magic
tech sky130A
magscale 1 2
timestamp 1607490450
<< locali >>
rect 75653 694195 75687 698309
rect 10793 676243 10827 685797
rect 140513 676243 140547 685797
rect 205557 684539 205591 694093
rect 270325 685899 270359 695453
rect 75561 656931 75595 666485
rect 85773 38675 85807 43469
rect 168757 38675 168791 48229
rect 109417 29019 109451 38573
rect 124321 29019 124355 38573
rect 197461 31603 197495 38573
rect 200497 31603 200531 42041
rect 203165 29019 203199 38573
rect 62313 19363 62347 28917
rect 291025 27659 291059 37145
rect 291393 29019 291427 38573
rect 293969 37315 294003 46869
rect 489653 38675 489687 48161
rect 487169 29019 487203 38573
rect 74733 19363 74767 22321
rect 147781 9707 147815 19261
rect 150817 9707 150851 22117
rect 203165 11747 203199 19261
rect 293969 18003 294003 27557
rect 438133 19363 438167 28917
rect 487169 9707 487203 19261
rect 499589 4743 499623 4981
rect 509157 4743 509191 4981
rect 518909 4743 518943 4981
rect 528477 4743 528511 4981
rect 59921 3179 59955 3417
rect 63509 3111 63543 3553
rect 95617 3383 95651 3689
rect 113833 3179 113867 3485
rect 121745 3179 121779 3553
rect 147873 3451 147907 3757
rect 162133 3383 162167 3757
rect 200773 3723 200807 4097
rect 171609 3247 171643 3621
rect 207213 3179 207247 4097
rect 209789 3791 209823 4097
rect 208501 3111 208535 3621
rect 213929 3519 213963 3893
rect 215401 3859 215435 3961
rect 221013 3791 221047 3961
rect 229109 3723 229143 3961
rect 231133 3587 231167 3689
rect 468987 3553 469321 3587
rect 495449 3383 495483 3893
<< viali >>
rect 75653 698309 75687 698343
rect 75653 694161 75687 694195
rect 270325 695453 270359 695487
rect 205557 694093 205591 694127
rect 10793 685797 10827 685831
rect 10793 676209 10827 676243
rect 140513 685797 140547 685831
rect 270325 685865 270359 685899
rect 205557 684505 205591 684539
rect 140513 676209 140547 676243
rect 75561 666485 75595 666519
rect 75561 656897 75595 656931
rect 168757 48229 168791 48263
rect 85773 43469 85807 43503
rect 85773 38641 85807 38675
rect 489653 48161 489687 48195
rect 293969 46869 294003 46903
rect 168757 38641 168791 38675
rect 200497 42041 200531 42075
rect 109417 38573 109451 38607
rect 109417 28985 109451 29019
rect 124321 38573 124355 38607
rect 197461 38573 197495 38607
rect 197461 31569 197495 31603
rect 200497 31569 200531 31603
rect 203165 38573 203199 38607
rect 124321 28985 124355 29019
rect 291393 38573 291427 38607
rect 203165 28985 203199 29019
rect 291025 37145 291059 37179
rect 62313 28917 62347 28951
rect 489653 38641 489687 38675
rect 293969 37281 294003 37315
rect 487169 38573 487203 38607
rect 291393 28985 291427 29019
rect 487169 28985 487203 29019
rect 291025 27625 291059 27659
rect 438133 28917 438167 28951
rect 293969 27557 294003 27591
rect 62313 19329 62347 19363
rect 74733 22321 74767 22355
rect 74733 19329 74767 19363
rect 150817 22117 150851 22151
rect 147781 19261 147815 19295
rect 147781 9673 147815 9707
rect 203165 19261 203199 19295
rect 438133 19329 438167 19363
rect 293969 17969 294003 18003
rect 487169 19261 487203 19295
rect 203165 11713 203199 11747
rect 150817 9673 150851 9707
rect 487169 9673 487203 9707
rect 499589 4981 499623 5015
rect 499589 4709 499623 4743
rect 509157 4981 509191 5015
rect 509157 4709 509191 4743
rect 518909 4981 518943 5015
rect 518909 4709 518943 4743
rect 528477 4981 528511 5015
rect 528477 4709 528511 4743
rect 200773 4097 200807 4131
rect 147873 3757 147907 3791
rect 95617 3689 95651 3723
rect 63509 3553 63543 3587
rect 59921 3417 59955 3451
rect 59921 3145 59955 3179
rect 121745 3553 121779 3587
rect 95617 3349 95651 3383
rect 113833 3485 113867 3519
rect 113833 3145 113867 3179
rect 147873 3417 147907 3451
rect 162133 3757 162167 3791
rect 200773 3689 200807 3723
rect 207213 4097 207247 4131
rect 162133 3349 162167 3383
rect 171609 3621 171643 3655
rect 171609 3213 171643 3247
rect 121745 3145 121779 3179
rect 209789 4097 209823 4131
rect 215401 3961 215435 3995
rect 209789 3757 209823 3791
rect 213929 3893 213963 3927
rect 207213 3145 207247 3179
rect 208501 3621 208535 3655
rect 63509 3077 63543 3111
rect 215401 3825 215435 3859
rect 221013 3961 221047 3995
rect 221013 3757 221047 3791
rect 229109 3961 229143 3995
rect 495449 3893 495483 3927
rect 229109 3689 229143 3723
rect 231133 3689 231167 3723
rect 231133 3553 231167 3587
rect 468953 3553 468987 3587
rect 469321 3553 469355 3587
rect 213929 3485 213963 3519
rect 495449 3349 495483 3383
rect 208501 3077 208535 3111
<< metal1 >>
rect 54018 700816 54024 700868
rect 54076 700856 54082 700868
rect 55122 700856 55128 700868
rect 54076 700828 55128 700856
rect 54076 700816 54082 700828
rect 55122 700816 55128 700828
rect 55180 700816 55186 700868
rect 429102 700408 429108 700460
rect 429160 700448 429166 700460
rect 464982 700448 464988 700460
rect 429160 700420 464988 700448
rect 429160 700408 429166 700420
rect 464982 700408 464988 700420
rect 465040 700408 465046 700460
rect 480162 700408 480168 700460
rect 480220 700448 480226 700460
rect 529842 700448 529848 700460
rect 480220 700420 529848 700448
rect 480220 700408 480226 700420
rect 529842 700408 529848 700420
rect 529900 700408 529906 700460
rect 360102 700340 360108 700392
rect 360160 700380 360166 700392
rect 378410 700380 378416 700392
rect 360160 700352 378416 700380
rect 360160 700340 360166 700352
rect 378410 700340 378416 700352
rect 378468 700340 378474 700392
rect 394602 700340 394608 700392
rect 394660 700380 394666 700392
rect 421742 700380 421748 700392
rect 394660 700352 421748 700380
rect 394660 700340 394666 700352
rect 421742 700340 421748 700352
rect 421800 700340 421806 700392
rect 445662 700340 445668 700392
rect 445720 700380 445726 700392
rect 486602 700380 486608 700392
rect 445720 700352 486608 700380
rect 445720 700340 445726 700352
rect 486602 700340 486608 700352
rect 486660 700340 486666 700392
rect 496722 700340 496728 700392
rect 496780 700380 496786 700392
rect 551462 700380 551468 700392
rect 496780 700352 551468 700380
rect 496780 700340 496786 700352
rect 551462 700340 551468 700352
rect 551520 700340 551526 700392
rect 343542 700272 343548 700324
rect 343600 700312 343606 700324
rect 356790 700312 356796 700324
rect 343600 700284 356796 700312
rect 343600 700272 343606 700284
rect 356790 700272 356796 700284
rect 356848 700272 356854 700324
rect 378042 700272 378048 700324
rect 378100 700312 378106 700324
rect 400122 700312 400128 700324
rect 378100 700284 400128 700312
rect 378100 700272 378106 700284
rect 400122 700272 400128 700284
rect 400180 700272 400186 700324
rect 411162 700272 411168 700324
rect 411220 700312 411226 700324
rect 443362 700312 443368 700324
rect 411220 700284 443368 700312
rect 411220 700272 411226 700284
rect 443362 700272 443368 700284
rect 443420 700272 443426 700324
rect 463602 700272 463608 700324
rect 463660 700312 463666 700324
rect 508222 700312 508228 700324
rect 463660 700284 508228 700312
rect 463660 700272 463666 700284
rect 508222 700272 508228 700284
rect 508280 700272 508286 700324
rect 514662 700272 514668 700324
rect 514720 700312 514726 700324
rect 573082 700312 573088 700324
rect 514720 700284 573088 700312
rect 514720 700272 514726 700284
rect 573082 700272 573088 700284
rect 573140 700272 573146 700324
rect 183738 700136 183744 700188
rect 183796 700176 183802 700188
rect 184842 700176 184848 700188
rect 183796 700148 184848 700176
rect 183796 700136 183802 700148
rect 184842 700136 184848 700148
rect 184900 700136 184906 700188
rect 32398 699660 32404 699712
rect 32456 699700 32462 699712
rect 33042 699700 33048 699712
rect 32456 699672 33048 699700
rect 32456 699660 32462 699672
rect 33042 699660 33048 699672
rect 33100 699660 33106 699712
rect 97258 699660 97264 699712
rect 97316 699700 97322 699712
rect 97902 699700 97908 699712
rect 97316 699672 97908 699700
rect 97316 699660 97322 699672
rect 97902 699660 97908 699672
rect 97960 699660 97966 699712
rect 118878 699660 118884 699712
rect 118936 699700 118942 699712
rect 119982 699700 119988 699712
rect 118936 699672 119988 699700
rect 118936 699660 118942 699672
rect 119982 699660 119988 699672
rect 120040 699660 120046 699712
rect 162118 699660 162124 699712
rect 162176 699700 162182 699712
rect 162762 699700 162768 699712
rect 162176 699672 162768 699700
rect 162176 699660 162182 699672
rect 162762 699660 162768 699672
rect 162820 699660 162826 699712
rect 227070 699660 227076 699712
rect 227128 699700 227134 699712
rect 227622 699700 227628 699712
rect 227128 699672 227628 699700
rect 227128 699660 227134 699672
rect 227622 699660 227628 699672
rect 227680 699660 227686 699712
rect 248690 699660 248696 699712
rect 248748 699700 248754 699712
rect 249702 699700 249708 699712
rect 248748 699672 249708 699700
rect 248748 699660 248754 699672
rect 249702 699660 249708 699672
rect 249760 699660 249766 699712
rect 291194 699660 291200 699712
rect 291252 699700 291258 699712
rect 291930 699700 291936 699712
rect 291252 699672 291936 699700
rect 291252 699660 291258 699672
rect 291930 699660 291936 699672
rect 291988 699660 291994 699712
rect 309042 699660 309048 699712
rect 309100 699700 309106 699712
rect 313550 699700 313556 699712
rect 309100 699672 313556 699700
rect 309100 699660 309106 699672
rect 313550 699660 313556 699672
rect 313608 699660 313614 699712
rect 326982 699660 326988 699712
rect 327040 699700 327046 699712
rect 335170 699700 335176 699712
rect 327040 699672 335176 699700
rect 327040 699660 327046 699672
rect 335170 699660 335176 699672
rect 335228 699660 335234 699712
rect 75638 698340 75644 698352
rect 75599 698312 75644 698340
rect 75638 698300 75644 698312
rect 75696 698300 75702 698352
rect 10686 695512 10692 695564
rect 10744 695552 10750 695564
rect 10778 695552 10784 695564
rect 10744 695524 10784 695552
rect 10744 695512 10750 695524
rect 10778 695512 10784 695524
rect 10836 695512 10842 695564
rect 140406 695512 140412 695564
rect 140464 695552 140470 695564
rect 140498 695552 140504 695564
rect 140464 695524 140504 695552
rect 140464 695512 140470 695524
rect 140498 695512 140504 695524
rect 140556 695512 140562 695564
rect 523678 695512 523684 695564
rect 523736 695552 523742 695564
rect 580166 695552 580172 695564
rect 523736 695524 580172 695552
rect 523736 695512 523742 695524
rect 580166 695512 580172 695524
rect 580224 695512 580230 695564
rect 270313 695487 270371 695493
rect 270313 695453 270325 695487
rect 270359 695484 270371 695487
rect 270402 695484 270408 695496
rect 270359 695456 270408 695484
rect 270359 695453 270371 695456
rect 270313 695447 270371 695453
rect 270402 695444 270408 695456
rect 270460 695444 270466 695496
rect 75638 694192 75644 694204
rect 75599 694164 75644 694192
rect 75638 694152 75644 694164
rect 75696 694152 75702 694204
rect 205545 694127 205603 694133
rect 205545 694093 205557 694127
rect 205591 694124 205603 694127
rect 205634 694124 205640 694136
rect 205591 694096 205640 694124
rect 205591 694093 205603 694096
rect 205545 694087 205603 694093
rect 205634 694084 205640 694096
rect 205692 694084 205698 694136
rect 75638 688684 75644 688696
rect 75564 688656 75644 688684
rect 75564 688628 75592 688656
rect 75638 688644 75644 688656
rect 75696 688644 75702 688696
rect 10686 688576 10692 688628
rect 10744 688616 10750 688628
rect 10870 688616 10876 688628
rect 10744 688588 10876 688616
rect 10744 688576 10750 688588
rect 10870 688576 10876 688588
rect 10928 688576 10934 688628
rect 75546 688576 75552 688628
rect 75604 688576 75610 688628
rect 140406 688576 140412 688628
rect 140464 688616 140470 688628
rect 140590 688616 140596 688628
rect 140464 688588 140596 688616
rect 140464 688576 140470 688588
rect 140590 688576 140596 688588
rect 140648 688576 140654 688628
rect 270310 685896 270316 685908
rect 270271 685868 270316 685896
rect 270310 685856 270316 685868
rect 270368 685856 270374 685908
rect 10781 685831 10839 685837
rect 10781 685797 10793 685831
rect 10827 685828 10839 685831
rect 10870 685828 10876 685840
rect 10827 685800 10876 685828
rect 10827 685797 10839 685800
rect 10781 685791 10839 685797
rect 10870 685788 10876 685800
rect 10928 685788 10934 685840
rect 140501 685831 140559 685837
rect 140501 685797 140513 685831
rect 140547 685828 140559 685831
rect 140590 685828 140596 685840
rect 140547 685800 140596 685828
rect 140547 685797 140559 685800
rect 140501 685791 140559 685797
rect 140590 685788 140596 685800
rect 140648 685788 140654 685840
rect 205542 684536 205548 684548
rect 205503 684508 205548 684536
rect 205542 684496 205548 684508
rect 205600 684496 205606 684548
rect 523770 680348 523776 680400
rect 523828 680388 523834 680400
rect 580166 680388 580172 680400
rect 523828 680360 580172 680388
rect 523828 680348 523834 680360
rect 580166 680348 580172 680360
rect 580224 680348 580230 680400
rect 75546 679028 75552 679040
rect 75472 679000 75552 679028
rect 75472 678972 75500 679000
rect 75546 678988 75552 679000
rect 75604 678988 75610 679040
rect 205542 679028 205548 679040
rect 205468 679000 205548 679028
rect 205468 678972 205496 679000
rect 205542 678988 205548 679000
rect 205600 678988 205606 679040
rect 270310 679028 270316 679040
rect 270236 679000 270316 679028
rect 270236 678972 270264 679000
rect 270310 678988 270316 679000
rect 270368 678988 270374 679040
rect 75454 678920 75460 678972
rect 75512 678920 75518 678972
rect 205450 678920 205456 678972
rect 205508 678920 205514 678972
rect 270218 678920 270224 678972
rect 270276 678920 270282 678972
rect 10778 676240 10784 676252
rect 10739 676212 10784 676240
rect 10778 676200 10784 676212
rect 10836 676200 10842 676252
rect 140498 676240 140504 676252
rect 140459 676212 140504 676240
rect 140498 676200 140504 676212
rect 140556 676200 140562 676252
rect 10778 673480 10784 673532
rect 10836 673520 10842 673532
rect 10962 673520 10968 673532
rect 10836 673492 10968 673520
rect 10836 673480 10842 673492
rect 10962 673480 10968 673492
rect 11020 673480 11026 673532
rect 140498 673480 140504 673532
rect 140556 673520 140562 673532
rect 140682 673520 140688 673532
rect 140556 673492 140688 673520
rect 140556 673480 140562 673492
rect 140682 673480 140688 673492
rect 140740 673480 140746 673532
rect 270218 673480 270224 673532
rect 270276 673520 270282 673532
rect 270402 673520 270408 673532
rect 270276 673492 270408 673520
rect 270276 673480 270282 673492
rect 270402 673480 270408 673492
rect 270460 673480 270466 673532
rect 205450 669372 205456 669384
rect 205376 669344 205456 669372
rect 205376 669316 205404 669344
rect 205450 669332 205456 669344
rect 205508 669332 205514 669384
rect 75454 669264 75460 669316
rect 75512 669304 75518 669316
rect 75638 669304 75644 669316
rect 75512 669276 75644 669304
rect 75512 669264 75518 669276
rect 75638 669264 75644 669276
rect 75696 669264 75702 669316
rect 205358 669264 205364 669316
rect 205416 669264 205422 669316
rect 75549 666519 75607 666525
rect 75549 666485 75561 666519
rect 75595 666516 75607 666519
rect 75638 666516 75644 666528
rect 75595 666488 75644 666516
rect 75595 666485 75607 666488
rect 75549 666479 75607 666485
rect 75638 666476 75644 666488
rect 75696 666476 75702 666528
rect 205358 659716 205364 659728
rect 205284 659688 205364 659716
rect 205284 659660 205312 659688
rect 205358 659676 205364 659688
rect 205416 659676 205422 659728
rect 205266 659608 205272 659660
rect 205324 659608 205330 659660
rect 75546 656928 75552 656940
rect 75507 656900 75552 656928
rect 75546 656888 75552 656900
rect 75604 656888 75610 656940
rect 249702 655460 249708 655512
rect 249760 655500 249766 655512
rect 257890 655500 257896 655512
rect 249760 655472 257896 655500
rect 249760 655460 249766 655472
rect 257890 655460 257896 655472
rect 257948 655460 257954 655512
rect 270218 655460 270224 655512
rect 270276 655500 270282 655512
rect 274910 655500 274916 655512
rect 270276 655472 274916 655500
rect 270276 655460 270282 655472
rect 274910 655460 274916 655472
rect 274968 655460 274974 655512
rect 377122 655460 377128 655512
rect 377180 655500 377186 655512
rect 378042 655500 378048 655512
rect 377180 655472 378048 655500
rect 377180 655460 377186 655472
rect 378042 655460 378048 655472
rect 378100 655460 378106 655512
rect 428182 655460 428188 655512
rect 428240 655500 428246 655512
rect 429102 655500 429108 655512
rect 428240 655472 429108 655500
rect 428240 655460 428246 655472
rect 429102 655460 429108 655472
rect 429160 655460 429166 655512
rect 462314 655460 462320 655512
rect 462372 655500 462378 655512
rect 463602 655500 463608 655512
rect 462372 655472 463608 655500
rect 462372 655460 462378 655472
rect 463602 655460 463608 655472
rect 463660 655460 463666 655512
rect 479334 655460 479340 655512
rect 479392 655500 479398 655512
rect 480162 655500 480168 655512
rect 479392 655472 480168 655500
rect 479392 655460 479398 655472
rect 480162 655460 480168 655472
rect 480220 655460 480226 655512
rect 513374 655256 513380 655308
rect 513432 655296 513438 655308
rect 514662 655296 514668 655308
rect 513432 655268 514668 655296
rect 513432 655256 513438 655268
rect 514662 655256 514668 655268
rect 514720 655256 514726 655308
rect 325970 655120 325976 655172
rect 326028 655160 326034 655172
rect 326982 655160 326988 655172
rect 326028 655132 326988 655160
rect 326028 655120 326034 655132
rect 326982 655120 326988 655132
rect 327040 655120 327046 655172
rect 55122 654916 55128 654968
rect 55180 654956 55186 654968
rect 104526 654956 104532 654968
rect 55180 654928 104532 654956
rect 55180 654916 55186 654928
rect 104526 654916 104532 654928
rect 104584 654916 104590 654968
rect 119982 654916 119988 654968
rect 120040 654956 120046 654968
rect 155586 654956 155592 654968
rect 120040 654928 155592 654956
rect 120040 654916 120046 654928
rect 155586 654916 155592 654928
rect 155644 654916 155650 654968
rect 33042 654848 33048 654900
rect 33100 654888 33106 654900
rect 87506 654888 87512 654900
rect 33100 654860 87512 654888
rect 33100 654848 33106 654860
rect 87506 654848 87512 654860
rect 87564 654848 87570 654900
rect 97902 654848 97908 654900
rect 97960 654888 97966 654900
rect 138566 654888 138572 654900
rect 97960 654860 138572 654888
rect 97960 654848 97966 654860
rect 138566 654848 138572 654860
rect 138624 654848 138630 654900
rect 162762 654848 162768 654900
rect 162820 654888 162826 654900
rect 189718 654888 189724 654900
rect 162820 654860 189724 654888
rect 162820 654848 162826 654860
rect 189718 654848 189724 654860
rect 189776 654848 189782 654900
rect 205266 654848 205272 654900
rect 205324 654888 205330 654900
rect 223758 654888 223764 654900
rect 205324 654860 223764 654888
rect 205324 654848 205330 654860
rect 223758 654848 223764 654860
rect 223816 654848 223822 654900
rect 10778 654780 10784 654832
rect 10836 654820 10842 654832
rect 70486 654820 70492 654832
rect 10836 654792 70492 654820
rect 10836 654780 10842 654792
rect 70486 654780 70492 654792
rect 70544 654780 70550 654832
rect 75546 654780 75552 654832
rect 75604 654820 75610 654832
rect 121546 654820 121552 654832
rect 75604 654792 121552 654820
rect 75604 654780 75610 654792
rect 121546 654780 121552 654792
rect 121604 654780 121610 654832
rect 140498 654780 140504 654832
rect 140556 654820 140562 654832
rect 172698 654820 172704 654832
rect 140556 654792 172704 654820
rect 140556 654780 140562 654792
rect 172698 654780 172704 654792
rect 172756 654780 172762 654832
rect 184842 654780 184848 654832
rect 184900 654820 184906 654832
rect 206738 654820 206744 654832
rect 184900 654792 206744 654820
rect 184900 654780 184906 654792
rect 206738 654780 206744 654792
rect 206796 654780 206802 654832
rect 227622 654780 227628 654832
rect 227680 654820 227686 654832
rect 240778 654820 240784 654832
rect 227680 654792 240784 654820
rect 227680 654780 227686 654792
rect 240778 654780 240784 654792
rect 240836 654780 240842 654832
rect 3418 645804 3424 645856
rect 3476 645844 3482 645856
rect 59354 645844 59360 645856
rect 3476 645816 59360 645844
rect 3476 645804 3482 645816
rect 59354 645804 59360 645816
rect 59412 645804 59418 645856
rect 523678 633428 523684 633480
rect 523736 633468 523742 633480
rect 580166 633468 580172 633480
rect 523736 633440 580172 633468
rect 523736 633428 523742 633440
rect 580166 633428 580172 633440
rect 580224 633428 580230 633480
rect 3510 630572 3516 630624
rect 3568 630612 3574 630624
rect 59354 630612 59360 630624
rect 3568 630584 59360 630612
rect 3568 630572 3574 630584
rect 59354 630572 59360 630584
rect 59412 630572 59418 630624
rect 524322 619556 524328 619608
rect 524380 619596 524386 619608
rect 580258 619596 580264 619608
rect 524380 619568 580264 619596
rect 524380 619556 524386 619568
rect 580258 619556 580264 619568
rect 580316 619556 580322 619608
rect 3602 616768 3608 616820
rect 3660 616808 3666 616820
rect 59354 616808 59360 616820
rect 3660 616780 59360 616808
rect 3660 616768 3666 616780
rect 59354 616768 59360 616780
rect 59412 616768 59418 616820
rect 523126 605752 523132 605804
rect 523184 605792 523190 605804
rect 580350 605792 580356 605804
rect 523184 605764 580356 605792
rect 523184 605752 523190 605764
rect 580350 605752 580356 605764
rect 580408 605752 580414 605804
rect 3694 603032 3700 603084
rect 3752 603072 3758 603084
rect 59354 603072 59360 603084
rect 3752 603044 59360 603072
rect 3752 603032 3758 603044
rect 59354 603032 59360 603044
rect 59412 603032 59418 603084
rect 523770 601672 523776 601724
rect 523828 601712 523834 601724
rect 580166 601712 580172 601724
rect 523828 601684 580172 601712
rect 523828 601672 523834 601684
rect 580166 601672 580172 601684
rect 580224 601672 580230 601724
rect 3418 587800 3424 587852
rect 3476 587840 3482 587852
rect 59354 587840 59360 587852
rect 3476 587812 59360 587840
rect 3476 587800 3482 587812
rect 59354 587800 59360 587812
rect 59412 587800 59418 587852
rect 523678 586508 523684 586560
rect 523736 586548 523742 586560
rect 580166 586548 580172 586560
rect 523736 586520 580172 586548
rect 523736 586508 523742 586520
rect 580166 586508 580172 586520
rect 580224 586508 580230 586560
rect 524322 579572 524328 579624
rect 524380 579612 524386 579624
rect 580258 579612 580264 579624
rect 524380 579584 580264 579612
rect 524380 579572 524386 579584
rect 580258 579572 580264 579584
rect 580316 579572 580322 579624
rect 3510 573996 3516 574048
rect 3568 574036 3574 574048
rect 59354 574036 59360 574048
rect 3568 574008 59360 574036
rect 3568 573996 3574 574008
rect 59354 573996 59360 574008
rect 59412 573996 59418 574048
rect 3602 560192 3608 560244
rect 3660 560232 3666 560244
rect 59354 560232 59360 560244
rect 3660 560204 59360 560232
rect 3660 560192 3666 560204
rect 59354 560192 59360 560204
rect 59412 560192 59418 560244
rect 523770 554752 523776 554804
rect 523828 554792 523834 554804
rect 580166 554792 580172 554804
rect 523828 554764 580172 554792
rect 523828 554752 523834 554764
rect 580166 554752 580172 554764
rect 580224 554752 580230 554804
rect 3418 545028 3424 545080
rect 3476 545068 3482 545080
rect 59354 545068 59360 545080
rect 3476 545040 59360 545068
rect 3476 545028 3482 545040
rect 59354 545028 59360 545040
rect 59412 545028 59418 545080
rect 523494 539588 523500 539640
rect 523552 539628 523558 539640
rect 580166 539628 580172 539640
rect 523552 539600 580172 539628
rect 523552 539588 523558 539600
rect 580166 539588 580172 539600
rect 580224 539588 580230 539640
rect 523678 539520 523684 539572
rect 523736 539560 523742 539572
rect 580258 539560 580264 539572
rect 523736 539532 580264 539560
rect 523736 539520 523742 539532
rect 580258 539520 580264 539532
rect 580316 539520 580322 539572
rect 3510 531224 3516 531276
rect 3568 531264 3574 531276
rect 59354 531264 59360 531276
rect 3568 531236 59360 531264
rect 3568 531224 3574 531236
rect 59354 531224 59360 531236
rect 59412 531224 59418 531276
rect 523770 522996 523776 523048
rect 523828 523036 523834 523048
rect 580166 523036 580172 523048
rect 523828 523008 580172 523036
rect 523828 522996 523834 523008
rect 580166 522996 580172 523008
rect 580224 522996 580230 523048
rect 3602 517420 3608 517472
rect 3660 517460 3666 517472
rect 59354 517460 59360 517472
rect 3660 517432 59360 517460
rect 3660 517420 3666 517432
rect 59354 517420 59360 517432
rect 59412 517420 59418 517472
rect 523678 507832 523684 507884
rect 523736 507872 523742 507884
rect 580166 507872 580172 507884
rect 523736 507844 580172 507872
rect 523736 507832 523742 507844
rect 580166 507832 580172 507844
rect 580224 507832 580230 507884
rect 3418 502256 3424 502308
rect 3476 502296 3482 502308
rect 59354 502296 59360 502308
rect 3476 502268 59360 502296
rect 3476 502256 3482 502268
rect 59354 502256 59360 502268
rect 59412 502256 59418 502308
rect 523770 492668 523776 492720
rect 523828 492708 523834 492720
rect 580166 492708 580172 492720
rect 523828 492680 580172 492708
rect 523828 492668 523834 492680
rect 580166 492668 580172 492680
rect 580224 492668 580230 492720
rect 3510 488452 3516 488504
rect 3568 488492 3574 488504
rect 59354 488492 59360 488504
rect 3568 488464 59360 488492
rect 3568 488452 3574 488464
rect 59354 488452 59360 488464
rect 59412 488452 59418 488504
rect 523678 476076 523684 476128
rect 523736 476116 523742 476128
rect 580166 476116 580172 476128
rect 523736 476088 580172 476116
rect 523736 476076 523742 476088
rect 580166 476076 580172 476088
rect 580224 476076 580230 476128
rect 3418 474648 3424 474700
rect 3476 474688 3482 474700
rect 59354 474688 59360 474700
rect 3476 474660 59360 474688
rect 3476 474648 3482 474660
rect 59354 474648 59360 474660
rect 59412 474648 59418 474700
rect 523770 460912 523776 460964
rect 523828 460952 523834 460964
rect 580166 460952 580172 460964
rect 523828 460924 580172 460952
rect 523828 460912 523834 460924
rect 580166 460912 580172 460924
rect 580224 460912 580230 460964
rect 3510 459484 3516 459536
rect 3568 459524 3574 459536
rect 59354 459524 59360 459536
rect 3568 459496 59360 459524
rect 3568 459484 3574 459496
rect 59354 459484 59360 459496
rect 59412 459484 59418 459536
rect 523678 445748 523684 445800
rect 523736 445788 523742 445800
rect 580166 445788 580172 445800
rect 523736 445760 580172 445788
rect 523736 445748 523742 445760
rect 580166 445748 580172 445760
rect 580224 445748 580230 445800
rect 3418 445680 3424 445732
rect 3476 445720 3482 445732
rect 59354 445720 59360 445732
rect 3476 445692 59360 445720
rect 3476 445680 3482 445692
rect 59354 445680 59360 445692
rect 59412 445680 59418 445732
rect 3418 430516 3424 430568
rect 3476 430556 3482 430568
rect 59354 430556 59360 430568
rect 3476 430528 59360 430556
rect 3476 430516 3482 430528
rect 59354 430516 59360 430528
rect 59412 430516 59418 430568
rect 523678 429156 523684 429208
rect 523736 429196 523742 429208
rect 580166 429196 580172 429208
rect 523736 429168 580172 429196
rect 523736 429156 523742 429168
rect 580166 429156 580172 429168
rect 580224 429156 580230 429208
rect 3418 416712 3424 416764
rect 3476 416752 3482 416764
rect 59354 416752 59360 416764
rect 3476 416724 59360 416752
rect 3476 416712 3482 416724
rect 59354 416712 59360 416724
rect 59412 416712 59418 416764
rect 523678 413992 523684 414044
rect 523736 414032 523742 414044
rect 580166 414032 580172 414044
rect 523736 414004 580172 414032
rect 523736 413992 523742 414004
rect 580166 413992 580172 414004
rect 580224 413992 580230 414044
rect 3418 402908 3424 402960
rect 3476 402948 3482 402960
rect 59354 402948 59360 402960
rect 3476 402920 59360 402948
rect 3476 402908 3482 402920
rect 59354 402908 59360 402920
rect 59412 402908 59418 402960
rect 523678 398828 523684 398880
rect 523736 398868 523742 398880
rect 580166 398868 580172 398880
rect 523736 398840 580172 398868
rect 523736 398828 523742 398840
rect 580166 398828 580172 398840
rect 580224 398828 580230 398880
rect 3878 387744 3884 387796
rect 3936 387784 3942 387796
rect 59354 387784 59360 387796
rect 3936 387756 59360 387784
rect 3936 387744 3942 387756
rect 59354 387744 59360 387756
rect 59412 387744 59418 387796
rect 523126 382236 523132 382288
rect 523184 382276 523190 382288
rect 580166 382276 580172 382288
rect 523184 382248 580172 382276
rect 523184 382236 523190 382248
rect 580166 382236 580172 382248
rect 580224 382236 580230 382288
rect 3418 373940 3424 373992
rect 3476 373980 3482 373992
rect 59354 373980 59360 373992
rect 3476 373952 59360 373980
rect 3476 373940 3482 373952
rect 59354 373940 59360 373952
rect 59412 373940 59418 373992
rect 523310 367072 523316 367124
rect 523368 367112 523374 367124
rect 580166 367112 580172 367124
rect 523368 367084 580172 367112
rect 523368 367072 523374 367084
rect 580166 367072 580172 367084
rect 580224 367072 580230 367124
rect 3418 360136 3424 360188
rect 3476 360176 3482 360188
rect 59354 360176 59360 360188
rect 3476 360148 59360 360176
rect 3476 360136 3482 360148
rect 59354 360136 59360 360148
rect 59412 360136 59418 360188
rect 524322 352520 524328 352572
rect 524380 352560 524386 352572
rect 580166 352560 580172 352572
rect 524380 352532 580172 352560
rect 524380 352520 524386 352532
rect 580166 352520 580172 352532
rect 580224 352520 580230 352572
rect 3418 343544 3424 343596
rect 3476 343584 3482 343596
rect 59354 343584 59360 343596
rect 3476 343556 59360 343584
rect 3476 343544 3482 343556
rect 59354 343544 59360 343556
rect 59412 343544 59418 343596
rect 523402 336676 523408 336728
rect 523460 336716 523466 336728
rect 580166 336716 580172 336728
rect 523460 336688 580172 336716
rect 523460 336676 523466 336688
rect 580166 336676 580172 336688
rect 580224 336676 580230 336728
rect 3326 327020 3332 327072
rect 3384 327060 3390 327072
rect 59354 327060 59360 327072
rect 3384 327032 59360 327060
rect 3384 327020 3390 327032
rect 59354 327020 59360 327032
rect 59412 327020 59418 327072
rect 523126 321512 523132 321564
rect 523184 321552 523190 321564
rect 580166 321552 580172 321564
rect 523184 321524 580172 321552
rect 523184 321512 523190 321524
rect 580166 321512 580172 321524
rect 580224 321512 580230 321564
rect 3418 310428 3424 310480
rect 3476 310468 3482 310480
rect 59998 310468 60004 310480
rect 3476 310440 60004 310468
rect 3476 310428 3482 310440
rect 59998 310428 60004 310440
rect 60056 310428 60062 310480
rect 523678 306280 523684 306332
rect 523736 306320 523742 306332
rect 580166 306320 580172 306332
rect 523736 306292 580172 306320
rect 523736 306280 523742 306292
rect 580166 306280 580172 306292
rect 580224 306280 580230 306332
rect 3142 293904 3148 293956
rect 3200 293944 3206 293956
rect 59998 293944 60004 293956
rect 3200 293916 60004 293944
rect 3200 293904 3206 293916
rect 59998 293904 60004 293916
rect 60056 293904 60062 293956
rect 523678 289756 523684 289808
rect 523736 289796 523742 289808
rect 580166 289796 580172 289808
rect 523736 289768 580172 289796
rect 523736 289756 523742 289768
rect 580166 289756 580172 289768
rect 580224 289756 580230 289808
rect 3418 277312 3424 277364
rect 3476 277352 3482 277364
rect 59998 277352 60004 277364
rect 3476 277324 60004 277352
rect 3476 277312 3482 277324
rect 59998 277312 60004 277324
rect 60056 277312 60062 277364
rect 523678 274592 523684 274644
rect 523736 274632 523742 274644
rect 580166 274632 580172 274644
rect 523736 274604 580172 274632
rect 523736 274592 523742 274604
rect 580166 274592 580172 274604
rect 580224 274592 580230 274644
rect 3418 260788 3424 260840
rect 3476 260828 3482 260840
rect 59998 260828 60004 260840
rect 3476 260800 60004 260828
rect 3476 260788 3482 260800
rect 59998 260788 60004 260800
rect 60056 260788 60062 260840
rect 523678 259360 523684 259412
rect 523736 259400 523742 259412
rect 580166 259400 580172 259412
rect 523736 259372 580172 259400
rect 523736 259360 523742 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3418 244196 3424 244248
rect 3476 244236 3482 244248
rect 59998 244236 60004 244248
rect 3476 244208 60004 244236
rect 3476 244196 3482 244208
rect 59998 244196 60004 244208
rect 60056 244196 60062 244248
rect 523770 242836 523776 242888
rect 523828 242876 523834 242888
rect 580166 242876 580172 242888
rect 523828 242848 580172 242876
rect 523828 242836 523834 242848
rect 580166 242836 580172 242848
rect 580224 242836 580230 242888
rect 523678 227672 523684 227724
rect 523736 227712 523742 227724
rect 580166 227712 580172 227724
rect 523736 227684 580172 227712
rect 523736 227672 523742 227684
rect 580166 227672 580172 227684
rect 580224 227672 580230 227724
rect 3418 226244 3424 226296
rect 3476 226284 3482 226296
rect 60090 226284 60096 226296
rect 3476 226256 60096 226284
rect 3476 226244 3482 226256
rect 60090 226244 60096 226256
rect 60148 226244 60154 226296
rect 523770 212440 523776 212492
rect 523828 212480 523834 212492
rect 580166 212480 580172 212492
rect 523828 212452 580172 212480
rect 523828 212440 523834 212452
rect 580166 212440 580172 212452
rect 580224 212440 580230 212492
rect 3418 209720 3424 209772
rect 3476 209760 3482 209772
rect 59998 209760 60004 209772
rect 3476 209732 60004 209760
rect 3476 209720 3482 209732
rect 59998 209720 60004 209732
rect 60056 209720 60062 209772
rect 523678 195916 523684 195968
rect 523736 195956 523742 195968
rect 580166 195956 580172 195968
rect 523736 195928 580172 195956
rect 523736 195916 523742 195928
rect 580166 195916 580172 195928
rect 580224 195916 580230 195968
rect 3510 193128 3516 193180
rect 3568 193168 3574 193180
rect 60090 193168 60096 193180
rect 3568 193140 60096 193168
rect 3568 193128 3574 193140
rect 60090 193128 60096 193140
rect 60148 193128 60154 193180
rect 523770 180752 523776 180804
rect 523828 180792 523834 180804
rect 580166 180792 580172 180804
rect 523828 180764 580172 180792
rect 523828 180752 523834 180764
rect 580166 180752 580172 180764
rect 580224 180752 580230 180804
rect 3418 176604 3424 176656
rect 3476 176644 3482 176656
rect 59998 176644 60004 176656
rect 3476 176616 60004 176644
rect 3476 176604 3482 176616
rect 59998 176604 60004 176616
rect 60056 176604 60062 176656
rect 523678 165520 523684 165572
rect 523736 165560 523742 165572
rect 580166 165560 580172 165572
rect 523736 165532 580172 165560
rect 523736 165520 523742 165532
rect 580166 165520 580172 165532
rect 580224 165520 580230 165572
rect 3142 160012 3148 160064
rect 3200 160052 3206 160064
rect 60182 160052 60188 160064
rect 3200 160024 60188 160052
rect 3200 160012 3206 160024
rect 60182 160012 60188 160024
rect 60240 160012 60246 160064
rect 523862 148996 523868 149048
rect 523920 149036 523926 149048
rect 580166 149036 580172 149048
rect 523920 149008 580172 149036
rect 523920 148996 523926 149008
rect 580166 148996 580172 149008
rect 580224 148996 580230 149048
rect 3234 143488 3240 143540
rect 3292 143528 3298 143540
rect 60090 143528 60096 143540
rect 3292 143500 60096 143528
rect 3292 143488 3298 143500
rect 60090 143488 60096 143500
rect 60148 143488 60154 143540
rect 523770 133832 523776 133884
rect 523828 133872 523834 133884
rect 580166 133872 580172 133884
rect 523828 133844 580172 133872
rect 523828 133832 523834 133844
rect 580166 133832 580172 133844
rect 580224 133832 580230 133884
rect 3234 126896 3240 126948
rect 3292 126936 3298 126948
rect 59998 126936 60004 126948
rect 3292 126908 60004 126936
rect 3292 126896 3298 126908
rect 59998 126896 60004 126908
rect 60056 126896 60062 126948
rect 523678 118600 523684 118652
rect 523736 118640 523742 118652
rect 580166 118640 580172 118652
rect 523736 118612 580172 118640
rect 523736 118600 523742 118612
rect 580166 118600 580172 118612
rect 580224 118600 580230 118652
rect 3418 108944 3424 108996
rect 3476 108984 3482 108996
rect 60182 108984 60188 108996
rect 3476 108956 60188 108984
rect 3476 108944 3482 108956
rect 60182 108944 60188 108956
rect 60240 108944 60246 108996
rect 523862 102076 523868 102128
rect 523920 102116 523926 102128
rect 580166 102116 580172 102128
rect 523920 102088 580172 102116
rect 523920 102076 523926 102088
rect 580166 102076 580172 102088
rect 580224 102076 580230 102128
rect 3326 92420 3332 92472
rect 3384 92460 3390 92472
rect 60090 92460 60096 92472
rect 3384 92432 60096 92460
rect 3384 92420 3390 92432
rect 60090 92420 60096 92432
rect 60148 92420 60154 92472
rect 523770 86912 523776 86964
rect 523828 86952 523834 86964
rect 580166 86952 580172 86964
rect 523828 86924 580172 86952
rect 523828 86912 523834 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3418 75828 3424 75880
rect 3476 75868 3482 75880
rect 59998 75868 60004 75880
rect 3476 75840 60004 75868
rect 3476 75828 3482 75840
rect 59998 75828 60004 75840
rect 60056 75828 60062 75880
rect 523678 71680 523684 71732
rect 523736 71720 523742 71732
rect 580166 71720 580172 71732
rect 523736 71692 580172 71720
rect 523736 71680 523742 71692
rect 580166 71680 580172 71692
rect 580224 71680 580230 71732
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 60274 59344 60280 59356
rect 3108 59316 60280 59344
rect 3108 59304 3114 59316
rect 60274 59304 60280 59316
rect 60332 59304 60338 59356
rect 523954 55156 523960 55208
rect 524012 55196 524018 55208
rect 580166 55196 580172 55208
rect 524012 55168 580172 55196
rect 524012 55156 524018 55168
rect 580166 55156 580172 55168
rect 580224 55156 580230 55208
rect 147766 51008 147772 51060
rect 147824 51048 147830 51060
rect 148042 51048 148048 51060
rect 147824 51020 148048 51048
rect 147824 51008 147830 51020
rect 148042 51008 148048 51020
rect 148100 51008 148106 51060
rect 209038 49648 209044 49700
rect 209096 49688 209102 49700
rect 209866 49688 209872 49700
rect 209096 49660 209872 49688
rect 209096 49648 209102 49660
rect 209866 49648 209872 49660
rect 209924 49648 209930 49700
rect 232498 49648 232504 49700
rect 232556 49688 232562 49700
rect 242710 49688 242716 49700
rect 232556 49660 242716 49688
rect 232556 49648 232562 49660
rect 242710 49648 242716 49660
rect 242768 49648 242774 49700
rect 245562 49648 245568 49700
rect 245620 49688 245626 49700
rect 254854 49688 254860 49700
rect 245620 49660 254860 49688
rect 245620 49648 245626 49660
rect 254854 49648 254860 49660
rect 254912 49648 254918 49700
rect 262122 49648 262128 49700
rect 262180 49688 262186 49700
rect 268010 49688 268016 49700
rect 262180 49660 268016 49688
rect 262180 49648 262186 49660
rect 268010 49648 268016 49660
rect 268068 49648 268074 49700
rect 275922 49648 275928 49700
rect 275980 49688 275986 49700
rect 279326 49688 279332 49700
rect 275980 49660 279332 49688
rect 275980 49648 275986 49660
rect 279326 49648 279332 49660
rect 279384 49648 279390 49700
rect 324314 49648 324320 49700
rect 324372 49688 324378 49700
rect 326338 49688 326344 49700
rect 324372 49660 326344 49688
rect 324372 49648 324378 49660
rect 326338 49648 326344 49660
rect 326396 49648 326402 49700
rect 450170 49648 450176 49700
rect 450228 49688 450234 49700
rect 451918 49688 451924 49700
rect 450228 49660 451924 49688
rect 450228 49648 450234 49660
rect 451918 49648 451924 49660
rect 451976 49648 451982 49700
rect 241422 49580 241428 49632
rect 241480 49620 241486 49632
rect 252094 49620 252100 49632
rect 241480 49592 252100 49620
rect 241480 49580 241486 49592
rect 252094 49580 252100 49592
rect 252152 49580 252158 49632
rect 257338 49580 257344 49632
rect 257396 49620 257402 49632
rect 262398 49620 262404 49632
rect 257396 49592 262404 49620
rect 257396 49580 257402 49592
rect 262398 49580 262404 49592
rect 262456 49580 262462 49632
rect 263410 49580 263416 49632
rect 263468 49620 263474 49632
rect 269942 49620 269948 49632
rect 263468 49592 269948 49620
rect 263468 49580 263474 49592
rect 269942 49580 269948 49592
rect 270000 49580 270006 49632
rect 274542 49580 274548 49632
rect 274600 49620 274606 49632
rect 278314 49620 278320 49632
rect 274600 49592 278320 49620
rect 274600 49580 274606 49592
rect 278314 49580 278320 49592
rect 278372 49580 278378 49632
rect 392854 49580 392860 49632
rect 392912 49620 392918 49632
rect 393958 49620 393964 49632
rect 392912 49592 393964 49620
rect 392912 49580 392918 49592
rect 393958 49580 393964 49592
rect 394016 49580 394022 49632
rect 237190 49512 237196 49564
rect 237248 49552 237254 49564
rect 248046 49552 248052 49564
rect 237248 49524 248052 49552
rect 237248 49512 237254 49524
rect 248046 49512 248052 49524
rect 248104 49512 248110 49564
rect 248322 49512 248328 49564
rect 248380 49552 248386 49564
rect 257706 49552 257712 49564
rect 248380 49524 257712 49552
rect 248380 49512 248386 49524
rect 257706 49512 257712 49524
rect 257764 49512 257770 49564
rect 219342 49444 219348 49496
rect 219400 49484 219406 49496
rect 234246 49484 234252 49496
rect 219400 49456 234252 49484
rect 219400 49444 219406 49456
rect 234246 49444 234252 49456
rect 234304 49444 234310 49496
rect 238662 49444 238668 49496
rect 238720 49484 238726 49496
rect 250162 49484 250168 49496
rect 238720 49456 250168 49484
rect 238720 49444 238726 49456
rect 250162 49444 250168 49456
rect 250220 49444 250226 49496
rect 255222 49444 255228 49496
rect 255280 49484 255286 49496
rect 263318 49484 263324 49496
rect 255280 49456 263324 49484
rect 255280 49444 255286 49456
rect 263318 49444 263324 49456
rect 263376 49444 263382 49496
rect 220722 49376 220728 49428
rect 220780 49416 220786 49428
rect 236086 49416 236092 49428
rect 220780 49388 236092 49416
rect 220780 49376 220786 49388
rect 236086 49376 236092 49388
rect 236144 49376 236150 49428
rect 237282 49376 237288 49428
rect 237340 49416 237346 49428
rect 249242 49416 249248 49428
rect 237340 49388 249248 49416
rect 237340 49376 237346 49388
rect 249242 49376 249248 49388
rect 249300 49376 249306 49428
rect 249702 49376 249708 49428
rect 249760 49416 249766 49428
rect 258626 49416 258632 49428
rect 249760 49388 258632 49416
rect 249760 49376 249766 49388
rect 258626 49376 258632 49388
rect 258684 49376 258690 49428
rect 64782 49308 64788 49360
rect 64840 49348 64846 49360
rect 113174 49348 113180 49360
rect 64840 49320 113180 49348
rect 64840 49308 64846 49320
rect 113174 49308 113180 49320
rect 113232 49308 113238 49360
rect 186222 49308 186228 49360
rect 186280 49348 186286 49360
rect 208854 49348 208860 49360
rect 186280 49320 208860 49348
rect 186280 49308 186286 49320
rect 208854 49308 208860 49320
rect 208912 49308 208918 49360
rect 217962 49308 217968 49360
rect 218020 49348 218026 49360
rect 233326 49348 233332 49360
rect 218020 49320 233332 49348
rect 218020 49308 218026 49320
rect 233326 49308 233332 49320
rect 233384 49308 233390 49360
rect 234522 49308 234528 49360
rect 234580 49348 234586 49360
rect 246482 49348 246488 49360
rect 234580 49320 246488 49348
rect 234580 49308 234586 49320
rect 246482 49308 246488 49320
rect 246540 49308 246546 49360
rect 251082 49308 251088 49360
rect 251140 49348 251146 49360
rect 259546 49348 259552 49360
rect 251140 49320 259552 49348
rect 251140 49308 251146 49320
rect 259546 49308 259552 49320
rect 259604 49308 259610 49360
rect 419166 49308 419172 49360
rect 419224 49348 419230 49360
rect 422938 49348 422944 49360
rect 419224 49320 422944 49348
rect 419224 49308 419230 49320
rect 422938 49308 422944 49320
rect 422996 49308 423002 49360
rect 465166 49308 465172 49360
rect 465224 49348 465230 49360
rect 510706 49348 510712 49360
rect 465224 49320 510712 49348
rect 465224 49308 465230 49320
rect 510706 49308 510712 49320
rect 510764 49308 510770 49360
rect 57882 49240 57888 49292
rect 57940 49280 57946 49292
rect 107470 49280 107476 49292
rect 57940 49252 107476 49280
rect 57940 49240 57946 49252
rect 107470 49240 107476 49252
rect 107528 49240 107534 49292
rect 122742 49240 122748 49292
rect 122800 49280 122806 49292
rect 158162 49280 158168 49292
rect 122800 49252 158168 49280
rect 122800 49240 122806 49252
rect 158162 49240 158168 49252
rect 158220 49240 158226 49292
rect 179322 49240 179328 49292
rect 179380 49280 179386 49292
rect 203242 49280 203248 49292
rect 179380 49252 203248 49280
rect 179380 49240 179386 49252
rect 203242 49240 203248 49252
rect 203300 49240 203306 49292
rect 215202 49240 215208 49292
rect 215260 49280 215266 49292
rect 231394 49280 231400 49292
rect 215260 49252 231400 49280
rect 215260 49240 215266 49252
rect 231394 49240 231400 49252
rect 231452 49240 231458 49292
rect 233142 49240 233148 49292
rect 233200 49280 233206 49292
rect 245470 49280 245476 49292
rect 233200 49252 245476 49280
rect 233200 49240 233206 49252
rect 245470 49240 245476 49252
rect 245528 49240 245534 49292
rect 246942 49240 246948 49292
rect 247000 49280 247006 49292
rect 256786 49280 256792 49292
rect 247000 49252 256792 49280
rect 247000 49240 247006 49252
rect 256786 49240 256792 49252
rect 256844 49240 256850 49292
rect 266262 49240 266268 49292
rect 266320 49280 266326 49292
rect 271782 49280 271788 49292
rect 266320 49252 271788 49280
rect 266320 49240 266326 49252
rect 271782 49240 271788 49252
rect 271840 49240 271846 49292
rect 476482 49240 476488 49292
rect 476540 49280 476546 49292
rect 524414 49280 524420 49292
rect 476540 49252 524420 49280
rect 476540 49240 476546 49252
rect 524414 49240 524420 49252
rect 524472 49240 524478 49292
rect 50982 49172 50988 49224
rect 51040 49212 51046 49224
rect 101858 49212 101864 49224
rect 51040 49184 101864 49212
rect 51040 49172 51046 49184
rect 101858 49172 101864 49184
rect 101916 49172 101922 49224
rect 115842 49172 115848 49224
rect 115900 49212 115906 49224
rect 152550 49212 152556 49224
rect 115900 49184 152556 49212
rect 115900 49172 115906 49184
rect 152550 49172 152556 49184
rect 152608 49172 152614 49224
rect 172422 49172 172428 49224
rect 172480 49212 172486 49224
rect 197630 49212 197636 49224
rect 172480 49184 197636 49212
rect 172480 49172 172486 49184
rect 197630 49172 197636 49184
rect 197688 49172 197694 49224
rect 208302 49172 208308 49224
rect 208360 49212 208366 49224
rect 225782 49212 225788 49224
rect 208360 49184 225788 49212
rect 208360 49172 208366 49184
rect 225782 49172 225788 49184
rect 225840 49172 225846 49224
rect 229002 49172 229008 49224
rect 229060 49212 229066 49224
rect 241698 49212 241704 49224
rect 229060 49184 241704 49212
rect 229060 49172 229066 49184
rect 241698 49172 241704 49184
rect 241756 49172 241762 49224
rect 242802 49172 242808 49224
rect 242860 49212 242866 49224
rect 253014 49212 253020 49224
rect 242860 49184 253020 49212
rect 242860 49172 242866 49184
rect 253014 49172 253020 49184
rect 253072 49172 253078 49224
rect 253842 49172 253848 49224
rect 253900 49212 253906 49224
rect 261478 49212 261484 49224
rect 253900 49184 261484 49212
rect 253900 49172 253906 49184
rect 261478 49172 261484 49184
rect 261536 49172 261542 49224
rect 482094 49172 482100 49224
rect 482152 49212 482158 49224
rect 531314 49212 531320 49224
rect 482152 49184 531320 49212
rect 482152 49172 482158 49184
rect 531314 49172 531320 49184
rect 531372 49172 531378 49224
rect 13078 49104 13084 49156
rect 13136 49144 13142 49156
rect 69934 49144 69940 49156
rect 13136 49116 69940 49144
rect 13136 49104 13142 49116
rect 69934 49104 69940 49116
rect 69992 49104 69998 49156
rect 107562 49104 107568 49156
rect 107620 49144 107626 49156
rect 146938 49144 146944 49156
rect 107620 49116 146944 49144
rect 107620 49104 107626 49116
rect 146938 49104 146944 49116
rect 146996 49104 147002 49156
rect 160002 49104 160008 49156
rect 160060 49144 160066 49156
rect 188246 49144 188252 49156
rect 160060 49116 188252 49144
rect 160060 49104 160066 49116
rect 188246 49104 188252 49116
rect 188304 49104 188310 49156
rect 206922 49104 206928 49156
rect 206980 49144 206986 49156
rect 224862 49144 224868 49156
rect 206980 49116 224868 49144
rect 206980 49104 206986 49116
rect 224862 49104 224868 49116
rect 224920 49104 224926 49156
rect 226242 49104 226248 49156
rect 226300 49144 226306 49156
rect 239858 49144 239864 49156
rect 226300 49116 239864 49144
rect 226300 49104 226306 49116
rect 239858 49104 239864 49116
rect 239916 49104 239922 49156
rect 244182 49104 244188 49156
rect 244240 49144 244246 49156
rect 253934 49144 253940 49156
rect 244240 49116 253940 49144
rect 244240 49104 244246 49116
rect 253934 49104 253940 49116
rect 253992 49104 253998 49156
rect 257982 49104 257988 49156
rect 258040 49144 258046 49156
rect 265250 49144 265256 49156
rect 258040 49116 265256 49144
rect 258040 49104 258046 49116
rect 265250 49104 265256 49116
rect 265308 49104 265314 49156
rect 267642 49104 267648 49156
rect 267700 49144 267706 49156
rect 272702 49144 272708 49156
rect 267700 49116 272708 49144
rect 267700 49104 267706 49116
rect 272702 49104 272708 49116
rect 272760 49104 272766 49156
rect 277302 49104 277308 49156
rect 277360 49144 277366 49156
rect 280246 49144 280252 49156
rect 277360 49116 280252 49144
rect 277360 49104 277366 49116
rect 280246 49104 280252 49116
rect 280304 49104 280310 49156
rect 426710 49104 426716 49156
rect 426768 49144 426774 49156
rect 438118 49144 438124 49156
rect 426768 49116 438124 49144
rect 426768 49104 426774 49116
rect 438118 49104 438124 49116
rect 438176 49104 438182 49156
rect 487706 49104 487712 49156
rect 487764 49144 487770 49156
rect 538214 49144 538220 49156
rect 487764 49116 538220 49144
rect 487764 49104 487770 49116
rect 538214 49104 538220 49116
rect 538272 49104 538278 49156
rect 8938 49036 8944 49088
rect 8996 49076 9002 49088
rect 66162 49076 66168 49088
rect 8996 49048 66168 49076
rect 8996 49036 9002 49048
rect 66162 49036 66168 49048
rect 66220 49036 66226 49088
rect 103422 49036 103428 49088
rect 103480 49076 103486 49088
rect 143166 49076 143172 49088
rect 103480 49048 143172 49076
rect 103480 49036 103486 49048
rect 143166 49036 143172 49048
rect 143224 49036 143230 49088
rect 158622 49036 158628 49088
rect 158680 49076 158686 49088
rect 186314 49076 186320 49088
rect 158680 49048 186320 49076
rect 158680 49036 158686 49048
rect 186314 49036 186320 49048
rect 186372 49036 186378 49088
rect 213822 49036 213828 49088
rect 213880 49076 213886 49088
rect 230474 49076 230480 49088
rect 213880 49048 230480 49076
rect 213880 49036 213886 49048
rect 230474 49036 230480 49048
rect 230532 49036 230538 49088
rect 231762 49036 231768 49088
rect 231820 49076 231826 49088
rect 244550 49076 244556 49088
rect 231820 49048 244556 49076
rect 231820 49036 231826 49048
rect 244550 49036 244556 49048
rect 244608 49036 244614 49088
rect 245562 49036 245568 49088
rect 245620 49076 245626 49088
rect 255866 49076 255872 49088
rect 245620 49048 255872 49076
rect 245620 49036 245626 49048
rect 255866 49036 255872 49048
rect 255924 49036 255930 49088
rect 256602 49036 256608 49088
rect 256660 49076 256666 49088
rect 264238 49076 264244 49088
rect 256660 49048 264244 49076
rect 256660 49036 256666 49048
rect 264238 49036 264244 49048
rect 264296 49036 264302 49088
rect 264882 49036 264888 49088
rect 264940 49076 264946 49088
rect 270862 49076 270868 49088
rect 264940 49048 270868 49076
rect 264940 49036 264946 49048
rect 270862 49036 270868 49048
rect 270920 49036 270926 49088
rect 273162 49036 273168 49088
rect 273220 49076 273226 49088
rect 277394 49076 277400 49088
rect 273220 49048 277400 49076
rect 273220 49036 273226 49048
rect 277394 49036 277400 49048
rect 277452 49036 277458 49088
rect 391014 49036 391020 49088
rect 391072 49076 391078 49088
rect 416866 49076 416872 49088
rect 391072 49048 416872 49076
rect 391072 49036 391078 49048
rect 416866 49036 416872 49048
rect 416924 49036 416930 49088
rect 435174 49036 435180 49088
rect 435232 49076 435238 49088
rect 457438 49076 457444 49088
rect 435232 49048 457444 49076
rect 435232 49036 435238 49048
rect 457438 49036 457444 49048
rect 457496 49036 457502 49088
rect 493318 49036 493324 49088
rect 493376 49076 493382 49088
rect 546494 49076 546500 49088
rect 493376 49048 546500 49076
rect 493376 49036 493382 49048
rect 546494 49036 546500 49048
rect 546552 49036 546558 49088
rect 17218 48968 17224 49020
rect 17276 49008 17282 49020
rect 74626 49008 74632 49020
rect 17276 48980 74632 49008
rect 17276 48968 17282 48980
rect 74626 48968 74632 48980
rect 74684 48968 74690 49020
rect 79962 48968 79968 49020
rect 80020 49008 80026 49020
rect 124398 49008 124404 49020
rect 80020 48980 124404 49008
rect 80020 48968 80026 48980
rect 124398 48968 124404 48980
rect 124456 48968 124462 49020
rect 125502 48968 125508 49020
rect 125560 49008 125566 49020
rect 160094 49008 160100 49020
rect 125560 48980 160100 49008
rect 125560 48968 125566 48980
rect 160094 48968 160100 48980
rect 160152 48968 160158 49020
rect 165522 48968 165528 49020
rect 165580 49008 165586 49020
rect 192018 49008 192024 49020
rect 165580 48980 192024 49008
rect 165580 48968 165586 48980
rect 192018 48968 192024 48980
rect 192076 48968 192082 49020
rect 202782 48968 202788 49020
rect 202840 49008 202846 49020
rect 222010 49008 222016 49020
rect 202840 48980 222016 49008
rect 202840 48968 202846 48980
rect 222010 48968 222016 48980
rect 222068 48968 222074 49020
rect 222102 48968 222108 49020
rect 222160 49008 222166 49020
rect 237006 49008 237012 49020
rect 222160 48980 237012 49008
rect 222160 48968 222166 48980
rect 237006 48968 237012 48980
rect 237064 48968 237070 49020
rect 240042 48968 240048 49020
rect 240100 49008 240106 49020
rect 251174 49008 251180 49020
rect 240100 48980 251180 49008
rect 240100 48968 240106 48980
rect 251174 48968 251180 48980
rect 251232 48968 251238 49020
rect 252462 48968 252468 49020
rect 252520 49008 252526 49020
rect 260558 49008 260564 49020
rect 252520 48980 260564 49008
rect 252520 48968 252526 48980
rect 260558 48968 260564 48980
rect 260616 48968 260622 49020
rect 350626 48968 350632 49020
rect 350684 49008 350690 49020
rect 365806 49008 365812 49020
rect 350684 48980 365812 49008
rect 350684 48968 350690 48980
rect 365806 48968 365812 48980
rect 365864 48968 365870 49020
rect 373166 48968 373172 49020
rect 373224 49008 373230 49020
rect 391198 49008 391204 49020
rect 373224 48980 391204 49008
rect 373224 48968 373230 48980
rect 391198 48968 391204 48980
rect 391256 48968 391262 49020
rect 406010 48968 406016 49020
rect 406068 49008 406074 49020
rect 434714 49008 434720 49020
rect 406068 48980 434720 49008
rect 406068 48968 406074 48980
rect 434714 48968 434720 48980
rect 434772 48968 434778 49020
rect 454862 48968 454868 49020
rect 454920 49008 454926 49020
rect 482278 49008 482284 49020
rect 454920 48980 482284 49008
rect 454920 48968 454926 48980
rect 482278 48968 482284 48980
rect 482336 48968 482342 49020
rect 498930 48968 498936 49020
rect 498988 49008 498994 49020
rect 553394 49008 553400 49020
rect 498988 48980 553400 49008
rect 498988 48968 498994 48980
rect 553394 48968 553400 48980
rect 553452 48968 553458 49020
rect 271782 48832 271788 48884
rect 271840 48872 271846 48884
rect 276474 48872 276480 48884
rect 271840 48844 276480 48872
rect 271840 48832 271846 48844
rect 276474 48832 276480 48844
rect 276532 48832 276538 48884
rect 79318 48764 79324 48816
rect 79376 48804 79382 48816
rect 80238 48804 80244 48816
rect 79376 48776 80244 48804
rect 79376 48764 79382 48776
rect 80238 48764 80244 48776
rect 80296 48764 80302 48816
rect 92474 48764 92480 48816
rect 92532 48804 92538 48816
rect 93118 48804 93124 48816
rect 92532 48776 93124 48804
rect 92532 48764 92538 48776
rect 93118 48764 93124 48776
rect 93176 48764 93182 48816
rect 95234 48764 95240 48816
rect 95292 48804 95298 48816
rect 95878 48804 95884 48816
rect 95292 48776 95884 48804
rect 95292 48764 95298 48776
rect 95878 48764 95884 48776
rect 95936 48764 95942 48816
rect 103514 48764 103520 48816
rect 103572 48804 103578 48816
rect 104342 48804 104348 48816
rect 103572 48776 104348 48804
rect 103572 48764 103578 48776
rect 104342 48764 104348 48776
rect 104400 48764 104406 48816
rect 108298 48764 108304 48816
rect 108356 48804 108362 48816
rect 109402 48804 109408 48816
rect 108356 48776 109408 48804
rect 108356 48764 108362 48776
rect 109402 48764 109408 48776
rect 109460 48764 109466 48816
rect 139394 48764 139400 48816
rect 139452 48804 139458 48816
rect 140038 48804 140044 48816
rect 139452 48776 140044 48804
rect 139452 48764 139458 48776
rect 140038 48764 140044 48776
rect 140096 48764 140102 48816
rect 144914 48764 144920 48816
rect 144972 48804 144978 48816
rect 145742 48804 145748 48816
rect 144972 48776 145748 48804
rect 144972 48764 144978 48776
rect 145742 48764 145748 48776
rect 145800 48764 145806 48816
rect 146938 48764 146944 48816
rect 146996 48804 147002 48816
rect 147858 48804 147864 48816
rect 146996 48776 147864 48804
rect 146996 48764 147002 48776
rect 147858 48764 147864 48776
rect 147916 48764 147922 48816
rect 162118 48764 162124 48816
rect 162176 48804 162182 48816
rect 162854 48804 162860 48816
rect 162176 48776 162860 48804
rect 162176 48764 162182 48776
rect 162854 48764 162860 48776
rect 162912 48764 162918 48816
rect 179414 48764 179420 48816
rect 179472 48804 179478 48816
rect 180334 48804 180340 48816
rect 179472 48776 180340 48804
rect 179472 48764 179478 48776
rect 180334 48764 180340 48776
rect 180392 48764 180398 48816
rect 212534 48764 212540 48816
rect 212592 48804 212598 48816
rect 213270 48804 213276 48816
rect 212592 48776 213276 48804
rect 212592 48764 212598 48776
rect 213270 48764 213276 48776
rect 213328 48764 213334 48816
rect 215294 48764 215300 48816
rect 215352 48804 215358 48816
rect 216030 48804 216036 48816
rect 215352 48776 216036 48804
rect 215352 48764 215358 48776
rect 216030 48764 216036 48776
rect 216088 48764 216094 48816
rect 226334 48764 226340 48816
rect 226392 48804 226398 48816
rect 227254 48804 227260 48816
rect 226392 48776 227260 48804
rect 226392 48764 226398 48776
rect 227254 48764 227260 48776
rect 227312 48764 227318 48816
rect 259362 48764 259368 48816
rect 259420 48804 259426 48816
rect 266170 48804 266176 48816
rect 259420 48776 266176 48804
rect 259420 48764 259426 48776
rect 266170 48764 266176 48776
rect 266228 48764 266234 48816
rect 272518 48764 272524 48816
rect 272576 48804 272582 48816
rect 275554 48804 275560 48816
rect 272576 48776 275560 48804
rect 272576 48764 272582 48776
rect 275554 48764 275560 48776
rect 275612 48764 275618 48816
rect 281442 48764 281448 48816
rect 281500 48804 281506 48816
rect 284018 48804 284024 48816
rect 281500 48776 284024 48804
rect 281500 48764 281506 48776
rect 284018 48764 284024 48776
rect 284076 48764 284082 48816
rect 296622 48764 296628 48816
rect 296680 48804 296686 48816
rect 296898 48804 296904 48816
rect 296680 48776 296904 48804
rect 296680 48764 296686 48776
rect 296898 48764 296904 48776
rect 296956 48764 296962 48816
rect 299934 48764 299940 48816
rect 299992 48804 299998 48816
rect 301038 48804 301044 48816
rect 299992 48776 301044 48804
rect 299992 48764 299998 48776
rect 301038 48764 301044 48776
rect 301096 48764 301102 48816
rect 309318 48764 309324 48816
rect 309376 48804 309382 48816
rect 310422 48804 310428 48816
rect 309376 48776 310428 48804
rect 309376 48764 309382 48776
rect 310422 48764 310428 48776
rect 310480 48764 310486 48816
rect 311250 48764 311256 48816
rect 311308 48804 311314 48816
rect 312538 48804 312544 48816
rect 311308 48776 312544 48804
rect 311308 48764 311314 48776
rect 312538 48764 312544 48776
rect 312596 48764 312602 48816
rect 314010 48764 314016 48816
rect 314068 48804 314074 48816
rect 315298 48804 315304 48816
rect 314068 48776 315304 48804
rect 314068 48764 314074 48776
rect 315298 48764 315304 48776
rect 315356 48764 315362 48816
rect 317782 48764 317788 48816
rect 317840 48804 317846 48816
rect 320818 48804 320824 48816
rect 317840 48776 320824 48804
rect 317840 48764 317846 48776
rect 320818 48764 320824 48776
rect 320876 48764 320882 48816
rect 321554 48764 321560 48816
rect 321612 48804 321618 48816
rect 322750 48804 322756 48816
rect 321612 48776 322756 48804
rect 321612 48764 321618 48776
rect 322750 48764 322756 48776
rect 322808 48764 322814 48816
rect 326246 48764 326252 48816
rect 326304 48804 326310 48816
rect 326982 48804 326988 48816
rect 326304 48776 326988 48804
rect 326304 48764 326310 48776
rect 326982 48764 326988 48776
rect 327040 48764 327046 48816
rect 327166 48764 327172 48816
rect 327224 48804 327230 48816
rect 328362 48804 328368 48816
rect 327224 48776 328368 48804
rect 327224 48764 327230 48776
rect 328362 48764 328368 48776
rect 328420 48764 328426 48816
rect 329006 48764 329012 48816
rect 329064 48804 329070 48816
rect 329742 48804 329748 48816
rect 329064 48776 329748 48804
rect 329064 48764 329070 48776
rect 329742 48764 329748 48776
rect 329800 48764 329806 48816
rect 330018 48764 330024 48816
rect 330076 48804 330082 48816
rect 331122 48804 331128 48816
rect 330076 48776 331128 48804
rect 330076 48764 330082 48776
rect 331122 48764 331128 48776
rect 331180 48764 331186 48816
rect 332778 48764 332784 48816
rect 332836 48804 332842 48816
rect 333882 48804 333888 48816
rect 332836 48776 333888 48804
rect 332836 48764 332842 48776
rect 333882 48764 333888 48776
rect 333940 48764 333946 48816
rect 335630 48764 335636 48816
rect 335688 48804 335694 48816
rect 336642 48804 336648 48816
rect 335688 48776 336648 48804
rect 335688 48764 335694 48776
rect 336642 48764 336648 48776
rect 336700 48764 336706 48816
rect 338482 48764 338488 48816
rect 338540 48804 338546 48816
rect 339402 48804 339408 48816
rect 338540 48776 339408 48804
rect 338540 48764 338546 48776
rect 339402 48764 339408 48776
rect 339460 48764 339466 48816
rect 341242 48764 341248 48816
rect 341300 48804 341306 48816
rect 342162 48804 342168 48816
rect 341300 48776 342168 48804
rect 341300 48764 341306 48776
rect 342162 48764 342168 48776
rect 342220 48764 342226 48816
rect 344094 48764 344100 48816
rect 344152 48804 344158 48816
rect 344922 48804 344928 48816
rect 344152 48776 344928 48804
rect 344152 48764 344158 48776
rect 344922 48764 344928 48776
rect 344980 48764 344986 48816
rect 345014 48764 345020 48816
rect 345072 48804 345078 48816
rect 346210 48804 346216 48816
rect 345072 48776 346216 48804
rect 345072 48764 345078 48776
rect 346210 48764 346216 48776
rect 346268 48764 346274 48816
rect 347866 48764 347872 48816
rect 347924 48804 347930 48816
rect 348970 48804 348976 48816
rect 347924 48776 348976 48804
rect 347924 48764 347930 48776
rect 348970 48764 348976 48776
rect 349028 48764 349034 48816
rect 353478 48764 353484 48816
rect 353536 48804 353542 48816
rect 354490 48804 354496 48816
rect 353536 48776 354496 48804
rect 353536 48764 353542 48776
rect 354490 48764 354496 48776
rect 354548 48764 354554 48816
rect 356238 48764 356244 48816
rect 356296 48804 356302 48816
rect 357250 48804 357256 48816
rect 356296 48776 357256 48804
rect 356296 48764 356302 48776
rect 357250 48764 357256 48776
rect 357308 48764 357314 48816
rect 359090 48764 359096 48816
rect 359148 48804 359154 48816
rect 360010 48804 360016 48816
rect 359148 48776 360016 48804
rect 359148 48764 359154 48776
rect 360010 48764 360016 48776
rect 360068 48764 360074 48816
rect 361942 48764 361948 48816
rect 362000 48804 362006 48816
rect 362770 48804 362776 48816
rect 362000 48776 362776 48804
rect 362000 48764 362006 48776
rect 362770 48764 362776 48776
rect 362828 48764 362834 48816
rect 367554 48764 367560 48816
rect 367612 48804 367618 48816
rect 368382 48804 368388 48816
rect 367612 48776 368388 48804
rect 367612 48764 367618 48776
rect 368382 48764 368388 48776
rect 368440 48764 368446 48816
rect 368474 48764 368480 48816
rect 368532 48804 368538 48816
rect 369670 48804 369676 48816
rect 368532 48776 369676 48804
rect 368532 48764 368538 48776
rect 369670 48764 369676 48776
rect 369728 48764 369734 48816
rect 370314 48764 370320 48816
rect 370372 48804 370378 48816
rect 371142 48804 371148 48816
rect 370372 48776 371148 48804
rect 370372 48764 370378 48776
rect 371142 48764 371148 48776
rect 371200 48764 371206 48816
rect 371326 48764 371332 48816
rect 371384 48804 371390 48816
rect 372430 48804 372436 48816
rect 371384 48776 372436 48804
rect 371384 48764 371390 48776
rect 372430 48764 372436 48776
rect 372488 48764 372494 48816
rect 374086 48764 374092 48816
rect 374144 48804 374150 48816
rect 375282 48804 375288 48816
rect 374144 48776 375288 48804
rect 374144 48764 374150 48776
rect 375282 48764 375288 48776
rect 375340 48764 375346 48816
rect 376938 48764 376944 48816
rect 376996 48804 377002 48816
rect 378042 48804 378048 48816
rect 376996 48776 378048 48804
rect 376996 48764 377002 48776
rect 378042 48764 378048 48776
rect 378100 48764 378106 48816
rect 379698 48764 379704 48816
rect 379756 48804 379762 48816
rect 380802 48804 380808 48816
rect 379756 48776 380808 48804
rect 379756 48764 379762 48776
rect 380802 48764 380808 48776
rect 380860 48764 380866 48816
rect 382550 48764 382556 48816
rect 382608 48804 382614 48816
rect 383470 48804 383476 48816
rect 382608 48776 383476 48804
rect 382608 48764 382614 48776
rect 383470 48764 383476 48776
rect 383528 48764 383534 48816
rect 385402 48764 385408 48816
rect 385460 48804 385466 48816
rect 386230 48804 386236 48816
rect 385460 48776 386236 48804
rect 385460 48764 385466 48776
rect 386230 48764 386236 48776
rect 386288 48764 386294 48816
rect 388162 48764 388168 48816
rect 388220 48804 388226 48816
rect 389082 48804 389088 48816
rect 388220 48776 389088 48804
rect 388220 48764 388226 48776
rect 389082 48764 389088 48776
rect 389140 48764 389146 48816
rect 389174 48764 389180 48816
rect 389232 48804 389238 48816
rect 390462 48804 390468 48816
rect 389232 48776 390468 48804
rect 389232 48764 389238 48776
rect 390462 48764 390468 48776
rect 390520 48764 390526 48816
rect 391934 48764 391940 48816
rect 391992 48804 391998 48816
rect 393222 48804 393228 48816
rect 391992 48776 393228 48804
rect 391992 48764 391998 48776
rect 393222 48764 393228 48776
rect 393280 48764 393286 48816
rect 394786 48764 394792 48816
rect 394844 48804 394850 48816
rect 395982 48804 395988 48816
rect 394844 48776 395988 48804
rect 394844 48764 394850 48776
rect 395982 48764 395988 48776
rect 396040 48764 396046 48816
rect 397546 48764 397552 48816
rect 397604 48804 397610 48816
rect 398742 48804 398748 48816
rect 397604 48776 398748 48804
rect 397604 48764 397610 48776
rect 398742 48764 398748 48776
rect 398800 48764 398806 48816
rect 400398 48764 400404 48816
rect 400456 48804 400462 48816
rect 401502 48804 401508 48816
rect 400456 48776 401508 48804
rect 400456 48764 400462 48776
rect 401502 48764 401508 48776
rect 401560 48764 401566 48816
rect 403250 48764 403256 48816
rect 403308 48804 403314 48816
rect 404262 48804 404268 48816
rect 403308 48776 404268 48804
rect 403308 48764 403314 48776
rect 404262 48764 404268 48776
rect 404320 48764 404326 48816
rect 408862 48764 408868 48816
rect 408920 48804 408926 48816
rect 409782 48804 409788 48816
rect 408920 48776 409788 48804
rect 408920 48764 408926 48776
rect 409782 48764 409788 48776
rect 409840 48764 409846 48816
rect 411622 48764 411628 48816
rect 411680 48804 411686 48816
rect 412542 48804 412548 48816
rect 411680 48776 412548 48804
rect 411680 48764 411686 48776
rect 412542 48764 412548 48776
rect 412600 48764 412606 48816
rect 412634 48764 412640 48816
rect 412692 48804 412698 48816
rect 413922 48804 413928 48816
rect 412692 48776 413928 48804
rect 412692 48764 412698 48776
rect 413922 48764 413928 48776
rect 413980 48764 413986 48816
rect 414474 48764 414480 48816
rect 414532 48804 414538 48816
rect 415302 48804 415308 48816
rect 414532 48776 415308 48804
rect 414532 48764 414538 48776
rect 415302 48764 415308 48776
rect 415360 48764 415366 48816
rect 415394 48764 415400 48816
rect 415452 48804 415458 48816
rect 416682 48804 416688 48816
rect 415452 48776 416688 48804
rect 415452 48764 415458 48776
rect 416682 48764 416688 48776
rect 416740 48764 416746 48816
rect 420086 48764 420092 48816
rect 420144 48804 420150 48816
rect 420822 48804 420828 48816
rect 420144 48776 420828 48804
rect 420144 48764 420150 48776
rect 420822 48764 420828 48776
rect 420880 48764 420886 48816
rect 421006 48764 421012 48816
rect 421064 48804 421070 48816
rect 422202 48804 422208 48816
rect 421064 48776 422208 48804
rect 421064 48764 421070 48776
rect 422202 48764 422208 48776
rect 422260 48764 422266 48816
rect 423858 48764 423864 48816
rect 423916 48804 423922 48816
rect 424870 48804 424876 48816
rect 423916 48776 424876 48804
rect 423916 48764 423922 48776
rect 424870 48764 424876 48776
rect 424928 48764 424934 48816
rect 432322 48764 432328 48816
rect 432380 48804 432386 48816
rect 433978 48804 433984 48816
rect 432380 48776 433984 48804
rect 432380 48764 432386 48776
rect 433978 48764 433984 48776
rect 434036 48764 434042 48816
rect 436094 48764 436100 48816
rect 436152 48804 436158 48816
rect 437290 48804 437296 48816
rect 436152 48776 437296 48804
rect 436152 48764 436158 48776
rect 437290 48764 437296 48776
rect 437348 48764 437354 48816
rect 437934 48764 437940 48816
rect 437992 48804 437998 48816
rect 438762 48804 438768 48816
rect 437992 48776 438768 48804
rect 437992 48764 437998 48776
rect 438762 48764 438768 48776
rect 438820 48764 438826 48816
rect 438854 48764 438860 48816
rect 438912 48804 438918 48816
rect 440142 48804 440148 48816
rect 438912 48776 440148 48804
rect 438912 48764 438918 48776
rect 440142 48764 440148 48776
rect 440200 48764 440206 48816
rect 441706 48764 441712 48816
rect 441764 48804 441770 48816
rect 442810 48804 442816 48816
rect 441764 48776 442816 48804
rect 441764 48764 441770 48776
rect 442810 48764 442816 48776
rect 442868 48764 442874 48816
rect 444558 48764 444564 48816
rect 444616 48804 444622 48816
rect 445570 48804 445576 48816
rect 444616 48776 445576 48804
rect 444616 48764 444622 48776
rect 445570 48764 445576 48776
rect 445628 48764 445634 48816
rect 452930 48764 452936 48816
rect 452988 48804 452994 48816
rect 453850 48804 453856 48816
rect 452988 48776 453856 48804
rect 452988 48764 452994 48776
rect 453850 48764 453856 48776
rect 453908 48764 453914 48816
rect 458634 48764 458640 48816
rect 458692 48804 458698 48816
rect 459462 48804 459468 48816
rect 458692 48776 459468 48804
rect 458692 48764 458698 48776
rect 459462 48764 459468 48776
rect 459520 48764 459526 48816
rect 459554 48764 459560 48816
rect 459612 48804 459618 48816
rect 460842 48804 460848 48816
rect 459612 48776 460848 48804
rect 459612 48764 459618 48776
rect 460842 48764 460848 48776
rect 460900 48764 460906 48816
rect 462314 48764 462320 48816
rect 462372 48804 462378 48816
rect 463602 48804 463608 48816
rect 462372 48776 463608 48804
rect 462372 48764 462378 48776
rect 463602 48764 463608 48776
rect 463660 48764 463666 48816
rect 464246 48764 464252 48816
rect 464304 48804 464310 48816
rect 464982 48804 464988 48816
rect 464304 48776 464988 48804
rect 464304 48764 464310 48776
rect 464982 48764 464988 48776
rect 465040 48764 465046 48816
rect 467006 48764 467012 48816
rect 467064 48804 467070 48816
rect 467742 48804 467748 48816
rect 467064 48776 467748 48804
rect 467064 48764 467070 48776
rect 467742 48764 467748 48776
rect 467800 48764 467806 48816
rect 468018 48764 468024 48816
rect 468076 48804 468082 48816
rect 469122 48804 469128 48816
rect 468076 48776 469128 48804
rect 468076 48764 468082 48776
rect 469122 48764 469128 48776
rect 469180 48764 469186 48816
rect 470778 48764 470784 48816
rect 470836 48804 470842 48816
rect 471882 48804 471888 48816
rect 470836 48776 471888 48804
rect 470836 48764 470842 48776
rect 471882 48764 471888 48776
rect 471940 48764 471946 48816
rect 473630 48764 473636 48816
rect 473688 48804 473694 48816
rect 474642 48804 474648 48816
rect 473688 48776 474648 48804
rect 473688 48764 473694 48776
rect 474642 48764 474648 48776
rect 474700 48764 474706 48816
rect 479242 48764 479248 48816
rect 479300 48804 479306 48816
rect 480162 48804 480168 48816
rect 479300 48776 480168 48804
rect 479300 48764 479306 48776
rect 480162 48764 480168 48776
rect 480220 48764 480226 48816
rect 483014 48764 483020 48816
rect 483072 48804 483078 48816
rect 484302 48804 484308 48816
rect 483072 48776 484308 48804
rect 483072 48764 483078 48776
rect 484302 48764 484308 48776
rect 484360 48764 484366 48816
rect 484854 48764 484860 48816
rect 484912 48804 484918 48816
rect 485682 48804 485688 48816
rect 484912 48776 485688 48804
rect 484912 48764 484918 48776
rect 485682 48764 485688 48776
rect 485740 48764 485746 48816
rect 506474 48764 506480 48816
rect 506532 48804 506538 48816
rect 507670 48804 507676 48816
rect 506532 48776 507676 48804
rect 506532 48764 506538 48776
rect 507670 48764 507676 48776
rect 507728 48764 507734 48816
rect 511166 48764 511172 48816
rect 511224 48804 511230 48816
rect 511902 48804 511908 48816
rect 511224 48776 511908 48804
rect 511224 48764 511230 48776
rect 511902 48764 511908 48776
rect 511960 48764 511966 48816
rect 514938 48764 514944 48816
rect 514996 48804 515002 48816
rect 516042 48804 516048 48816
rect 514996 48776 516048 48804
rect 514996 48764 515002 48776
rect 516042 48764 516048 48776
rect 516100 48764 516106 48816
rect 517698 48764 517704 48816
rect 517756 48804 517762 48816
rect 518802 48804 518808 48816
rect 517756 48776 518808 48804
rect 517756 48764 517762 48776
rect 518802 48764 518808 48776
rect 518860 48764 518866 48816
rect 520550 48764 520556 48816
rect 520608 48804 520614 48816
rect 521470 48804 521476 48816
rect 520608 48776 521476 48804
rect 520608 48764 520614 48776
rect 521470 48764 521476 48776
rect 521528 48764 521534 48816
rect 204898 48696 204904 48748
rect 204956 48736 204962 48748
rect 207014 48736 207020 48748
rect 204956 48708 207020 48736
rect 204956 48696 204962 48708
rect 207014 48696 207020 48708
rect 207072 48696 207078 48748
rect 269022 48696 269028 48748
rect 269080 48736 269086 48748
rect 273622 48736 273628 48748
rect 269080 48708 273628 48736
rect 269080 48696 269086 48708
rect 273622 48696 273628 48708
rect 273680 48696 273686 48748
rect 280062 48696 280068 48748
rect 280120 48736 280126 48748
rect 282086 48736 282092 48748
rect 280120 48708 282092 48736
rect 280120 48696 280126 48708
rect 282086 48696 282092 48708
rect 282144 48696 282150 48748
rect 312170 48696 312176 48748
rect 312228 48736 312234 48748
rect 313182 48736 313188 48748
rect 312228 48708 313188 48736
rect 312228 48696 312234 48708
rect 313182 48696 313188 48708
rect 313240 48696 313246 48748
rect 314930 48696 314936 48748
rect 314988 48736 314994 48748
rect 315942 48736 315948 48748
rect 314988 48708 315948 48736
rect 314988 48696 314994 48708
rect 315942 48696 315948 48708
rect 316000 48696 316006 48748
rect 378778 48696 378784 48748
rect 378836 48736 378842 48748
rect 381538 48736 381544 48748
rect 378836 48708 381544 48736
rect 378836 48696 378842 48708
rect 381538 48696 381544 48708
rect 381596 48696 381602 48748
rect 390094 48696 390100 48748
rect 390152 48736 390158 48748
rect 391290 48736 391296 48748
rect 390152 48708 391296 48736
rect 390152 48696 390158 48708
rect 391290 48696 391296 48708
rect 391348 48696 391354 48748
rect 401318 48696 401324 48748
rect 401376 48736 401382 48748
rect 402238 48736 402244 48748
rect 401376 48708 402244 48736
rect 401376 48696 401382 48708
rect 402238 48696 402244 48708
rect 402296 48696 402302 48748
rect 407942 48696 407948 48748
rect 408000 48736 408006 48748
rect 410518 48736 410524 48748
rect 408000 48708 410524 48736
rect 408000 48696 408006 48708
rect 410518 48696 410524 48708
rect 410576 48696 410582 48748
rect 443546 48696 443552 48748
rect 443604 48736 443610 48748
rect 446398 48736 446404 48748
rect 443604 48708 446404 48736
rect 443604 48696 443610 48708
rect 446398 48696 446404 48708
rect 446456 48696 446462 48748
rect 461394 48696 461400 48748
rect 461452 48736 461458 48748
rect 464338 48736 464344 48748
rect 461452 48708 464344 48736
rect 461452 48696 461458 48708
rect 464338 48696 464344 48708
rect 464396 48696 464402 48748
rect 468938 48696 468944 48748
rect 468996 48736 469002 48748
rect 469858 48736 469864 48748
rect 468996 48708 469864 48736
rect 468996 48696 469002 48708
rect 469858 48696 469864 48708
rect 469916 48696 469922 48748
rect 472710 48696 472716 48748
rect 472768 48736 472774 48748
rect 475378 48736 475384 48748
rect 472768 48708 475384 48736
rect 472768 48696 472774 48708
rect 475378 48696 475384 48708
rect 475436 48696 475442 48748
rect 306558 48628 306564 48680
rect 306616 48668 306622 48680
rect 309318 48668 309324 48680
rect 306616 48640 309324 48668
rect 306616 48628 306622 48640
rect 309318 48628 309324 48640
rect 309376 48628 309382 48680
rect 396626 48628 396632 48680
rect 396684 48668 396690 48680
rect 399478 48668 399484 48680
rect 396684 48640 399484 48668
rect 396684 48628 396690 48640
rect 399478 48628 399484 48640
rect 399536 48628 399542 48680
rect 509326 48628 509332 48680
rect 509384 48668 509390 48680
rect 510430 48668 510436 48680
rect 509384 48640 510436 48668
rect 509384 48628 509390 48640
rect 510430 48628 510436 48640
rect 510488 48628 510494 48680
rect 512086 48628 512092 48680
rect 512144 48668 512150 48680
rect 513190 48668 513196 48680
rect 512144 48640 513196 48668
rect 512144 48628 512150 48640
rect 513190 48628 513196 48640
rect 513248 48628 513254 48680
rect 270402 48560 270408 48612
rect 270460 48600 270466 48612
rect 274634 48600 274640 48612
rect 270460 48572 274640 48600
rect 270460 48560 270466 48572
rect 274634 48560 274640 48572
rect 274692 48560 274698 48612
rect 279970 48560 279976 48612
rect 280028 48600 280034 48612
rect 283006 48600 283012 48612
rect 280028 48572 283012 48600
rect 280028 48560 280034 48572
rect 283006 48560 283012 48572
rect 283064 48560 283070 48612
rect 320634 48560 320640 48612
rect 320692 48600 320698 48612
rect 321462 48600 321468 48612
rect 320692 48572 321468 48600
rect 320692 48560 320698 48572
rect 321462 48560 321468 48572
rect 321520 48560 321526 48612
rect 323394 48560 323400 48612
rect 323452 48600 323458 48612
rect 324222 48600 324228 48612
rect 323452 48572 324228 48600
rect 323452 48560 323458 48572
rect 324222 48560 324228 48572
rect 324280 48560 324286 48612
rect 263502 48492 263508 48544
rect 263560 48532 263566 48544
rect 268930 48532 268936 48544
rect 263560 48504 268936 48532
rect 263560 48492 263566 48504
rect 268930 48492 268936 48504
rect 268988 48492 268994 48544
rect 346854 48492 346860 48544
rect 346912 48532 346918 48544
rect 347682 48532 347688 48544
rect 346912 48504 347688 48532
rect 346912 48492 346918 48504
rect 347682 48492 347688 48504
rect 347740 48492 347746 48544
rect 364702 48492 364708 48544
rect 364760 48532 364766 48544
rect 373258 48532 373264 48544
rect 364760 48504 373264 48532
rect 364760 48492 364766 48504
rect 373258 48492 373264 48504
rect 373316 48492 373322 48544
rect 418246 48492 418252 48544
rect 418304 48532 418310 48544
rect 420178 48532 420184 48544
rect 418304 48504 420184 48532
rect 418304 48492 418310 48504
rect 420178 48492 420184 48504
rect 420236 48492 420242 48544
rect 485866 48492 485872 48544
rect 485924 48532 485930 48544
rect 487062 48532 487068 48544
rect 485924 48504 487068 48532
rect 485924 48492 485930 48504
rect 487062 48492 487068 48504
rect 487120 48492 487126 48544
rect 491478 48492 491484 48544
rect 491536 48532 491542 48544
rect 492582 48532 492588 48544
rect 491536 48504 492588 48532
rect 491536 48492 491542 48504
rect 492582 48492 492588 48504
rect 492640 48492 492646 48544
rect 303706 48424 303712 48476
rect 303764 48464 303770 48476
rect 304902 48464 304908 48476
rect 303764 48436 304908 48464
rect 303764 48424 303770 48436
rect 304902 48424 304908 48436
rect 304960 48424 304966 48476
rect 417326 48424 417332 48476
rect 417384 48464 417390 48476
rect 418062 48464 418068 48476
rect 417384 48436 418068 48464
rect 417384 48424 417390 48436
rect 418062 48424 418068 48436
rect 418120 48424 418126 48476
rect 261478 48356 261484 48408
rect 261536 48396 261542 48408
rect 267090 48396 267096 48408
rect 261536 48368 267096 48396
rect 261536 48356 261542 48368
rect 267090 48356 267096 48368
rect 267148 48356 267154 48408
rect 429470 48356 429476 48408
rect 429528 48396 429534 48408
rect 430482 48396 430488 48408
rect 429528 48368 430488 48396
rect 429528 48356 429534 48368
rect 430482 48356 430488 48368
rect 430540 48356 430546 48408
rect 61378 48288 61384 48340
rect 61436 48328 61442 48340
rect 62482 48328 62488 48340
rect 61436 48300 62488 48328
rect 61436 48288 61442 48300
rect 62482 48288 62488 48300
rect 62540 48288 62546 48340
rect 111058 48288 111064 48340
rect 111116 48328 111122 48340
rect 112162 48328 112168 48340
rect 111116 48300 112168 48328
rect 111116 48288 111122 48300
rect 112162 48288 112168 48300
rect 112220 48288 112226 48340
rect 120718 48288 120724 48340
rect 120776 48328 120782 48340
rect 122558 48328 122564 48340
rect 120776 48300 122564 48328
rect 120776 48288 120782 48300
rect 122558 48288 122564 48300
rect 122616 48288 122622 48340
rect 126238 48288 126244 48340
rect 126296 48328 126302 48340
rect 128170 48328 128176 48340
rect 126296 48300 128176 48328
rect 126296 48288 126302 48300
rect 128170 48288 128176 48300
rect 128228 48288 128234 48340
rect 167638 48288 167644 48340
rect 167696 48328 167702 48340
rect 170398 48328 170404 48340
rect 167696 48300 170404 48328
rect 167696 48288 167702 48300
rect 170398 48288 170404 48300
rect 170456 48288 170462 48340
rect 284202 48288 284208 48340
rect 284260 48328 284266 48340
rect 285858 48328 285864 48340
rect 284260 48300 285864 48328
rect 284260 48288 284266 48300
rect 285858 48288 285864 48300
rect 285916 48288 285922 48340
rect 286962 48288 286968 48340
rect 287020 48328 287026 48340
rect 287698 48328 287704 48340
rect 287020 48300 287704 48328
rect 287020 48288 287026 48300
rect 287698 48288 287704 48300
rect 287756 48288 287762 48340
rect 289630 48328 289636 48340
rect 288268 48300 289636 48328
rect 288268 48272 288296 48300
rect 289630 48288 289636 48300
rect 289688 48288 289694 48340
rect 290918 48288 290924 48340
rect 290976 48328 290982 48340
rect 291470 48328 291476 48340
rect 290976 48300 291476 48328
rect 290976 48288 290982 48300
rect 291470 48288 291476 48300
rect 291528 48288 291534 48340
rect 300854 48288 300860 48340
rect 300912 48328 300918 48340
rect 302142 48328 302148 48340
rect 300912 48300 302148 48328
rect 300912 48288 300918 48300
rect 302142 48288 302148 48300
rect 302200 48288 302206 48340
rect 488994 48288 489000 48340
rect 489052 48328 489058 48340
rect 489638 48328 489644 48340
rect 489052 48300 489644 48328
rect 489052 48288 489058 48300
rect 489638 48288 489644 48300
rect 489696 48288 489702 48340
rect 494238 48288 494244 48340
rect 494296 48328 494302 48340
rect 495066 48328 495072 48340
rect 494296 48300 495072 48328
rect 494296 48288 494302 48300
rect 495066 48288 495072 48300
rect 495124 48288 495130 48340
rect 495158 48288 495164 48340
rect 495216 48328 495222 48340
rect 496078 48328 496084 48340
rect 495216 48300 496084 48328
rect 495216 48288 495222 48300
rect 496078 48288 496084 48300
rect 496136 48288 496142 48340
rect 505554 48288 505560 48340
rect 505612 48328 505618 48340
rect 506382 48328 506388 48340
rect 505612 48300 506388 48328
rect 505612 48288 505618 48300
rect 506382 48288 506388 48300
rect 506440 48288 506446 48340
rect 508314 48288 508320 48340
rect 508372 48328 508378 48340
rect 509142 48328 509148 48340
rect 508372 48300 509148 48328
rect 508372 48288 508378 48300
rect 509142 48288 509148 48300
rect 509200 48288 509206 48340
rect 168742 48260 168748 48272
rect 168703 48232 168748 48260
rect 168742 48220 168748 48232
rect 168800 48220 168806 48272
rect 288250 48220 288256 48272
rect 288308 48220 288314 48272
rect 489638 48192 489644 48204
rect 489599 48164 489644 48192
rect 489638 48152 489644 48164
rect 489696 48152 489702 48204
rect 10318 47540 10324 47592
rect 10376 47580 10382 47592
rect 65242 47580 65248 47592
rect 10376 47552 65248 47580
rect 10376 47540 10382 47552
rect 65242 47540 65248 47552
rect 65300 47540 65306 47592
rect 70302 47540 70308 47592
rect 70360 47580 70366 47592
rect 116854 47580 116860 47592
rect 70360 47552 116860 47580
rect 70360 47540 70366 47552
rect 116854 47540 116860 47552
rect 116912 47540 116918 47592
rect 155862 47540 155868 47592
rect 155920 47580 155926 47592
rect 184474 47580 184480 47592
rect 155920 47552 184480 47580
rect 155920 47540 155926 47552
rect 184474 47540 184480 47552
rect 184532 47540 184538 47592
rect 447318 47540 447324 47592
rect 447376 47580 447382 47592
rect 487154 47580 487160 47592
rect 447376 47552 487160 47580
rect 447376 47540 447382 47552
rect 487154 47540 487160 47552
rect 487212 47540 487218 47592
rect 497090 47540 497096 47592
rect 497148 47580 497154 47592
rect 550634 47580 550640 47592
rect 497148 47552 550640 47580
rect 497148 47540 497154 47552
rect 550634 47540 550640 47552
rect 550692 47540 550698 47592
rect 176654 46860 176660 46912
rect 176712 46900 176718 46912
rect 177574 46900 177580 46912
rect 176712 46872 177580 46900
rect 176712 46860 176718 46872
rect 177574 46860 177580 46872
rect 177632 46860 177638 46912
rect 293954 46900 293960 46912
rect 293915 46872 293960 46900
rect 293954 46860 293960 46872
rect 294012 46860 294018 46912
rect 118786 46248 118792 46300
rect 118844 46288 118850 46300
rect 119430 46288 119436 46300
rect 118844 46260 119436 46288
rect 118844 46248 118850 46260
rect 119430 46248 119436 46260
rect 119488 46248 119494 46300
rect 153194 46248 153200 46300
rect 153252 46288 153258 46300
rect 154206 46288 154212 46300
rect 153252 46260 154212 46288
rect 153252 46248 153258 46260
rect 154206 46248 154212 46260
rect 154264 46248 154270 46300
rect 155954 46248 155960 46300
rect 156012 46288 156018 46300
rect 156966 46288 156972 46300
rect 156012 46260 156972 46288
rect 156012 46248 156018 46260
rect 156966 46248 156972 46260
rect 157024 46248 157030 46300
rect 22002 46180 22008 46232
rect 22060 46220 22066 46232
rect 22060 46192 74028 46220
rect 22060 46180 22066 46192
rect 74000 46152 74028 46192
rect 77386 46180 77392 46232
rect 77444 46220 77450 46232
rect 78030 46220 78036 46232
rect 77444 46192 78036 46220
rect 77444 46180 77450 46192
rect 78030 46180 78036 46192
rect 78088 46180 78094 46232
rect 88242 46180 88248 46232
rect 88300 46220 88306 46232
rect 130930 46220 130936 46232
rect 88300 46192 130936 46220
rect 88300 46180 88306 46192
rect 130930 46180 130936 46192
rect 130988 46180 130994 46232
rect 132402 46180 132408 46232
rect 132460 46220 132466 46232
rect 165706 46220 165712 46232
rect 132460 46192 165712 46220
rect 132460 46180 132466 46192
rect 165706 46180 165712 46192
rect 165764 46180 165770 46232
rect 173894 46180 173900 46232
rect 173952 46220 173958 46232
rect 174814 46220 174820 46232
rect 173952 46192 174820 46220
rect 173952 46180 173958 46192
rect 174814 46180 174820 46192
rect 174872 46180 174878 46232
rect 455782 46180 455788 46232
rect 455840 46220 455846 46232
rect 498194 46220 498200 46232
rect 455840 46192 498200 46220
rect 455840 46180 455846 46192
rect 498194 46180 498200 46192
rect 498252 46180 498258 46232
rect 499942 46180 499948 46232
rect 500000 46220 500006 46232
rect 554774 46220 554780 46232
rect 500000 46192 554780 46220
rect 500000 46180 500006 46192
rect 554774 46180 554780 46192
rect 554832 46180 554838 46232
rect 78950 46152 78956 46164
rect 74000 46124 78956 46152
rect 78950 46112 78956 46124
rect 79008 46112 79014 46164
rect 27522 44820 27528 44872
rect 27580 44860 27586 44872
rect 82906 44860 82912 44872
rect 27580 44832 82912 44860
rect 27580 44820 27586 44832
rect 82906 44820 82912 44832
rect 82964 44820 82970 44872
rect 92382 44820 92388 44872
rect 92440 44860 92446 44872
rect 133874 44860 133880 44872
rect 92440 44832 133880 44860
rect 92440 44820 92446 44832
rect 133874 44820 133880 44832
rect 133932 44820 133938 44872
rect 139302 44820 139308 44872
rect 139360 44860 139366 44872
rect 171226 44860 171232 44872
rect 139360 44832 171232 44860
rect 139360 44820 139366 44832
rect 171226 44820 171232 44832
rect 171284 44820 171290 44872
rect 502702 44820 502708 44872
rect 502760 44860 502766 44872
rect 557534 44860 557540 44872
rect 502760 44832 557540 44860
rect 502760 44820 502766 44832
rect 557534 44820 557540 44832
rect 557592 44820 557598 44872
rect 85761 43503 85819 43509
rect 85761 43469 85773 43503
rect 85807 43500 85819 43503
rect 86494 43500 86500 43512
rect 85807 43472 86500 43500
rect 85807 43469 85819 43472
rect 85761 43463 85819 43469
rect 86494 43460 86500 43472
rect 86552 43460 86558 43512
rect 34422 43392 34428 43444
rect 34480 43432 34486 43444
rect 88426 43432 88432 43444
rect 34480 43404 88432 43432
rect 34480 43392 34486 43404
rect 88426 43392 88432 43404
rect 88484 43392 88490 43444
rect 129642 43392 129648 43444
rect 129700 43432 129706 43444
rect 162946 43432 162952 43444
rect 129700 43404 162952 43432
rect 129700 43392 129706 43404
rect 162946 43392 162952 43404
rect 163004 43392 163010 43444
rect 509142 43392 509148 43444
rect 509200 43432 509206 43444
rect 564434 43432 564440 43444
rect 509200 43404 564440 43432
rect 509200 43392 509206 43404
rect 564434 43392 564440 43404
rect 564492 43392 564498 43444
rect 3418 42712 3424 42764
rect 3476 42752 3482 42764
rect 60182 42752 60188 42764
rect 3476 42724 60188 42752
rect 3476 42712 3482 42724
rect 60182 42712 60188 42724
rect 60240 42712 60246 42764
rect 42702 42032 42708 42084
rect 42760 42072 42766 42084
rect 95326 42072 95332 42084
rect 42760 42044 95332 42072
rect 42760 42032 42766 42044
rect 95326 42032 95332 42044
rect 95384 42032 95390 42084
rect 106182 42032 106188 42084
rect 106240 42072 106246 42084
rect 145006 42072 145012 42084
rect 106240 42044 145012 42072
rect 106240 42032 106246 42044
rect 145006 42032 145012 42044
rect 145064 42032 145070 42084
rect 200485 42075 200543 42081
rect 200485 42041 200497 42075
rect 200531 42072 200543 42075
rect 201126 42072 201132 42084
rect 200531 42044 201132 42072
rect 200531 42041 200543 42044
rect 200485 42035 200543 42041
rect 201126 42032 201132 42044
rect 201184 42032 201190 42084
rect 511902 42032 511908 42084
rect 511960 42072 511966 42084
rect 568574 42072 568580 42084
rect 511960 42044 568580 42072
rect 511960 42032 511966 42044
rect 568574 42032 568580 42044
rect 568632 42032 568638 42084
rect 194778 41420 194784 41472
rect 194836 41460 194842 41472
rect 195422 41460 195428 41472
rect 194836 41432 195428 41460
rect 194836 41420 194842 41432
rect 195422 41420 195428 41432
rect 195480 41420 195486 41472
rect 489730 41420 489736 41472
rect 489788 41420 489794 41472
rect 62390 41352 62396 41404
rect 62448 41392 62454 41404
rect 63126 41392 63132 41404
rect 62448 41364 63132 41392
rect 62448 41352 62454 41364
rect 63126 41352 63132 41364
rect 63184 41352 63190 41404
rect 124214 41352 124220 41404
rect 124272 41392 124278 41404
rect 124398 41392 124404 41404
rect 124272 41364 124404 41392
rect 124272 41352 124278 41364
rect 124398 41352 124404 41364
rect 124456 41352 124462 41404
rect 296898 41352 296904 41404
rect 296956 41392 296962 41404
rect 297082 41392 297088 41404
rect 296956 41364 297088 41392
rect 296956 41352 296962 41364
rect 297082 41352 297088 41364
rect 297140 41352 297146 41404
rect 489748 41336 489776 41420
rect 489730 41284 489736 41336
rect 489788 41284 489794 41336
rect 49602 40672 49608 40724
rect 49660 40712 49666 40724
rect 100846 40712 100852 40724
rect 49660 40684 100852 40712
rect 49660 40672 49666 40684
rect 100846 40672 100852 40684
rect 100904 40672 100910 40724
rect 484210 40672 484216 40724
rect 484268 40712 484274 40724
rect 534074 40712 534080 40724
rect 484268 40684 534080 40712
rect 484268 40672 484274 40684
rect 534074 40672 534080 40684
rect 534132 40672 534138 40724
rect 523862 39992 523868 40044
rect 523920 40032 523926 40044
rect 580166 40032 580172 40044
rect 523920 40004 580172 40032
rect 523920 39992 523926 40004
rect 580166 39992 580172 40004
rect 580224 39992 580230 40044
rect 53742 39312 53748 39364
rect 53800 39352 53806 39364
rect 103606 39352 103612 39364
rect 53800 39324 103612 39352
rect 53800 39312 53806 39324
rect 103606 39312 103612 39324
rect 103664 39312 103670 39364
rect 74718 38632 74724 38684
rect 74776 38672 74782 38684
rect 74902 38672 74908 38684
rect 74776 38644 74908 38672
rect 74776 38632 74782 38644
rect 74902 38632 74908 38644
rect 74960 38632 74966 38684
rect 82814 38632 82820 38684
rect 82872 38672 82878 38684
rect 83734 38672 83740 38684
rect 82872 38644 83740 38672
rect 82872 38632 82878 38644
rect 83734 38632 83740 38644
rect 83792 38632 83798 38684
rect 85758 38672 85764 38684
rect 85719 38644 85764 38672
rect 85758 38632 85764 38644
rect 85816 38632 85822 38684
rect 132862 38632 132868 38684
rect 132920 38672 132926 38684
rect 133414 38672 133420 38684
rect 132920 38644 133420 38672
rect 132920 38632 132926 38644
rect 133414 38632 133420 38644
rect 133472 38632 133478 38684
rect 168745 38675 168803 38681
rect 168745 38641 168757 38675
rect 168791 38672 168803 38675
rect 168834 38672 168840 38684
rect 168791 38644 168840 38672
rect 168791 38641 168803 38644
rect 168745 38635 168803 38641
rect 168834 38632 168840 38644
rect 168892 38632 168898 38684
rect 489641 38675 489699 38681
rect 489641 38641 489653 38675
rect 489687 38672 489699 38675
rect 489822 38672 489828 38684
rect 489687 38644 489828 38672
rect 489687 38641 489699 38644
rect 489641 38635 489699 38641
rect 489822 38632 489828 38644
rect 489880 38632 489886 38684
rect 109402 38604 109408 38616
rect 109363 38576 109408 38604
rect 109402 38564 109408 38576
rect 109460 38564 109466 38616
rect 124309 38607 124367 38613
rect 124309 38573 124321 38607
rect 124355 38604 124367 38607
rect 124398 38604 124404 38616
rect 124355 38576 124404 38604
rect 124355 38573 124367 38576
rect 124309 38567 124367 38573
rect 124398 38564 124404 38576
rect 124456 38564 124462 38616
rect 197446 38604 197452 38616
rect 197407 38576 197452 38604
rect 197446 38564 197452 38576
rect 197504 38564 197510 38616
rect 203153 38607 203211 38613
rect 203153 38573 203165 38607
rect 203199 38604 203211 38607
rect 203242 38604 203248 38616
rect 203199 38576 203248 38604
rect 203199 38573 203211 38576
rect 203153 38567 203211 38573
rect 203242 38564 203248 38576
rect 203300 38564 203306 38616
rect 291378 38604 291384 38616
rect 291339 38576 291384 38604
rect 291378 38564 291384 38576
rect 291436 38564 291442 38616
rect 487154 38604 487160 38616
rect 487115 38576 487160 38604
rect 487154 38564 487160 38576
rect 487212 38564 487218 38616
rect 56410 37884 56416 37936
rect 56468 37924 56474 37936
rect 106366 37924 106372 37936
rect 56468 37896 106372 37924
rect 56468 37884 56474 37896
rect 106366 37884 106372 37896
rect 106424 37884 106430 37936
rect 486970 37884 486976 37936
rect 487028 37924 487034 37936
rect 536834 37924 536840 37936
rect 487028 37896 536840 37924
rect 487028 37884 487034 37896
rect 536834 37884 536840 37896
rect 536892 37884 536898 37936
rect 293954 37312 293960 37324
rect 293915 37284 293960 37312
rect 293954 37272 293960 37284
rect 294012 37272 294018 37324
rect 290826 37136 290832 37188
rect 290884 37176 290890 37188
rect 291013 37179 291071 37185
rect 291013 37176 291025 37179
rect 290884 37148 291025 37176
rect 290884 37136 290890 37148
rect 291013 37145 291025 37148
rect 291059 37145 291071 37179
rect 291013 37139 291071 37145
rect 14458 36524 14464 36576
rect 14516 36564 14522 36576
rect 72050 36564 72056 36576
rect 14516 36536 72056 36564
rect 14516 36524 14522 36536
rect 72050 36524 72056 36536
rect 72108 36524 72114 36576
rect 288158 36524 288164 36576
rect 288216 36564 288222 36576
rect 288342 36564 288348 36576
rect 288216 36536 288348 36564
rect 288216 36524 288222 36536
rect 288342 36524 288348 36536
rect 288400 36524 288406 36576
rect 492490 36524 492496 36576
rect 492548 36564 492554 36576
rect 545114 36564 545120 36576
rect 492548 36536 545120 36564
rect 492548 36524 492554 36536
rect 545114 36524 545120 36536
rect 545172 36524 545178 36576
rect 98086 35912 98092 35964
rect 98144 35952 98150 35964
rect 98270 35952 98276 35964
rect 98144 35924 98276 35952
rect 98144 35912 98150 35924
rect 98270 35912 98276 35924
rect 98328 35912 98334 35964
rect 19978 35164 19984 35216
rect 20036 35204 20042 35216
rect 75914 35204 75920 35216
rect 20036 35176 75920 35204
rect 20036 35164 20042 35176
rect 75914 35164 75920 35176
rect 75972 35164 75978 35216
rect 498010 35164 498016 35216
rect 498068 35204 498074 35216
rect 552014 35204 552020 35216
rect 498068 35176 552020 35204
rect 498068 35164 498074 35176
rect 552014 35164 552020 35176
rect 552072 35164 552078 35216
rect 28902 33736 28908 33788
rect 28960 33776 28966 33788
rect 82814 33776 82820 33788
rect 28960 33748 82820 33776
rect 28960 33736 28966 33748
rect 82814 33736 82820 33748
rect 82872 33736 82878 33788
rect 433242 33736 433248 33788
rect 433300 33776 433306 33788
rect 469214 33776 469220 33788
rect 433300 33748 469220 33776
rect 433300 33736 433306 33748
rect 469214 33736 469220 33748
rect 469272 33736 469278 33788
rect 507670 33736 507676 33788
rect 507728 33776 507734 33788
rect 563146 33776 563152 33788
rect 507728 33748 563152 33776
rect 507728 33736 507734 33748
rect 563146 33736 563152 33748
rect 563204 33736 563210 33788
rect 31662 32376 31668 32428
rect 31720 32416 31726 32428
rect 85758 32416 85764 32428
rect 31720 32388 85764 32416
rect 31720 32376 31726 32388
rect 85758 32376 85764 32388
rect 85816 32376 85822 32428
rect 96522 32376 96528 32428
rect 96580 32416 96586 32428
rect 136726 32416 136732 32428
rect 96580 32388 136732 32416
rect 96580 32376 96586 32388
rect 136726 32376 136732 32388
rect 136784 32376 136790 32428
rect 430390 32376 430396 32428
rect 430448 32416 430454 32428
rect 466454 32416 466460 32428
rect 430448 32388 466460 32416
rect 430448 32376 430454 32388
rect 466454 32376 466460 32388
rect 466512 32376 466518 32428
rect 489638 31696 489644 31748
rect 489696 31736 489702 31748
rect 489822 31736 489828 31748
rect 489696 31708 489828 31736
rect 489696 31696 489702 31708
rect 489822 31696 489828 31708
rect 489880 31696 489886 31748
rect 495066 31696 495072 31748
rect 495124 31736 495130 31748
rect 495250 31736 495256 31748
rect 495124 31708 495256 31736
rect 495124 31696 495130 31708
rect 495250 31696 495256 31708
rect 495308 31696 495314 31748
rect 197446 31600 197452 31612
rect 197407 31572 197452 31600
rect 197446 31560 197452 31572
rect 197504 31560 197510 31612
rect 200482 31600 200488 31612
rect 200443 31572 200488 31600
rect 200482 31560 200488 31572
rect 200540 31560 200546 31612
rect 35802 31016 35808 31068
rect 35860 31056 35866 31068
rect 88334 31056 88340 31068
rect 35860 31028 88340 31056
rect 35860 31016 35866 31028
rect 88334 31016 88340 31028
rect 88392 31016 88398 31068
rect 89622 31016 89628 31068
rect 89680 31056 89686 31068
rect 131114 31056 131120 31068
rect 89680 31028 131120 31056
rect 89680 31016 89686 31028
rect 131114 31016 131120 31028
rect 131172 31016 131178 31068
rect 427722 31016 427728 31068
rect 427780 31056 427786 31068
rect 462314 31056 462320 31068
rect 427780 31028 462320 31056
rect 427780 31016 427786 31028
rect 462314 31016 462320 31028
rect 462372 31016 462378 31068
rect 478782 31016 478788 31068
rect 478840 31056 478846 31068
rect 527174 31056 527180 31068
rect 478840 31028 527180 31056
rect 478840 31016 478846 31028
rect 527174 31016 527180 31028
rect 527232 31016 527238 31068
rect 85482 29656 85488 29708
rect 85540 29696 85546 29708
rect 128354 29696 128360 29708
rect 85540 29668 128360 29696
rect 85540 29656 85546 29668
rect 128354 29656 128360 29668
rect 128412 29656 128418 29708
rect 38562 29588 38568 29640
rect 38620 29628 38626 29640
rect 92566 29628 92572 29640
rect 38620 29600 92572 29628
rect 38620 29588 38626 29600
rect 92566 29588 92572 29600
rect 92624 29588 92630 29640
rect 422110 29588 422116 29640
rect 422168 29628 422174 29640
rect 455414 29628 455420 29640
rect 422168 29600 455420 29628
rect 422168 29588 422174 29600
rect 455414 29588 455420 29600
rect 455472 29588 455478 29640
rect 489730 29588 489736 29640
rect 489788 29628 489794 29640
rect 540974 29628 540980 29640
rect 489788 29600 540980 29628
rect 489788 29588 489794 29600
rect 540974 29588 540980 29600
rect 541032 29588 541038 29640
rect 109405 29019 109463 29025
rect 109405 28985 109417 29019
rect 109451 29016 109463 29019
rect 109494 29016 109500 29028
rect 109451 28988 109500 29016
rect 109451 28985 109463 28988
rect 109405 28979 109463 28985
rect 109494 28976 109500 28988
rect 109552 28976 109558 29028
rect 124306 29016 124312 29028
rect 124267 28988 124312 29016
rect 124306 28976 124312 28988
rect 124364 28976 124370 29028
rect 203150 29016 203156 29028
rect 203111 28988 203156 29016
rect 203150 28976 203156 28988
rect 203208 28976 203214 29028
rect 291381 29019 291439 29025
rect 291381 28985 291393 29019
rect 291427 29016 291439 29019
rect 291470 29016 291476 29028
rect 291427 28988 291476 29016
rect 291427 28985 291439 28988
rect 291381 28979 291439 28985
rect 291470 28976 291476 28988
rect 291528 28976 291534 29028
rect 296990 28976 296996 29028
rect 297048 29016 297054 29028
rect 297082 29016 297088 29028
rect 297048 28988 297088 29016
rect 297048 28976 297054 28988
rect 297082 28976 297088 28988
rect 297140 28976 297146 29028
rect 487154 29016 487160 29028
rect 487115 28988 487160 29016
rect 487154 28976 487160 28988
rect 487212 28976 487218 29028
rect 62298 28948 62304 28960
rect 62259 28920 62304 28948
rect 62298 28908 62304 28920
rect 62356 28908 62362 28960
rect 438118 28948 438124 28960
rect 438079 28920 438124 28948
rect 438118 28908 438124 28920
rect 438176 28908 438182 28960
rect 82722 28228 82728 28280
rect 82780 28268 82786 28280
rect 125594 28268 125600 28280
rect 82780 28240 125600 28268
rect 82780 28228 82786 28240
rect 125594 28228 125600 28240
rect 125652 28228 125658 28280
rect 422938 28228 422944 28280
rect 422996 28268 423002 28280
rect 451274 28268 451280 28280
rect 422996 28240 451280 28268
rect 422996 28228 423002 28240
rect 451274 28228 451280 28240
rect 451332 28228 451338 28280
rect 470502 28228 470508 28280
rect 470560 28268 470566 28280
rect 516134 28268 516140 28280
rect 470560 28240 516140 28268
rect 470560 28228 470566 28240
rect 516134 28228 516140 28240
rect 516192 28228 516198 28280
rect 80146 27616 80152 27668
rect 80204 27656 80210 27668
rect 80238 27656 80244 27668
rect 80204 27628 80244 27656
rect 80204 27616 80210 27628
rect 80238 27616 80244 27628
rect 80296 27616 80302 27668
rect 291010 27656 291016 27668
rect 290971 27628 291016 27656
rect 291010 27616 291016 27628
rect 291068 27616 291074 27668
rect 293954 27588 293960 27600
rect 293915 27560 293960 27588
rect 293954 27548 293960 27560
rect 294012 27548 294018 27600
rect 296990 27548 296996 27600
rect 297048 27588 297054 27600
rect 297082 27588 297088 27600
rect 297048 27560 297088 27588
rect 297048 27548 297054 27560
rect 297082 27548 297088 27560
rect 297140 27548 297146 27600
rect 78582 26868 78588 26920
rect 78640 26908 78646 26920
rect 122834 26908 122840 26920
rect 78640 26880 122840 26908
rect 78640 26868 78646 26880
rect 122834 26868 122840 26880
rect 122892 26868 122898 26920
rect 124122 26868 124128 26920
rect 124180 26908 124186 26920
rect 158714 26908 158720 26920
rect 124180 26880 158720 26908
rect 124180 26868 124186 26880
rect 158714 26868 158720 26880
rect 158772 26868 158778 26920
rect 416590 26868 416596 26920
rect 416648 26908 416654 26920
rect 448514 26908 448520 26920
rect 416648 26880 448520 26908
rect 416648 26868 416654 26880
rect 448514 26868 448520 26880
rect 448572 26868 448578 26920
rect 464338 26868 464344 26920
rect 464396 26908 464402 26920
rect 505094 26908 505100 26920
rect 464396 26880 505100 26908
rect 464396 26868 464402 26880
rect 505094 26868 505100 26880
rect 505152 26868 505158 26920
rect 150802 26256 150808 26308
rect 150860 26296 150866 26308
rect 150894 26296 150900 26308
rect 150860 26268 150900 26296
rect 150860 26256 150866 26268
rect 150894 26256 150900 26268
rect 150952 26256 150958 26308
rect 3418 26188 3424 26240
rect 3476 26228 3482 26240
rect 60090 26228 60096 26240
rect 3476 26200 60096 26228
rect 3476 26188 3482 26200
rect 60090 26188 60096 26200
rect 60148 26188 60154 26240
rect 74442 25508 74448 25560
rect 74500 25548 74506 25560
rect 120074 25548 120080 25560
rect 74500 25520 120080 25548
rect 74500 25508 74506 25520
rect 120074 25508 120080 25520
rect 120132 25508 120138 25560
rect 140682 25508 140688 25560
rect 140740 25548 140746 25560
rect 171134 25548 171140 25560
rect 140740 25520 171140 25548
rect 140740 25508 140746 25520
rect 171134 25508 171140 25520
rect 171192 25508 171198 25560
rect 413830 25508 413836 25560
rect 413888 25548 413894 25560
rect 444374 25548 444380 25560
rect 413888 25520 444380 25548
rect 413888 25508 413894 25520
rect 444374 25508 444380 25520
rect 444432 25508 444438 25560
rect 459462 25508 459468 25560
rect 459520 25548 459526 25560
rect 502426 25548 502432 25560
rect 459520 25520 502432 25548
rect 459520 25508 459526 25520
rect 502426 25508 502432 25520
rect 502484 25508 502490 25560
rect 503622 25508 503628 25560
rect 503680 25548 503686 25560
rect 558914 25548 558920 25560
rect 503680 25520 558920 25548
rect 503680 25508 503686 25520
rect 558914 25508 558920 25520
rect 558972 25508 558978 25560
rect 523770 24760 523776 24812
rect 523828 24800 523834 24812
rect 580166 24800 580172 24812
rect 523828 24772 580172 24800
rect 523828 24760 523834 24772
rect 580166 24760 580172 24772
rect 580224 24760 580230 24812
rect 200298 24148 200304 24200
rect 200356 24188 200362 24200
rect 200482 24188 200488 24200
rect 200356 24160 200488 24188
rect 200356 24148 200362 24160
rect 200482 24148 200488 24160
rect 200540 24148 200546 24200
rect 67542 24080 67548 24132
rect 67600 24120 67606 24132
rect 114554 24120 114560 24132
rect 67600 24092 114560 24120
rect 67600 24080 67606 24092
rect 114554 24080 114560 24092
rect 114612 24080 114618 24132
rect 136542 24080 136548 24132
rect 136600 24120 136606 24132
rect 168834 24120 168840 24132
rect 136600 24092 168840 24120
rect 136600 24080 136606 24092
rect 168834 24080 168840 24092
rect 168892 24080 168898 24132
rect 411162 24080 411168 24132
rect 411220 24120 411226 24132
rect 441614 24120 441620 24132
rect 411220 24092 441620 24120
rect 411220 24080 411226 24092
rect 441614 24080 441620 24092
rect 441672 24080 441678 24132
rect 451918 24080 451924 24132
rect 451976 24120 451982 24132
rect 491294 24120 491300 24132
rect 451976 24092 491300 24120
rect 451976 24080 451982 24092
rect 491294 24080 491300 24092
rect 491352 24080 491358 24132
rect 445570 22788 445576 22840
rect 445628 22828 445634 22840
rect 484394 22828 484400 22840
rect 445628 22800 484400 22828
rect 445628 22788 445634 22800
rect 484394 22788 484400 22800
rect 484452 22788 484458 22840
rect 23382 22720 23388 22772
rect 23440 22760 23446 22772
rect 79318 22760 79324 22772
rect 23440 22732 79324 22760
rect 23440 22720 23446 22732
rect 79318 22720 79324 22732
rect 79376 22720 79382 22772
rect 91002 22720 91008 22772
rect 91060 22760 91066 22772
rect 132862 22760 132868 22772
rect 91060 22732 132868 22760
rect 91060 22720 91066 22732
rect 132862 22720 132868 22732
rect 132920 22720 132926 22772
rect 133782 22720 133788 22772
rect 133840 22760 133846 22772
rect 165614 22760 165620 22772
rect 133840 22732 165620 22760
rect 133840 22720 133846 22732
rect 165614 22720 165620 22732
rect 165672 22720 165678 22772
rect 368382 22720 368388 22772
rect 368440 22760 368446 22772
rect 386414 22760 386420 22772
rect 368440 22732 386420 22760
rect 368440 22720 368446 22732
rect 386414 22720 386420 22732
rect 386472 22720 386478 22772
rect 402882 22720 402888 22772
rect 402940 22760 402946 22772
rect 430574 22760 430580 22772
rect 402940 22732 430580 22760
rect 402940 22720 402946 22732
rect 430574 22720 430580 22732
rect 430632 22720 430638 22772
rect 481542 22720 481548 22772
rect 481600 22760 481606 22772
rect 529934 22760 529940 22772
rect 481600 22732 529940 22760
rect 481600 22720 481606 22732
rect 529934 22720 529940 22732
rect 529992 22720 529998 22772
rect 74718 22352 74724 22364
rect 74679 22324 74724 22352
rect 74718 22312 74724 22324
rect 74776 22312 74782 22364
rect 124306 22108 124312 22160
rect 124364 22108 124370 22160
rect 150618 22108 150624 22160
rect 150676 22148 150682 22160
rect 150805 22151 150863 22157
rect 150805 22148 150817 22151
rect 150676 22120 150817 22148
rect 150676 22108 150682 22120
rect 150805 22117 150817 22120
rect 150851 22117 150863 22151
rect 150805 22111 150863 22117
rect 495250 22108 495256 22160
rect 495308 22108 495314 22160
rect 124324 22024 124352 22108
rect 202966 22040 202972 22092
rect 203024 22080 203030 22092
rect 203150 22080 203156 22092
rect 203024 22052 203156 22080
rect 203024 22040 203030 22052
rect 203150 22040 203156 22052
rect 203208 22040 203214 22092
rect 291286 22040 291292 22092
rect 291344 22080 291350 22092
rect 291470 22080 291476 22092
rect 291344 22052 291476 22080
rect 291344 22040 291350 22052
rect 291470 22040 291476 22052
rect 291528 22040 291534 22092
rect 495268 22024 495296 22108
rect 124306 21972 124312 22024
rect 124364 21972 124370 22024
rect 495250 21972 495256 22024
rect 495308 21972 495314 22024
rect 146202 21428 146208 21480
rect 146260 21468 146266 21480
rect 176746 21468 176752 21480
rect 146260 21440 176752 21468
rect 146260 21428 146266 21440
rect 176746 21428 176752 21440
rect 176804 21428 176810 21480
rect 438762 21428 438768 21480
rect 438820 21468 438826 21480
rect 476114 21468 476120 21480
rect 438820 21440 476120 21468
rect 438820 21428 438826 21440
rect 476114 21428 476120 21440
rect 476172 21428 476178 21480
rect 60642 21360 60648 21412
rect 60700 21400 60706 21412
rect 108298 21400 108304 21412
rect 60700 21372 108304 21400
rect 60700 21360 60706 21372
rect 108298 21360 108304 21372
rect 108356 21360 108362 21412
rect 108942 21360 108948 21412
rect 109000 21400 109006 21412
rect 146938 21400 146944 21412
rect 109000 21372 146944 21400
rect 109000 21360 109006 21372
rect 146938 21360 146944 21372
rect 146996 21360 147002 21412
rect 410518 21360 410524 21412
rect 410576 21400 410582 21412
rect 437474 21400 437480 21412
rect 410576 21372 437480 21400
rect 410576 21360 410582 21372
rect 437474 21360 437480 21372
rect 437532 21360 437538 21412
rect 476022 21360 476028 21412
rect 476080 21400 476086 21412
rect 523034 21400 523040 21412
rect 476080 21372 523040 21400
rect 476080 21360 476086 21372
rect 523034 21360 523040 21372
rect 523092 21360 523098 21412
rect 64690 19932 64696 19984
rect 64748 19972 64754 19984
rect 111058 19972 111064 19984
rect 64748 19944 111064 19972
rect 64748 19932 64754 19944
rect 111058 19932 111064 19944
rect 111116 19932 111122 19984
rect 142062 19932 142068 19984
rect 142120 19972 142126 19984
rect 173986 19972 173992 19984
rect 142120 19944 173992 19972
rect 142120 19932 142126 19944
rect 173986 19932 173992 19944
rect 174044 19932 174050 19984
rect 405642 19932 405648 19984
rect 405700 19972 405706 19984
rect 433334 19972 433340 19984
rect 405700 19944 433340 19972
rect 405700 19932 405706 19944
rect 433334 19932 433340 19944
rect 433392 19932 433398 19984
rect 433978 19932 433984 19984
rect 434036 19972 434042 19984
rect 467926 19972 467932 19984
rect 434036 19944 467932 19972
rect 434036 19932 434042 19944
rect 467926 19932 467932 19944
rect 467984 19932 467990 19984
rect 475378 19932 475384 19984
rect 475436 19972 475442 19984
rect 520366 19972 520372 19984
rect 475436 19944 520372 19972
rect 475436 19932 475442 19944
rect 520366 19932 520372 19944
rect 520424 19932 520430 19984
rect 62301 19363 62359 19369
rect 62301 19329 62313 19363
rect 62347 19360 62359 19363
rect 62482 19360 62488 19372
rect 62347 19332 62488 19360
rect 62347 19329 62359 19332
rect 62301 19323 62359 19329
rect 62482 19320 62488 19332
rect 62540 19320 62546 19372
rect 74718 19360 74724 19372
rect 74679 19332 74724 19360
rect 74718 19320 74724 19332
rect 74776 19320 74782 19372
rect 109310 19320 109316 19372
rect 109368 19360 109374 19372
rect 109402 19360 109408 19372
rect 109368 19332 109408 19360
rect 109368 19320 109374 19332
rect 109402 19320 109408 19332
rect 109460 19320 109466 19372
rect 438121 19363 438179 19369
rect 438121 19329 438133 19363
rect 438167 19360 438179 19363
rect 438302 19360 438308 19372
rect 438167 19332 438308 19360
rect 438167 19329 438179 19332
rect 438121 19323 438179 19329
rect 438302 19320 438308 19332
rect 438360 19320 438366 19372
rect 147769 19295 147827 19301
rect 147769 19261 147781 19295
rect 147815 19292 147827 19295
rect 147858 19292 147864 19304
rect 147815 19264 147864 19292
rect 147815 19261 147827 19264
rect 147769 19255 147827 19261
rect 147858 19252 147864 19264
rect 147916 19252 147922 19304
rect 203150 19292 203156 19304
rect 203111 19264 203156 19292
rect 203150 19252 203156 19264
rect 203208 19252 203214 19304
rect 487154 19292 487160 19304
rect 487115 19264 487160 19292
rect 487154 19252 487160 19264
rect 487212 19252 487218 19304
rect 430482 18640 430488 18692
rect 430540 18680 430546 18692
rect 465074 18680 465080 18692
rect 430540 18652 465080 18680
rect 430540 18640 430546 18652
rect 465074 18640 465080 18652
rect 465132 18640 465138 18692
rect 10410 18572 10416 18624
rect 10468 18612 10474 18624
rect 69106 18612 69112 18624
rect 10468 18584 69112 18612
rect 10468 18572 10474 18584
rect 69106 18572 69112 18584
rect 69164 18572 69170 18624
rect 71682 18572 71688 18624
rect 71740 18612 71746 18624
rect 117314 18612 117320 18624
rect 71740 18584 117320 18612
rect 71740 18572 71746 18584
rect 117314 18572 117320 18584
rect 117372 18572 117378 18624
rect 135162 18572 135168 18624
rect 135220 18612 135226 18624
rect 168374 18612 168380 18624
rect 135220 18584 168380 18612
rect 135220 18572 135226 18584
rect 168374 18572 168380 18584
rect 168432 18572 168438 18624
rect 290642 18572 290648 18624
rect 290700 18612 290706 18624
rect 291102 18612 291108 18624
rect 290700 18584 291108 18612
rect 290700 18572 290706 18584
rect 291102 18572 291108 18584
rect 291160 18572 291166 18624
rect 400122 18572 400128 18624
rect 400180 18612 400186 18624
rect 426434 18612 426440 18624
rect 400180 18584 426440 18612
rect 400180 18572 400186 18584
rect 426434 18572 426440 18584
rect 426492 18572 426498 18624
rect 464982 18572 464988 18624
rect 465040 18612 465046 18624
rect 509234 18612 509240 18624
rect 465040 18584 509240 18612
rect 465040 18572 465046 18584
rect 509234 18572 509240 18584
rect 509292 18572 509298 18624
rect 293954 18000 293960 18012
rect 293915 17972 293960 18000
rect 293954 17960 293960 17972
rect 294012 17960 294018 18012
rect 424870 17280 424876 17332
rect 424928 17320 424934 17332
rect 458174 17320 458180 17332
rect 424928 17292 458180 17320
rect 424928 17280 424934 17292
rect 458174 17280 458180 17292
rect 458232 17280 458238 17332
rect 45462 17212 45468 17264
rect 45520 17252 45526 17264
rect 96614 17252 96620 17264
rect 45520 17224 96620 17252
rect 45520 17212 45526 17224
rect 96614 17212 96620 17224
rect 96672 17212 96678 17264
rect 128262 17212 128268 17264
rect 128320 17252 128326 17264
rect 162118 17252 162124 17264
rect 128320 17224 162124 17252
rect 128320 17212 128326 17224
rect 162118 17212 162124 17224
rect 162176 17212 162182 17264
rect 164142 17212 164148 17264
rect 164200 17252 164206 17264
rect 190454 17252 190460 17264
rect 164200 17224 190460 17252
rect 164200 17212 164206 17224
rect 190454 17212 190460 17224
rect 190512 17212 190518 17264
rect 399478 17212 399484 17264
rect 399536 17252 399542 17264
rect 423674 17252 423680 17264
rect 399536 17224 423680 17252
rect 399536 17212 399542 17224
rect 423674 17212 423680 17224
rect 423732 17212 423738 17264
rect 453850 17212 453856 17264
rect 453908 17252 453914 17264
rect 494054 17252 494060 17264
rect 453908 17224 494060 17252
rect 453908 17212 453914 17224
rect 494054 17212 494060 17224
rect 494112 17212 494118 17264
rect 496078 17212 496084 17264
rect 496136 17252 496142 17264
rect 547874 17252 547880 17264
rect 496136 17224 547880 17252
rect 496136 17212 496142 17224
rect 547874 17212 547880 17224
rect 547932 17212 547938 17264
rect 98086 16600 98092 16652
rect 98144 16640 98150 16652
rect 98270 16640 98276 16652
rect 98144 16612 98276 16640
rect 98144 16600 98150 16612
rect 98270 16600 98276 16612
rect 98328 16600 98334 16652
rect 41322 15852 41328 15904
rect 41380 15892 41386 15904
rect 93854 15892 93860 15904
rect 41380 15864 93860 15892
rect 41380 15852 41386 15864
rect 93854 15852 93860 15864
rect 93912 15852 93918 15904
rect 102042 15852 102048 15904
rect 102100 15892 102106 15904
rect 142246 15892 142252 15904
rect 102100 15864 142252 15892
rect 102100 15852 102106 15864
rect 142246 15852 142252 15864
rect 142304 15852 142310 15904
rect 159910 15852 159916 15904
rect 159968 15892 159974 15904
rect 186406 15892 186412 15904
rect 159968 15864 186412 15892
rect 159968 15852 159974 15864
rect 186406 15852 186412 15864
rect 186464 15852 186470 15904
rect 394602 15852 394608 15904
rect 394660 15892 394666 15904
rect 419534 15892 419540 15904
rect 394660 15864 419540 15892
rect 394660 15852 394666 15864
rect 419534 15852 419540 15864
rect 419592 15852 419598 15904
rect 420178 15852 420184 15904
rect 420236 15892 420242 15904
rect 451366 15892 451372 15904
rect 420236 15864 451372 15892
rect 420236 15852 420242 15864
rect 451366 15852 451372 15864
rect 451424 15852 451430 15904
rect 469858 15852 469864 15904
rect 469916 15892 469922 15904
rect 514754 15892 514760 15904
rect 469916 15864 514760 15892
rect 469916 15852 469922 15864
rect 514754 15852 514760 15864
rect 514812 15852 514818 15904
rect 404170 14492 404176 14544
rect 404228 14532 404234 14544
rect 433426 14532 433432 14544
rect 404228 14504 433432 14532
rect 404228 14492 404234 14504
rect 433426 14492 433432 14504
rect 433484 14492 433490 14544
rect 38470 14424 38476 14476
rect 38528 14464 38534 14476
rect 91094 14464 91100 14476
rect 38528 14436 91100 14464
rect 38528 14424 38534 14436
rect 91094 14424 91100 14436
rect 91152 14424 91158 14476
rect 99282 14424 99288 14476
rect 99340 14464 99346 14476
rect 139486 14464 139492 14476
rect 99340 14436 139492 14464
rect 99340 14424 99346 14436
rect 139486 14424 139492 14436
rect 139544 14424 139550 14476
rect 151722 14424 151728 14476
rect 151780 14464 151786 14476
rect 180794 14464 180800 14476
rect 151780 14436 180800 14464
rect 151780 14424 151786 14436
rect 180794 14424 180800 14436
rect 180852 14424 180858 14476
rect 424962 14424 424968 14476
rect 425020 14464 425026 14476
rect 459646 14464 459652 14476
rect 425020 14436 459652 14464
rect 425020 14424 425026 14436
rect 459646 14424 459652 14436
rect 459704 14424 459710 14476
rect 463510 14424 463516 14476
rect 463568 14464 463574 14476
rect 507854 14464 507860 14476
rect 463568 14436 507860 14464
rect 463568 14424 463574 14436
rect 507854 14424 507860 14436
rect 507912 14424 507918 14476
rect 510430 14424 510436 14476
rect 510488 14464 510494 14476
rect 565814 14464 565820 14476
rect 510488 14436 565820 14464
rect 510488 14424 510494 14436
rect 565814 14424 565820 14436
rect 565872 14424 565878 14476
rect 395890 13132 395896 13184
rect 395948 13172 395954 13184
rect 422294 13172 422300 13184
rect 395948 13144 422300 13172
rect 395948 13132 395954 13144
rect 422294 13132 422300 13144
rect 422352 13132 422358 13184
rect 460750 13132 460756 13184
rect 460808 13172 460814 13184
rect 503714 13172 503720 13184
rect 460808 13144 503720 13172
rect 460808 13132 460814 13144
rect 503714 13132 503720 13144
rect 503772 13132 503778 13184
rect 30282 13064 30288 13116
rect 30340 13104 30346 13116
rect 85574 13104 85580 13116
rect 30340 13076 85580 13104
rect 30340 13064 30346 13076
rect 85574 13064 85580 13076
rect 85632 13064 85638 13116
rect 95142 13064 95148 13116
rect 95200 13104 95206 13116
rect 136634 13104 136640 13116
rect 95200 13076 136640 13104
rect 95200 13064 95206 13076
rect 136634 13064 136640 13076
rect 136692 13064 136698 13116
rect 148962 13064 148968 13116
rect 149020 13104 149026 13116
rect 178034 13104 178040 13116
rect 149020 13076 178040 13104
rect 149020 13064 149026 13076
rect 178034 13064 178040 13076
rect 178092 13064 178098 13116
rect 187602 13064 187608 13116
rect 187660 13104 187666 13116
rect 209038 13104 209044 13116
rect 187660 13076 209044 13104
rect 187660 13064 187666 13076
rect 209038 13064 209044 13076
rect 209096 13064 209102 13116
rect 422202 13064 422208 13116
rect 422260 13104 422266 13116
rect 454034 13104 454040 13116
rect 422260 13076 454040 13104
rect 422260 13064 422266 13076
rect 454034 13064 454040 13076
rect 454092 13064 454098 13116
rect 500862 13064 500868 13116
rect 500920 13104 500926 13116
rect 554866 13104 554872 13116
rect 500920 13076 554872 13104
rect 500920 13064 500926 13076
rect 554866 13064 554872 13076
rect 554924 13064 554930 13116
rect 80054 12384 80060 12436
rect 80112 12424 80118 12436
rect 80422 12424 80428 12436
rect 80112 12396 80428 12424
rect 80112 12384 80118 12396
rect 80422 12384 80428 12396
rect 80480 12384 80486 12436
rect 300946 12248 300952 12300
rect 301004 12288 301010 12300
rect 301406 12288 301412 12300
rect 301004 12260 301412 12288
rect 301004 12248 301010 12260
rect 301406 12248 301412 12260
rect 301464 12248 301470 12300
rect 513190 11976 513196 12028
rect 513248 11976 513254 12028
rect 513208 11812 513236 11976
rect 513282 11812 513288 11824
rect 513208 11784 513288 11812
rect 513282 11772 513288 11784
rect 513340 11772 513346 11824
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 67634 11744 67640 11756
rect 9088 11716 67640 11744
rect 9088 11704 9094 11716
rect 67634 11704 67640 11716
rect 67692 11704 67698 11756
rect 84102 11704 84108 11756
rect 84160 11744 84166 11756
rect 126238 11744 126244 11756
rect 84160 11716 126244 11744
rect 84160 11704 84166 11716
rect 126238 11704 126244 11716
rect 126296 11704 126302 11756
rect 144822 11704 144828 11756
rect 144880 11744 144886 11756
rect 175274 11744 175280 11756
rect 144880 11716 175280 11744
rect 144880 11704 144886 11716
rect 175274 11704 175280 11716
rect 175332 11704 175338 11756
rect 180702 11704 180708 11756
rect 180760 11744 180766 11756
rect 203153 11747 203211 11753
rect 203153 11744 203165 11747
rect 180760 11716 203165 11744
rect 180760 11704 180766 11716
rect 203153 11713 203165 11716
rect 203199 11713 203211 11747
rect 203153 11707 203211 11713
rect 387702 11704 387708 11756
rect 387760 11744 387766 11756
rect 411254 11744 411260 11756
rect 387760 11716 411260 11744
rect 387760 11704 387766 11716
rect 411254 11704 411260 11716
rect 411312 11704 411318 11756
rect 413922 11704 413928 11756
rect 413980 11744 413986 11756
rect 443086 11744 443092 11756
rect 413980 11716 443092 11744
rect 413980 11704 413986 11716
rect 443086 11704 443092 11716
rect 443144 11704 443150 11756
rect 458082 11704 458088 11756
rect 458140 11744 458146 11756
rect 500954 11744 500960 11756
rect 458140 11716 500960 11744
rect 458140 11704 458146 11716
rect 500954 11704 500960 11716
rect 501012 11704 501018 11756
rect 517422 11704 517428 11756
rect 517480 11744 517486 11756
rect 574738 11744 574744 11756
rect 517480 11716 574744 11744
rect 517480 11704 517486 11716
rect 574738 11704 574744 11716
rect 574796 11704 574802 11756
rect 4062 10276 4068 10328
rect 4120 10316 4126 10328
rect 63494 10316 63500 10328
rect 4120 10288 63500 10316
rect 4120 10276 4126 10288
rect 63494 10276 63500 10288
rect 63552 10276 63558 10328
rect 80238 10276 80244 10328
rect 80296 10316 80302 10328
rect 124398 10316 124404 10328
rect 80296 10288 124404 10316
rect 80296 10276 80302 10288
rect 124398 10276 124404 10288
rect 124456 10276 124462 10328
rect 141970 10276 141976 10328
rect 142028 10316 142034 10328
rect 172514 10316 172520 10328
rect 142028 10288 172520 10316
rect 142028 10276 142034 10288
rect 172514 10276 172520 10288
rect 172572 10276 172578 10328
rect 176562 10276 176568 10328
rect 176620 10316 176626 10328
rect 200390 10316 200396 10328
rect 176620 10288 200396 10316
rect 176620 10276 176626 10288
rect 200390 10276 200396 10288
rect 200448 10276 200454 10328
rect 384942 10276 384948 10328
rect 385000 10316 385006 10328
rect 408586 10316 408592 10328
rect 385000 10288 408592 10316
rect 385000 10276 385006 10288
rect 408586 10276 408592 10288
rect 408644 10276 408650 10328
rect 409690 10276 409696 10328
rect 409748 10316 409754 10328
rect 440234 10316 440240 10328
rect 409748 10288 440240 10316
rect 409748 10276 409754 10288
rect 440234 10276 440240 10288
rect 440292 10276 440298 10328
rect 452562 10276 452568 10328
rect 452620 10316 452626 10328
rect 494146 10316 494152 10328
rect 452620 10288 494152 10316
rect 452620 10276 452626 10288
rect 494146 10276 494152 10288
rect 494204 10276 494210 10328
rect 520182 10276 520188 10328
rect 520240 10316 520246 10328
rect 579614 10316 579620 10328
rect 520240 10288 579620 10316
rect 520240 10276 520246 10288
rect 579614 10276 579620 10288
rect 579672 10276 579678 10328
rect 147766 9704 147772 9716
rect 147727 9676 147772 9704
rect 147766 9664 147772 9676
rect 147824 9664 147830 9716
rect 150802 9704 150808 9716
rect 150763 9676 150808 9704
rect 150802 9664 150808 9676
rect 150860 9664 150866 9716
rect 487154 9704 487160 9716
rect 487115 9676 487160 9704
rect 487154 9664 487160 9676
rect 487212 9664 487218 9716
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 59998 9636 60004 9648
rect 3476 9608 60004 9636
rect 3476 9596 3482 9608
rect 59998 9596 60004 9608
rect 60056 9596 60062 9648
rect 119430 8984 119436 9036
rect 119488 9024 119494 9036
rect 156046 9024 156052 9036
rect 119488 8996 156052 9024
rect 119488 8984 119494 8996
rect 156046 8984 156052 8996
rect 156104 8984 156110 9036
rect 449802 8984 449808 9036
rect 449860 9024 449866 9036
rect 490558 9024 490564 9036
rect 449860 8996 490564 9024
rect 449860 8984 449866 8996
rect 490558 8984 490564 8996
rect 490616 8984 490622 9036
rect 76650 8916 76656 8968
rect 76708 8956 76714 8968
rect 120718 8956 120724 8968
rect 76708 8928 120724 8956
rect 76708 8916 76714 8928
rect 120718 8916 120724 8928
rect 120776 8916 120782 8968
rect 137278 8916 137284 8968
rect 137336 8956 137342 8968
rect 167638 8956 167644 8968
rect 137336 8928 167644 8956
rect 137336 8916 137342 8928
rect 167638 8916 167644 8928
rect 167696 8916 167702 8968
rect 172974 8916 172980 8968
rect 173032 8956 173038 8968
rect 197446 8956 197452 8968
rect 173032 8928 197452 8956
rect 173032 8916 173038 8928
rect 197446 8916 197452 8928
rect 197504 8916 197510 8968
rect 371142 8916 371148 8968
rect 371200 8956 371206 8968
rect 390646 8956 390652 8968
rect 371200 8928 390652 8956
rect 371200 8916 371206 8928
rect 390646 8916 390652 8928
rect 390704 8916 390710 8968
rect 391290 8916 391296 8968
rect 391348 8956 391354 8968
rect 415670 8956 415676 8968
rect 391348 8928 415676 8956
rect 391348 8916 391354 8928
rect 415670 8916 415676 8928
rect 415728 8916 415734 8968
rect 416682 8916 416688 8968
rect 416740 8956 416746 8968
rect 447778 8956 447784 8968
rect 416740 8928 447784 8956
rect 416740 8916 416746 8928
rect 447778 8916 447784 8928
rect 447836 8916 447842 8968
rect 467742 8916 467748 8968
rect 467800 8956 467806 8968
rect 513190 8956 513196 8968
rect 467800 8928 513196 8956
rect 467800 8916 467806 8928
rect 513190 8916 513196 8928
rect 513248 8916 513254 8968
rect 514662 8916 514668 8968
rect 514720 8956 514726 8968
rect 572622 8956 572628 8968
rect 514720 8928 572628 8956
rect 514720 8916 514726 8928
rect 572622 8916 572628 8928
rect 572680 8916 572686 8968
rect 523678 8236 523684 8288
rect 523736 8276 523742 8288
rect 580166 8276 580172 8288
rect 523736 8248 580172 8276
rect 523736 8236 523742 8248
rect 580166 8236 580172 8248
rect 580224 8236 580230 8288
rect 133690 7624 133696 7676
rect 133748 7664 133754 7676
rect 166994 7664 167000 7676
rect 133748 7636 167000 7664
rect 133748 7624 133754 7636
rect 166994 7624 167000 7636
rect 167052 7624 167058 7676
rect 382182 7624 382188 7676
rect 382240 7664 382246 7676
rect 404906 7664 404912 7676
rect 382240 7636 404912 7664
rect 382240 7624 382246 7636
rect 404906 7624 404912 7636
rect 404964 7624 404970 7676
rect 447042 7624 447048 7676
rect 447100 7664 447106 7676
rect 486970 7664 486976 7676
rect 447100 7636 486976 7664
rect 447100 7624 447106 7636
rect 486970 7624 486976 7636
rect 487028 7624 487034 7676
rect 494054 7624 494060 7676
rect 494112 7664 494118 7676
rect 495342 7664 495348 7676
rect 494112 7636 495348 7664
rect 494112 7624 494118 7636
rect 495342 7624 495348 7636
rect 495400 7624 495406 7676
rect 1670 7556 1676 7608
rect 1728 7596 1734 7608
rect 62482 7596 62488 7608
rect 1728 7568 62488 7596
rect 1728 7556 1734 7568
rect 62482 7556 62488 7568
rect 62540 7556 62546 7608
rect 65978 7556 65984 7608
rect 66036 7596 66042 7608
rect 113266 7596 113272 7608
rect 66036 7568 113272 7596
rect 66036 7556 66042 7568
rect 113266 7556 113272 7568
rect 113324 7556 113330 7608
rect 115934 7556 115940 7608
rect 115992 7596 115998 7608
rect 153286 7596 153292 7608
rect 115992 7568 153292 7596
rect 115992 7556 115998 7568
rect 153286 7556 153292 7568
rect 153344 7556 153350 7608
rect 169386 7556 169392 7608
rect 169444 7596 169450 7608
rect 194686 7596 194692 7608
rect 169444 7568 194692 7596
rect 169444 7556 169450 7568
rect 194686 7556 194692 7568
rect 194744 7556 194750 7608
rect 362770 7556 362776 7608
rect 362828 7596 362834 7608
rect 379974 7596 379980 7608
rect 362828 7568 379980 7596
rect 362828 7556 362834 7568
rect 379974 7556 379980 7568
rect 380032 7556 380038 7608
rect 402238 7556 402244 7608
rect 402296 7596 402302 7608
rect 429930 7596 429936 7608
rect 402296 7568 429936 7596
rect 402296 7556 402302 7568
rect 429930 7556 429936 7568
rect 429988 7556 429994 7608
rect 466362 7556 466368 7608
rect 466420 7596 466426 7608
rect 511994 7596 512000 7608
rect 466420 7568 512000 7596
rect 466420 7556 466426 7568
rect 511994 7556 512000 7568
rect 512052 7556 512058 7608
rect 130194 6196 130200 6248
rect 130252 6236 130258 6248
rect 164234 6236 164240 6248
rect 130252 6208 164240 6236
rect 130252 6196 130258 6208
rect 164234 6196 164240 6208
rect 164292 6196 164298 6248
rect 446398 6196 446404 6248
rect 446456 6236 446462 6248
rect 483474 6236 483480 6248
rect 446456 6208 483480 6236
rect 446456 6196 446462 6208
rect 483474 6196 483480 6208
rect 483532 6196 483538 6248
rect 566 6128 572 6180
rect 624 6168 630 6180
rect 61378 6168 61384 6180
rect 624 6140 61384 6168
rect 624 6128 630 6140
rect 61378 6128 61384 6140
rect 61436 6128 61442 6180
rect 62390 6128 62396 6180
rect 62448 6168 62454 6180
rect 110414 6168 110420 6180
rect 62448 6140 110420 6168
rect 62448 6128 62454 6140
rect 110414 6128 110420 6140
rect 110472 6128 110478 6180
rect 112346 6128 112352 6180
rect 112404 6168 112410 6180
rect 150526 6168 150532 6180
rect 112404 6140 150532 6168
rect 112404 6128 112410 6140
rect 150526 6128 150532 6140
rect 150584 6128 150590 6180
rect 165890 6128 165896 6180
rect 165948 6168 165954 6180
rect 191926 6168 191932 6180
rect 165948 6140 191932 6168
rect 165948 6128 165954 6140
rect 191926 6128 191932 6140
rect 191984 6128 191990 6180
rect 360010 6128 360016 6180
rect 360068 6168 360074 6180
rect 376386 6168 376392 6180
rect 360068 6140 376392 6168
rect 360068 6128 360074 6140
rect 376386 6128 376392 6140
rect 376444 6128 376450 6180
rect 376662 6128 376668 6180
rect 376720 6168 376726 6180
rect 397822 6168 397828 6180
rect 376720 6140 397828 6168
rect 376720 6128 376726 6140
rect 397822 6128 397828 6140
rect 397880 6128 397886 6180
rect 398650 6128 398656 6180
rect 398708 6168 398714 6180
rect 426250 6168 426256 6180
rect 398708 6140 426256 6168
rect 398708 6128 398714 6140
rect 426250 6128 426256 6140
rect 426308 6128 426314 6180
rect 441522 6128 441528 6180
rect 441580 6168 441586 6180
rect 479886 6168 479892 6180
rect 441580 6140 479892 6168
rect 441580 6128 441586 6140
rect 479886 6128 479892 6140
rect 479944 6128 479950 6180
rect 482278 6128 482284 6180
rect 482336 6168 482342 6180
rect 497734 6168 497740 6180
rect 482336 6140 497740 6168
rect 482336 6128 482342 6140
rect 497734 6128 497740 6140
rect 497792 6128 497798 6180
rect 506382 6128 506388 6180
rect 506440 6168 506446 6180
rect 561950 6168 561956 6180
rect 506440 6140 561956 6168
rect 506440 6128 506446 6140
rect 561950 6128 561956 6140
rect 562008 6128 562014 6180
rect 471790 5312 471796 5364
rect 471848 5352 471854 5364
rect 519078 5352 519084 5364
rect 471848 5324 519084 5352
rect 471848 5312 471854 5324
rect 519078 5312 519084 5324
rect 519136 5312 519142 5364
rect 474550 5244 474556 5296
rect 474608 5284 474614 5296
rect 522666 5284 522672 5296
rect 474608 5256 522672 5284
rect 474608 5244 474614 5256
rect 522666 5244 522672 5256
rect 522724 5244 522730 5296
rect 484302 5176 484308 5228
rect 484360 5216 484366 5228
rect 533430 5216 533436 5228
rect 484360 5188 533436 5216
rect 484360 5176 484366 5188
rect 533430 5176 533436 5188
rect 533488 5176 533494 5228
rect 55214 5108 55220 5160
rect 55272 5148 55278 5160
rect 104894 5148 104900 5160
rect 55272 5120 104900 5148
rect 55272 5108 55278 5120
rect 104894 5108 104900 5120
rect 104952 5108 104958 5160
rect 477402 5108 477408 5160
rect 477460 5148 477466 5160
rect 526254 5148 526260 5160
rect 477460 5120 526260 5148
rect 477460 5108 477466 5120
rect 526254 5108 526260 5120
rect 526312 5108 526318 5160
rect 540514 5148 540520 5160
rect 533356 5120 540520 5148
rect 58802 5040 58808 5092
rect 58860 5080 58866 5092
rect 107654 5080 107660 5092
rect 58860 5052 107660 5080
rect 58860 5040 58866 5052
rect 107654 5040 107660 5052
rect 107712 5040 107718 5092
rect 480070 5040 480076 5092
rect 480128 5080 480134 5092
rect 529842 5080 529848 5092
rect 480128 5052 529848 5080
rect 480128 5040 480134 5052
rect 529842 5040 529848 5052
rect 529900 5040 529906 5092
rect 51626 4972 51632 5024
rect 51684 5012 51690 5024
rect 102134 5012 102140 5024
rect 51684 4984 102140 5012
rect 51684 4972 51690 4984
rect 102134 4972 102140 4984
rect 102192 4972 102198 5024
rect 489638 4972 489644 5024
rect 489696 5012 489702 5024
rect 499577 5015 499635 5021
rect 499577 5012 499589 5015
rect 489696 4984 499589 5012
rect 489696 4972 489702 4984
rect 499577 4981 499589 4984
rect 499623 4981 499635 5015
rect 499577 4975 499635 4981
rect 509145 5015 509203 5021
rect 509145 4981 509157 5015
rect 509191 5012 509203 5015
rect 518897 5015 518955 5021
rect 518897 5012 518909 5015
rect 509191 4984 518909 5012
rect 509191 4981 509203 4984
rect 509145 4975 509203 4981
rect 518897 4981 518909 4984
rect 518943 4981 518955 5015
rect 518897 4975 518955 4981
rect 528465 5015 528523 5021
rect 528465 4981 528477 5015
rect 528511 5012 528523 5015
rect 533356 5012 533384 5120
rect 540514 5108 540520 5120
rect 540572 5108 540578 5160
rect 528511 4984 533384 5012
rect 528511 4981 528523 4984
rect 528465 4975 528523 4981
rect 48130 4904 48136 4956
rect 48188 4944 48194 4956
rect 99374 4944 99380 4956
rect 48188 4916 99380 4944
rect 48188 4904 48194 4916
rect 99374 4904 99380 4916
rect 99432 4904 99438 4956
rect 279878 4904 279884 4956
rect 279936 4944 279942 4956
rect 280062 4944 280068 4956
rect 279936 4916 280068 4944
rect 279936 4904 279942 4916
rect 280062 4904 280068 4916
rect 280120 4904 280126 4956
rect 487062 4904 487068 4956
rect 487120 4944 487126 4956
rect 536926 4944 536932 4956
rect 487120 4916 536932 4944
rect 487120 4904 487126 4916
rect 536926 4904 536932 4916
rect 536984 4904 536990 4956
rect 17310 4836 17316 4888
rect 17368 4876 17374 4888
rect 74718 4876 74724 4888
rect 17368 4848 74724 4876
rect 17368 4836 17374 4848
rect 74718 4836 74724 4848
rect 74776 4836 74782 4888
rect 183738 4836 183744 4888
rect 183796 4876 183802 4888
rect 204898 4876 204904 4888
rect 183796 4848 204904 4876
rect 183796 4836 183802 4848
rect 204898 4836 204904 4848
rect 204956 4836 204962 4888
rect 373258 4836 373264 4888
rect 373316 4876 373322 4888
rect 383378 4876 383384 4888
rect 373316 4848 383384 4876
rect 373316 4836 373322 4848
rect 383378 4836 383384 4848
rect 383436 4836 383442 4888
rect 393958 4836 393964 4888
rect 394016 4876 394022 4888
rect 419166 4876 419172 4888
rect 394016 4848 419172 4876
rect 394016 4836 394022 4848
rect 419166 4836 419172 4848
rect 419224 4836 419230 4888
rect 457438 4836 457444 4888
rect 457496 4876 457502 4888
rect 457496 4848 462268 4876
rect 457496 4836 457502 4848
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 71774 4808 71780 4820
rect 12492 4780 71780 4808
rect 12492 4768 12498 4780
rect 71774 4768 71780 4780
rect 71832 4768 71838 4820
rect 73062 4768 73068 4820
rect 73120 4808 73126 4820
rect 118786 4808 118792 4820
rect 73120 4780 118792 4808
rect 73120 4768 73126 4780
rect 118786 4768 118792 4780
rect 118844 4768 118850 4820
rect 126606 4768 126612 4820
rect 126664 4808 126670 4820
rect 161474 4808 161480 4820
rect 126664 4780 161480 4808
rect 126664 4768 126670 4780
rect 161474 4768 161480 4780
rect 161532 4768 161538 4820
rect 162302 4768 162308 4820
rect 162360 4808 162366 4820
rect 189166 4808 189172 4820
rect 162360 4780 189172 4808
rect 162360 4768 162366 4780
rect 189166 4768 189172 4780
rect 189224 4768 189230 4820
rect 357250 4768 357256 4820
rect 357308 4808 357314 4820
rect 372798 4808 372804 4820
rect 357308 4780 372804 4808
rect 357308 4768 357314 4780
rect 372798 4768 372804 4780
rect 372856 4768 372862 4820
rect 381538 4768 381544 4820
rect 381596 4808 381602 4820
rect 401318 4808 401324 4820
rect 381596 4780 401324 4808
rect 381596 4768 381602 4780
rect 401318 4768 401324 4780
rect 401376 4768 401382 4820
rect 407022 4768 407028 4820
rect 407080 4808 407086 4820
rect 437014 4808 437020 4820
rect 407080 4780 437020 4808
rect 407080 4768 407086 4780
rect 437014 4768 437020 4780
rect 437072 4768 437078 4820
rect 438302 4768 438308 4820
rect 438360 4808 438366 4820
rect 462038 4808 462044 4820
rect 438360 4780 462044 4808
rect 438360 4768 438366 4780
rect 462038 4768 462044 4780
rect 462096 4768 462102 4820
rect 462240 4808 462268 4848
rect 492582 4836 492588 4888
rect 492640 4876 492646 4888
rect 544102 4876 544108 4888
rect 492640 4848 544108 4876
rect 492640 4836 492646 4848
rect 544102 4836 544108 4848
rect 544160 4836 544166 4888
rect 472710 4808 472716 4820
rect 462240 4780 472716 4808
rect 472710 4768 472716 4780
rect 472768 4768 472774 4820
rect 495158 4768 495164 4820
rect 495216 4808 495222 4820
rect 547690 4808 547696 4820
rect 495216 4780 547696 4808
rect 495216 4768 495222 4780
rect 547690 4768 547696 4780
rect 547748 4768 547754 4820
rect 499577 4743 499635 4749
rect 499577 4709 499589 4743
rect 499623 4740 499635 4743
rect 509145 4743 509203 4749
rect 509145 4740 509157 4743
rect 499623 4712 509157 4740
rect 499623 4709 499635 4712
rect 499577 4703 499635 4709
rect 509145 4709 509157 4712
rect 509191 4709 509203 4743
rect 509145 4703 509203 4709
rect 518897 4743 518955 4749
rect 518897 4709 518909 4743
rect 518943 4740 518955 4743
rect 528465 4743 528523 4749
rect 528465 4740 528477 4743
rect 518943 4712 528477 4740
rect 518943 4709 518955 4712
rect 518897 4703 518955 4709
rect 528465 4709 528477 4712
rect 528511 4709 528523 4743
rect 528465 4703 528523 4709
rect 391198 4632 391204 4684
rect 391256 4672 391262 4684
rect 394234 4672 394240 4684
rect 391256 4644 394240 4672
rect 391256 4632 391262 4644
rect 394234 4632 394240 4644
rect 394292 4632 394298 4684
rect 296714 4360 296720 4412
rect 296772 4400 296778 4412
rect 297082 4400 297088 4412
rect 296772 4372 297088 4400
rect 296772 4360 296778 4372
rect 297082 4360 297088 4372
rect 297140 4360 297146 4412
rect 45738 4088 45744 4140
rect 45796 4128 45802 4140
rect 97994 4128 98000 4140
rect 45796 4100 98000 4128
rect 45796 4088 45802 4100
rect 97994 4088 98000 4100
rect 98052 4088 98058 4140
rect 106366 4088 106372 4140
rect 106424 4128 106430 4140
rect 144914 4128 144920 4140
rect 106424 4100 144920 4128
rect 106424 4088 106430 4100
rect 144914 4088 144920 4100
rect 144972 4088 144978 4140
rect 155126 4088 155132 4140
rect 155184 4128 155190 4140
rect 155862 4128 155868 4140
rect 155184 4100 155868 4128
rect 155184 4088 155190 4100
rect 155862 4088 155868 4100
rect 155920 4088 155926 4140
rect 158714 4088 158720 4140
rect 158772 4128 158778 4140
rect 159910 4128 159916 4140
rect 158772 4100 159916 4128
rect 158772 4088 158778 4100
rect 159910 4088 159916 4100
rect 159968 4088 159974 4140
rect 163498 4088 163504 4140
rect 163556 4128 163562 4140
rect 164142 4128 164148 4140
rect 163556 4100 164148 4128
rect 163556 4088 163562 4100
rect 164142 4088 164148 4100
rect 164200 4088 164206 4140
rect 170582 4088 170588 4140
rect 170640 4128 170646 4140
rect 195974 4128 195980 4140
rect 170640 4100 195980 4128
rect 170640 4088 170646 4100
rect 195974 4088 195980 4100
rect 196032 4088 196038 4140
rect 200761 4131 200819 4137
rect 200761 4097 200773 4131
rect 200807 4128 200819 4131
rect 207106 4128 207112 4140
rect 200807 4100 207112 4128
rect 200807 4097 200819 4100
rect 200761 4091 200819 4097
rect 207106 4088 207112 4100
rect 207164 4088 207170 4140
rect 207201 4131 207259 4137
rect 207201 4097 207213 4131
rect 207247 4128 207259 4131
rect 209777 4131 209835 4137
rect 209777 4128 209789 4131
rect 207247 4100 209789 4128
rect 207247 4097 207259 4100
rect 207201 4091 207259 4097
rect 209777 4097 209789 4100
rect 209823 4097 209835 4131
rect 209777 4091 209835 4097
rect 278866 4088 278872 4140
rect 278924 4128 278930 4140
rect 279878 4128 279884 4140
rect 278924 4100 279884 4128
rect 278924 4088 278930 4100
rect 279878 4088 279884 4100
rect 279936 4088 279942 4140
rect 287146 4088 287152 4140
rect 287204 4128 287210 4140
rect 288342 4128 288348 4140
rect 287204 4100 288348 4128
rect 287204 4088 287210 4100
rect 288342 4088 288348 4100
rect 288400 4088 288406 4140
rect 289538 4088 289544 4140
rect 289596 4128 289602 4140
rect 289906 4128 289912 4140
rect 289596 4100 289912 4128
rect 289596 4088 289602 4100
rect 289906 4088 289912 4100
rect 289964 4088 289970 4140
rect 291470 4088 291476 4140
rect 291528 4128 291534 4140
rect 291930 4128 291936 4140
rect 291528 4100 291936 4128
rect 291528 4088 291534 4100
rect 291930 4088 291936 4100
rect 291988 4088 291994 4140
rect 292574 4088 292580 4140
rect 292632 4128 292638 4140
rect 293126 4128 293132 4140
rect 292632 4100 293132 4128
rect 292632 4088 292638 4100
rect 293126 4088 293132 4100
rect 293184 4088 293190 4140
rect 296806 4088 296812 4140
rect 296864 4128 296870 4140
rect 297910 4128 297916 4140
rect 296864 4100 297916 4128
rect 296864 4088 296870 4100
rect 297910 4088 297916 4100
rect 297968 4088 297974 4140
rect 298094 4088 298100 4140
rect 298152 4128 298158 4140
rect 299106 4128 299112 4140
rect 298152 4100 299112 4128
rect 298152 4088 298158 4100
rect 299106 4088 299112 4100
rect 299164 4088 299170 4140
rect 299382 4088 299388 4140
rect 299440 4128 299446 4140
rect 300302 4128 300308 4140
rect 299440 4100 300308 4128
rect 299440 4088 299446 4100
rect 300302 4088 300308 4100
rect 300360 4088 300366 4140
rect 306282 4088 306288 4140
rect 306340 4128 306346 4140
rect 308582 4128 308588 4140
rect 306340 4100 308588 4128
rect 306340 4088 306346 4100
rect 308582 4088 308588 4100
rect 308640 4088 308646 4140
rect 338022 4088 338028 4140
rect 338080 4128 338086 4140
rect 348878 4128 348884 4140
rect 338080 4100 348884 4128
rect 338080 4088 338086 4100
rect 348878 4088 348884 4100
rect 348936 4088 348942 4140
rect 350442 4088 350448 4140
rect 350500 4128 350506 4140
rect 364518 4128 364524 4140
rect 350500 4100 364524 4128
rect 350500 4088 350506 4100
rect 364518 4088 364524 4100
rect 364576 4088 364582 4140
rect 367002 4088 367008 4140
rect 367060 4128 367066 4140
rect 385862 4128 385868 4140
rect 367060 4100 385868 4128
rect 367060 4088 367066 4100
rect 385862 4088 385868 4100
rect 385920 4088 385926 4140
rect 386230 4088 386236 4140
rect 386288 4128 386294 4140
rect 409690 4128 409696 4140
rect 386288 4100 409696 4128
rect 386288 4088 386294 4100
rect 409690 4088 409696 4100
rect 409748 4088 409754 4140
rect 442810 4088 442816 4140
rect 442868 4128 442874 4140
rect 481082 4128 481088 4140
rect 442868 4100 481088 4128
rect 442868 4088 442874 4100
rect 481082 4088 481088 4100
rect 481140 4088 481146 4140
rect 496722 4088 496728 4140
rect 496780 4128 496786 4140
rect 550082 4128 550088 4140
rect 496780 4100 550088 4128
rect 496780 4088 496786 4100
rect 550082 4088 550088 4100
rect 550140 4088 550146 4140
rect 43346 4020 43352 4072
rect 43404 4060 43410 4072
rect 43404 4032 92612 4060
rect 43404 4020 43410 4032
rect 36170 3952 36176 4004
rect 36228 3992 36234 4004
rect 89714 3992 89720 4004
rect 36228 3964 89720 3992
rect 36228 3952 36234 3964
rect 89714 3952 89720 3964
rect 89772 3952 89778 4004
rect 39758 3884 39764 3936
rect 39816 3924 39822 3936
rect 92474 3924 92480 3936
rect 39816 3896 92480 3924
rect 39816 3884 39822 3896
rect 92474 3884 92480 3896
rect 92532 3884 92538 3936
rect 32674 3816 32680 3868
rect 32732 3856 32738 3868
rect 32732 3828 84332 3856
rect 32732 3816 32738 3828
rect 5258 3748 5264 3800
rect 5316 3788 5322 3800
rect 8938 3788 8944 3800
rect 5316 3760 8944 3788
rect 5316 3748 5322 3760
rect 8938 3748 8944 3760
rect 8996 3748 9002 3800
rect 29086 3748 29092 3800
rect 29144 3788 29150 3800
rect 84194 3788 84200 3800
rect 29144 3760 84200 3788
rect 29144 3748 29150 3760
rect 84194 3748 84200 3760
rect 84252 3748 84258 3800
rect 84304 3788 84332 3828
rect 84930 3816 84936 3868
rect 84988 3856 84994 3868
rect 85482 3856 85488 3868
rect 84988 3828 85488 3856
rect 84988 3816 84994 3828
rect 85482 3816 85488 3828
rect 85540 3816 85546 3868
rect 88518 3816 88524 3868
rect 88576 3856 88582 3868
rect 89622 3856 89628 3868
rect 88576 3828 89628 3856
rect 88576 3816 88582 3828
rect 89622 3816 89628 3828
rect 89680 3816 89686 3868
rect 92584 3856 92612 4032
rect 109954 4020 109960 4072
rect 110012 4060 110018 4072
rect 147766 4060 147772 4072
rect 110012 4032 147772 4060
rect 110012 4020 110018 4032
rect 147766 4020 147772 4032
rect 147824 4020 147830 4072
rect 167086 4020 167092 4072
rect 167144 4060 167150 4072
rect 193214 4060 193220 4072
rect 167144 4032 193220 4060
rect 167144 4020 167150 4032
rect 193214 4020 193220 4032
rect 193272 4020 193278 4072
rect 196802 4020 196808 4072
rect 196860 4060 196866 4072
rect 216674 4060 216680 4072
rect 196860 4032 216680 4060
rect 196860 4020 196866 4032
rect 216674 4020 216680 4032
rect 216732 4020 216738 4072
rect 218238 4020 218244 4072
rect 218296 4060 218302 4072
rect 219342 4060 219348 4072
rect 218296 4032 219348 4060
rect 218296 4020 218302 4032
rect 219342 4020 219348 4032
rect 219400 4020 219406 4072
rect 304810 4020 304816 4072
rect 304868 4060 304874 4072
rect 307386 4060 307392 4072
rect 304868 4032 307392 4060
rect 304868 4020 304874 4032
rect 307386 4020 307392 4032
rect 307444 4020 307450 4072
rect 331122 4020 331128 4072
rect 331180 4060 331186 4072
rect 339494 4060 339500 4072
rect 331180 4032 339500 4060
rect 331180 4020 331186 4032
rect 339494 4020 339500 4032
rect 339552 4020 339558 4072
rect 342162 4020 342168 4072
rect 342220 4060 342226 4072
rect 353754 4060 353760 4072
rect 342220 4032 353760 4060
rect 342220 4020 342226 4032
rect 353754 4020 353760 4032
rect 353812 4020 353818 4072
rect 354582 4020 354588 4072
rect 354640 4060 354646 4072
rect 370406 4060 370412 4072
rect 354640 4032 370412 4060
rect 354640 4020 354646 4032
rect 370406 4020 370412 4032
rect 370464 4020 370470 4072
rect 372522 4020 372528 4072
rect 372580 4060 372586 4072
rect 393038 4060 393044 4072
rect 372580 4032 393044 4060
rect 372580 4020 372586 4032
rect 393038 4020 393044 4032
rect 393096 4020 393102 4072
rect 393222 4020 393228 4072
rect 393280 4060 393286 4072
rect 417970 4060 417976 4072
rect 393280 4032 417976 4060
rect 393280 4020 393286 4032
rect 417970 4020 417976 4032
rect 418028 4020 418034 4072
rect 440050 4020 440056 4072
rect 440108 4060 440114 4072
rect 478690 4060 478696 4072
rect 440108 4032 478696 4060
rect 440108 4020 440114 4032
rect 478690 4020 478696 4032
rect 478748 4020 478754 4072
rect 502242 4020 502248 4072
rect 502300 4060 502306 4072
rect 557166 4060 557172 4072
rect 502300 4032 557172 4060
rect 502300 4020 502306 4032
rect 557166 4020 557172 4032
rect 557224 4020 557230 4072
rect 111150 3952 111156 4004
rect 111208 3992 111214 4004
rect 149054 3992 149060 4004
rect 111208 3964 149060 3992
rect 111208 3952 111214 3964
rect 149054 3952 149060 3964
rect 149112 3952 149118 4004
rect 156322 3952 156328 4004
rect 156380 3992 156386 4004
rect 184934 3992 184940 4004
rect 156380 3964 184940 3992
rect 156380 3952 156386 3964
rect 184934 3952 184940 3964
rect 184992 3952 184998 4004
rect 195606 3952 195612 4004
rect 195664 3992 195670 4004
rect 215294 3992 215300 4004
rect 195664 3964 215300 3992
rect 195664 3952 195670 3964
rect 215294 3952 215300 3964
rect 215352 3952 215358 4004
rect 215389 3995 215447 4001
rect 215389 3961 215401 3995
rect 215435 3992 215447 3995
rect 221001 3995 221059 4001
rect 215435 3964 218284 3992
rect 215435 3961 215447 3964
rect 215389 3955 215447 3961
rect 103974 3884 103980 3936
rect 104032 3924 104038 3936
rect 104032 3896 140912 3924
rect 104032 3884 104038 3896
rect 95234 3856 95240 3868
rect 92584 3828 95240 3856
rect 95234 3816 95240 3828
rect 95292 3816 95298 3868
rect 99190 3816 99196 3868
rect 99248 3856 99254 3868
rect 139394 3856 139400 3868
rect 99248 3828 139400 3856
rect 99248 3816 99254 3828
rect 139394 3816 139400 3828
rect 139452 3816 139458 3868
rect 86954 3788 86960 3800
rect 84304 3760 86960 3788
rect 86954 3748 86960 3760
rect 87012 3748 87018 3800
rect 96890 3748 96896 3800
rect 96948 3788 96954 3800
rect 138014 3788 138020 3800
rect 96948 3760 138020 3788
rect 96948 3748 96954 3760
rect 138014 3748 138020 3760
rect 138072 3748 138078 3800
rect 24302 3680 24308 3732
rect 24360 3720 24366 3732
rect 80146 3720 80152 3732
rect 24360 3692 80152 3720
rect 24360 3680 24366 3692
rect 80146 3680 80152 3692
rect 80204 3680 80210 3732
rect 95605 3723 95663 3729
rect 95605 3689 95617 3723
rect 95651 3720 95663 3723
rect 98270 3720 98276 3732
rect 95651 3692 98276 3720
rect 95651 3689 95663 3692
rect 95605 3683 95663 3689
rect 98270 3680 98276 3692
rect 98328 3680 98334 3732
rect 100478 3680 100484 3732
rect 100536 3720 100542 3732
rect 140774 3720 140780 3732
rect 100536 3692 140780 3720
rect 100536 3680 100542 3692
rect 140774 3680 140780 3692
rect 140832 3680 140838 3732
rect 10318 3652 10324 3664
rect 7576 3624 10324 3652
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4062 3516 4068 3528
rect 2924 3488 4068 3516
rect 2924 3476 2930 3488
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 7576 3516 7604 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 20772 3624 70624 3652
rect 20772 3612 20778 3624
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11296 3556 14596 3584
rect 11296 3544 11302 3556
rect 4172 3488 7604 3516
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 4172 3380 4200 3488
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 9030 3516 9036 3528
rect 7708 3488 9036 3516
rect 7708 3476 7714 3488
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 14458 3516 14464 3528
rect 13688 3488 14464 3516
rect 13688 3476 13694 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14568 3516 14596 3556
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 63497 3587 63555 3593
rect 63497 3584 63509 3587
rect 14884 3556 63509 3584
rect 14884 3544 14890 3556
rect 63497 3553 63509 3556
rect 63543 3553 63555 3587
rect 63497 3547 63555 3553
rect 63586 3544 63592 3596
rect 63644 3584 63650 3596
rect 64690 3584 64696 3596
rect 63644 3556 64696 3584
rect 63644 3544 63650 3556
rect 64690 3544 64696 3556
rect 64748 3544 64754 3596
rect 70486 3584 70492 3596
rect 65536 3556 70492 3584
rect 65536 3516 65564 3556
rect 70486 3544 70492 3556
rect 70544 3544 70550 3596
rect 70596 3584 70624 3624
rect 70670 3612 70676 3664
rect 70728 3652 70734 3664
rect 71682 3652 71688 3664
rect 70728 3624 71688 3652
rect 70728 3612 70734 3624
rect 71682 3612 71688 3624
rect 71740 3612 71746 3664
rect 77386 3652 77392 3664
rect 71792 3624 77392 3652
rect 71792 3584 71820 3624
rect 77386 3612 77392 3624
rect 77444 3612 77450 3664
rect 77846 3612 77852 3664
rect 77904 3652 77910 3664
rect 78582 3652 78588 3664
rect 77904 3624 78588 3652
rect 77904 3612 77910 3624
rect 78582 3612 78588 3624
rect 78640 3612 78646 3664
rect 93302 3612 93308 3664
rect 93360 3652 93366 3664
rect 135254 3652 135260 3664
rect 93360 3624 135260 3652
rect 93360 3612 93366 3624
rect 135254 3612 135260 3624
rect 135312 3612 135318 3664
rect 140884 3652 140912 3896
rect 150434 3884 150440 3936
rect 150492 3924 150498 3936
rect 179414 3924 179420 3936
rect 150492 3896 179420 3924
rect 150492 3884 150498 3896
rect 179414 3884 179420 3896
rect 179472 3884 179478 3936
rect 192018 3884 192024 3936
rect 192076 3924 192082 3936
rect 212534 3924 212540 3936
rect 192076 3896 212540 3924
rect 192076 3884 192082 3896
rect 212534 3884 212540 3896
rect 212592 3884 212598 3936
rect 213917 3927 213975 3933
rect 213917 3893 213929 3927
rect 213963 3924 213975 3927
rect 218146 3924 218152 3936
rect 213963 3896 218152 3924
rect 213963 3893 213975 3896
rect 213917 3887 213975 3893
rect 218146 3884 218152 3896
rect 218204 3884 218210 3936
rect 218256 3924 218284 3964
rect 221001 3961 221013 3995
rect 221047 3992 221059 3995
rect 227714 3992 227720 4004
rect 221047 3964 227720 3992
rect 221047 3961 221059 3964
rect 221001 3955 221059 3961
rect 227714 3952 227720 3964
rect 227772 3952 227778 4004
rect 229097 3995 229155 4001
rect 229097 3961 229109 3995
rect 229143 3992 229155 3995
rect 240134 3992 240140 4004
rect 229143 3964 240140 3992
rect 229143 3961 229155 3964
rect 229097 3955 229155 3961
rect 240134 3952 240140 3964
rect 240192 3952 240198 4004
rect 284754 3952 284760 4004
rect 284812 3992 284818 4004
rect 285766 3992 285772 4004
rect 284812 3964 285772 3992
rect 284812 3952 284818 3964
rect 285766 3952 285772 3964
rect 285824 3952 285830 4004
rect 320082 3952 320088 4004
rect 320140 3992 320146 4004
rect 326430 3992 326436 4004
rect 320140 3964 326436 3992
rect 320140 3952 320146 3964
rect 326430 3952 326436 3964
rect 326488 3952 326494 4004
rect 332502 3952 332508 4004
rect 332560 3992 332566 4004
rect 341886 3992 341892 4004
rect 332560 3964 341892 3992
rect 332560 3952 332566 3964
rect 341886 3952 341892 3964
rect 341944 3952 341950 4004
rect 346302 3952 346308 4004
rect 346360 3992 346366 4004
rect 359734 3992 359740 4004
rect 346360 3964 359740 3992
rect 346360 3952 346366 3964
rect 359734 3952 359740 3964
rect 359792 3952 359798 4004
rect 361482 3952 361488 4004
rect 361540 3992 361546 4004
rect 378778 3992 378784 4004
rect 361540 3964 378784 3992
rect 361540 3952 361546 3964
rect 378778 3952 378784 3964
rect 378836 3952 378842 4004
rect 383470 3952 383476 4004
rect 383528 3992 383534 4004
rect 406102 3992 406108 4004
rect 383528 3964 406108 3992
rect 383528 3952 383534 3964
rect 406102 3952 406108 3964
rect 406160 3952 406166 4004
rect 409782 3952 409788 4004
rect 409840 3992 409846 4004
rect 439406 3992 439412 4004
rect 409840 3964 439412 3992
rect 409840 3952 409846 3964
rect 439406 3952 439412 3964
rect 439464 3952 439470 4004
rect 448330 3952 448336 4004
rect 448388 3992 448394 4004
rect 489362 3992 489368 4004
rect 448388 3964 489368 3992
rect 448388 3952 448394 3964
rect 489362 3952 489368 3964
rect 489420 3952 489426 4004
rect 505002 3952 505008 4004
rect 505060 3992 505066 4004
rect 560754 3992 560760 4004
rect 505060 3964 560760 3992
rect 505060 3952 505066 3964
rect 560754 3952 560760 3964
rect 560812 3952 560818 4004
rect 220906 3924 220912 3936
rect 218256 3896 220912 3924
rect 220906 3884 220912 3896
rect 220964 3884 220970 3936
rect 224126 3884 224132 3936
rect 224184 3924 224190 3936
rect 238846 3924 238852 3936
rect 224184 3896 238852 3924
rect 224184 3884 224190 3896
rect 238846 3884 238852 3896
rect 238904 3884 238910 3936
rect 335262 3884 335268 3936
rect 335320 3924 335326 3936
rect 345474 3924 345480 3936
rect 335320 3896 345480 3924
rect 335320 3884 335326 3896
rect 345474 3884 345480 3896
rect 345532 3884 345538 3936
rect 347682 3884 347688 3936
rect 347740 3924 347746 3936
rect 360930 3924 360936 3936
rect 347740 3896 360936 3924
rect 347740 3884 347746 3896
rect 360930 3884 360936 3896
rect 360988 3884 360994 3936
rect 364242 3884 364248 3936
rect 364300 3924 364306 3936
rect 382366 3924 382372 3936
rect 364300 3896 382372 3924
rect 364300 3884 364306 3896
rect 382366 3884 382372 3896
rect 382424 3884 382430 3936
rect 386322 3884 386328 3936
rect 386380 3924 386386 3936
rect 410886 3924 410892 3936
rect 386380 3896 410892 3924
rect 386380 3884 386386 3896
rect 410886 3884 410892 3896
rect 410944 3884 410950 3936
rect 412542 3884 412548 3936
rect 412600 3924 412606 3936
rect 442994 3924 443000 3936
rect 412600 3896 443000 3924
rect 412600 3884 412606 3896
rect 442994 3884 443000 3896
rect 443052 3884 443058 3936
rect 445662 3884 445668 3936
rect 445720 3924 445726 3936
rect 485774 3924 485780 3936
rect 445720 3896 485780 3924
rect 445720 3884 445726 3896
rect 485774 3884 485780 3896
rect 485832 3884 485838 3936
rect 491202 3884 491208 3936
rect 491260 3924 491266 3936
rect 495437 3927 495495 3933
rect 495437 3924 495449 3927
rect 491260 3896 495449 3924
rect 491260 3884 491266 3896
rect 495437 3893 495449 3896
rect 495483 3893 495495 3927
rect 495437 3887 495495 3893
rect 507762 3884 507768 3936
rect 507820 3924 507826 3936
rect 564342 3924 564348 3936
rect 507820 3896 564348 3924
rect 507820 3884 507826 3896
rect 564342 3884 564348 3896
rect 564400 3884 564406 3936
rect 153930 3816 153936 3868
rect 153988 3856 153994 3868
rect 183554 3856 183560 3868
rect 153988 3828 183560 3856
rect 153988 3816 153994 3828
rect 183554 3816 183560 3828
rect 183612 3816 183618 3868
rect 188430 3816 188436 3868
rect 188488 3856 188494 3868
rect 209958 3856 209964 3868
rect 188488 3828 209964 3856
rect 188488 3816 188494 3828
rect 209958 3816 209964 3828
rect 210016 3816 210022 3868
rect 215389 3859 215447 3865
rect 215389 3856 215401 3859
rect 210068 3828 215401 3856
rect 147861 3791 147919 3797
rect 147861 3757 147873 3791
rect 147907 3788 147919 3791
rect 154666 3788 154672 3800
rect 147907 3760 154672 3788
rect 147907 3757 147919 3760
rect 147861 3751 147919 3757
rect 154666 3748 154672 3760
rect 154724 3748 154730 3800
rect 162121 3791 162179 3797
rect 162121 3757 162133 3791
rect 162167 3788 162179 3791
rect 182174 3788 182180 3800
rect 162167 3760 182180 3788
rect 162167 3757 162179 3760
rect 162121 3751 162179 3757
rect 182174 3748 182180 3760
rect 182232 3748 182238 3800
rect 182542 3748 182548 3800
rect 182600 3788 182606 3800
rect 205634 3788 205640 3800
rect 182600 3760 205640 3788
rect 182600 3748 182606 3760
rect 205634 3748 205640 3760
rect 205692 3748 205698 3800
rect 209777 3791 209835 3797
rect 209777 3757 209789 3791
rect 209823 3788 209835 3791
rect 210068 3788 210096 3828
rect 215389 3825 215401 3828
rect 215435 3825 215447 3859
rect 215389 3819 215447 3825
rect 215846 3816 215852 3868
rect 215904 3856 215910 3868
rect 231854 3856 231860 3868
rect 215904 3828 231860 3856
rect 215904 3816 215910 3828
rect 231854 3816 231860 3828
rect 231912 3816 231918 3868
rect 328362 3816 328368 3868
rect 328420 3856 328426 3868
rect 335906 3856 335912 3868
rect 328420 3828 335912 3856
rect 328420 3816 328426 3828
rect 335906 3816 335912 3828
rect 335964 3816 335970 3868
rect 336642 3816 336648 3868
rect 336700 3856 336706 3868
rect 346670 3856 346676 3868
rect 336700 3828 346676 3856
rect 336700 3816 336706 3828
rect 346670 3816 346676 3828
rect 346728 3816 346734 3868
rect 349062 3816 349068 3868
rect 349120 3856 349126 3868
rect 363322 3856 363328 3868
rect 349120 3828 363328 3856
rect 349120 3816 349126 3828
rect 363322 3816 363328 3828
rect 363380 3816 363386 3868
rect 365622 3816 365628 3868
rect 365680 3856 365686 3868
rect 384666 3856 384672 3868
rect 365680 3828 384672 3856
rect 365680 3816 365686 3828
rect 384666 3816 384672 3828
rect 384724 3816 384730 3868
rect 389082 3816 389088 3868
rect 389140 3856 389146 3868
rect 413278 3856 413284 3868
rect 389140 3828 413284 3856
rect 389140 3816 389146 3828
rect 413278 3816 413284 3828
rect 413336 3816 413342 3868
rect 415302 3816 415308 3868
rect 415360 3856 415366 3868
rect 446582 3856 446588 3868
rect 415360 3828 446588 3856
rect 415360 3816 415366 3828
rect 446582 3816 446588 3828
rect 446640 3816 446646 3868
rect 451182 3816 451188 3868
rect 451240 3856 451246 3868
rect 492950 3856 492956 3868
rect 451240 3828 492956 3856
rect 451240 3816 451246 3828
rect 492950 3816 492956 3828
rect 493008 3816 493014 3868
rect 510522 3816 510528 3868
rect 510580 3856 510586 3868
rect 567838 3856 567844 3868
rect 510580 3828 567844 3856
rect 510580 3816 510586 3828
rect 567838 3816 567844 3828
rect 567896 3816 567902 3868
rect 209823 3760 210096 3788
rect 209823 3757 209835 3760
rect 209777 3751 209835 3757
rect 211062 3748 211068 3800
rect 211120 3788 211126 3800
rect 221001 3791 221059 3797
rect 221001 3788 221013 3791
rect 211120 3760 221013 3788
rect 211120 3748 211126 3760
rect 221001 3757 221013 3760
rect 221047 3757 221059 3791
rect 226426 3788 226432 3800
rect 221001 3751 221059 3757
rect 221108 3760 226432 3788
rect 146846 3680 146852 3732
rect 146904 3720 146910 3732
rect 176654 3720 176660 3732
rect 146904 3692 176660 3720
rect 146904 3680 146910 3692
rect 176654 3680 176660 3692
rect 176712 3680 176718 3732
rect 184842 3680 184848 3732
rect 184900 3720 184906 3732
rect 200761 3723 200819 3729
rect 200761 3720 200773 3723
rect 184900 3692 200773 3720
rect 184900 3680 184906 3692
rect 200761 3689 200773 3692
rect 200807 3689 200819 3723
rect 200761 3683 200819 3689
rect 203886 3680 203892 3732
rect 203944 3720 203950 3732
rect 203944 3692 208440 3720
rect 203944 3680 203950 3692
rect 143534 3652 143540 3664
rect 140884 3624 143540 3652
rect 143534 3612 143540 3624
rect 143592 3612 143598 3664
rect 143644 3624 149192 3652
rect 70596 3556 71820 3584
rect 75454 3544 75460 3596
rect 75512 3584 75518 3596
rect 75512 3556 89668 3584
rect 75512 3544 75518 3556
rect 14568 3488 65564 3516
rect 69474 3476 69480 3528
rect 69532 3516 69538 3528
rect 70302 3516 70308 3528
rect 69532 3488 70308 3516
rect 69532 3476 69538 3488
rect 70302 3476 70308 3488
rect 70360 3476 70366 3528
rect 89640 3516 89668 3556
rect 89714 3544 89720 3596
rect 89772 3584 89778 3596
rect 121733 3587 121791 3593
rect 121733 3584 121745 3587
rect 89772 3556 121745 3584
rect 89772 3544 89778 3556
rect 121733 3553 121745 3556
rect 121779 3553 121791 3587
rect 121733 3547 121791 3553
rect 121822 3544 121828 3596
rect 121880 3584 121886 3596
rect 122742 3584 122748 3596
rect 121880 3556 122748 3584
rect 121880 3544 121886 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 123018 3544 123024 3596
rect 123076 3584 123082 3596
rect 124122 3584 124128 3596
rect 123076 3556 124128 3584
rect 123076 3544 123082 3556
rect 124122 3544 124128 3556
rect 124180 3544 124186 3596
rect 124214 3544 124220 3596
rect 124272 3584 124278 3596
rect 125502 3584 125508 3596
rect 124272 3556 125508 3584
rect 124272 3544 124278 3556
rect 125502 3544 125508 3556
rect 125560 3544 125566 3596
rect 125612 3556 129780 3584
rect 113821 3519 113879 3525
rect 113821 3516 113833 3519
rect 89640 3488 113833 3516
rect 113821 3485 113833 3488
rect 113867 3485 113879 3519
rect 113821 3479 113879 3485
rect 125410 3476 125416 3528
rect 125468 3516 125474 3528
rect 125612 3516 125640 3556
rect 125468 3488 125640 3516
rect 125468 3476 125474 3488
rect 127802 3476 127808 3528
rect 127860 3516 127866 3528
rect 128262 3516 128268 3528
rect 127860 3488 128268 3516
rect 127860 3476 127866 3488
rect 128262 3476 128268 3488
rect 128320 3476 128326 3528
rect 128998 3476 129004 3528
rect 129056 3516 129062 3528
rect 129642 3516 129648 3528
rect 129056 3488 129648 3516
rect 129056 3476 129062 3488
rect 129642 3476 129648 3488
rect 129700 3476 129706 3528
rect 129752 3516 129780 3556
rect 131390 3544 131396 3596
rect 131448 3584 131454 3596
rect 132402 3584 132408 3596
rect 131448 3556 132408 3584
rect 131448 3544 131454 3556
rect 132402 3544 132408 3556
rect 132460 3544 132466 3596
rect 132586 3544 132592 3596
rect 132644 3584 132650 3596
rect 133782 3584 133788 3596
rect 132644 3556 133788 3584
rect 132644 3544 132650 3556
rect 133782 3544 133788 3556
rect 133840 3544 133846 3596
rect 136082 3544 136088 3596
rect 136140 3584 136146 3596
rect 136542 3584 136548 3596
rect 136140 3556 136548 3584
rect 136140 3544 136146 3556
rect 136542 3544 136548 3556
rect 136600 3544 136606 3596
rect 139670 3544 139676 3596
rect 139728 3584 139734 3596
rect 140682 3584 140688 3596
rect 139728 3556 140688 3584
rect 139728 3544 139734 3556
rect 140682 3544 140688 3556
rect 140740 3544 140746 3596
rect 140866 3544 140872 3596
rect 140924 3584 140930 3596
rect 141970 3584 141976 3596
rect 140924 3556 141976 3584
rect 140924 3544 140930 3556
rect 141970 3544 141976 3556
rect 142028 3544 142034 3596
rect 143258 3544 143264 3596
rect 143316 3584 143322 3596
rect 143644 3584 143672 3624
rect 143316 3556 143672 3584
rect 143316 3544 143322 3556
rect 145650 3544 145656 3596
rect 145708 3584 145714 3596
rect 146202 3584 146208 3596
rect 145708 3556 146208 3584
rect 145708 3544 145714 3556
rect 146202 3544 146208 3556
rect 146260 3544 146266 3596
rect 129752 3488 147996 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 59909 3451 59967 3457
rect 59909 3448 59921 3451
rect 6512 3420 59921 3448
rect 6512 3408 6518 3420
rect 59909 3417 59921 3420
rect 59955 3417 59967 3451
rect 59909 3411 59967 3417
rect 59998 3408 60004 3460
rect 60056 3448 60062 3460
rect 60642 3448 60648 3460
rect 60056 3420 60648 3448
rect 60056 3408 60062 3420
rect 60642 3408 60648 3420
rect 60700 3408 60706 3460
rect 68278 3408 68284 3460
rect 68336 3448 68342 3460
rect 116118 3448 116124 3460
rect 68336 3420 116124 3448
rect 68336 3408 68342 3420
rect 116118 3408 116124 3420
rect 116176 3408 116182 3460
rect 118234 3408 118240 3460
rect 118292 3448 118298 3460
rect 147861 3451 147919 3457
rect 147861 3448 147873 3451
rect 118292 3420 147873 3448
rect 118292 3408 118298 3420
rect 147861 3417 147873 3420
rect 147907 3417 147919 3451
rect 147968 3448 147996 3488
rect 148042 3476 148048 3528
rect 148100 3516 148106 3528
rect 148962 3516 148968 3528
rect 148100 3488 148968 3516
rect 148100 3476 148106 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149164 3516 149192 3624
rect 149238 3612 149244 3664
rect 149296 3652 149302 3664
rect 171597 3655 171655 3661
rect 171597 3652 171609 3655
rect 149296 3624 171609 3652
rect 149296 3612 149302 3624
rect 171597 3621 171609 3624
rect 171643 3621 171655 3655
rect 173894 3652 173900 3664
rect 171597 3615 171655 3621
rect 171704 3624 173900 3652
rect 171704 3584 171732 3624
rect 173894 3612 173900 3624
rect 173952 3612 173958 3664
rect 180150 3612 180156 3664
rect 180208 3652 180214 3664
rect 180702 3652 180708 3664
rect 180208 3624 180708 3652
rect 180208 3612 180214 3624
rect 180702 3612 180708 3624
rect 180760 3612 180766 3664
rect 181346 3612 181352 3664
rect 181404 3652 181410 3664
rect 204254 3652 204260 3664
rect 181404 3624 204260 3652
rect 181404 3612 181410 3624
rect 204254 3612 204260 3624
rect 204312 3612 204318 3664
rect 157352 3556 171732 3584
rect 157352 3516 157380 3556
rect 171778 3544 171784 3596
rect 171836 3584 171842 3596
rect 172422 3584 172428 3596
rect 171836 3556 172428 3584
rect 171836 3544 171842 3556
rect 172422 3544 172428 3556
rect 172480 3544 172486 3596
rect 177758 3544 177764 3596
rect 177816 3584 177822 3596
rect 201494 3584 201500 3596
rect 177816 3556 201500 3584
rect 177816 3544 177822 3556
rect 201494 3544 201500 3556
rect 201552 3544 201558 3596
rect 206278 3544 206284 3596
rect 206336 3584 206342 3596
rect 206922 3584 206928 3596
rect 206336 3556 206928 3584
rect 206336 3544 206342 3556
rect 206922 3544 206928 3556
rect 206980 3544 206986 3596
rect 207474 3544 207480 3596
rect 207532 3584 207538 3596
rect 208302 3584 208308 3596
rect 207532 3556 208308 3584
rect 207532 3544 207538 3556
rect 208302 3544 208308 3556
rect 208360 3544 208366 3596
rect 208412 3584 208440 3692
rect 208670 3680 208676 3732
rect 208728 3720 208734 3732
rect 221108 3720 221136 3760
rect 226426 3748 226432 3760
rect 226484 3748 226490 3800
rect 228910 3748 228916 3800
rect 228968 3788 228974 3800
rect 232498 3788 232504 3800
rect 228968 3760 232504 3788
rect 228968 3748 228974 3760
rect 232498 3748 232504 3760
rect 232556 3748 232562 3800
rect 315298 3748 315304 3800
rect 315356 3788 315362 3800
rect 319254 3788 319260 3800
rect 315356 3760 319260 3788
rect 315356 3748 315362 3760
rect 319254 3748 319260 3760
rect 319312 3748 319318 3800
rect 339402 3748 339408 3800
rect 339460 3788 339466 3800
rect 350258 3788 350264 3800
rect 339460 3760 350264 3788
rect 339460 3748 339466 3760
rect 350258 3748 350264 3760
rect 350316 3748 350322 3800
rect 351822 3748 351828 3800
rect 351880 3788 351886 3800
rect 366910 3788 366916 3800
rect 351880 3760 366916 3788
rect 351880 3748 351886 3760
rect 366910 3748 366916 3760
rect 366968 3748 366974 3800
rect 369670 3748 369676 3800
rect 369728 3788 369734 3800
rect 388254 3788 388260 3800
rect 369728 3760 388260 3788
rect 369728 3748 369734 3760
rect 388254 3748 388260 3760
rect 388312 3748 388318 3800
rect 390462 3748 390468 3800
rect 390520 3788 390526 3800
rect 414474 3788 414480 3800
rect 390520 3760 414480 3788
rect 390520 3748 390526 3760
rect 414474 3748 414480 3760
rect 414532 3748 414538 3800
rect 423582 3748 423588 3800
rect 423640 3788 423646 3800
rect 457254 3788 457260 3800
rect 423640 3760 457260 3788
rect 423640 3748 423646 3760
rect 457254 3748 457260 3760
rect 457312 3748 457318 3800
rect 460842 3748 460848 3800
rect 460900 3788 460906 3800
rect 503622 3788 503628 3800
rect 460900 3760 503628 3788
rect 460900 3748 460906 3760
rect 503622 3748 503628 3760
rect 503680 3748 503686 3800
rect 516042 3748 516048 3800
rect 516100 3788 516106 3800
rect 573818 3788 573824 3800
rect 516100 3760 573824 3788
rect 516100 3748 516106 3760
rect 573818 3748 573824 3760
rect 573876 3748 573882 3800
rect 223758 3720 223764 3732
rect 208728 3692 221136 3720
rect 221200 3692 223764 3720
rect 208728 3680 208734 3692
rect 208489 3655 208547 3661
rect 208489 3621 208501 3655
rect 208535 3652 208547 3655
rect 221200 3652 221228 3692
rect 223758 3680 223764 3692
rect 223816 3680 223822 3732
rect 226518 3680 226524 3732
rect 226576 3720 226582 3732
rect 229097 3723 229155 3729
rect 229097 3720 229109 3723
rect 226576 3692 229109 3720
rect 226576 3680 226582 3692
rect 229097 3689 229109 3692
rect 229143 3689 229155 3723
rect 229097 3683 229155 3689
rect 231121 3723 231179 3729
rect 231121 3689 231133 3723
rect 231167 3720 231179 3723
rect 237374 3720 237380 3732
rect 231167 3692 237380 3720
rect 231167 3689 231179 3692
rect 231121 3683 231179 3689
rect 237374 3680 237380 3692
rect 237432 3680 237438 3732
rect 313090 3680 313096 3732
rect 313148 3720 313154 3732
rect 318058 3720 318064 3732
rect 313148 3692 318064 3720
rect 313148 3680 313154 3692
rect 318058 3680 318064 3692
rect 318116 3680 318122 3732
rect 325602 3680 325608 3732
rect 325660 3720 325666 3732
rect 333606 3720 333612 3732
rect 325660 3692 333612 3720
rect 325660 3680 325666 3692
rect 333606 3680 333612 3692
rect 333664 3680 333670 3732
rect 333790 3680 333796 3732
rect 333848 3720 333854 3732
rect 344278 3720 344284 3732
rect 333848 3692 344284 3720
rect 333848 3680 333854 3692
rect 344278 3680 344284 3692
rect 344336 3680 344342 3732
rect 348970 3680 348976 3732
rect 349028 3720 349034 3732
rect 362126 3720 362132 3732
rect 349028 3692 362132 3720
rect 349028 3680 349034 3692
rect 362126 3680 362132 3692
rect 362184 3680 362190 3732
rect 362862 3680 362868 3732
rect 362920 3720 362926 3732
rect 381170 3720 381176 3732
rect 362920 3692 381176 3720
rect 362920 3680 362926 3692
rect 381170 3680 381176 3692
rect 381228 3680 381234 3732
rect 383562 3680 383568 3732
rect 383620 3720 383626 3732
rect 407298 3720 407304 3732
rect 383620 3692 407304 3720
rect 383620 3680 383626 3692
rect 407298 3680 407304 3692
rect 407356 3680 407362 3732
rect 418062 3680 418068 3732
rect 418120 3720 418126 3732
rect 450170 3720 450176 3732
rect 418120 3692 450176 3720
rect 418120 3680 418126 3692
rect 450170 3680 450176 3692
rect 450228 3680 450234 3732
rect 451274 3680 451280 3732
rect 451332 3720 451338 3732
rect 452470 3720 452476 3732
rect 451332 3692 452476 3720
rect 451332 3680 451338 3692
rect 452470 3680 452476 3692
rect 452528 3680 452534 3732
rect 453942 3680 453948 3732
rect 454000 3720 454006 3732
rect 496538 3720 496544 3732
rect 454000 3692 496544 3720
rect 454000 3680 454006 3692
rect 496538 3680 496544 3692
rect 496596 3680 496602 3732
rect 513282 3680 513288 3732
rect 513340 3720 513346 3732
rect 570230 3720 570236 3732
rect 513340 3692 570236 3720
rect 513340 3680 513346 3692
rect 570230 3680 570236 3692
rect 570288 3680 570294 3732
rect 208535 3624 221228 3652
rect 208535 3621 208547 3624
rect 208489 3615 208547 3621
rect 222930 3612 222936 3664
rect 222988 3652 222994 3664
rect 247126 3652 247132 3664
rect 222988 3624 226380 3652
rect 222988 3612 222994 3624
rect 222194 3584 222200 3596
rect 208412 3556 222200 3584
rect 222194 3544 222200 3556
rect 222252 3544 222258 3596
rect 225322 3544 225328 3596
rect 225380 3584 225386 3596
rect 226242 3584 226248 3596
rect 225380 3556 226248 3584
rect 225380 3544 225386 3556
rect 226242 3544 226248 3556
rect 226300 3544 226306 3596
rect 226352 3584 226380 3624
rect 239508 3624 247132 3652
rect 231121 3587 231179 3593
rect 231121 3584 231133 3587
rect 226352 3556 231133 3584
rect 231121 3553 231133 3556
rect 231167 3553 231179 3587
rect 234614 3584 234620 3596
rect 231121 3547 231179 3553
rect 231228 3556 234620 3584
rect 160278 3516 160284 3528
rect 149164 3488 157380 3516
rect 157444 3488 160284 3516
rect 157444 3448 157472 3488
rect 160278 3476 160284 3488
rect 160336 3476 160342 3528
rect 168190 3476 168196 3528
rect 168248 3516 168254 3528
rect 194594 3516 194600 3528
rect 168248 3488 194600 3516
rect 168248 3476 168254 3488
rect 194594 3476 194600 3488
rect 194652 3476 194658 3528
rect 197998 3476 198004 3528
rect 198056 3516 198062 3528
rect 213917 3519 213975 3525
rect 213917 3516 213929 3519
rect 198056 3488 213929 3516
rect 198056 3476 198062 3488
rect 213917 3485 213929 3488
rect 213963 3485 213975 3519
rect 213917 3479 213975 3485
rect 214650 3476 214656 3528
rect 214708 3516 214714 3528
rect 215202 3516 215208 3528
rect 214708 3488 215208 3516
rect 214708 3476 214714 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 217042 3476 217048 3528
rect 217100 3516 217106 3528
rect 217962 3516 217968 3528
rect 217100 3488 217968 3516
rect 217100 3476 217106 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 219342 3476 219348 3528
rect 219400 3516 219406 3528
rect 231228 3516 231256 3556
rect 234614 3544 234620 3556
rect 234672 3544 234678 3596
rect 235994 3544 236000 3596
rect 236052 3584 236058 3596
rect 237190 3584 237196 3596
rect 236052 3556 237196 3584
rect 236052 3544 236058 3556
rect 237190 3544 237196 3556
rect 237248 3544 237254 3596
rect 219400 3488 231256 3516
rect 219400 3476 219406 3488
rect 231302 3476 231308 3528
rect 231360 3516 231366 3528
rect 231762 3516 231768 3528
rect 231360 3488 231768 3516
rect 231360 3476 231366 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232498 3476 232504 3528
rect 232556 3516 232562 3528
rect 233142 3516 233148 3528
rect 232556 3488 233148 3516
rect 232556 3476 232562 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233694 3476 233700 3528
rect 233752 3516 233758 3528
rect 234522 3516 234528 3528
rect 233752 3488 234528 3516
rect 233752 3476 233758 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234798 3476 234804 3528
rect 234856 3516 234862 3528
rect 239508 3516 239536 3624
rect 247126 3612 247132 3624
rect 247184 3612 247190 3664
rect 285950 3612 285956 3664
rect 286008 3652 286014 3664
rect 286962 3652 286968 3664
rect 286008 3624 286968 3652
rect 286008 3612 286014 3624
rect 286962 3612 286968 3624
rect 287020 3612 287026 3664
rect 315942 3612 315948 3664
rect 316000 3652 316006 3664
rect 320450 3652 320456 3664
rect 316000 3624 320456 3652
rect 316000 3612 316006 3624
rect 320450 3612 320456 3624
rect 320508 3612 320514 3664
rect 324222 3612 324228 3664
rect 324280 3652 324286 3664
rect 331214 3652 331220 3664
rect 324280 3624 331220 3652
rect 324280 3612 324286 3624
rect 331214 3612 331220 3624
rect 331272 3612 331278 3664
rect 336550 3612 336556 3664
rect 336608 3652 336614 3664
rect 347866 3652 347872 3664
rect 336608 3624 347872 3652
rect 336608 3612 336614 3624
rect 347866 3612 347872 3624
rect 347924 3612 347930 3664
rect 355962 3612 355968 3664
rect 356020 3652 356026 3664
rect 371602 3652 371608 3664
rect 356020 3624 371608 3652
rect 356020 3612 356026 3624
rect 371602 3612 371608 3624
rect 371660 3612 371666 3664
rect 377950 3612 377956 3664
rect 378008 3652 378014 3664
rect 400214 3652 400220 3664
rect 378008 3624 400220 3652
rect 378008 3612 378014 3624
rect 400214 3612 400220 3624
rect 400272 3612 400278 3664
rect 401502 3612 401508 3664
rect 401560 3652 401566 3664
rect 428734 3652 428740 3664
rect 401560 3624 428740 3652
rect 401560 3612 401566 3624
rect 428734 3612 428740 3624
rect 428792 3612 428798 3664
rect 434622 3612 434628 3664
rect 434680 3652 434686 3664
rect 471514 3652 471520 3664
rect 434680 3624 471520 3652
rect 434680 3612 434686 3624
rect 471514 3612 471520 3624
rect 471572 3612 471578 3664
rect 471882 3612 471888 3664
rect 471940 3652 471946 3664
rect 517882 3652 517888 3664
rect 471940 3624 517888 3652
rect 471940 3612 471946 3624
rect 517882 3612 517888 3624
rect 517940 3612 517946 3664
rect 518802 3612 518808 3664
rect 518860 3652 518866 3664
rect 577406 3652 577412 3664
rect 518860 3624 577412 3652
rect 518860 3612 518866 3624
rect 577406 3612 577412 3624
rect 577464 3612 577470 3664
rect 302050 3544 302056 3596
rect 302108 3584 302114 3596
rect 303798 3584 303804 3596
rect 302108 3556 303804 3584
rect 302108 3544 302114 3556
rect 303798 3544 303804 3556
rect 303856 3544 303862 3596
rect 309042 3544 309048 3596
rect 309100 3584 309106 3596
rect 312170 3584 312176 3596
rect 309100 3556 312176 3584
rect 309100 3544 309106 3556
rect 312170 3544 312176 3556
rect 312228 3544 312234 3596
rect 322750 3544 322756 3596
rect 322808 3584 322814 3596
rect 328822 3584 328828 3596
rect 322808 3556 328828 3584
rect 322808 3544 322814 3556
rect 328822 3544 328828 3556
rect 328880 3544 328886 3596
rect 329742 3544 329748 3596
rect 329800 3584 329806 3596
rect 338298 3584 338304 3596
rect 329800 3556 338304 3584
rect 329800 3544 329806 3556
rect 338298 3544 338304 3556
rect 338356 3544 338362 3596
rect 339310 3544 339316 3596
rect 339368 3584 339374 3596
rect 351362 3584 351368 3596
rect 339368 3556 351368 3584
rect 339368 3544 339374 3556
rect 351362 3544 351368 3556
rect 351420 3544 351426 3596
rect 354490 3544 354496 3596
rect 354548 3584 354554 3596
rect 369210 3584 369216 3596
rect 354548 3556 369216 3584
rect 354548 3544 354554 3556
rect 369210 3544 369216 3556
rect 369268 3544 369274 3596
rect 369762 3544 369768 3596
rect 369820 3584 369826 3596
rect 389450 3584 389456 3596
rect 369820 3556 389456 3584
rect 369820 3544 369826 3556
rect 389450 3544 389456 3556
rect 389508 3544 389514 3596
rect 395982 3544 395988 3596
rect 396040 3584 396046 3596
rect 421558 3584 421564 3596
rect 396040 3556 421564 3584
rect 396040 3544 396046 3556
rect 421558 3544 421564 3556
rect 421616 3544 421622 3596
rect 426342 3544 426348 3596
rect 426400 3584 426406 3596
rect 460842 3584 460848 3596
rect 426400 3556 460848 3584
rect 426400 3544 426406 3556
rect 460842 3544 460848 3556
rect 460900 3544 460906 3596
rect 463602 3544 463608 3596
rect 463660 3584 463666 3596
rect 468941 3587 468999 3593
rect 468941 3584 468953 3587
rect 463660 3556 468953 3584
rect 463660 3544 463666 3556
rect 468941 3553 468953 3556
rect 468987 3553 468999 3587
rect 468941 3547 468999 3553
rect 469030 3544 469036 3596
rect 469088 3584 469094 3596
rect 469309 3587 469367 3593
rect 469088 3556 469260 3584
rect 469088 3544 469094 3556
rect 234856 3488 239536 3516
rect 234856 3476 234862 3488
rect 239582 3476 239588 3528
rect 239640 3516 239646 3528
rect 240042 3516 240048 3528
rect 239640 3488 240048 3516
rect 239640 3476 239646 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 240778 3476 240784 3528
rect 240836 3516 240842 3528
rect 241422 3516 241428 3528
rect 240836 3488 241428 3516
rect 240836 3476 240842 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 241974 3476 241980 3528
rect 242032 3516 242038 3528
rect 242802 3516 242808 3528
rect 242032 3488 242808 3516
rect 242032 3476 242038 3488
rect 242802 3476 242808 3488
rect 242860 3476 242866 3528
rect 243170 3476 243176 3528
rect 243228 3516 243234 3528
rect 244182 3516 244188 3528
rect 243228 3488 244188 3516
rect 243228 3476 243234 3488
rect 244182 3476 244188 3488
rect 244240 3476 244246 3528
rect 244366 3476 244372 3528
rect 244424 3516 244430 3528
rect 245470 3516 245476 3528
rect 244424 3488 245476 3516
rect 244424 3476 244430 3488
rect 245470 3476 245476 3488
rect 245528 3476 245534 3528
rect 249150 3476 249156 3528
rect 249208 3516 249214 3528
rect 249702 3516 249708 3528
rect 249208 3488 249708 3516
rect 249208 3476 249214 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 250346 3476 250352 3528
rect 250404 3516 250410 3528
rect 251082 3516 251088 3528
rect 250404 3488 251088 3516
rect 250404 3476 250410 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251450 3476 251456 3528
rect 251508 3516 251514 3528
rect 252462 3516 252468 3528
rect 251508 3488 252468 3516
rect 251508 3476 251514 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 252646 3476 252652 3528
rect 252704 3516 252710 3528
rect 253842 3516 253848 3528
rect 252704 3488 253848 3516
rect 252704 3476 252710 3488
rect 253842 3476 253848 3488
rect 253900 3476 253906 3528
rect 257430 3476 257436 3528
rect 257488 3516 257494 3528
rect 257982 3516 257988 3528
rect 257488 3488 257988 3516
rect 257488 3476 257494 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 259822 3476 259828 3528
rect 259880 3516 259886 3528
rect 261478 3516 261484 3528
rect 259880 3488 261484 3516
rect 259880 3476 259886 3488
rect 261478 3476 261484 3488
rect 261536 3476 261542 3528
rect 262214 3476 262220 3528
rect 262272 3516 262278 3528
rect 263502 3516 263508 3528
rect 262272 3488 263508 3516
rect 262272 3476 262278 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 265802 3476 265808 3528
rect 265860 3516 265866 3528
rect 266262 3516 266268 3528
rect 265860 3488 266268 3516
rect 265860 3476 265866 3488
rect 266262 3476 266268 3488
rect 266320 3476 266326 3528
rect 268102 3476 268108 3528
rect 268160 3516 268166 3528
rect 269022 3516 269028 3528
rect 268160 3488 269028 3516
rect 268160 3476 268166 3488
rect 269022 3476 269028 3488
rect 269080 3476 269086 3528
rect 270494 3476 270500 3528
rect 270552 3516 270558 3528
rect 272518 3516 272524 3528
rect 270552 3488 272524 3516
rect 270552 3476 270558 3488
rect 272518 3476 272524 3488
rect 272576 3476 272582 3528
rect 274082 3476 274088 3528
rect 274140 3516 274146 3528
rect 274542 3516 274548 3528
rect 274140 3488 274548 3516
rect 274140 3476 274146 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 275278 3476 275284 3528
rect 275336 3516 275342 3528
rect 275922 3516 275928 3528
rect 275336 3488 275928 3516
rect 275336 3476 275342 3488
rect 275922 3476 275928 3488
rect 275980 3476 275986 3528
rect 276474 3476 276480 3528
rect 276532 3516 276538 3528
rect 277302 3516 277308 3528
rect 276532 3488 277308 3516
rect 276532 3476 276538 3488
rect 277302 3476 277308 3488
rect 277360 3476 277366 3528
rect 302142 3476 302148 3528
rect 302200 3516 302206 3528
rect 302602 3516 302608 3528
rect 302200 3488 302608 3516
rect 302200 3476 302206 3488
rect 302602 3476 302608 3488
rect 302660 3476 302666 3528
rect 304902 3476 304908 3528
rect 304960 3516 304966 3528
rect 306190 3516 306196 3528
rect 304960 3488 306196 3516
rect 304960 3476 304966 3488
rect 306190 3476 306196 3488
rect 306248 3476 306254 3528
rect 310422 3476 310428 3528
rect 310480 3516 310486 3528
rect 313366 3516 313372 3528
rect 310480 3488 313372 3516
rect 310480 3476 310486 3488
rect 313366 3476 313372 3488
rect 313424 3476 313430 3528
rect 316954 3516 316960 3528
rect 313476 3488 316960 3516
rect 147968 3420 157472 3448
rect 147861 3411 147919 3417
rect 157518 3408 157524 3460
rect 157576 3448 157582 3460
rect 158622 3448 158628 3460
rect 157576 3420 158628 3448
rect 157576 3408 157582 3420
rect 158622 3408 158628 3420
rect 158680 3408 158686 3460
rect 161106 3408 161112 3460
rect 161164 3448 161170 3460
rect 189074 3448 189080 3460
rect 161164 3420 189080 3448
rect 161164 3408 161170 3420
rect 189074 3408 189080 3420
rect 189132 3408 189138 3460
rect 189626 3408 189632 3460
rect 189684 3448 189690 3460
rect 211154 3448 211160 3460
rect 189684 3420 211160 3448
rect 189684 3408 189690 3420
rect 211154 3408 211160 3420
rect 211212 3408 211218 3460
rect 212258 3408 212264 3460
rect 212316 3448 212322 3460
rect 229094 3448 229100 3460
rect 212316 3420 229100 3448
rect 212316 3408 212322 3420
rect 229094 3408 229100 3420
rect 229152 3408 229158 3460
rect 230106 3408 230112 3460
rect 230164 3448 230170 3460
rect 242986 3448 242992 3460
rect 230164 3420 242992 3448
rect 230164 3408 230170 3420
rect 242986 3408 242992 3420
rect 243044 3408 243050 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 267642 3448 267648 3460
rect 267056 3420 267648 3448
rect 267056 3408 267062 3420
rect 267642 3408 267648 3420
rect 267700 3408 267706 3460
rect 277670 3408 277676 3460
rect 277728 3448 277734 3460
rect 280246 3448 280252 3460
rect 277728 3420 280252 3448
rect 277728 3408 277734 3420
rect 280246 3408 280252 3420
rect 280304 3408 280310 3460
rect 303522 3408 303528 3460
rect 303580 3448 303586 3460
rect 304994 3448 305000 3460
rect 303580 3420 305000 3448
rect 303580 3408 303586 3420
rect 304994 3408 305000 3420
rect 305052 3408 305058 3460
rect 307662 3408 307668 3460
rect 307720 3448 307726 3460
rect 310974 3448 310980 3460
rect 307720 3420 310980 3448
rect 307720 3408 307726 3420
rect 310974 3408 310980 3420
rect 311032 3408 311038 3460
rect 313182 3408 313188 3460
rect 313240 3448 313246 3460
rect 313476 3448 313504 3488
rect 316954 3476 316960 3488
rect 317012 3476 317018 3528
rect 318702 3476 318708 3528
rect 318760 3516 318766 3528
rect 325234 3516 325240 3528
rect 318760 3488 325240 3516
rect 318760 3476 318766 3488
rect 325234 3476 325240 3488
rect 325292 3476 325298 3528
rect 326338 3476 326344 3528
rect 326396 3516 326402 3528
rect 332410 3516 332416 3528
rect 326396 3488 332416 3516
rect 326396 3476 326402 3488
rect 332410 3476 332416 3488
rect 332468 3476 332474 3528
rect 337102 3516 337108 3528
rect 332520 3488 337108 3516
rect 313240 3420 313504 3448
rect 313240 3408 313246 3420
rect 315850 3408 315856 3460
rect 315908 3448 315914 3460
rect 321646 3448 321652 3460
rect 315908 3420 321652 3448
rect 315908 3408 315914 3420
rect 321646 3408 321652 3420
rect 321704 3408 321710 3460
rect 322842 3408 322848 3460
rect 322900 3448 322906 3460
rect 330018 3448 330024 3460
rect 322900 3420 330024 3448
rect 322900 3408 322906 3420
rect 330018 3408 330024 3420
rect 330076 3408 330082 3460
rect 4120 3352 4200 3380
rect 4120 3340 4126 3352
rect 18322 3340 18328 3392
rect 18380 3380 18386 3392
rect 19978 3380 19984 3392
rect 18380 3352 19984 3380
rect 18380 3340 18386 3352
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 26694 3340 26700 3392
rect 26752 3380 26758 3392
rect 27522 3380 27528 3392
rect 26752 3352 27528 3380
rect 26752 3340 26758 3352
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28902 3380 28908 3392
rect 27948 3352 28908 3380
rect 27948 3340 27954 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 33870 3340 33876 3392
rect 33928 3380 33934 3392
rect 34422 3380 34428 3392
rect 33928 3352 34428 3380
rect 33928 3340 33934 3352
rect 34422 3340 34428 3352
rect 34480 3340 34486 3392
rect 34974 3340 34980 3392
rect 35032 3380 35038 3392
rect 35802 3380 35808 3392
rect 35032 3352 35808 3380
rect 35032 3340 35038 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 37366 3340 37372 3392
rect 37424 3380 37430 3392
rect 38470 3380 38476 3392
rect 37424 3352 38476 3380
rect 37424 3340 37430 3352
rect 38470 3340 38476 3352
rect 38528 3340 38534 3392
rect 42150 3340 42156 3392
rect 42208 3380 42214 3392
rect 42702 3380 42708 3392
rect 42208 3352 42708 3380
rect 42208 3340 42214 3352
rect 42702 3340 42708 3352
rect 42760 3340 42766 3392
rect 50522 3340 50528 3392
rect 50580 3380 50586 3392
rect 50982 3380 50988 3392
rect 50580 3352 50988 3380
rect 50580 3340 50586 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 52822 3340 52828 3392
rect 52880 3380 52886 3392
rect 53742 3380 53748 3392
rect 52880 3352 53748 3380
rect 52880 3340 52886 3352
rect 53742 3340 53748 3352
rect 53800 3340 53806 3392
rect 95605 3383 95663 3389
rect 95605 3380 95617 3383
rect 53852 3352 95617 3380
rect 44542 3272 44548 3324
rect 44600 3312 44606 3324
rect 45462 3312 45468 3324
rect 44600 3284 45468 3312
rect 44600 3272 44606 3284
rect 45462 3272 45468 3284
rect 45520 3272 45526 3324
rect 46934 3272 46940 3324
rect 46992 3312 46998 3324
rect 53852 3312 53880 3352
rect 95605 3349 95617 3352
rect 95651 3349 95663 3383
rect 95605 3343 95663 3349
rect 95694 3340 95700 3392
rect 95752 3380 95758 3392
rect 96522 3380 96528 3392
rect 95752 3352 96528 3380
rect 95752 3340 95758 3352
rect 96522 3340 96528 3352
rect 96580 3340 96586 3392
rect 98086 3340 98092 3392
rect 98144 3380 98150 3392
rect 99282 3380 99288 3392
rect 98144 3352 99288 3380
rect 98144 3340 98150 3352
rect 99282 3340 99288 3352
rect 99340 3340 99346 3392
rect 101582 3340 101588 3392
rect 101640 3380 101646 3392
rect 102042 3380 102048 3392
rect 101640 3352 102048 3380
rect 101640 3340 101646 3352
rect 102042 3340 102048 3352
rect 102100 3340 102106 3392
rect 102778 3340 102784 3392
rect 102836 3380 102842 3392
rect 103422 3380 103428 3392
rect 102836 3352 103428 3380
rect 102836 3340 102842 3352
rect 103422 3340 103428 3352
rect 103480 3340 103486 3392
rect 105170 3340 105176 3392
rect 105228 3380 105234 3392
rect 106182 3380 106188 3392
rect 105228 3352 106188 3380
rect 105228 3340 105234 3352
rect 106182 3340 106188 3352
rect 106240 3340 106246 3392
rect 113542 3340 113548 3392
rect 113600 3380 113606 3392
rect 150802 3380 150808 3392
rect 113600 3352 150808 3380
rect 113600 3340 113606 3352
rect 150802 3340 150808 3352
rect 150860 3340 150866 3392
rect 152734 3340 152740 3392
rect 152792 3380 152798 3392
rect 162121 3383 162179 3389
rect 162121 3380 162133 3383
rect 152792 3352 162133 3380
rect 152792 3340 152798 3352
rect 162121 3349 162133 3352
rect 162167 3349 162179 3383
rect 162121 3343 162179 3349
rect 175366 3340 175372 3392
rect 175424 3380 175430 3392
rect 200114 3380 200120 3392
rect 175424 3352 200120 3380
rect 175424 3340 175430 3352
rect 200114 3340 200120 3352
rect 200172 3340 200178 3392
rect 200390 3340 200396 3392
rect 200448 3380 200454 3392
rect 219526 3380 219532 3392
rect 200448 3352 219532 3380
rect 200448 3340 200454 3352
rect 219526 3340 219532 3352
rect 219584 3340 219590 3392
rect 227714 3340 227720 3392
rect 227772 3380 227778 3392
rect 229002 3380 229008 3392
rect 227772 3352 229008 3380
rect 227772 3340 227778 3352
rect 229002 3340 229008 3352
rect 229060 3340 229066 3392
rect 310330 3340 310336 3392
rect 310388 3380 310394 3392
rect 314562 3380 314568 3392
rect 310388 3352 314568 3380
rect 310388 3340 310394 3352
rect 314562 3340 314568 3352
rect 314620 3340 314626 3392
rect 328270 3340 328276 3392
rect 328328 3380 328334 3392
rect 332520 3380 332548 3488
rect 337102 3476 337108 3488
rect 337160 3476 337166 3528
rect 343542 3476 343548 3528
rect 343600 3516 343606 3528
rect 356146 3516 356152 3528
rect 343600 3488 356152 3516
rect 343600 3476 343606 3488
rect 356146 3476 356152 3488
rect 356204 3476 356210 3528
rect 357342 3476 357348 3528
rect 357400 3516 357406 3528
rect 373994 3516 374000 3528
rect 357400 3488 374000 3516
rect 357400 3476 357406 3488
rect 373994 3476 374000 3488
rect 374052 3476 374058 3528
rect 375190 3476 375196 3528
rect 375248 3516 375254 3528
rect 396626 3516 396632 3528
rect 375248 3488 396632 3516
rect 375248 3476 375254 3488
rect 396626 3476 396632 3488
rect 396684 3476 396690 3528
rect 398742 3476 398748 3528
rect 398800 3516 398806 3528
rect 425146 3516 425152 3528
rect 398800 3488 425152 3516
rect 398800 3476 398806 3488
rect 425146 3476 425152 3488
rect 425204 3476 425210 3528
rect 431862 3476 431868 3528
rect 431920 3516 431926 3528
rect 467834 3516 467840 3528
rect 431920 3488 467840 3516
rect 431920 3476 431926 3488
rect 467834 3476 467840 3488
rect 467892 3476 467898 3528
rect 467926 3476 467932 3528
rect 467984 3516 467990 3528
rect 469122 3516 469128 3528
rect 467984 3488 469128 3516
rect 467984 3476 467990 3488
rect 469122 3476 469128 3488
rect 469180 3476 469186 3528
rect 469232 3516 469260 3556
rect 469309 3553 469321 3587
rect 469355 3584 469367 3587
rect 507210 3584 507216 3596
rect 469355 3556 507216 3584
rect 469355 3553 469367 3556
rect 469309 3547 469367 3553
rect 507210 3544 507216 3556
rect 507268 3544 507274 3596
rect 513098 3544 513104 3596
rect 513156 3584 513162 3596
rect 571426 3584 571432 3596
rect 513156 3556 571432 3584
rect 513156 3544 513162 3556
rect 571426 3544 571432 3556
rect 571484 3544 571490 3596
rect 575014 3584 575020 3596
rect 571536 3556 575020 3584
rect 514386 3516 514392 3528
rect 469232 3488 514392 3516
rect 514386 3476 514392 3488
rect 514444 3476 514450 3528
rect 515950 3476 515956 3528
rect 516008 3516 516014 3528
rect 571536 3516 571564 3556
rect 575014 3544 575020 3556
rect 575072 3544 575078 3596
rect 516008 3488 571564 3516
rect 516008 3476 516014 3488
rect 574738 3476 574744 3528
rect 574796 3516 574802 3528
rect 576210 3516 576216 3528
rect 574796 3488 576216 3516
rect 574796 3476 574802 3488
rect 576210 3476 576216 3488
rect 576268 3476 576274 3528
rect 340690 3448 340696 3460
rect 328328 3352 332548 3380
rect 332612 3420 340696 3448
rect 328328 3340 328334 3352
rect 46992 3284 53880 3312
rect 46992 3272 46998 3284
rect 54018 3272 54024 3324
rect 54076 3312 54082 3324
rect 103514 3312 103520 3324
rect 54076 3284 103520 3312
rect 54076 3272 54082 3284
rect 103514 3272 103520 3284
rect 103572 3272 103578 3324
rect 117130 3272 117136 3324
rect 117188 3312 117194 3324
rect 153194 3312 153200 3324
rect 117188 3284 153200 3312
rect 117188 3272 117194 3284
rect 153194 3272 153200 3284
rect 153252 3272 153258 3324
rect 174170 3272 174176 3324
rect 174228 3312 174234 3324
rect 198734 3312 198740 3324
rect 174228 3284 198740 3312
rect 174228 3272 174234 3284
rect 198734 3272 198740 3284
rect 198792 3272 198798 3324
rect 199194 3272 199200 3324
rect 199252 3312 199258 3324
rect 218330 3312 218336 3324
rect 199252 3284 218336 3312
rect 199252 3272 199258 3284
rect 218330 3272 218336 3284
rect 218388 3272 218394 3324
rect 253842 3272 253848 3324
rect 253900 3312 253906 3324
rect 257338 3312 257344 3324
rect 253900 3284 257344 3312
rect 253900 3272 253906 3284
rect 257338 3272 257344 3284
rect 257396 3272 257402 3324
rect 320818 3272 320824 3324
rect 320876 3312 320882 3324
rect 324038 3312 324044 3324
rect 320876 3284 324044 3312
rect 320876 3272 320882 3284
rect 324038 3272 324044 3284
rect 324096 3272 324102 3324
rect 331030 3272 331036 3324
rect 331088 3312 331094 3324
rect 332612 3312 332640 3420
rect 340690 3408 340696 3420
rect 340748 3408 340754 3460
rect 342070 3408 342076 3460
rect 342128 3448 342134 3460
rect 354950 3448 354956 3460
rect 342128 3420 354956 3448
rect 342128 3408 342134 3420
rect 354950 3408 354956 3420
rect 355008 3408 355014 3460
rect 360102 3408 360108 3460
rect 360160 3448 360166 3460
rect 377582 3448 377588 3460
rect 360160 3420 377588 3448
rect 360160 3408 360166 3420
rect 377582 3408 377588 3420
rect 377640 3408 377646 3460
rect 380710 3408 380716 3460
rect 380768 3448 380774 3460
rect 403710 3448 403716 3460
rect 380768 3420 403716 3448
rect 380768 3408 380774 3420
rect 403710 3408 403716 3420
rect 403768 3408 403774 3460
rect 404262 3408 404268 3460
rect 404320 3448 404326 3460
rect 432322 3448 432328 3460
rect 404320 3420 432328 3448
rect 404320 3408 404326 3420
rect 432322 3408 432328 3420
rect 432380 3408 432386 3460
rect 433334 3408 433340 3460
rect 433392 3448 433398 3460
rect 434622 3448 434628 3460
rect 433392 3420 434628 3448
rect 433392 3408 433398 3420
rect 434622 3408 434628 3420
rect 434680 3408 434686 3460
rect 437290 3408 437296 3460
rect 437348 3448 437354 3460
rect 473906 3448 473912 3460
rect 437348 3420 473912 3448
rect 437348 3408 437354 3420
rect 473906 3408 473912 3420
rect 473964 3408 473970 3460
rect 474642 3408 474648 3460
rect 474700 3448 474706 3460
rect 521378 3448 521384 3460
rect 474700 3420 521384 3448
rect 474700 3408 474706 3420
rect 521378 3408 521384 3420
rect 521436 3408 521442 3460
rect 521562 3408 521568 3460
rect 521620 3448 521626 3460
rect 580994 3448 581000 3460
rect 521620 3420 581000 3448
rect 521620 3408 521626 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 333882 3340 333888 3392
rect 333940 3380 333946 3392
rect 343082 3380 343088 3392
rect 333940 3352 343088 3380
rect 333940 3340 333946 3352
rect 343082 3340 343088 3352
rect 343140 3340 343146 3392
rect 346210 3340 346216 3392
rect 346268 3380 346274 3392
rect 358538 3380 358544 3392
rect 346268 3352 358544 3380
rect 346268 3340 346274 3352
rect 358538 3340 358544 3352
rect 358596 3340 358602 3392
rect 358722 3340 358728 3392
rect 358780 3380 358786 3392
rect 375190 3380 375196 3392
rect 358780 3352 375196 3380
rect 358780 3340 358786 3352
rect 375190 3340 375196 3352
rect 375248 3340 375254 3392
rect 378042 3340 378048 3392
rect 378100 3380 378106 3392
rect 399018 3380 399024 3392
rect 378100 3352 399024 3380
rect 378100 3340 378106 3352
rect 399018 3340 399024 3352
rect 399076 3340 399082 3392
rect 437382 3340 437388 3392
rect 437440 3380 437446 3392
rect 475102 3380 475108 3392
rect 437440 3352 475108 3380
rect 437440 3340 437446 3352
rect 475102 3340 475108 3352
rect 475160 3340 475166 3392
rect 495437 3383 495495 3389
rect 495437 3349 495449 3383
rect 495483 3380 495495 3383
rect 542906 3380 542912 3392
rect 495483 3352 542912 3380
rect 495483 3349 495495 3352
rect 495437 3343 495495 3349
rect 542906 3340 542912 3352
rect 542964 3340 542970 3392
rect 331088 3284 332640 3312
rect 331088 3272 331094 3284
rect 340782 3272 340788 3324
rect 340840 3312 340846 3324
rect 352558 3312 352564 3324
rect 340840 3284 352564 3312
rect 340840 3272 340846 3284
rect 352558 3272 352564 3284
rect 352616 3272 352622 3324
rect 353202 3272 353208 3324
rect 353260 3312 353266 3324
rect 368014 3312 368020 3324
rect 353260 3284 368020 3312
rect 353260 3272 353266 3284
rect 368014 3272 368020 3284
rect 368072 3272 368078 3324
rect 380802 3272 380808 3324
rect 380860 3312 380866 3324
rect 402514 3312 402520 3324
rect 380860 3284 402520 3312
rect 380860 3272 380866 3284
rect 402514 3272 402520 3284
rect 402572 3272 402578 3324
rect 440142 3272 440148 3324
rect 440200 3312 440206 3324
rect 477494 3312 477500 3324
rect 440200 3284 477500 3312
rect 440200 3272 440206 3284
rect 477494 3272 477500 3284
rect 477552 3272 477558 3324
rect 485682 3272 485688 3324
rect 485740 3312 485746 3324
rect 535730 3312 535736 3324
rect 485740 3284 535736 3312
rect 485740 3272 485746 3284
rect 535730 3272 535736 3284
rect 535788 3272 535794 3324
rect 536834 3272 536840 3324
rect 536892 3312 536898 3324
rect 538122 3312 538128 3324
rect 536892 3284 538128 3312
rect 536892 3272 536898 3284
rect 538122 3272 538128 3284
rect 538180 3272 538186 3324
rect 10042 3204 10048 3256
rect 10100 3244 10106 3256
rect 13078 3244 13084 3256
rect 10100 3216 13084 3244
rect 10100 3204 10106 3216
rect 13078 3204 13084 3216
rect 13136 3204 13142 3256
rect 61194 3204 61200 3256
rect 61252 3244 61258 3256
rect 109402 3244 109408 3256
rect 61252 3216 109408 3244
rect 61252 3204 61258 3216
rect 109402 3204 109408 3216
rect 109460 3204 109466 3256
rect 114738 3204 114744 3256
rect 114796 3244 114802 3256
rect 115842 3244 115848 3256
rect 114796 3216 115848 3244
rect 114796 3204 114802 3216
rect 115842 3204 115848 3216
rect 115900 3204 115906 3256
rect 120626 3204 120632 3256
rect 120684 3244 120690 3256
rect 155954 3244 155960 3256
rect 120684 3216 155960 3244
rect 120684 3204 120690 3216
rect 155954 3204 155960 3216
rect 156012 3204 156018 3256
rect 171597 3247 171655 3253
rect 171597 3213 171609 3247
rect 171643 3244 171655 3247
rect 179506 3244 179512 3256
rect 171643 3216 179512 3244
rect 171643 3213 171655 3216
rect 171597 3207 171655 3213
rect 179506 3204 179512 3216
rect 179564 3204 179570 3256
rect 193214 3204 193220 3256
rect 193272 3244 193278 3256
rect 214006 3244 214012 3256
rect 193272 3216 214012 3244
rect 193272 3204 193278 3216
rect 214006 3204 214012 3216
rect 214064 3204 214070 3256
rect 261018 3204 261024 3256
rect 261076 3244 261082 3256
rect 262122 3244 262128 3256
rect 261076 3216 262128 3244
rect 261076 3204 261082 3216
rect 262122 3204 262128 3216
rect 262180 3204 262186 3256
rect 312538 3204 312544 3256
rect 312596 3244 312602 3256
rect 315758 3244 315764 3256
rect 312596 3216 315764 3244
rect 312596 3204 312602 3216
rect 315758 3204 315764 3216
rect 315816 3204 315822 3256
rect 317322 3204 317328 3256
rect 317380 3244 317386 3256
rect 322842 3244 322848 3256
rect 317380 3216 322848 3244
rect 317380 3204 317386 3216
rect 322842 3204 322848 3216
rect 322900 3204 322906 3256
rect 344922 3204 344928 3256
rect 344980 3244 344986 3256
rect 357342 3244 357348 3256
rect 344980 3216 357348 3244
rect 344980 3204 344986 3216
rect 357342 3204 357348 3216
rect 357400 3204 357406 3256
rect 375282 3204 375288 3256
rect 375340 3244 375346 3256
rect 395430 3244 395436 3256
rect 375340 3216 395436 3244
rect 375340 3204 375346 3216
rect 395430 3204 395436 3216
rect 395488 3204 395494 3256
rect 429102 3204 429108 3256
rect 429160 3244 429166 3256
rect 464430 3244 464436 3256
rect 429160 3216 464436 3244
rect 429160 3204 429166 3216
rect 464430 3204 464436 3216
rect 464488 3204 464494 3256
rect 480162 3204 480168 3256
rect 480220 3244 480226 3256
rect 528646 3244 528652 3256
rect 480220 3216 528652 3244
rect 480220 3204 480226 3216
rect 528646 3204 528652 3216
rect 528704 3204 528710 3256
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 17218 3176 17224 3188
rect 16080 3148 17224 3176
rect 16080 3136 16086 3148
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 59909 3179 59967 3185
rect 59909 3145 59921 3179
rect 59955 3176 59967 3179
rect 66346 3176 66352 3188
rect 59955 3148 66352 3176
rect 59955 3145 59967 3148
rect 59909 3139 59967 3145
rect 66346 3136 66352 3148
rect 66404 3136 66410 3188
rect 71866 3136 71872 3188
rect 71924 3176 71930 3188
rect 113821 3179 113879 3185
rect 71924 3148 113404 3176
rect 71924 3136 71930 3148
rect 63497 3111 63555 3117
rect 63497 3077 63509 3111
rect 63543 3108 63555 3111
rect 73154 3108 73160 3120
rect 63543 3080 73160 3108
rect 63543 3077 63555 3080
rect 63497 3071 63555 3077
rect 73154 3068 73160 3080
rect 73212 3068 73218 3120
rect 81434 3068 81440 3120
rect 81492 3108 81498 3120
rect 82722 3108 82728 3120
rect 81492 3080 82728 3108
rect 81492 3068 81498 3080
rect 82722 3068 82728 3080
rect 82780 3068 82786 3120
rect 113376 3108 113404 3148
rect 113821 3145 113833 3179
rect 113867 3176 113879 3179
rect 121546 3176 121552 3188
rect 113867 3148 121552 3176
rect 113867 3145 113879 3148
rect 113821 3139 113879 3145
rect 121546 3136 121552 3148
rect 121604 3136 121610 3188
rect 121733 3179 121791 3185
rect 121733 3145 121745 3179
rect 121779 3176 121791 3179
rect 132494 3176 132500 3188
rect 121779 3148 132500 3176
rect 121779 3145 121791 3148
rect 121733 3139 121791 3145
rect 132494 3136 132500 3148
rect 132552 3136 132558 3188
rect 201494 3136 201500 3188
rect 201552 3176 201558 3188
rect 207201 3179 207259 3185
rect 207201 3176 207213 3179
rect 201552 3148 207213 3176
rect 201552 3136 201558 3148
rect 207201 3145 207213 3148
rect 207247 3145 207259 3179
rect 207201 3139 207259 3145
rect 209866 3136 209872 3188
rect 209924 3176 209930 3188
rect 226334 3176 226340 3188
rect 209924 3148 226340 3176
rect 209924 3136 209930 3148
rect 226334 3136 226340 3148
rect 226392 3136 226398 3188
rect 282454 3136 282460 3188
rect 282512 3176 282518 3188
rect 284294 3176 284300 3188
rect 282512 3148 284300 3176
rect 282512 3136 282518 3148
rect 284294 3136 284300 3148
rect 284352 3136 284358 3188
rect 372430 3136 372436 3188
rect 372488 3176 372494 3188
rect 391842 3176 391848 3188
rect 372488 3148 391848 3176
rect 372488 3136 372494 3148
rect 391842 3136 391848 3148
rect 391900 3136 391906 3188
rect 420822 3136 420828 3188
rect 420880 3176 420886 3188
rect 453666 3176 453672 3188
rect 420880 3148 453672 3176
rect 420880 3136 420886 3148
rect 453666 3136 453672 3148
rect 453724 3136 453730 3188
rect 118878 3108 118884 3120
rect 113376 3080 118884 3108
rect 118878 3068 118884 3080
rect 118936 3068 118942 3120
rect 164694 3068 164700 3120
rect 164752 3108 164758 3120
rect 165522 3108 165528 3120
rect 164752 3080 165528 3108
rect 164752 3068 164758 3080
rect 165522 3068 165528 3080
rect 165580 3068 165586 3120
rect 205082 3068 205088 3120
rect 205140 3108 205146 3120
rect 208489 3111 208547 3117
rect 208489 3108 208501 3111
rect 205140 3080 208501 3108
rect 205140 3068 205146 3080
rect 208489 3077 208501 3080
rect 208535 3077 208547 3111
rect 208489 3071 208547 3077
rect 258626 3068 258632 3120
rect 258684 3108 258690 3120
rect 259362 3108 259368 3120
rect 258684 3080 259368 3108
rect 258684 3068 258690 3080
rect 259362 3068 259368 3080
rect 259420 3068 259426 3120
rect 283650 3068 283656 3120
rect 283708 3108 283714 3120
rect 284202 3108 284208 3120
rect 283708 3080 284208 3108
rect 283708 3068 283714 3080
rect 284202 3068 284208 3080
rect 284260 3068 284266 3120
rect 138474 3000 138480 3052
rect 138532 3040 138538 3052
rect 139302 3040 139308 3052
rect 138532 3012 139308 3040
rect 138532 3000 138538 3012
rect 139302 3000 139308 3012
rect 139360 3000 139366 3052
rect 269298 3000 269304 3052
rect 269356 3040 269362 3052
rect 270402 3040 270408 3052
rect 269356 3012 270408 3040
rect 269356 3000 269362 3012
rect 270402 3000 270408 3012
rect 270460 3000 270466 3052
rect 321462 3000 321468 3052
rect 321520 3040 321526 3052
rect 327626 3040 327632 3052
rect 321520 3012 327632 3040
rect 321520 3000 321526 3012
rect 327626 3000 327632 3012
rect 327684 3000 327690 3052
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 10410 2972 10416 2984
rect 8904 2944 10416 2972
rect 8904 2932 8910 2944
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 87322 2864 87328 2916
rect 87380 2904 87386 2916
rect 88242 2904 88248 2916
rect 87380 2876 88248 2904
rect 87380 2864 87386 2876
rect 88242 2864 88248 2876
rect 88300 2864 88306 2916
rect 94498 2864 94504 2916
rect 94556 2904 94562 2916
rect 95142 2904 95148 2916
rect 94556 2876 95148 2904
rect 94556 2864 94562 2876
rect 95142 2864 95148 2876
rect 95200 2864 95206 2916
rect 326982 2864 326988 2916
rect 327040 2904 327046 2916
rect 334710 2904 334716 2916
rect 327040 2876 334716 2904
rect 327040 2864 327046 2876
rect 334710 2864 334716 2876
rect 334768 2864 334774 2916
rect 79042 824 79048 876
rect 79100 864 79106 876
rect 79962 864 79968 876
rect 79100 836 79968 864
rect 79100 824 79106 836
rect 79962 824 79968 836
rect 80020 824 80026 876
rect 74258 552 74264 604
rect 74316 592 74322 604
rect 74442 592 74448 604
rect 74316 564 74448 592
rect 74316 552 74322 564
rect 74442 552 74448 564
rect 74500 552 74506 604
rect 83826 552 83832 604
rect 83884 592 83890 604
rect 84102 592 84108 604
rect 83884 564 84108 592
rect 83884 552 83890 564
rect 84102 552 84108 564
rect 84160 552 84166 604
rect 151538 552 151544 604
rect 151596 592 151602 604
rect 151722 592 151728 604
rect 151596 564 151728 592
rect 151596 552 151602 564
rect 151722 552 151728 564
rect 151780 552 151786 604
rect 187234 552 187240 604
rect 187292 592 187298 604
rect 187602 592 187608 604
rect 187292 564 187608 592
rect 187292 552 187298 564
rect 187602 552 187608 564
rect 187660 552 187666 604
rect 220538 552 220544 604
rect 220596 592 220602 604
rect 220722 592 220728 604
rect 220596 564 220728 592
rect 220596 552 220602 564
rect 220722 552 220728 564
rect 220780 552 220786 604
rect 238386 552 238392 604
rect 238444 592 238450 604
rect 238662 592 238668 604
rect 238444 564 238668 592
rect 238444 552 238450 564
rect 238662 552 238668 564
rect 238720 552 238726 604
rect 386414 552 386420 604
rect 386472 592 386478 604
rect 387058 592 387064 604
rect 386472 564 387064 592
rect 386472 552 386478 564
rect 387058 552 387064 564
rect 387116 552 387122 604
rect 434714 552 434720 604
rect 434772 592 434778 604
rect 435818 592 435824 604
rect 434772 564 435824 592
rect 434772 552 434778 564
rect 435818 552 435824 564
rect 435876 552 435882 604
rect 437474 552 437480 604
rect 437532 592 437538 604
rect 438210 592 438216 604
rect 437532 564 438216 592
rect 437532 552 437538 564
rect 438210 552 438216 564
rect 438268 552 438274 604
rect 441614 552 441620 604
rect 441672 592 441678 604
rect 441798 592 441804 604
rect 441672 564 441804 592
rect 441672 552 441678 564
rect 441798 552 441804 564
rect 441856 552 441862 604
rect 443086 552 443092 604
rect 443144 592 443150 604
rect 444190 592 444196 604
rect 443144 564 444196 592
rect 443144 552 443150 564
rect 444190 552 444196 564
rect 444248 552 444254 604
rect 444374 552 444380 604
rect 444432 592 444438 604
rect 445386 592 445392 604
rect 444432 564 445392 592
rect 444432 552 444438 564
rect 445386 552 445392 564
rect 445444 552 445450 604
rect 448514 552 448520 604
rect 448572 592 448578 604
rect 448974 592 448980 604
rect 448572 564 448980 592
rect 448572 552 448578 564
rect 448974 552 448980 564
rect 449032 552 449038 604
rect 487062 552 487068 604
rect 487120 592 487126 604
rect 488166 592 488172 604
rect 487120 564 488172 592
rect 487120 552 487126 564
rect 488166 552 488172 564
rect 488224 552 488230 604
rect 491202 552 491208 604
rect 491260 592 491266 604
rect 491754 592 491760 604
rect 491260 564 491760 592
rect 491260 552 491266 564
rect 491754 552 491760 564
rect 491812 552 491818 604
rect 579614 552 579620 604
rect 579672 592 579678 604
rect 579798 592 579804 604
rect 579672 564 579804 592
rect 579672 552 579678 564
rect 579798 552 579804 564
rect 579856 552 579862 604
<< via1 >>
rect 54024 700816 54076 700868
rect 55128 700816 55180 700868
rect 429108 700408 429160 700460
rect 464988 700408 465040 700460
rect 480168 700408 480220 700460
rect 529848 700408 529900 700460
rect 360108 700340 360160 700392
rect 378416 700340 378468 700392
rect 394608 700340 394660 700392
rect 421748 700340 421800 700392
rect 445668 700340 445720 700392
rect 486608 700340 486660 700392
rect 496728 700340 496780 700392
rect 551468 700340 551520 700392
rect 343548 700272 343600 700324
rect 356796 700272 356848 700324
rect 378048 700272 378100 700324
rect 400128 700272 400180 700324
rect 411168 700272 411220 700324
rect 443368 700272 443420 700324
rect 463608 700272 463660 700324
rect 508228 700272 508280 700324
rect 514668 700272 514720 700324
rect 573088 700272 573140 700324
rect 183744 700136 183796 700188
rect 184848 700136 184900 700188
rect 32404 699660 32456 699712
rect 33048 699660 33100 699712
rect 97264 699660 97316 699712
rect 97908 699660 97960 699712
rect 118884 699660 118936 699712
rect 119988 699660 120040 699712
rect 162124 699660 162176 699712
rect 162768 699660 162820 699712
rect 227076 699660 227128 699712
rect 227628 699660 227680 699712
rect 248696 699660 248748 699712
rect 249708 699660 249760 699712
rect 291200 699660 291252 699712
rect 291936 699660 291988 699712
rect 309048 699660 309100 699712
rect 313556 699660 313608 699712
rect 326988 699660 327040 699712
rect 335176 699660 335228 699712
rect 75644 698343 75696 698352
rect 75644 698309 75653 698343
rect 75653 698309 75687 698343
rect 75687 698309 75696 698343
rect 75644 698300 75696 698309
rect 10692 695512 10744 695564
rect 10784 695512 10836 695564
rect 140412 695512 140464 695564
rect 140504 695512 140556 695564
rect 523684 695512 523736 695564
rect 580172 695512 580224 695564
rect 270408 695444 270460 695496
rect 75644 694195 75696 694204
rect 75644 694161 75653 694195
rect 75653 694161 75687 694195
rect 75687 694161 75696 694195
rect 75644 694152 75696 694161
rect 205640 694084 205692 694136
rect 75644 688644 75696 688696
rect 10692 688576 10744 688628
rect 10876 688576 10928 688628
rect 75552 688576 75604 688628
rect 140412 688576 140464 688628
rect 140596 688576 140648 688628
rect 270316 685899 270368 685908
rect 270316 685865 270325 685899
rect 270325 685865 270359 685899
rect 270359 685865 270368 685899
rect 270316 685856 270368 685865
rect 10876 685788 10928 685840
rect 140596 685788 140648 685840
rect 205548 684539 205600 684548
rect 205548 684505 205557 684539
rect 205557 684505 205591 684539
rect 205591 684505 205600 684539
rect 205548 684496 205600 684505
rect 523776 680348 523828 680400
rect 580172 680348 580224 680400
rect 75552 678988 75604 679040
rect 205548 678988 205600 679040
rect 270316 678988 270368 679040
rect 75460 678920 75512 678972
rect 205456 678920 205508 678972
rect 270224 678920 270276 678972
rect 10784 676243 10836 676252
rect 10784 676209 10793 676243
rect 10793 676209 10827 676243
rect 10827 676209 10836 676243
rect 10784 676200 10836 676209
rect 140504 676243 140556 676252
rect 140504 676209 140513 676243
rect 140513 676209 140547 676243
rect 140547 676209 140556 676243
rect 140504 676200 140556 676209
rect 10784 673480 10836 673532
rect 10968 673480 11020 673532
rect 140504 673480 140556 673532
rect 140688 673480 140740 673532
rect 270224 673480 270276 673532
rect 270408 673480 270460 673532
rect 205456 669332 205508 669384
rect 75460 669264 75512 669316
rect 75644 669264 75696 669316
rect 205364 669264 205416 669316
rect 75644 666476 75696 666528
rect 205364 659676 205416 659728
rect 205272 659608 205324 659660
rect 75552 656931 75604 656940
rect 75552 656897 75561 656931
rect 75561 656897 75595 656931
rect 75595 656897 75604 656931
rect 75552 656888 75604 656897
rect 249708 655460 249760 655512
rect 257896 655460 257948 655512
rect 270224 655460 270276 655512
rect 274916 655460 274968 655512
rect 377128 655460 377180 655512
rect 378048 655460 378100 655512
rect 428188 655460 428240 655512
rect 429108 655460 429160 655512
rect 462320 655460 462372 655512
rect 463608 655460 463660 655512
rect 479340 655460 479392 655512
rect 480168 655460 480220 655512
rect 513380 655256 513432 655308
rect 514668 655256 514720 655308
rect 325976 655120 326028 655172
rect 326988 655120 327040 655172
rect 55128 654916 55180 654968
rect 104532 654916 104584 654968
rect 119988 654916 120040 654968
rect 155592 654916 155644 654968
rect 33048 654848 33100 654900
rect 87512 654848 87564 654900
rect 97908 654848 97960 654900
rect 138572 654848 138624 654900
rect 162768 654848 162820 654900
rect 189724 654848 189776 654900
rect 205272 654848 205324 654900
rect 223764 654848 223816 654900
rect 10784 654780 10836 654832
rect 70492 654780 70544 654832
rect 75552 654780 75604 654832
rect 121552 654780 121604 654832
rect 140504 654780 140556 654832
rect 172704 654780 172756 654832
rect 184848 654780 184900 654832
rect 206744 654780 206796 654832
rect 227628 654780 227680 654832
rect 240784 654780 240836 654832
rect 3424 645804 3476 645856
rect 59360 645804 59412 645856
rect 523684 633428 523736 633480
rect 580172 633428 580224 633480
rect 3516 630572 3568 630624
rect 59360 630572 59412 630624
rect 524328 619556 524380 619608
rect 580264 619556 580316 619608
rect 3608 616768 3660 616820
rect 59360 616768 59412 616820
rect 523132 605752 523184 605804
rect 580356 605752 580408 605804
rect 3700 603032 3752 603084
rect 59360 603032 59412 603084
rect 523776 601672 523828 601724
rect 580172 601672 580224 601724
rect 3424 587800 3476 587852
rect 59360 587800 59412 587852
rect 523684 586508 523736 586560
rect 580172 586508 580224 586560
rect 524328 579572 524380 579624
rect 580264 579572 580316 579624
rect 3516 573996 3568 574048
rect 59360 573996 59412 574048
rect 3608 560192 3660 560244
rect 59360 560192 59412 560244
rect 523776 554752 523828 554804
rect 580172 554752 580224 554804
rect 3424 545028 3476 545080
rect 59360 545028 59412 545080
rect 523500 539588 523552 539640
rect 580172 539588 580224 539640
rect 523684 539520 523736 539572
rect 580264 539520 580316 539572
rect 3516 531224 3568 531276
rect 59360 531224 59412 531276
rect 523776 522996 523828 523048
rect 580172 522996 580224 523048
rect 3608 517420 3660 517472
rect 59360 517420 59412 517472
rect 523684 507832 523736 507884
rect 580172 507832 580224 507884
rect 3424 502256 3476 502308
rect 59360 502256 59412 502308
rect 523776 492668 523828 492720
rect 580172 492668 580224 492720
rect 3516 488452 3568 488504
rect 59360 488452 59412 488504
rect 523684 476076 523736 476128
rect 580172 476076 580224 476128
rect 3424 474648 3476 474700
rect 59360 474648 59412 474700
rect 523776 460912 523828 460964
rect 580172 460912 580224 460964
rect 3516 459484 3568 459536
rect 59360 459484 59412 459536
rect 523684 445748 523736 445800
rect 580172 445748 580224 445800
rect 3424 445680 3476 445732
rect 59360 445680 59412 445732
rect 3424 430516 3476 430568
rect 59360 430516 59412 430568
rect 523684 429156 523736 429208
rect 580172 429156 580224 429208
rect 3424 416712 3476 416764
rect 59360 416712 59412 416764
rect 523684 413992 523736 414044
rect 580172 413992 580224 414044
rect 3424 402908 3476 402960
rect 59360 402908 59412 402960
rect 523684 398828 523736 398880
rect 580172 398828 580224 398880
rect 3884 387744 3936 387796
rect 59360 387744 59412 387796
rect 523132 382236 523184 382288
rect 580172 382236 580224 382288
rect 3424 373940 3476 373992
rect 59360 373940 59412 373992
rect 523316 367072 523368 367124
rect 580172 367072 580224 367124
rect 3424 360136 3476 360188
rect 59360 360136 59412 360188
rect 524328 352520 524380 352572
rect 580172 352520 580224 352572
rect 3424 343544 3476 343596
rect 59360 343544 59412 343596
rect 523408 336676 523460 336728
rect 580172 336676 580224 336728
rect 3332 327020 3384 327072
rect 59360 327020 59412 327072
rect 523132 321512 523184 321564
rect 580172 321512 580224 321564
rect 3424 310428 3476 310480
rect 60004 310428 60056 310480
rect 523684 306280 523736 306332
rect 580172 306280 580224 306332
rect 3148 293904 3200 293956
rect 60004 293904 60056 293956
rect 523684 289756 523736 289808
rect 580172 289756 580224 289808
rect 3424 277312 3476 277364
rect 60004 277312 60056 277364
rect 523684 274592 523736 274644
rect 580172 274592 580224 274644
rect 3424 260788 3476 260840
rect 60004 260788 60056 260840
rect 523684 259360 523736 259412
rect 580172 259360 580224 259412
rect 3424 244196 3476 244248
rect 60004 244196 60056 244248
rect 523776 242836 523828 242888
rect 580172 242836 580224 242888
rect 523684 227672 523736 227724
rect 580172 227672 580224 227724
rect 3424 226244 3476 226296
rect 60096 226244 60148 226296
rect 523776 212440 523828 212492
rect 580172 212440 580224 212492
rect 3424 209720 3476 209772
rect 60004 209720 60056 209772
rect 523684 195916 523736 195968
rect 580172 195916 580224 195968
rect 3516 193128 3568 193180
rect 60096 193128 60148 193180
rect 523776 180752 523828 180804
rect 580172 180752 580224 180804
rect 3424 176604 3476 176656
rect 60004 176604 60056 176656
rect 523684 165520 523736 165572
rect 580172 165520 580224 165572
rect 3148 160012 3200 160064
rect 60188 160012 60240 160064
rect 523868 148996 523920 149048
rect 580172 148996 580224 149048
rect 3240 143488 3292 143540
rect 60096 143488 60148 143540
rect 523776 133832 523828 133884
rect 580172 133832 580224 133884
rect 3240 126896 3292 126948
rect 60004 126896 60056 126948
rect 523684 118600 523736 118652
rect 580172 118600 580224 118652
rect 3424 108944 3476 108996
rect 60188 108944 60240 108996
rect 523868 102076 523920 102128
rect 580172 102076 580224 102128
rect 3332 92420 3384 92472
rect 60096 92420 60148 92472
rect 523776 86912 523828 86964
rect 580172 86912 580224 86964
rect 3424 75828 3476 75880
rect 60004 75828 60056 75880
rect 523684 71680 523736 71732
rect 580172 71680 580224 71732
rect 3056 59304 3108 59356
rect 60280 59304 60332 59356
rect 523960 55156 524012 55208
rect 580172 55156 580224 55208
rect 147772 51008 147824 51060
rect 148048 51008 148100 51060
rect 209044 49648 209096 49700
rect 209872 49648 209924 49700
rect 232504 49648 232556 49700
rect 242716 49648 242768 49700
rect 245568 49648 245620 49700
rect 254860 49648 254912 49700
rect 262128 49648 262180 49700
rect 268016 49648 268068 49700
rect 275928 49648 275980 49700
rect 279332 49648 279384 49700
rect 324320 49648 324372 49700
rect 326344 49648 326396 49700
rect 450176 49648 450228 49700
rect 451924 49648 451976 49700
rect 241428 49580 241480 49632
rect 252100 49580 252152 49632
rect 257344 49580 257396 49632
rect 262404 49580 262456 49632
rect 263416 49580 263468 49632
rect 269948 49580 270000 49632
rect 274548 49580 274600 49632
rect 278320 49580 278372 49632
rect 392860 49580 392912 49632
rect 393964 49580 394016 49632
rect 237196 49512 237248 49564
rect 248052 49512 248104 49564
rect 248328 49512 248380 49564
rect 257712 49512 257764 49564
rect 219348 49444 219400 49496
rect 234252 49444 234304 49496
rect 238668 49444 238720 49496
rect 250168 49444 250220 49496
rect 255228 49444 255280 49496
rect 263324 49444 263376 49496
rect 220728 49376 220780 49428
rect 236092 49376 236144 49428
rect 237288 49376 237340 49428
rect 249248 49376 249300 49428
rect 249708 49376 249760 49428
rect 258632 49376 258684 49428
rect 64788 49308 64840 49360
rect 113180 49308 113232 49360
rect 186228 49308 186280 49360
rect 208860 49308 208912 49360
rect 217968 49308 218020 49360
rect 233332 49308 233384 49360
rect 234528 49308 234580 49360
rect 246488 49308 246540 49360
rect 251088 49308 251140 49360
rect 259552 49308 259604 49360
rect 419172 49308 419224 49360
rect 422944 49308 422996 49360
rect 465172 49308 465224 49360
rect 510712 49308 510764 49360
rect 57888 49240 57940 49292
rect 107476 49240 107528 49292
rect 122748 49240 122800 49292
rect 158168 49240 158220 49292
rect 179328 49240 179380 49292
rect 203248 49240 203300 49292
rect 215208 49240 215260 49292
rect 231400 49240 231452 49292
rect 233148 49240 233200 49292
rect 245476 49240 245528 49292
rect 246948 49240 247000 49292
rect 256792 49240 256844 49292
rect 266268 49240 266320 49292
rect 271788 49240 271840 49292
rect 476488 49240 476540 49292
rect 524420 49240 524472 49292
rect 50988 49172 51040 49224
rect 101864 49172 101916 49224
rect 115848 49172 115900 49224
rect 152556 49172 152608 49224
rect 172428 49172 172480 49224
rect 197636 49172 197688 49224
rect 208308 49172 208360 49224
rect 225788 49172 225840 49224
rect 229008 49172 229060 49224
rect 241704 49172 241756 49224
rect 242808 49172 242860 49224
rect 253020 49172 253072 49224
rect 253848 49172 253900 49224
rect 261484 49172 261536 49224
rect 482100 49172 482152 49224
rect 531320 49172 531372 49224
rect 13084 49104 13136 49156
rect 69940 49104 69992 49156
rect 107568 49104 107620 49156
rect 146944 49104 146996 49156
rect 160008 49104 160060 49156
rect 188252 49104 188304 49156
rect 206928 49104 206980 49156
rect 224868 49104 224920 49156
rect 226248 49104 226300 49156
rect 239864 49104 239916 49156
rect 244188 49104 244240 49156
rect 253940 49104 253992 49156
rect 257988 49104 258040 49156
rect 265256 49104 265308 49156
rect 267648 49104 267700 49156
rect 272708 49104 272760 49156
rect 277308 49104 277360 49156
rect 280252 49104 280304 49156
rect 426716 49104 426768 49156
rect 438124 49104 438176 49156
rect 487712 49104 487764 49156
rect 538220 49104 538272 49156
rect 8944 49036 8996 49088
rect 66168 49036 66220 49088
rect 103428 49036 103480 49088
rect 143172 49036 143224 49088
rect 158628 49036 158680 49088
rect 186320 49036 186372 49088
rect 213828 49036 213880 49088
rect 230480 49036 230532 49088
rect 231768 49036 231820 49088
rect 244556 49036 244608 49088
rect 245568 49036 245620 49088
rect 255872 49036 255924 49088
rect 256608 49036 256660 49088
rect 264244 49036 264296 49088
rect 264888 49036 264940 49088
rect 270868 49036 270920 49088
rect 273168 49036 273220 49088
rect 277400 49036 277452 49088
rect 391020 49036 391072 49088
rect 416872 49036 416924 49088
rect 435180 49036 435232 49088
rect 457444 49036 457496 49088
rect 493324 49036 493376 49088
rect 546500 49036 546552 49088
rect 17224 48968 17276 49020
rect 74632 48968 74684 49020
rect 79968 48968 80020 49020
rect 124404 48968 124456 49020
rect 125508 48968 125560 49020
rect 160100 48968 160152 49020
rect 165528 48968 165580 49020
rect 192024 48968 192076 49020
rect 202788 48968 202840 49020
rect 222016 48968 222068 49020
rect 222108 48968 222160 49020
rect 237012 48968 237064 49020
rect 240048 48968 240100 49020
rect 251180 48968 251232 49020
rect 252468 48968 252520 49020
rect 260564 48968 260616 49020
rect 350632 48968 350684 49020
rect 365812 48968 365864 49020
rect 373172 48968 373224 49020
rect 391204 48968 391256 49020
rect 406016 48968 406068 49020
rect 434720 48968 434772 49020
rect 454868 48968 454920 49020
rect 482284 48968 482336 49020
rect 498936 48968 498988 49020
rect 553400 48968 553452 49020
rect 271788 48832 271840 48884
rect 276480 48832 276532 48884
rect 79324 48764 79376 48816
rect 80244 48764 80296 48816
rect 92480 48764 92532 48816
rect 93124 48764 93176 48816
rect 95240 48764 95292 48816
rect 95884 48764 95936 48816
rect 103520 48764 103572 48816
rect 104348 48764 104400 48816
rect 108304 48764 108356 48816
rect 109408 48764 109460 48816
rect 139400 48764 139452 48816
rect 140044 48764 140096 48816
rect 144920 48764 144972 48816
rect 145748 48764 145800 48816
rect 146944 48764 146996 48816
rect 147864 48764 147916 48816
rect 162124 48764 162176 48816
rect 162860 48764 162912 48816
rect 179420 48764 179472 48816
rect 180340 48764 180392 48816
rect 212540 48764 212592 48816
rect 213276 48764 213328 48816
rect 215300 48764 215352 48816
rect 216036 48764 216088 48816
rect 226340 48764 226392 48816
rect 227260 48764 227312 48816
rect 259368 48764 259420 48816
rect 266176 48764 266228 48816
rect 272524 48764 272576 48816
rect 275560 48764 275612 48816
rect 281448 48764 281500 48816
rect 284024 48764 284076 48816
rect 296628 48764 296680 48816
rect 296904 48764 296956 48816
rect 299940 48764 299992 48816
rect 301044 48764 301096 48816
rect 309324 48764 309376 48816
rect 310428 48764 310480 48816
rect 311256 48764 311308 48816
rect 312544 48764 312596 48816
rect 314016 48764 314068 48816
rect 315304 48764 315356 48816
rect 317788 48764 317840 48816
rect 320824 48764 320876 48816
rect 321560 48764 321612 48816
rect 322756 48764 322808 48816
rect 326252 48764 326304 48816
rect 326988 48764 327040 48816
rect 327172 48764 327224 48816
rect 328368 48764 328420 48816
rect 329012 48764 329064 48816
rect 329748 48764 329800 48816
rect 330024 48764 330076 48816
rect 331128 48764 331180 48816
rect 332784 48764 332836 48816
rect 333888 48764 333940 48816
rect 335636 48764 335688 48816
rect 336648 48764 336700 48816
rect 338488 48764 338540 48816
rect 339408 48764 339460 48816
rect 341248 48764 341300 48816
rect 342168 48764 342220 48816
rect 344100 48764 344152 48816
rect 344928 48764 344980 48816
rect 345020 48764 345072 48816
rect 346216 48764 346268 48816
rect 347872 48764 347924 48816
rect 348976 48764 349028 48816
rect 353484 48764 353536 48816
rect 354496 48764 354548 48816
rect 356244 48764 356296 48816
rect 357256 48764 357308 48816
rect 359096 48764 359148 48816
rect 360016 48764 360068 48816
rect 361948 48764 362000 48816
rect 362776 48764 362828 48816
rect 367560 48764 367612 48816
rect 368388 48764 368440 48816
rect 368480 48764 368532 48816
rect 369676 48764 369728 48816
rect 370320 48764 370372 48816
rect 371148 48764 371200 48816
rect 371332 48764 371384 48816
rect 372436 48764 372488 48816
rect 374092 48764 374144 48816
rect 375288 48764 375340 48816
rect 376944 48764 376996 48816
rect 378048 48764 378100 48816
rect 379704 48764 379756 48816
rect 380808 48764 380860 48816
rect 382556 48764 382608 48816
rect 383476 48764 383528 48816
rect 385408 48764 385460 48816
rect 386236 48764 386288 48816
rect 388168 48764 388220 48816
rect 389088 48764 389140 48816
rect 389180 48764 389232 48816
rect 390468 48764 390520 48816
rect 391940 48764 391992 48816
rect 393228 48764 393280 48816
rect 394792 48764 394844 48816
rect 395988 48764 396040 48816
rect 397552 48764 397604 48816
rect 398748 48764 398800 48816
rect 400404 48764 400456 48816
rect 401508 48764 401560 48816
rect 403256 48764 403308 48816
rect 404268 48764 404320 48816
rect 408868 48764 408920 48816
rect 409788 48764 409840 48816
rect 411628 48764 411680 48816
rect 412548 48764 412600 48816
rect 412640 48764 412692 48816
rect 413928 48764 413980 48816
rect 414480 48764 414532 48816
rect 415308 48764 415360 48816
rect 415400 48764 415452 48816
rect 416688 48764 416740 48816
rect 420092 48764 420144 48816
rect 420828 48764 420880 48816
rect 421012 48764 421064 48816
rect 422208 48764 422260 48816
rect 423864 48764 423916 48816
rect 424876 48764 424928 48816
rect 432328 48764 432380 48816
rect 433984 48764 434036 48816
rect 436100 48764 436152 48816
rect 437296 48764 437348 48816
rect 437940 48764 437992 48816
rect 438768 48764 438820 48816
rect 438860 48764 438912 48816
rect 440148 48764 440200 48816
rect 441712 48764 441764 48816
rect 442816 48764 442868 48816
rect 444564 48764 444616 48816
rect 445576 48764 445628 48816
rect 452936 48764 452988 48816
rect 453856 48764 453908 48816
rect 458640 48764 458692 48816
rect 459468 48764 459520 48816
rect 459560 48764 459612 48816
rect 460848 48764 460900 48816
rect 462320 48764 462372 48816
rect 463608 48764 463660 48816
rect 464252 48764 464304 48816
rect 464988 48764 465040 48816
rect 467012 48764 467064 48816
rect 467748 48764 467800 48816
rect 468024 48764 468076 48816
rect 469128 48764 469180 48816
rect 470784 48764 470836 48816
rect 471888 48764 471940 48816
rect 473636 48764 473688 48816
rect 474648 48764 474700 48816
rect 479248 48764 479300 48816
rect 480168 48764 480220 48816
rect 483020 48764 483072 48816
rect 484308 48764 484360 48816
rect 484860 48764 484912 48816
rect 485688 48764 485740 48816
rect 506480 48764 506532 48816
rect 507676 48764 507728 48816
rect 511172 48764 511224 48816
rect 511908 48764 511960 48816
rect 514944 48764 514996 48816
rect 516048 48764 516100 48816
rect 517704 48764 517756 48816
rect 518808 48764 518860 48816
rect 520556 48764 520608 48816
rect 521476 48764 521528 48816
rect 204904 48696 204956 48748
rect 207020 48696 207072 48748
rect 269028 48696 269080 48748
rect 273628 48696 273680 48748
rect 280068 48696 280120 48748
rect 282092 48696 282144 48748
rect 312176 48696 312228 48748
rect 313188 48696 313240 48748
rect 314936 48696 314988 48748
rect 315948 48696 316000 48748
rect 378784 48696 378836 48748
rect 381544 48696 381596 48748
rect 390100 48696 390152 48748
rect 391296 48696 391348 48748
rect 401324 48696 401376 48748
rect 402244 48696 402296 48748
rect 407948 48696 408000 48748
rect 410524 48696 410576 48748
rect 443552 48696 443604 48748
rect 446404 48696 446456 48748
rect 461400 48696 461452 48748
rect 464344 48696 464396 48748
rect 468944 48696 468996 48748
rect 469864 48696 469916 48748
rect 472716 48696 472768 48748
rect 475384 48696 475436 48748
rect 306564 48628 306616 48680
rect 309324 48628 309376 48680
rect 396632 48628 396684 48680
rect 399484 48628 399536 48680
rect 509332 48628 509384 48680
rect 510436 48628 510488 48680
rect 512092 48628 512144 48680
rect 513196 48628 513248 48680
rect 270408 48560 270460 48612
rect 274640 48560 274692 48612
rect 279976 48560 280028 48612
rect 283012 48560 283064 48612
rect 320640 48560 320692 48612
rect 321468 48560 321520 48612
rect 323400 48560 323452 48612
rect 324228 48560 324280 48612
rect 263508 48492 263560 48544
rect 268936 48492 268988 48544
rect 346860 48492 346912 48544
rect 347688 48492 347740 48544
rect 364708 48492 364760 48544
rect 373264 48492 373316 48544
rect 418252 48492 418304 48544
rect 420184 48492 420236 48544
rect 485872 48492 485924 48544
rect 487068 48492 487120 48544
rect 491484 48492 491536 48544
rect 492588 48492 492640 48544
rect 303712 48424 303764 48476
rect 304908 48424 304960 48476
rect 417332 48424 417384 48476
rect 418068 48424 418120 48476
rect 261484 48356 261536 48408
rect 267096 48356 267148 48408
rect 429476 48356 429528 48408
rect 430488 48356 430540 48408
rect 61384 48288 61436 48340
rect 62488 48288 62540 48340
rect 111064 48288 111116 48340
rect 112168 48288 112220 48340
rect 120724 48288 120776 48340
rect 122564 48288 122616 48340
rect 126244 48288 126296 48340
rect 128176 48288 128228 48340
rect 167644 48288 167696 48340
rect 170404 48288 170456 48340
rect 284208 48288 284260 48340
rect 285864 48288 285916 48340
rect 286968 48288 287020 48340
rect 287704 48288 287756 48340
rect 289636 48288 289688 48340
rect 290924 48288 290976 48340
rect 291476 48288 291528 48340
rect 300860 48288 300912 48340
rect 302148 48288 302200 48340
rect 489000 48288 489052 48340
rect 489644 48288 489696 48340
rect 494244 48288 494296 48340
rect 495072 48288 495124 48340
rect 495164 48288 495216 48340
rect 496084 48288 496136 48340
rect 505560 48288 505612 48340
rect 506388 48288 506440 48340
rect 508320 48288 508372 48340
rect 509148 48288 509200 48340
rect 168748 48263 168800 48272
rect 168748 48229 168757 48263
rect 168757 48229 168791 48263
rect 168791 48229 168800 48263
rect 168748 48220 168800 48229
rect 288256 48220 288308 48272
rect 489644 48195 489696 48204
rect 489644 48161 489653 48195
rect 489653 48161 489687 48195
rect 489687 48161 489696 48195
rect 489644 48152 489696 48161
rect 10324 47540 10376 47592
rect 65248 47540 65300 47592
rect 70308 47540 70360 47592
rect 116860 47540 116912 47592
rect 155868 47540 155920 47592
rect 184480 47540 184532 47592
rect 447324 47540 447376 47592
rect 487160 47540 487212 47592
rect 497096 47540 497148 47592
rect 550640 47540 550692 47592
rect 176660 46860 176712 46912
rect 177580 46860 177632 46912
rect 293960 46903 294012 46912
rect 293960 46869 293969 46903
rect 293969 46869 294003 46903
rect 294003 46869 294012 46903
rect 293960 46860 294012 46869
rect 118792 46248 118844 46300
rect 119436 46248 119488 46300
rect 153200 46248 153252 46300
rect 154212 46248 154264 46300
rect 155960 46248 156012 46300
rect 156972 46248 157024 46300
rect 22008 46180 22060 46232
rect 77392 46180 77444 46232
rect 78036 46180 78088 46232
rect 88248 46180 88300 46232
rect 130936 46180 130988 46232
rect 132408 46180 132460 46232
rect 165712 46180 165764 46232
rect 173900 46180 173952 46232
rect 174820 46180 174872 46232
rect 455788 46180 455840 46232
rect 498200 46180 498252 46232
rect 499948 46180 500000 46232
rect 554780 46180 554832 46232
rect 78956 46112 79008 46164
rect 27528 44820 27580 44872
rect 82912 44820 82964 44872
rect 92388 44820 92440 44872
rect 133880 44820 133932 44872
rect 139308 44820 139360 44872
rect 171232 44820 171284 44872
rect 502708 44820 502760 44872
rect 557540 44820 557592 44872
rect 86500 43460 86552 43512
rect 34428 43392 34480 43444
rect 88432 43392 88484 43444
rect 129648 43392 129700 43444
rect 162952 43392 163004 43444
rect 509148 43392 509200 43444
rect 564440 43392 564492 43444
rect 3424 42712 3476 42764
rect 60188 42712 60240 42764
rect 42708 42032 42760 42084
rect 95332 42032 95384 42084
rect 106188 42032 106240 42084
rect 145012 42032 145064 42084
rect 201132 42032 201184 42084
rect 511908 42032 511960 42084
rect 568580 42032 568632 42084
rect 194784 41420 194836 41472
rect 195428 41420 195480 41472
rect 489736 41420 489788 41472
rect 62396 41352 62448 41404
rect 63132 41352 63184 41404
rect 124220 41352 124272 41404
rect 124404 41352 124456 41404
rect 296904 41352 296956 41404
rect 297088 41352 297140 41404
rect 489736 41284 489788 41336
rect 49608 40672 49660 40724
rect 100852 40672 100904 40724
rect 484216 40672 484268 40724
rect 534080 40672 534132 40724
rect 523868 39992 523920 40044
rect 580172 39992 580224 40044
rect 53748 39312 53800 39364
rect 103612 39312 103664 39364
rect 74724 38632 74776 38684
rect 74908 38632 74960 38684
rect 82820 38632 82872 38684
rect 83740 38632 83792 38684
rect 85764 38675 85816 38684
rect 85764 38641 85773 38675
rect 85773 38641 85807 38675
rect 85807 38641 85816 38675
rect 85764 38632 85816 38641
rect 132868 38632 132920 38684
rect 133420 38632 133472 38684
rect 168840 38632 168892 38684
rect 489828 38632 489880 38684
rect 109408 38607 109460 38616
rect 109408 38573 109417 38607
rect 109417 38573 109451 38607
rect 109451 38573 109460 38607
rect 109408 38564 109460 38573
rect 124404 38564 124456 38616
rect 197452 38607 197504 38616
rect 197452 38573 197461 38607
rect 197461 38573 197495 38607
rect 197495 38573 197504 38607
rect 197452 38564 197504 38573
rect 203248 38564 203300 38616
rect 291384 38607 291436 38616
rect 291384 38573 291393 38607
rect 291393 38573 291427 38607
rect 291427 38573 291436 38607
rect 291384 38564 291436 38573
rect 487160 38607 487212 38616
rect 487160 38573 487169 38607
rect 487169 38573 487203 38607
rect 487203 38573 487212 38607
rect 487160 38564 487212 38573
rect 56416 37884 56468 37936
rect 106372 37884 106424 37936
rect 486976 37884 487028 37936
rect 536840 37884 536892 37936
rect 293960 37315 294012 37324
rect 293960 37281 293969 37315
rect 293969 37281 294003 37315
rect 294003 37281 294012 37315
rect 293960 37272 294012 37281
rect 290832 37136 290884 37188
rect 14464 36524 14516 36576
rect 72056 36524 72108 36576
rect 288164 36524 288216 36576
rect 288348 36524 288400 36576
rect 492496 36524 492548 36576
rect 545120 36524 545172 36576
rect 98092 35912 98144 35964
rect 98276 35912 98328 35964
rect 19984 35164 20036 35216
rect 75920 35164 75972 35216
rect 498016 35164 498068 35216
rect 552020 35164 552072 35216
rect 28908 33736 28960 33788
rect 82820 33736 82872 33788
rect 433248 33736 433300 33788
rect 469220 33736 469272 33788
rect 507676 33736 507728 33788
rect 563152 33736 563204 33788
rect 31668 32376 31720 32428
rect 85764 32376 85816 32428
rect 96528 32376 96580 32428
rect 136732 32376 136784 32428
rect 430396 32376 430448 32428
rect 466460 32376 466512 32428
rect 489644 31696 489696 31748
rect 489828 31696 489880 31748
rect 495072 31696 495124 31748
rect 495256 31696 495308 31748
rect 197452 31603 197504 31612
rect 197452 31569 197461 31603
rect 197461 31569 197495 31603
rect 197495 31569 197504 31603
rect 197452 31560 197504 31569
rect 200488 31603 200540 31612
rect 200488 31569 200497 31603
rect 200497 31569 200531 31603
rect 200531 31569 200540 31603
rect 200488 31560 200540 31569
rect 35808 31016 35860 31068
rect 88340 31016 88392 31068
rect 89628 31016 89680 31068
rect 131120 31016 131172 31068
rect 427728 31016 427780 31068
rect 462320 31016 462372 31068
rect 478788 31016 478840 31068
rect 527180 31016 527232 31068
rect 85488 29656 85540 29708
rect 128360 29656 128412 29708
rect 38568 29588 38620 29640
rect 92572 29588 92624 29640
rect 422116 29588 422168 29640
rect 455420 29588 455472 29640
rect 489736 29588 489788 29640
rect 540980 29588 541032 29640
rect 109500 28976 109552 29028
rect 124312 29019 124364 29028
rect 124312 28985 124321 29019
rect 124321 28985 124355 29019
rect 124355 28985 124364 29019
rect 124312 28976 124364 28985
rect 203156 29019 203208 29028
rect 203156 28985 203165 29019
rect 203165 28985 203199 29019
rect 203199 28985 203208 29019
rect 203156 28976 203208 28985
rect 291476 28976 291528 29028
rect 296996 28976 297048 29028
rect 297088 28976 297140 29028
rect 487160 29019 487212 29028
rect 487160 28985 487169 29019
rect 487169 28985 487203 29019
rect 487203 28985 487212 29019
rect 487160 28976 487212 28985
rect 62304 28951 62356 28960
rect 62304 28917 62313 28951
rect 62313 28917 62347 28951
rect 62347 28917 62356 28951
rect 62304 28908 62356 28917
rect 438124 28951 438176 28960
rect 438124 28917 438133 28951
rect 438133 28917 438167 28951
rect 438167 28917 438176 28951
rect 438124 28908 438176 28917
rect 82728 28228 82780 28280
rect 125600 28228 125652 28280
rect 422944 28228 422996 28280
rect 451280 28228 451332 28280
rect 470508 28228 470560 28280
rect 516140 28228 516192 28280
rect 80152 27616 80204 27668
rect 80244 27616 80296 27668
rect 291016 27659 291068 27668
rect 291016 27625 291025 27659
rect 291025 27625 291059 27659
rect 291059 27625 291068 27659
rect 291016 27616 291068 27625
rect 293960 27591 294012 27600
rect 293960 27557 293969 27591
rect 293969 27557 294003 27591
rect 294003 27557 294012 27591
rect 293960 27548 294012 27557
rect 296996 27548 297048 27600
rect 297088 27548 297140 27600
rect 78588 26868 78640 26920
rect 122840 26868 122892 26920
rect 124128 26868 124180 26920
rect 158720 26868 158772 26920
rect 416596 26868 416648 26920
rect 448520 26868 448572 26920
rect 464344 26868 464396 26920
rect 505100 26868 505152 26920
rect 150808 26256 150860 26308
rect 150900 26256 150952 26308
rect 3424 26188 3476 26240
rect 60096 26188 60148 26240
rect 74448 25508 74500 25560
rect 120080 25508 120132 25560
rect 140688 25508 140740 25560
rect 171140 25508 171192 25560
rect 413836 25508 413888 25560
rect 444380 25508 444432 25560
rect 459468 25508 459520 25560
rect 502432 25508 502484 25560
rect 503628 25508 503680 25560
rect 558920 25508 558972 25560
rect 523776 24760 523828 24812
rect 580172 24760 580224 24812
rect 200304 24148 200356 24200
rect 200488 24148 200540 24200
rect 67548 24080 67600 24132
rect 114560 24080 114612 24132
rect 136548 24080 136600 24132
rect 168840 24080 168892 24132
rect 411168 24080 411220 24132
rect 441620 24080 441672 24132
rect 451924 24080 451976 24132
rect 491300 24080 491352 24132
rect 445576 22788 445628 22840
rect 484400 22788 484452 22840
rect 23388 22720 23440 22772
rect 79324 22720 79376 22772
rect 91008 22720 91060 22772
rect 132868 22720 132920 22772
rect 133788 22720 133840 22772
rect 165620 22720 165672 22772
rect 368388 22720 368440 22772
rect 386420 22720 386472 22772
rect 402888 22720 402940 22772
rect 430580 22720 430632 22772
rect 481548 22720 481600 22772
rect 529940 22720 529992 22772
rect 74724 22355 74776 22364
rect 74724 22321 74733 22355
rect 74733 22321 74767 22355
rect 74767 22321 74776 22355
rect 74724 22312 74776 22321
rect 124312 22108 124364 22160
rect 150624 22108 150676 22160
rect 495256 22108 495308 22160
rect 202972 22040 203024 22092
rect 203156 22040 203208 22092
rect 291292 22040 291344 22092
rect 291476 22040 291528 22092
rect 124312 21972 124364 22024
rect 495256 21972 495308 22024
rect 146208 21428 146260 21480
rect 176752 21428 176804 21480
rect 438768 21428 438820 21480
rect 476120 21428 476172 21480
rect 60648 21360 60700 21412
rect 108304 21360 108356 21412
rect 108948 21360 109000 21412
rect 146944 21360 146996 21412
rect 410524 21360 410576 21412
rect 437480 21360 437532 21412
rect 476028 21360 476080 21412
rect 523040 21360 523092 21412
rect 64696 19932 64748 19984
rect 111064 19932 111116 19984
rect 142068 19932 142120 19984
rect 173992 19932 174044 19984
rect 405648 19932 405700 19984
rect 433340 19932 433392 19984
rect 433984 19932 434036 19984
rect 467932 19932 467984 19984
rect 475384 19932 475436 19984
rect 520372 19932 520424 19984
rect 62488 19320 62540 19372
rect 74724 19363 74776 19372
rect 74724 19329 74733 19363
rect 74733 19329 74767 19363
rect 74767 19329 74776 19363
rect 74724 19320 74776 19329
rect 109316 19320 109368 19372
rect 109408 19320 109460 19372
rect 438308 19320 438360 19372
rect 147864 19252 147916 19304
rect 203156 19295 203208 19304
rect 203156 19261 203165 19295
rect 203165 19261 203199 19295
rect 203199 19261 203208 19295
rect 203156 19252 203208 19261
rect 487160 19295 487212 19304
rect 487160 19261 487169 19295
rect 487169 19261 487203 19295
rect 487203 19261 487212 19295
rect 487160 19252 487212 19261
rect 430488 18640 430540 18692
rect 465080 18640 465132 18692
rect 10416 18572 10468 18624
rect 69112 18572 69164 18624
rect 71688 18572 71740 18624
rect 117320 18572 117372 18624
rect 135168 18572 135220 18624
rect 168380 18572 168432 18624
rect 290648 18572 290700 18624
rect 291108 18572 291160 18624
rect 400128 18572 400180 18624
rect 426440 18572 426492 18624
rect 464988 18572 465040 18624
rect 509240 18572 509292 18624
rect 293960 18003 294012 18012
rect 293960 17969 293969 18003
rect 293969 17969 294003 18003
rect 294003 17969 294012 18003
rect 293960 17960 294012 17969
rect 424876 17280 424928 17332
rect 458180 17280 458232 17332
rect 45468 17212 45520 17264
rect 96620 17212 96672 17264
rect 128268 17212 128320 17264
rect 162124 17212 162176 17264
rect 164148 17212 164200 17264
rect 190460 17212 190512 17264
rect 399484 17212 399536 17264
rect 423680 17212 423732 17264
rect 453856 17212 453908 17264
rect 494060 17212 494112 17264
rect 496084 17212 496136 17264
rect 547880 17212 547932 17264
rect 98092 16600 98144 16652
rect 98276 16600 98328 16652
rect 41328 15852 41380 15904
rect 93860 15852 93912 15904
rect 102048 15852 102100 15904
rect 142252 15852 142304 15904
rect 159916 15852 159968 15904
rect 186412 15852 186464 15904
rect 394608 15852 394660 15904
rect 419540 15852 419592 15904
rect 420184 15852 420236 15904
rect 451372 15852 451424 15904
rect 469864 15852 469916 15904
rect 514760 15852 514812 15904
rect 404176 14492 404228 14544
rect 433432 14492 433484 14544
rect 38476 14424 38528 14476
rect 91100 14424 91152 14476
rect 99288 14424 99340 14476
rect 139492 14424 139544 14476
rect 151728 14424 151780 14476
rect 180800 14424 180852 14476
rect 424968 14424 425020 14476
rect 459652 14424 459704 14476
rect 463516 14424 463568 14476
rect 507860 14424 507912 14476
rect 510436 14424 510488 14476
rect 565820 14424 565872 14476
rect 395896 13132 395948 13184
rect 422300 13132 422352 13184
rect 460756 13132 460808 13184
rect 503720 13132 503772 13184
rect 30288 13064 30340 13116
rect 85580 13064 85632 13116
rect 95148 13064 95200 13116
rect 136640 13064 136692 13116
rect 148968 13064 149020 13116
rect 178040 13064 178092 13116
rect 187608 13064 187660 13116
rect 209044 13064 209096 13116
rect 422208 13064 422260 13116
rect 454040 13064 454092 13116
rect 500868 13064 500920 13116
rect 554872 13064 554924 13116
rect 80060 12384 80112 12436
rect 80428 12384 80480 12436
rect 300952 12248 301004 12300
rect 301412 12248 301464 12300
rect 513196 11976 513248 12028
rect 513288 11772 513340 11824
rect 9036 11704 9088 11756
rect 67640 11704 67692 11756
rect 84108 11704 84160 11756
rect 126244 11704 126296 11756
rect 144828 11704 144880 11756
rect 175280 11704 175332 11756
rect 180708 11704 180760 11756
rect 387708 11704 387760 11756
rect 411260 11704 411312 11756
rect 413928 11704 413980 11756
rect 443092 11704 443144 11756
rect 458088 11704 458140 11756
rect 500960 11704 501012 11756
rect 517428 11704 517480 11756
rect 574744 11704 574796 11756
rect 4068 10276 4120 10328
rect 63500 10276 63552 10328
rect 80244 10276 80296 10328
rect 124404 10276 124456 10328
rect 141976 10276 142028 10328
rect 172520 10276 172572 10328
rect 176568 10276 176620 10328
rect 200396 10276 200448 10328
rect 384948 10276 385000 10328
rect 408592 10276 408644 10328
rect 409696 10276 409748 10328
rect 440240 10276 440292 10328
rect 452568 10276 452620 10328
rect 494152 10276 494204 10328
rect 520188 10276 520240 10328
rect 579620 10276 579672 10328
rect 147772 9707 147824 9716
rect 147772 9673 147781 9707
rect 147781 9673 147815 9707
rect 147815 9673 147824 9707
rect 147772 9664 147824 9673
rect 150808 9707 150860 9716
rect 150808 9673 150817 9707
rect 150817 9673 150851 9707
rect 150851 9673 150860 9707
rect 150808 9664 150860 9673
rect 487160 9707 487212 9716
rect 487160 9673 487169 9707
rect 487169 9673 487203 9707
rect 487203 9673 487212 9707
rect 487160 9664 487212 9673
rect 3424 9596 3476 9648
rect 60004 9596 60056 9648
rect 119436 8984 119488 9036
rect 156052 8984 156104 9036
rect 449808 8984 449860 9036
rect 490564 8984 490616 9036
rect 76656 8916 76708 8968
rect 120724 8916 120776 8968
rect 137284 8916 137336 8968
rect 167644 8916 167696 8968
rect 172980 8916 173032 8968
rect 197452 8916 197504 8968
rect 371148 8916 371200 8968
rect 390652 8916 390704 8968
rect 391296 8916 391348 8968
rect 415676 8916 415728 8968
rect 416688 8916 416740 8968
rect 447784 8916 447836 8968
rect 467748 8916 467800 8968
rect 513196 8916 513248 8968
rect 514668 8916 514720 8968
rect 572628 8916 572680 8968
rect 523684 8236 523736 8288
rect 580172 8236 580224 8288
rect 133696 7624 133748 7676
rect 167000 7624 167052 7676
rect 382188 7624 382240 7676
rect 404912 7624 404964 7676
rect 447048 7624 447100 7676
rect 486976 7624 487028 7676
rect 494060 7624 494112 7676
rect 495348 7624 495400 7676
rect 1676 7556 1728 7608
rect 62488 7556 62540 7608
rect 65984 7556 66036 7608
rect 113272 7556 113324 7608
rect 115940 7556 115992 7608
rect 153292 7556 153344 7608
rect 169392 7556 169444 7608
rect 194692 7556 194744 7608
rect 362776 7556 362828 7608
rect 379980 7556 380032 7608
rect 402244 7556 402296 7608
rect 429936 7556 429988 7608
rect 466368 7556 466420 7608
rect 512000 7556 512052 7608
rect 130200 6196 130252 6248
rect 164240 6196 164292 6248
rect 446404 6196 446456 6248
rect 483480 6196 483532 6248
rect 572 6128 624 6180
rect 61384 6128 61436 6180
rect 62396 6128 62448 6180
rect 110420 6128 110472 6180
rect 112352 6128 112404 6180
rect 150532 6128 150584 6180
rect 165896 6128 165948 6180
rect 191932 6128 191984 6180
rect 360016 6128 360068 6180
rect 376392 6128 376444 6180
rect 376668 6128 376720 6180
rect 397828 6128 397880 6180
rect 398656 6128 398708 6180
rect 426256 6128 426308 6180
rect 441528 6128 441580 6180
rect 479892 6128 479944 6180
rect 482284 6128 482336 6180
rect 497740 6128 497792 6180
rect 506388 6128 506440 6180
rect 561956 6128 562008 6180
rect 471796 5312 471848 5364
rect 519084 5312 519136 5364
rect 474556 5244 474608 5296
rect 522672 5244 522724 5296
rect 484308 5176 484360 5228
rect 533436 5176 533488 5228
rect 55220 5108 55272 5160
rect 104900 5108 104952 5160
rect 477408 5108 477460 5160
rect 526260 5108 526312 5160
rect 58808 5040 58860 5092
rect 107660 5040 107712 5092
rect 480076 5040 480128 5092
rect 529848 5040 529900 5092
rect 51632 4972 51684 5024
rect 102140 4972 102192 5024
rect 489644 4972 489696 5024
rect 540520 5108 540572 5160
rect 48136 4904 48188 4956
rect 99380 4904 99432 4956
rect 279884 4904 279936 4956
rect 280068 4904 280120 4956
rect 487068 4904 487120 4956
rect 536932 4904 536984 4956
rect 17316 4836 17368 4888
rect 74724 4836 74776 4888
rect 183744 4836 183796 4888
rect 204904 4836 204956 4888
rect 373264 4836 373316 4888
rect 383384 4836 383436 4888
rect 393964 4836 394016 4888
rect 419172 4836 419224 4888
rect 457444 4836 457496 4888
rect 12440 4768 12492 4820
rect 71780 4768 71832 4820
rect 73068 4768 73120 4820
rect 118792 4768 118844 4820
rect 126612 4768 126664 4820
rect 161480 4768 161532 4820
rect 162308 4768 162360 4820
rect 189172 4768 189224 4820
rect 357256 4768 357308 4820
rect 372804 4768 372856 4820
rect 381544 4768 381596 4820
rect 401324 4768 401376 4820
rect 407028 4768 407080 4820
rect 437020 4768 437072 4820
rect 438308 4768 438360 4820
rect 462044 4768 462096 4820
rect 492588 4836 492640 4888
rect 544108 4836 544160 4888
rect 472716 4768 472768 4820
rect 495164 4768 495216 4820
rect 547696 4768 547748 4820
rect 391204 4632 391256 4684
rect 394240 4632 394292 4684
rect 296720 4360 296772 4412
rect 297088 4360 297140 4412
rect 45744 4088 45796 4140
rect 98000 4088 98052 4140
rect 106372 4088 106424 4140
rect 144920 4088 144972 4140
rect 155132 4088 155184 4140
rect 155868 4088 155920 4140
rect 158720 4088 158772 4140
rect 159916 4088 159968 4140
rect 163504 4088 163556 4140
rect 164148 4088 164200 4140
rect 170588 4088 170640 4140
rect 195980 4088 196032 4140
rect 207112 4088 207164 4140
rect 278872 4088 278924 4140
rect 279884 4088 279936 4140
rect 287152 4088 287204 4140
rect 288348 4088 288400 4140
rect 289544 4088 289596 4140
rect 289912 4088 289964 4140
rect 291476 4088 291528 4140
rect 291936 4088 291988 4140
rect 292580 4088 292632 4140
rect 293132 4088 293184 4140
rect 296812 4088 296864 4140
rect 297916 4088 297968 4140
rect 298100 4088 298152 4140
rect 299112 4088 299164 4140
rect 299388 4088 299440 4140
rect 300308 4088 300360 4140
rect 306288 4088 306340 4140
rect 308588 4088 308640 4140
rect 338028 4088 338080 4140
rect 348884 4088 348936 4140
rect 350448 4088 350500 4140
rect 364524 4088 364576 4140
rect 367008 4088 367060 4140
rect 385868 4088 385920 4140
rect 386236 4088 386288 4140
rect 409696 4088 409748 4140
rect 442816 4088 442868 4140
rect 481088 4088 481140 4140
rect 496728 4088 496780 4140
rect 550088 4088 550140 4140
rect 43352 4020 43404 4072
rect 36176 3952 36228 4004
rect 89720 3952 89772 4004
rect 39764 3884 39816 3936
rect 92480 3884 92532 3936
rect 32680 3816 32732 3868
rect 5264 3748 5316 3800
rect 8944 3748 8996 3800
rect 29092 3748 29144 3800
rect 84200 3748 84252 3800
rect 84936 3816 84988 3868
rect 85488 3816 85540 3868
rect 88524 3816 88576 3868
rect 89628 3816 89680 3868
rect 109960 4020 110012 4072
rect 147772 4020 147824 4072
rect 167092 4020 167144 4072
rect 193220 4020 193272 4072
rect 196808 4020 196860 4072
rect 216680 4020 216732 4072
rect 218244 4020 218296 4072
rect 219348 4020 219400 4072
rect 304816 4020 304868 4072
rect 307392 4020 307444 4072
rect 331128 4020 331180 4072
rect 339500 4020 339552 4072
rect 342168 4020 342220 4072
rect 353760 4020 353812 4072
rect 354588 4020 354640 4072
rect 370412 4020 370464 4072
rect 372528 4020 372580 4072
rect 393044 4020 393096 4072
rect 393228 4020 393280 4072
rect 417976 4020 418028 4072
rect 440056 4020 440108 4072
rect 478696 4020 478748 4072
rect 502248 4020 502300 4072
rect 557172 4020 557224 4072
rect 111156 3952 111208 4004
rect 149060 3952 149112 4004
rect 156328 3952 156380 4004
rect 184940 3952 184992 4004
rect 195612 3952 195664 4004
rect 215300 3952 215352 4004
rect 103980 3884 104032 3936
rect 95240 3816 95292 3868
rect 99196 3816 99248 3868
rect 139400 3816 139452 3868
rect 86960 3748 87012 3800
rect 96896 3748 96948 3800
rect 138020 3748 138072 3800
rect 24308 3680 24360 3732
rect 80152 3680 80204 3732
rect 98276 3680 98328 3732
rect 100484 3680 100536 3732
rect 140780 3680 140832 3732
rect 2872 3476 2924 3528
rect 4068 3476 4120 3528
rect 10324 3612 10376 3664
rect 20720 3612 20772 3664
rect 11244 3544 11296 3596
rect 4068 3340 4120 3392
rect 7656 3476 7708 3528
rect 9036 3476 9088 3528
rect 13636 3476 13688 3528
rect 14464 3476 14516 3528
rect 14832 3544 14884 3596
rect 63592 3544 63644 3596
rect 64696 3544 64748 3596
rect 70492 3544 70544 3596
rect 70676 3612 70728 3664
rect 71688 3612 71740 3664
rect 77392 3612 77444 3664
rect 77852 3612 77904 3664
rect 78588 3612 78640 3664
rect 93308 3612 93360 3664
rect 135260 3612 135312 3664
rect 150440 3884 150492 3936
rect 179420 3884 179472 3936
rect 192024 3884 192076 3936
rect 212540 3884 212592 3936
rect 218152 3884 218204 3936
rect 227720 3952 227772 4004
rect 240140 3952 240192 4004
rect 284760 3952 284812 4004
rect 285772 3952 285824 4004
rect 320088 3952 320140 4004
rect 326436 3952 326488 4004
rect 332508 3952 332560 4004
rect 341892 3952 341944 4004
rect 346308 3952 346360 4004
rect 359740 3952 359792 4004
rect 361488 3952 361540 4004
rect 378784 3952 378836 4004
rect 383476 3952 383528 4004
rect 406108 3952 406160 4004
rect 409788 3952 409840 4004
rect 439412 3952 439464 4004
rect 448336 3952 448388 4004
rect 489368 3952 489420 4004
rect 505008 3952 505060 4004
rect 560760 3952 560812 4004
rect 220912 3884 220964 3936
rect 224132 3884 224184 3936
rect 238852 3884 238904 3936
rect 335268 3884 335320 3936
rect 345480 3884 345532 3936
rect 347688 3884 347740 3936
rect 360936 3884 360988 3936
rect 364248 3884 364300 3936
rect 382372 3884 382424 3936
rect 386328 3884 386380 3936
rect 410892 3884 410944 3936
rect 412548 3884 412600 3936
rect 443000 3884 443052 3936
rect 445668 3884 445720 3936
rect 485780 3884 485832 3936
rect 491208 3884 491260 3936
rect 507768 3884 507820 3936
rect 564348 3884 564400 3936
rect 153936 3816 153988 3868
rect 183560 3816 183612 3868
rect 188436 3816 188488 3868
rect 209964 3816 210016 3868
rect 154672 3748 154724 3800
rect 182180 3748 182232 3800
rect 182548 3748 182600 3800
rect 205640 3748 205692 3800
rect 215852 3816 215904 3868
rect 231860 3816 231912 3868
rect 328368 3816 328420 3868
rect 335912 3816 335964 3868
rect 336648 3816 336700 3868
rect 346676 3816 346728 3868
rect 349068 3816 349120 3868
rect 363328 3816 363380 3868
rect 365628 3816 365680 3868
rect 384672 3816 384724 3868
rect 389088 3816 389140 3868
rect 413284 3816 413336 3868
rect 415308 3816 415360 3868
rect 446588 3816 446640 3868
rect 451188 3816 451240 3868
rect 492956 3816 493008 3868
rect 510528 3816 510580 3868
rect 567844 3816 567896 3868
rect 211068 3748 211120 3800
rect 146852 3680 146904 3732
rect 176660 3680 176712 3732
rect 184848 3680 184900 3732
rect 203892 3680 203944 3732
rect 143540 3612 143592 3664
rect 75460 3544 75512 3596
rect 69480 3476 69532 3528
rect 70308 3476 70360 3528
rect 89720 3544 89772 3596
rect 121828 3544 121880 3596
rect 122748 3544 122800 3596
rect 123024 3544 123076 3596
rect 124128 3544 124180 3596
rect 124220 3544 124272 3596
rect 125508 3544 125560 3596
rect 125416 3476 125468 3528
rect 127808 3476 127860 3528
rect 128268 3476 128320 3528
rect 129004 3476 129056 3528
rect 129648 3476 129700 3528
rect 131396 3544 131448 3596
rect 132408 3544 132460 3596
rect 132592 3544 132644 3596
rect 133788 3544 133840 3596
rect 136088 3544 136140 3596
rect 136548 3544 136600 3596
rect 139676 3544 139728 3596
rect 140688 3544 140740 3596
rect 140872 3544 140924 3596
rect 141976 3544 142028 3596
rect 143264 3544 143316 3596
rect 145656 3544 145708 3596
rect 146208 3544 146260 3596
rect 6460 3408 6512 3460
rect 60004 3408 60056 3460
rect 60648 3408 60700 3460
rect 68284 3408 68336 3460
rect 116124 3408 116176 3460
rect 118240 3408 118292 3460
rect 148048 3476 148100 3528
rect 148968 3476 149020 3528
rect 149244 3612 149296 3664
rect 173900 3612 173952 3664
rect 180156 3612 180208 3664
rect 180708 3612 180760 3664
rect 181352 3612 181404 3664
rect 204260 3612 204312 3664
rect 171784 3544 171836 3596
rect 172428 3544 172480 3596
rect 177764 3544 177816 3596
rect 201500 3544 201552 3596
rect 206284 3544 206336 3596
rect 206928 3544 206980 3596
rect 207480 3544 207532 3596
rect 208308 3544 208360 3596
rect 208676 3680 208728 3732
rect 226432 3748 226484 3800
rect 228916 3748 228968 3800
rect 232504 3748 232556 3800
rect 315304 3748 315356 3800
rect 319260 3748 319312 3800
rect 339408 3748 339460 3800
rect 350264 3748 350316 3800
rect 351828 3748 351880 3800
rect 366916 3748 366968 3800
rect 369676 3748 369728 3800
rect 388260 3748 388312 3800
rect 390468 3748 390520 3800
rect 414480 3748 414532 3800
rect 423588 3748 423640 3800
rect 457260 3748 457312 3800
rect 460848 3748 460900 3800
rect 503628 3748 503680 3800
rect 516048 3748 516100 3800
rect 573824 3748 573876 3800
rect 223764 3680 223816 3732
rect 226524 3680 226576 3732
rect 237380 3680 237432 3732
rect 313096 3680 313148 3732
rect 318064 3680 318116 3732
rect 325608 3680 325660 3732
rect 333612 3680 333664 3732
rect 333796 3680 333848 3732
rect 344284 3680 344336 3732
rect 348976 3680 349028 3732
rect 362132 3680 362184 3732
rect 362868 3680 362920 3732
rect 381176 3680 381228 3732
rect 383568 3680 383620 3732
rect 407304 3680 407356 3732
rect 418068 3680 418120 3732
rect 450176 3680 450228 3732
rect 451280 3680 451332 3732
rect 452476 3680 452528 3732
rect 453948 3680 454000 3732
rect 496544 3680 496596 3732
rect 513288 3680 513340 3732
rect 570236 3680 570288 3732
rect 222936 3612 222988 3664
rect 222200 3544 222252 3596
rect 225328 3544 225380 3596
rect 226248 3544 226300 3596
rect 160284 3476 160336 3528
rect 168196 3476 168248 3528
rect 194600 3476 194652 3528
rect 198004 3476 198056 3528
rect 214656 3476 214708 3528
rect 215208 3476 215260 3528
rect 217048 3476 217100 3528
rect 217968 3476 218020 3528
rect 219348 3476 219400 3528
rect 234620 3544 234672 3596
rect 236000 3544 236052 3596
rect 237196 3544 237248 3596
rect 231308 3476 231360 3528
rect 231768 3476 231820 3528
rect 232504 3476 232556 3528
rect 233148 3476 233200 3528
rect 233700 3476 233752 3528
rect 234528 3476 234580 3528
rect 234804 3476 234856 3528
rect 247132 3612 247184 3664
rect 285956 3612 286008 3664
rect 286968 3612 287020 3664
rect 315948 3612 316000 3664
rect 320456 3612 320508 3664
rect 324228 3612 324280 3664
rect 331220 3612 331272 3664
rect 336556 3612 336608 3664
rect 347872 3612 347924 3664
rect 355968 3612 356020 3664
rect 371608 3612 371660 3664
rect 377956 3612 378008 3664
rect 400220 3612 400272 3664
rect 401508 3612 401560 3664
rect 428740 3612 428792 3664
rect 434628 3612 434680 3664
rect 471520 3612 471572 3664
rect 471888 3612 471940 3664
rect 517888 3612 517940 3664
rect 518808 3612 518860 3664
rect 577412 3612 577464 3664
rect 302056 3544 302108 3596
rect 303804 3544 303856 3596
rect 309048 3544 309100 3596
rect 312176 3544 312228 3596
rect 322756 3544 322808 3596
rect 328828 3544 328880 3596
rect 329748 3544 329800 3596
rect 338304 3544 338356 3596
rect 339316 3544 339368 3596
rect 351368 3544 351420 3596
rect 354496 3544 354548 3596
rect 369216 3544 369268 3596
rect 369768 3544 369820 3596
rect 389456 3544 389508 3596
rect 395988 3544 396040 3596
rect 421564 3544 421616 3596
rect 426348 3544 426400 3596
rect 460848 3544 460900 3596
rect 463608 3544 463660 3596
rect 469036 3544 469088 3596
rect 239588 3476 239640 3528
rect 240048 3476 240100 3528
rect 240784 3476 240836 3528
rect 241428 3476 241480 3528
rect 241980 3476 242032 3528
rect 242808 3476 242860 3528
rect 243176 3476 243228 3528
rect 244188 3476 244240 3528
rect 244372 3476 244424 3528
rect 245476 3476 245528 3528
rect 249156 3476 249208 3528
rect 249708 3476 249760 3528
rect 250352 3476 250404 3528
rect 251088 3476 251140 3528
rect 251456 3476 251508 3528
rect 252468 3476 252520 3528
rect 252652 3476 252704 3528
rect 253848 3476 253900 3528
rect 257436 3476 257488 3528
rect 257988 3476 258040 3528
rect 259828 3476 259880 3528
rect 261484 3476 261536 3528
rect 262220 3476 262272 3528
rect 263508 3476 263560 3528
rect 265808 3476 265860 3528
rect 266268 3476 266320 3528
rect 268108 3476 268160 3528
rect 269028 3476 269080 3528
rect 270500 3476 270552 3528
rect 272524 3476 272576 3528
rect 274088 3476 274140 3528
rect 274548 3476 274600 3528
rect 275284 3476 275336 3528
rect 275928 3476 275980 3528
rect 276480 3476 276532 3528
rect 277308 3476 277360 3528
rect 302148 3476 302200 3528
rect 302608 3476 302660 3528
rect 304908 3476 304960 3528
rect 306196 3476 306248 3528
rect 310428 3476 310480 3528
rect 313372 3476 313424 3528
rect 157524 3408 157576 3460
rect 158628 3408 158680 3460
rect 161112 3408 161164 3460
rect 189080 3408 189132 3460
rect 189632 3408 189684 3460
rect 211160 3408 211212 3460
rect 212264 3408 212316 3460
rect 229100 3408 229152 3460
rect 230112 3408 230164 3460
rect 242992 3408 243044 3460
rect 267004 3408 267056 3460
rect 267648 3408 267700 3460
rect 277676 3408 277728 3460
rect 280252 3408 280304 3460
rect 303528 3408 303580 3460
rect 305000 3408 305052 3460
rect 307668 3408 307720 3460
rect 310980 3408 311032 3460
rect 313188 3408 313240 3460
rect 316960 3476 317012 3528
rect 318708 3476 318760 3528
rect 325240 3476 325292 3528
rect 326344 3476 326396 3528
rect 332416 3476 332468 3528
rect 315856 3408 315908 3460
rect 321652 3408 321704 3460
rect 322848 3408 322900 3460
rect 330024 3408 330076 3460
rect 18328 3340 18380 3392
rect 19984 3340 20036 3392
rect 26700 3340 26752 3392
rect 27528 3340 27580 3392
rect 27896 3340 27948 3392
rect 28908 3340 28960 3392
rect 33876 3340 33928 3392
rect 34428 3340 34480 3392
rect 34980 3340 35032 3392
rect 35808 3340 35860 3392
rect 37372 3340 37424 3392
rect 38476 3340 38528 3392
rect 42156 3340 42208 3392
rect 42708 3340 42760 3392
rect 50528 3340 50580 3392
rect 50988 3340 51040 3392
rect 52828 3340 52880 3392
rect 53748 3340 53800 3392
rect 44548 3272 44600 3324
rect 45468 3272 45520 3324
rect 46940 3272 46992 3324
rect 95700 3340 95752 3392
rect 96528 3340 96580 3392
rect 98092 3340 98144 3392
rect 99288 3340 99340 3392
rect 101588 3340 101640 3392
rect 102048 3340 102100 3392
rect 102784 3340 102836 3392
rect 103428 3340 103480 3392
rect 105176 3340 105228 3392
rect 106188 3340 106240 3392
rect 113548 3340 113600 3392
rect 150808 3340 150860 3392
rect 152740 3340 152792 3392
rect 175372 3340 175424 3392
rect 200120 3340 200172 3392
rect 200396 3340 200448 3392
rect 219532 3340 219584 3392
rect 227720 3340 227772 3392
rect 229008 3340 229060 3392
rect 310336 3340 310388 3392
rect 314568 3340 314620 3392
rect 328276 3340 328328 3392
rect 337108 3476 337160 3528
rect 343548 3476 343600 3528
rect 356152 3476 356204 3528
rect 357348 3476 357400 3528
rect 374000 3476 374052 3528
rect 375196 3476 375248 3528
rect 396632 3476 396684 3528
rect 398748 3476 398800 3528
rect 425152 3476 425204 3528
rect 431868 3476 431920 3528
rect 467840 3476 467892 3528
rect 467932 3476 467984 3528
rect 469128 3476 469180 3528
rect 507216 3544 507268 3596
rect 513104 3544 513156 3596
rect 571432 3544 571484 3596
rect 514392 3476 514444 3528
rect 515956 3476 516008 3528
rect 575020 3544 575072 3596
rect 574744 3476 574796 3528
rect 576216 3476 576268 3528
rect 54024 3272 54076 3324
rect 103520 3272 103572 3324
rect 117136 3272 117188 3324
rect 153200 3272 153252 3324
rect 174176 3272 174228 3324
rect 198740 3272 198792 3324
rect 199200 3272 199252 3324
rect 218336 3272 218388 3324
rect 253848 3272 253900 3324
rect 257344 3272 257396 3324
rect 320824 3272 320876 3324
rect 324044 3272 324096 3324
rect 331036 3272 331088 3324
rect 340696 3408 340748 3460
rect 342076 3408 342128 3460
rect 354956 3408 355008 3460
rect 360108 3408 360160 3460
rect 377588 3408 377640 3460
rect 380716 3408 380768 3460
rect 403716 3408 403768 3460
rect 404268 3408 404320 3460
rect 432328 3408 432380 3460
rect 433340 3408 433392 3460
rect 434628 3408 434680 3460
rect 437296 3408 437348 3460
rect 473912 3408 473964 3460
rect 474648 3408 474700 3460
rect 521384 3408 521436 3460
rect 521568 3408 521620 3460
rect 581000 3408 581052 3460
rect 333888 3340 333940 3392
rect 343088 3340 343140 3392
rect 346216 3340 346268 3392
rect 358544 3340 358596 3392
rect 358728 3340 358780 3392
rect 375196 3340 375248 3392
rect 378048 3340 378100 3392
rect 399024 3340 399076 3392
rect 437388 3340 437440 3392
rect 475108 3340 475160 3392
rect 542912 3340 542964 3392
rect 340788 3272 340840 3324
rect 352564 3272 352616 3324
rect 353208 3272 353260 3324
rect 368020 3272 368072 3324
rect 380808 3272 380860 3324
rect 402520 3272 402572 3324
rect 440148 3272 440200 3324
rect 477500 3272 477552 3324
rect 485688 3272 485740 3324
rect 535736 3272 535788 3324
rect 536840 3272 536892 3324
rect 538128 3272 538180 3324
rect 10048 3204 10100 3256
rect 13084 3204 13136 3256
rect 61200 3204 61252 3256
rect 109408 3204 109460 3256
rect 114744 3204 114796 3256
rect 115848 3204 115900 3256
rect 120632 3204 120684 3256
rect 155960 3204 156012 3256
rect 179512 3204 179564 3256
rect 193220 3204 193272 3256
rect 214012 3204 214064 3256
rect 261024 3204 261076 3256
rect 262128 3204 262180 3256
rect 312544 3204 312596 3256
rect 315764 3204 315816 3256
rect 317328 3204 317380 3256
rect 322848 3204 322900 3256
rect 344928 3204 344980 3256
rect 357348 3204 357400 3256
rect 375288 3204 375340 3256
rect 395436 3204 395488 3256
rect 429108 3204 429160 3256
rect 464436 3204 464488 3256
rect 480168 3204 480220 3256
rect 528652 3204 528704 3256
rect 16028 3136 16080 3188
rect 17224 3136 17276 3188
rect 66352 3136 66404 3188
rect 71872 3136 71924 3188
rect 73160 3068 73212 3120
rect 81440 3068 81492 3120
rect 82728 3068 82780 3120
rect 121552 3136 121604 3188
rect 132500 3136 132552 3188
rect 201500 3136 201552 3188
rect 209872 3136 209924 3188
rect 226340 3136 226392 3188
rect 282460 3136 282512 3188
rect 284300 3136 284352 3188
rect 372436 3136 372488 3188
rect 391848 3136 391900 3188
rect 420828 3136 420880 3188
rect 453672 3136 453724 3188
rect 118884 3068 118936 3120
rect 164700 3068 164752 3120
rect 165528 3068 165580 3120
rect 205088 3068 205140 3120
rect 258632 3068 258684 3120
rect 259368 3068 259420 3120
rect 283656 3068 283708 3120
rect 284208 3068 284260 3120
rect 138480 3000 138532 3052
rect 139308 3000 139360 3052
rect 269304 3000 269356 3052
rect 270408 3000 270460 3052
rect 321468 3000 321520 3052
rect 327632 3000 327684 3052
rect 8852 2932 8904 2984
rect 10416 2932 10468 2984
rect 87328 2864 87380 2916
rect 88248 2864 88300 2916
rect 94504 2864 94556 2916
rect 95148 2864 95200 2916
rect 326988 2864 327040 2916
rect 334716 2864 334768 2916
rect 79048 824 79100 876
rect 79968 824 80020 876
rect 74264 552 74316 604
rect 74448 552 74500 604
rect 83832 552 83884 604
rect 84108 552 84160 604
rect 151544 552 151596 604
rect 151728 552 151780 604
rect 187240 552 187292 604
rect 187608 552 187660 604
rect 220544 552 220596 604
rect 220728 552 220780 604
rect 238392 552 238444 604
rect 238668 552 238720 604
rect 386420 552 386472 604
rect 387064 552 387116 604
rect 434720 552 434772 604
rect 435824 552 435876 604
rect 437480 552 437532 604
rect 438216 552 438268 604
rect 441620 552 441672 604
rect 441804 552 441856 604
rect 443092 552 443144 604
rect 444196 552 444248 604
rect 444380 552 444432 604
rect 445392 552 445444 604
rect 448520 552 448572 604
rect 448980 552 449032 604
rect 487068 552 487120 604
rect 488172 552 488224 604
rect 491208 552 491260 604
rect 491760 552 491812 604
rect 579620 552 579672 604
rect 579804 552 579856 604
<< metal2 >>
rect 10754 703520 10866 704960
rect 32374 703520 32486 704960
rect 53994 703520 54106 704960
rect 75614 703520 75726 704960
rect 97234 703520 97346 704960
rect 118854 703520 118966 704960
rect 140474 703520 140586 704960
rect 162094 703520 162206 704960
rect 183714 703520 183826 704960
rect 205426 703520 205538 704960
rect 227046 703520 227158 704960
rect 248666 703520 248778 704960
rect 270286 703520 270398 704960
rect 291906 703520 292018 704960
rect 313526 703520 313638 704960
rect 335146 703520 335258 704960
rect 356766 703520 356878 704960
rect 378386 703520 378498 704960
rect 400098 703520 400210 704960
rect 421718 703520 421830 704960
rect 443338 703520 443450 704960
rect 464958 703520 465070 704960
rect 486578 703520 486690 704960
rect 508198 703520 508310 704960
rect 529818 703520 529930 704960
rect 551438 703520 551550 704960
rect 573058 703520 573170 704960
rect 10796 695570 10824 703520
rect 32416 699718 32444 703520
rect 54036 700874 54064 703520
rect 54024 700868 54076 700874
rect 54024 700810 54076 700816
rect 55128 700868 55180 700874
rect 55128 700810 55180 700816
rect 32404 699712 32456 699718
rect 32404 699654 32456 699660
rect 33048 699712 33100 699718
rect 33048 699654 33100 699660
rect 10692 695564 10744 695570
rect 10692 695506 10744 695512
rect 10784 695564 10836 695570
rect 10784 695506 10836 695512
rect 3422 695464 3478 695473
rect 3422 695399 3478 695408
rect 3436 645862 3464 695399
rect 10704 688634 10732 695506
rect 10692 688628 10744 688634
rect 10692 688570 10744 688576
rect 10876 688628 10928 688634
rect 10876 688570 10928 688576
rect 10888 685846 10916 688570
rect 10876 685840 10928 685846
rect 10876 685782 10928 685788
rect 3514 678736 3570 678745
rect 3514 678671 3570 678680
rect 3424 645856 3476 645862
rect 3424 645798 3476 645804
rect 3528 630630 3556 678671
rect 10784 676252 10836 676258
rect 10784 676194 10836 676200
rect 10796 673538 10824 676194
rect 10784 673532 10836 673538
rect 10784 673474 10836 673480
rect 10968 673532 11020 673538
rect 10968 673474 11020 673480
rect 10980 663762 11008 673474
rect 10796 663734 11008 663762
rect 3606 662008 3662 662017
rect 3606 661943 3662 661952
rect 3516 630624 3568 630630
rect 3516 630566 3568 630572
rect 3422 628416 3478 628425
rect 3422 628351 3478 628360
rect 3436 587858 3464 628351
rect 3620 616826 3648 661943
rect 10796 654838 10824 663734
rect 33060 654906 33088 699654
rect 55140 654974 55168 700810
rect 75656 698358 75684 703520
rect 97276 699718 97304 703520
rect 118896 699718 118924 703520
rect 97264 699712 97316 699718
rect 97264 699654 97316 699660
rect 97908 699712 97960 699718
rect 97908 699654 97960 699660
rect 118884 699712 118936 699718
rect 118884 699654 118936 699660
rect 119988 699712 120040 699718
rect 119988 699654 120040 699660
rect 75644 698352 75696 698358
rect 75644 698294 75696 698300
rect 75644 694204 75696 694210
rect 75644 694146 75696 694152
rect 75656 688702 75684 694146
rect 75644 688696 75696 688702
rect 75644 688638 75696 688644
rect 75552 688628 75604 688634
rect 75552 688570 75604 688576
rect 75564 679046 75592 688570
rect 75552 679040 75604 679046
rect 75552 678982 75604 678988
rect 75460 678972 75512 678978
rect 75460 678914 75512 678920
rect 75472 669322 75500 678914
rect 75460 669316 75512 669322
rect 75460 669258 75512 669264
rect 75644 669316 75696 669322
rect 75644 669258 75696 669264
rect 75656 666534 75684 669258
rect 75644 666528 75696 666534
rect 75644 666470 75696 666476
rect 75552 656940 75604 656946
rect 75552 656882 75604 656888
rect 55128 654968 55180 654974
rect 55128 654910 55180 654916
rect 33048 654900 33100 654906
rect 33048 654842 33100 654848
rect 75564 654838 75592 656882
rect 97920 654906 97948 699654
rect 120000 654974 120028 699654
rect 140516 695570 140544 703520
rect 162136 699718 162164 703520
rect 183756 700194 183784 703520
rect 183744 700188 183796 700194
rect 183744 700130 183796 700136
rect 184848 700188 184900 700194
rect 184848 700130 184900 700136
rect 162124 699712 162176 699718
rect 162124 699654 162176 699660
rect 162768 699712 162820 699718
rect 162768 699654 162820 699660
rect 140412 695564 140464 695570
rect 140412 695506 140464 695512
rect 140504 695564 140556 695570
rect 140504 695506 140556 695512
rect 140424 688634 140452 695506
rect 140412 688628 140464 688634
rect 140412 688570 140464 688576
rect 140596 688628 140648 688634
rect 140596 688570 140648 688576
rect 140608 685846 140636 688570
rect 140596 685840 140648 685846
rect 140596 685782 140648 685788
rect 140504 676252 140556 676258
rect 140504 676194 140556 676200
rect 140516 673538 140544 676194
rect 140504 673532 140556 673538
rect 140504 673474 140556 673480
rect 140688 673532 140740 673538
rect 140688 673474 140740 673480
rect 140700 663762 140728 673474
rect 140516 663734 140728 663762
rect 104532 654968 104584 654974
rect 104532 654910 104584 654916
rect 119988 654968 120040 654974
rect 119988 654910 120040 654916
rect 87512 654900 87564 654906
rect 87512 654842 87564 654848
rect 97908 654900 97960 654906
rect 97908 654842 97960 654848
rect 10784 654832 10836 654838
rect 10784 654774 10836 654780
rect 70492 654832 70544 654838
rect 70492 654774 70544 654780
rect 75552 654832 75604 654838
rect 75552 654774 75604 654780
rect 70504 651916 70532 654774
rect 87524 651916 87552 654842
rect 104544 651916 104572 654910
rect 138572 654900 138624 654906
rect 138572 654842 138624 654848
rect 121552 654832 121604 654838
rect 121552 654774 121604 654780
rect 121564 651916 121592 654774
rect 138584 651916 138612 654842
rect 140516 654838 140544 663734
rect 155592 654968 155644 654974
rect 155592 654910 155644 654916
rect 140504 654832 140556 654838
rect 140504 654774 140556 654780
rect 155604 651916 155632 654910
rect 162780 654906 162808 699654
rect 162768 654900 162820 654906
rect 162768 654842 162820 654848
rect 184860 654838 184888 700130
rect 205468 698442 205496 703520
rect 227088 699718 227116 703520
rect 248708 699718 248736 703520
rect 270328 703474 270356 703520
rect 270328 703446 270448 703474
rect 227076 699712 227128 699718
rect 227076 699654 227128 699660
rect 227628 699712 227680 699718
rect 227628 699654 227680 699660
rect 248696 699712 248748 699718
rect 248696 699654 248748 699660
rect 249708 699712 249760 699718
rect 249708 699654 249760 699660
rect 205468 698414 205680 698442
rect 205652 694142 205680 698414
rect 205640 694136 205692 694142
rect 205640 694078 205692 694084
rect 205548 684548 205600 684554
rect 205548 684490 205600 684496
rect 205560 679046 205588 684490
rect 205548 679040 205600 679046
rect 205548 678982 205600 678988
rect 205456 678972 205508 678978
rect 205456 678914 205508 678920
rect 205468 669390 205496 678914
rect 205456 669384 205508 669390
rect 205456 669326 205508 669332
rect 205364 669316 205416 669322
rect 205364 669258 205416 669264
rect 205376 659734 205404 669258
rect 205364 659728 205416 659734
rect 205364 659670 205416 659676
rect 205272 659660 205324 659666
rect 205272 659602 205324 659608
rect 205284 654906 205312 659602
rect 189724 654900 189776 654906
rect 189724 654842 189776 654848
rect 205272 654900 205324 654906
rect 205272 654842 205324 654848
rect 223764 654900 223816 654906
rect 223764 654842 223816 654848
rect 172704 654832 172756 654838
rect 172704 654774 172756 654780
rect 184848 654832 184900 654838
rect 184848 654774 184900 654780
rect 172716 651916 172744 654774
rect 189736 651916 189764 654842
rect 206744 654832 206796 654838
rect 206744 654774 206796 654780
rect 206756 651916 206784 654774
rect 223776 651916 223804 654842
rect 227640 654838 227668 699654
rect 249720 655518 249748 699654
rect 270420 695502 270448 703446
rect 291948 699718 291976 703520
rect 313568 699718 313596 703520
rect 335188 699718 335216 703520
rect 356808 700330 356836 703520
rect 378428 700398 378456 703520
rect 360108 700392 360160 700398
rect 360108 700334 360160 700340
rect 378416 700392 378468 700398
rect 378416 700334 378468 700340
rect 394608 700392 394660 700398
rect 394608 700334 394660 700340
rect 343548 700324 343600 700330
rect 343548 700266 343600 700272
rect 356796 700324 356848 700330
rect 356796 700266 356848 700272
rect 291200 699712 291252 699718
rect 291200 699654 291252 699660
rect 291936 699712 291988 699718
rect 291936 699654 291988 699660
rect 309048 699712 309100 699718
rect 309048 699654 309100 699660
rect 313556 699712 313608 699718
rect 313556 699654 313608 699660
rect 326988 699712 327040 699718
rect 326988 699654 327040 699660
rect 335176 699712 335228 699718
rect 335176 699654 335228 699660
rect 270408 695496 270460 695502
rect 270408 695438 270460 695444
rect 270316 685908 270368 685914
rect 270316 685850 270368 685856
rect 270328 679046 270356 685850
rect 270316 679040 270368 679046
rect 270316 678982 270368 678988
rect 270224 678972 270276 678978
rect 270224 678914 270276 678920
rect 270236 673538 270264 678914
rect 270224 673532 270276 673538
rect 270224 673474 270276 673480
rect 270408 673532 270460 673538
rect 270408 673474 270460 673480
rect 270420 663762 270448 673474
rect 270236 663734 270448 663762
rect 270236 655518 270264 663734
rect 249708 655512 249760 655518
rect 249708 655454 249760 655460
rect 257896 655512 257948 655518
rect 257896 655454 257948 655460
rect 270224 655512 270276 655518
rect 270224 655454 270276 655460
rect 274916 655512 274968 655518
rect 274916 655454 274968 655460
rect 227628 654832 227680 654838
rect 227628 654774 227680 654780
rect 240784 654832 240836 654838
rect 240784 654774 240836 654780
rect 240796 651916 240824 654774
rect 257908 651916 257936 655454
rect 274928 651916 274956 655454
rect 291212 651794 291240 699654
rect 309060 651930 309088 699654
rect 327000 655178 327028 699654
rect 325976 655172 326028 655178
rect 325976 655114 326028 655120
rect 326988 655172 327040 655178
rect 326988 655114 327040 655120
rect 308982 651902 309088 651930
rect 325988 651916 326016 655114
rect 343560 651794 343588 700266
rect 360120 651916 360148 700334
rect 378048 700324 378100 700330
rect 378048 700266 378100 700272
rect 378060 655518 378088 700266
rect 377128 655512 377180 655518
rect 377128 655454 377180 655460
rect 378048 655512 378100 655518
rect 378048 655454 378100 655460
rect 377140 651916 377168 655454
rect 394620 651794 394648 700334
rect 400140 700330 400168 703520
rect 421760 700398 421788 703520
rect 429108 700460 429160 700466
rect 429108 700402 429160 700408
rect 421748 700392 421800 700398
rect 421748 700334 421800 700340
rect 400128 700324 400180 700330
rect 400128 700266 400180 700272
rect 411168 700324 411220 700330
rect 411168 700266 411220 700272
rect 411180 651916 411208 700266
rect 429120 655518 429148 700402
rect 443380 700330 443408 703520
rect 465000 700466 465028 703520
rect 464988 700460 465040 700466
rect 464988 700402 465040 700408
rect 480168 700460 480220 700466
rect 480168 700402 480220 700408
rect 445668 700392 445720 700398
rect 445668 700334 445720 700340
rect 443368 700324 443420 700330
rect 443368 700266 443420 700272
rect 428188 655512 428240 655518
rect 428188 655454 428240 655460
rect 429108 655512 429160 655518
rect 429108 655454 429160 655460
rect 428200 651916 428228 655454
rect 445680 651930 445708 700334
rect 463608 700324 463660 700330
rect 463608 700266 463660 700272
rect 463620 655518 463648 700266
rect 480180 655518 480208 700402
rect 486620 700398 486648 703520
rect 486608 700392 486660 700398
rect 486608 700334 486660 700340
rect 496728 700392 496780 700398
rect 496728 700334 496780 700340
rect 462320 655512 462372 655518
rect 462320 655454 462372 655460
rect 463608 655512 463660 655518
rect 463608 655454 463660 655460
rect 479340 655512 479392 655518
rect 479340 655454 479392 655460
rect 480168 655512 480220 655518
rect 480168 655454 480220 655460
rect 445326 651902 445708 651930
rect 462332 651916 462360 655454
rect 479352 651916 479380 655454
rect 496740 651930 496768 700334
rect 508240 700330 508268 703520
rect 529860 700466 529888 703520
rect 529848 700460 529900 700466
rect 529848 700402 529900 700408
rect 551480 700398 551508 703520
rect 551468 700392 551520 700398
rect 551468 700334 551520 700340
rect 573100 700330 573128 703520
rect 508228 700324 508280 700330
rect 508228 700266 508280 700272
rect 514668 700324 514720 700330
rect 514668 700266 514720 700272
rect 573088 700324 573140 700330
rect 573088 700266 573140 700272
rect 514680 655314 514708 700266
rect 580170 696008 580226 696017
rect 580170 695943 580226 695952
rect 580184 695570 580212 695943
rect 523684 695564 523736 695570
rect 523684 695506 523736 695512
rect 580172 695564 580224 695570
rect 580172 695506 580224 695512
rect 513380 655308 513432 655314
rect 513380 655250 513432 655256
rect 514668 655308 514720 655314
rect 514668 655250 514720 655256
rect 496386 651902 496768 651930
rect 513392 651916 513420 655250
rect 291212 651766 291962 651794
rect 343022 651766 343588 651794
rect 394174 651766 394648 651794
rect 59360 645856 59412 645862
rect 59360 645798 59412 645804
rect 3698 645280 3754 645289
rect 3698 645215 3754 645224
rect 3608 616820 3660 616826
rect 3608 616762 3660 616768
rect 3514 611688 3570 611697
rect 3514 611623 3570 611632
rect 3424 587852 3476 587858
rect 3424 587794 3476 587800
rect 3422 578232 3478 578241
rect 3422 578167 3478 578176
rect 3436 545086 3464 578167
rect 3528 574054 3556 611623
rect 3712 603090 3740 645215
rect 59372 644745 59400 645798
rect 523696 645289 523724 695506
rect 523776 680400 523828 680406
rect 580172 680400 580224 680406
rect 523776 680342 523828 680348
rect 580170 680368 580172 680377
rect 580224 680368 580226 680377
rect 523682 645280 523738 645289
rect 523682 645215 523738 645224
rect 59358 644736 59414 644745
rect 59358 644671 59414 644680
rect 523684 633480 523736 633486
rect 523684 633422 523736 633428
rect 59360 630624 59412 630630
rect 59360 630566 59412 630572
rect 59372 630465 59400 630566
rect 59358 630456 59414 630465
rect 59358 630391 59414 630400
rect 59360 616820 59412 616826
rect 59360 616762 59412 616768
rect 59372 616185 59400 616762
rect 59358 616176 59414 616185
rect 59358 616111 59414 616120
rect 523132 605804 523184 605810
rect 523132 605746 523184 605752
rect 523144 605305 523172 605746
rect 523130 605296 523186 605305
rect 523130 605231 523186 605240
rect 3700 603084 3752 603090
rect 3700 603026 3752 603032
rect 59360 603084 59412 603090
rect 59360 603026 59412 603032
rect 59372 601905 59400 603026
rect 59358 601896 59414 601905
rect 59358 601831 59414 601840
rect 3606 594960 3662 594969
rect 3606 594895 3662 594904
rect 3516 574048 3568 574054
rect 3516 573990 3568 573996
rect 3514 561368 3570 561377
rect 3514 561303 3570 561312
rect 3424 545080 3476 545086
rect 3424 545022 3476 545028
rect 3528 531282 3556 561303
rect 3620 560250 3648 594895
rect 523696 591977 523724 633422
rect 523788 631961 523816 680342
rect 580170 680303 580226 680312
rect 580262 664728 580318 664737
rect 580262 664663 580318 664672
rect 580172 633480 580224 633486
rect 580170 633448 580172 633457
rect 580224 633448 580226 633457
rect 580170 633383 580226 633392
rect 523774 631952 523830 631961
rect 523774 631887 523830 631896
rect 580276 619614 580304 664663
rect 580354 649088 580410 649097
rect 580354 649023 580410 649032
rect 524328 619608 524380 619614
rect 524328 619550 524380 619556
rect 580264 619608 580316 619614
rect 580264 619550 580316 619556
rect 524340 618633 524368 619550
rect 524326 618624 524382 618633
rect 524326 618559 524382 618568
rect 580262 617808 580318 617817
rect 580262 617743 580318 617752
rect 580170 602168 580226 602177
rect 580170 602103 580226 602112
rect 580184 601730 580212 602103
rect 523776 601724 523828 601730
rect 523776 601666 523828 601672
rect 580172 601724 580224 601730
rect 580172 601666 580224 601672
rect 523682 591968 523738 591977
rect 523682 591903 523738 591912
rect 59360 587852 59412 587858
rect 59360 587794 59412 587800
rect 59372 587625 59400 587794
rect 59358 587616 59414 587625
rect 59358 587551 59414 587560
rect 523684 586560 523736 586566
rect 523684 586502 523736 586508
rect 59360 574048 59412 574054
rect 59360 573990 59412 573996
rect 59372 573345 59400 573990
rect 59358 573336 59414 573345
rect 59358 573271 59414 573280
rect 3608 560244 3660 560250
rect 3608 560186 3660 560192
rect 59360 560244 59412 560250
rect 59360 560186 59412 560192
rect 59372 559065 59400 560186
rect 59358 559056 59414 559065
rect 59358 558991 59414 559000
rect 523696 551993 523724 586502
rect 523788 565321 523816 601666
rect 580172 586560 580224 586566
rect 580170 586528 580172 586537
rect 580224 586528 580226 586537
rect 580170 586463 580226 586472
rect 580276 579630 580304 617743
rect 580368 605810 580396 649023
rect 580356 605804 580408 605810
rect 580356 605746 580408 605752
rect 524328 579624 524380 579630
rect 524328 579566 524380 579572
rect 580264 579624 580316 579630
rect 580264 579566 580316 579572
rect 524340 578649 524368 579566
rect 524326 578640 524382 578649
rect 524326 578575 524382 578584
rect 580262 570888 580318 570897
rect 580262 570823 580318 570832
rect 523774 565312 523830 565321
rect 523774 565247 523830 565256
rect 580170 555248 580226 555257
rect 580170 555183 580226 555192
rect 580184 554810 580212 555183
rect 523776 554804 523828 554810
rect 523776 554746 523828 554752
rect 580172 554804 580224 554810
rect 580172 554746 580224 554752
rect 523682 551984 523738 551993
rect 523682 551919 523738 551928
rect 59360 545080 59412 545086
rect 59360 545022 59412 545028
rect 59372 544785 59400 545022
rect 59358 544776 59414 544785
rect 59358 544711 59414 544720
rect 3606 544640 3662 544649
rect 3606 544575 3662 544584
rect 3516 531276 3568 531282
rect 3516 531218 3568 531224
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 502314 3464 527847
rect 3620 517478 3648 544575
rect 523500 539640 523552 539646
rect 523500 539582 523552 539588
rect 523512 538234 523540 539582
rect 523684 539572 523736 539578
rect 523684 539514 523736 539520
rect 523696 538665 523724 539514
rect 523682 538656 523738 538665
rect 523682 538591 523738 538600
rect 523512 538206 523724 538234
rect 59360 531276 59412 531282
rect 59360 531218 59412 531224
rect 59372 530505 59400 531218
rect 59358 530496 59414 530505
rect 59358 530431 59414 530440
rect 3608 517472 3660 517478
rect 3608 517414 3660 517420
rect 59360 517472 59412 517478
rect 59360 517414 59412 517420
rect 59372 516225 59400 517414
rect 59358 516216 59414 516225
rect 59358 516151 59414 516160
rect 523696 512009 523724 538206
rect 523788 525337 523816 554746
rect 580172 539640 580224 539646
rect 580170 539608 580172 539617
rect 580224 539608 580226 539617
rect 580276 539578 580304 570823
rect 580170 539543 580226 539552
rect 580264 539572 580316 539578
rect 580264 539514 580316 539520
rect 523774 525328 523830 525337
rect 523774 525263 523830 525272
rect 580170 523968 580226 523977
rect 580170 523903 580226 523912
rect 580184 523054 580212 523903
rect 523776 523048 523828 523054
rect 523776 522990 523828 522996
rect 580172 523048 580224 523054
rect 580172 522990 580224 522996
rect 523682 512000 523738 512009
rect 523682 511935 523738 511944
rect 3514 511184 3570 511193
rect 3514 511119 3570 511128
rect 3424 502308 3476 502314
rect 3424 502250 3476 502256
rect 3422 494320 3478 494329
rect 3422 494255 3478 494264
rect 3436 474706 3464 494255
rect 3528 488510 3556 511119
rect 523684 507884 523736 507890
rect 523684 507826 523736 507832
rect 59360 502308 59412 502314
rect 59360 502250 59412 502256
rect 59372 501945 59400 502250
rect 59358 501936 59414 501945
rect 59358 501871 59414 501880
rect 3516 488504 3568 488510
rect 3516 488446 3568 488452
rect 59360 488504 59412 488510
rect 59360 488446 59412 488452
rect 59372 487665 59400 488446
rect 59358 487656 59414 487665
rect 59358 487591 59414 487600
rect 523696 485353 523724 507826
rect 523788 498681 523816 522990
rect 580170 508328 580226 508337
rect 580170 508263 580226 508272
rect 580184 507890 580212 508263
rect 580172 507884 580224 507890
rect 580172 507826 580224 507832
rect 523774 498672 523830 498681
rect 523774 498607 523830 498616
rect 523776 492720 523828 492726
rect 580172 492720 580224 492726
rect 523776 492662 523828 492668
rect 580170 492688 580172 492697
rect 580224 492688 580226 492697
rect 523682 485344 523738 485353
rect 523682 485279 523738 485288
rect 3514 477592 3570 477601
rect 3514 477527 3570 477536
rect 3424 474700 3476 474706
rect 3424 474642 3476 474648
rect 3422 460864 3478 460873
rect 3422 460799 3478 460808
rect 3436 445738 3464 460799
rect 3528 459542 3556 477527
rect 523684 476128 523736 476134
rect 523684 476070 523736 476076
rect 59360 474700 59412 474706
rect 59360 474642 59412 474648
rect 59372 473385 59400 474642
rect 59358 473376 59414 473385
rect 59358 473311 59414 473320
rect 3516 459536 3568 459542
rect 3516 459478 3568 459484
rect 59360 459536 59412 459542
rect 59360 459478 59412 459484
rect 59372 459105 59400 459478
rect 59358 459096 59414 459105
rect 59358 459031 59414 459040
rect 523696 458697 523724 476070
rect 523788 472025 523816 492662
rect 580170 492623 580226 492632
rect 580170 477048 580226 477057
rect 580170 476983 580226 476992
rect 580184 476134 580212 476983
rect 580172 476128 580224 476134
rect 580172 476070 580224 476076
rect 523774 472016 523830 472025
rect 523774 471951 523830 471960
rect 580170 461408 580226 461417
rect 580170 461343 580226 461352
rect 580184 460970 580212 461343
rect 523776 460964 523828 460970
rect 523776 460906 523828 460912
rect 580172 460964 580224 460970
rect 580172 460906 580224 460912
rect 523682 458688 523738 458697
rect 523682 458623 523738 458632
rect 523684 445800 523736 445806
rect 523684 445742 523736 445748
rect 3424 445732 3476 445738
rect 3424 445674 3476 445680
rect 59360 445732 59412 445738
rect 59360 445674 59412 445680
rect 59372 444825 59400 445674
rect 59358 444816 59414 444825
rect 59358 444751 59414 444760
rect 3422 444136 3478 444145
rect 3422 444071 3478 444080
rect 3436 430574 3464 444071
rect 523696 432041 523724 445742
rect 523788 445369 523816 460906
rect 580172 445800 580224 445806
rect 580170 445768 580172 445777
rect 580224 445768 580226 445777
rect 580170 445703 580226 445712
rect 523774 445360 523830 445369
rect 523774 445295 523830 445304
rect 523682 432032 523738 432041
rect 523682 431967 523738 431976
rect 3424 430568 3476 430574
rect 59360 430568 59412 430574
rect 3424 430510 3476 430516
rect 59358 430536 59360 430545
rect 59412 430536 59414 430545
rect 59358 430471 59414 430480
rect 580170 430128 580226 430137
rect 580170 430063 580226 430072
rect 580184 429214 580212 430063
rect 523684 429208 523736 429214
rect 523684 429150 523736 429156
rect 580172 429208 580224 429214
rect 580172 429150 580224 429156
rect 3422 427272 3478 427281
rect 3422 427207 3478 427216
rect 3436 416770 3464 427207
rect 523696 418713 523724 429150
rect 523682 418704 523738 418713
rect 523682 418639 523738 418648
rect 3424 416764 3476 416770
rect 3424 416706 3476 416712
rect 59360 416764 59412 416770
rect 59360 416706 59412 416712
rect 59372 416265 59400 416706
rect 59358 416256 59414 416265
rect 59358 416191 59414 416200
rect 580170 414488 580226 414497
rect 580170 414423 580226 414432
rect 580184 414050 580212 414423
rect 523684 414044 523736 414050
rect 523684 413986 523736 413992
rect 580172 414044 580224 414050
rect 580172 413986 580224 413992
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 402966 3464 410479
rect 523696 405385 523724 413986
rect 523682 405376 523738 405385
rect 523682 405311 523738 405320
rect 3424 402960 3476 402966
rect 3424 402902 3476 402908
rect 59360 402960 59412 402966
rect 59360 402902 59412 402908
rect 59372 401985 59400 402902
rect 59358 401976 59414 401985
rect 59358 401911 59414 401920
rect 523684 398880 523736 398886
rect 580172 398880 580224 398886
rect 523684 398822 523736 398828
rect 580170 398848 580172 398857
rect 580224 398848 580226 398857
rect 3882 393816 3938 393825
rect 3882 393751 3938 393760
rect 3896 387802 3924 393751
rect 523696 392057 523724 398822
rect 580170 398783 580226 398792
rect 523682 392048 523738 392057
rect 523682 391983 523738 391992
rect 3884 387796 3936 387802
rect 3884 387738 3936 387744
rect 59360 387796 59412 387802
rect 59360 387738 59412 387744
rect 59372 387705 59400 387738
rect 59358 387696 59414 387705
rect 59358 387631 59414 387640
rect 580170 383208 580226 383217
rect 580170 383143 580226 383152
rect 580184 382294 580212 383143
rect 523132 382288 523184 382294
rect 523132 382230 523184 382236
rect 580172 382288 580224 382294
rect 580172 382230 580224 382236
rect 523144 378729 523172 382230
rect 523130 378720 523186 378729
rect 523130 378655 523186 378664
rect 3422 377088 3478 377097
rect 3422 377023 3478 377032
rect 3436 373998 3464 377023
rect 3424 373992 3476 373998
rect 3424 373934 3476 373940
rect 59360 373992 59412 373998
rect 59360 373934 59412 373940
rect 59372 373425 59400 373934
rect 59358 373416 59414 373425
rect 59358 373351 59414 373360
rect 580170 367568 580226 367577
rect 580170 367503 580226 367512
rect 580184 367130 580212 367503
rect 523316 367124 523368 367130
rect 523316 367066 523368 367072
rect 580172 367124 580224 367130
rect 580172 367066 580224 367072
rect 523328 365401 523356 367066
rect 523314 365392 523370 365401
rect 523314 365327 523370 365336
rect 3422 360360 3478 360369
rect 3422 360295 3478 360304
rect 3436 360194 3464 360295
rect 3424 360188 3476 360194
rect 3424 360130 3476 360136
rect 59360 360188 59412 360194
rect 59360 360130 59412 360136
rect 59372 359145 59400 360130
rect 59358 359136 59414 359145
rect 59358 359071 59414 359080
rect 524328 352572 524380 352578
rect 524328 352514 524380 352520
rect 580172 352572 580224 352578
rect 580172 352514 580224 352520
rect 524340 351937 524368 352514
rect 580184 351937 580212 352514
rect 524326 351928 524382 351937
rect 524326 351863 524382 351872
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 59358 344720 59414 344729
rect 59358 344655 59414 344664
rect 59372 343602 59400 344655
rect 3424 343596 3476 343602
rect 3424 343538 3476 343544
rect 59360 343596 59412 343602
rect 59360 343538 59412 343544
rect 3436 343505 3464 343538
rect 3422 343496 3478 343505
rect 3422 343431 3478 343440
rect 523406 338600 523462 338609
rect 523406 338535 523462 338544
rect 523420 336734 523448 338535
rect 523408 336728 523460 336734
rect 523408 336670 523460 336676
rect 580172 336728 580224 336734
rect 580172 336670 580224 336676
rect 580184 336297 580212 336670
rect 580170 336288 580226 336297
rect 580170 336223 580226 336232
rect 59358 330440 59414 330449
rect 59358 330375 59414 330384
rect 59372 327078 59400 330375
rect 3332 327072 3384 327078
rect 3332 327014 3384 327020
rect 59360 327072 59412 327078
rect 59360 327014 59412 327020
rect 3344 326777 3372 327014
rect 3330 326768 3386 326777
rect 3330 326703 3386 326712
rect 523130 325272 523186 325281
rect 523130 325207 523186 325216
rect 523144 321570 523172 325207
rect 523132 321564 523184 321570
rect 523132 321506 523184 321512
rect 580172 321564 580224 321570
rect 580172 321506 580224 321512
rect 580184 320657 580212 321506
rect 580170 320648 580226 320657
rect 580170 320583 580226 320592
rect 60002 316160 60058 316169
rect 60002 316095 60058 316104
rect 60016 310486 60044 316095
rect 523682 311944 523738 311953
rect 523682 311879 523738 311888
rect 3424 310480 3476 310486
rect 3424 310422 3476 310428
rect 60004 310480 60056 310486
rect 60004 310422 60056 310428
rect 3436 310049 3464 310422
rect 3422 310040 3478 310049
rect 3422 309975 3478 309984
rect 523696 306338 523724 311879
rect 523684 306332 523736 306338
rect 523684 306274 523736 306280
rect 580172 306332 580224 306338
rect 580172 306274 580224 306280
rect 580184 305017 580212 306274
rect 580170 305008 580226 305017
rect 580170 304943 580226 304952
rect 60002 301880 60058 301889
rect 60002 301815 60058 301824
rect 60016 293962 60044 301815
rect 523682 298616 523738 298625
rect 523682 298551 523738 298560
rect 3148 293956 3200 293962
rect 3148 293898 3200 293904
rect 60004 293956 60056 293962
rect 60004 293898 60056 293904
rect 3160 293321 3188 293898
rect 3146 293312 3202 293321
rect 3146 293247 3202 293256
rect 523696 289814 523724 298551
rect 523684 289808 523736 289814
rect 523684 289750 523736 289756
rect 580172 289808 580224 289814
rect 580172 289750 580224 289756
rect 580184 289377 580212 289750
rect 580170 289368 580226 289377
rect 580170 289303 580226 289312
rect 60002 287600 60058 287609
rect 60002 287535 60058 287544
rect 60016 277370 60044 287535
rect 523682 285288 523738 285297
rect 523682 285223 523738 285232
rect 3424 277364 3476 277370
rect 3424 277306 3476 277312
rect 60004 277364 60056 277370
rect 60004 277306 60056 277312
rect 3436 276457 3464 277306
rect 3422 276448 3478 276457
rect 3422 276383 3478 276392
rect 523696 274650 523724 285223
rect 523684 274644 523736 274650
rect 523684 274586 523736 274592
rect 580172 274644 580224 274650
rect 580172 274586 580224 274592
rect 580184 273737 580212 274586
rect 580170 273728 580226 273737
rect 580170 273663 580226 273672
rect 60002 273320 60058 273329
rect 60002 273255 60058 273264
rect 60016 260846 60044 273255
rect 523682 271960 523738 271969
rect 523682 271895 523738 271904
rect 3424 260840 3476 260846
rect 3424 260782 3476 260788
rect 60004 260840 60056 260846
rect 60004 260782 60056 260788
rect 3436 259729 3464 260782
rect 3422 259720 3478 259729
rect 3422 259655 3478 259664
rect 523696 259418 523724 271895
rect 523684 259412 523736 259418
rect 523684 259354 523736 259360
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 60002 259040 60058 259049
rect 60002 258975 60058 258984
rect 60016 244254 60044 258975
rect 523774 258632 523830 258641
rect 523774 258567 523830 258576
rect 523682 245304 523738 245313
rect 523682 245239 523738 245248
rect 60094 244760 60150 244769
rect 60094 244695 60150 244704
rect 3424 244248 3476 244254
rect 3424 244190 3476 244196
rect 60004 244248 60056 244254
rect 60004 244190 60056 244196
rect 3436 243001 3464 244190
rect 3422 242992 3478 243001
rect 3422 242927 3478 242936
rect 60002 230480 60058 230489
rect 60002 230415 60058 230424
rect 3424 226296 3476 226302
rect 3422 226264 3424 226273
rect 3476 226264 3478 226273
rect 3422 226199 3478 226208
rect 60016 209778 60044 230415
rect 60108 226302 60136 244695
rect 523696 227730 523724 245239
rect 523788 242894 523816 258567
rect 580184 258097 580212 259354
rect 580170 258088 580226 258097
rect 580170 258023 580226 258032
rect 523776 242888 523828 242894
rect 523776 242830 523828 242836
rect 580172 242888 580224 242894
rect 580172 242830 580224 242836
rect 580184 242457 580212 242830
rect 580170 242448 580226 242457
rect 580170 242383 580226 242392
rect 523774 231976 523830 231985
rect 523774 231911 523830 231920
rect 523684 227724 523736 227730
rect 523684 227666 523736 227672
rect 60096 226296 60148 226302
rect 60096 226238 60148 226244
rect 523682 218648 523738 218657
rect 523682 218583 523738 218592
rect 60094 216200 60150 216209
rect 60094 216135 60150 216144
rect 3424 209772 3476 209778
rect 3424 209714 3476 209720
rect 60004 209772 60056 209778
rect 60004 209714 60056 209720
rect 3436 209409 3464 209714
rect 3422 209400 3478 209409
rect 3422 209335 3478 209344
rect 60002 201920 60058 201929
rect 60002 201855 60058 201864
rect 3516 193180 3568 193186
rect 3516 193122 3568 193128
rect 3528 192681 3556 193122
rect 3514 192672 3570 192681
rect 3514 192607 3570 192616
rect 60016 176662 60044 201855
rect 60108 193186 60136 216135
rect 523696 195974 523724 218583
rect 523788 212498 523816 231911
rect 580172 227724 580224 227730
rect 580172 227666 580224 227672
rect 580184 226817 580212 227666
rect 580170 226808 580226 226817
rect 580170 226743 580226 226752
rect 523776 212492 523828 212498
rect 523776 212434 523828 212440
rect 580172 212492 580224 212498
rect 580172 212434 580224 212440
rect 580184 211177 580212 212434
rect 580170 211168 580226 211177
rect 580170 211103 580226 211112
rect 523774 205320 523830 205329
rect 523774 205255 523830 205264
rect 523684 195968 523736 195974
rect 523684 195910 523736 195916
rect 60096 193180 60148 193186
rect 60096 193122 60148 193128
rect 523682 191992 523738 192001
rect 523682 191927 523738 191936
rect 60186 187640 60242 187649
rect 60186 187575 60242 187584
rect 3424 176656 3476 176662
rect 3424 176598 3476 176604
rect 60004 176656 60056 176662
rect 60004 176598 60056 176604
rect 3436 175953 3464 176598
rect 3422 175944 3478 175953
rect 3422 175879 3478 175888
rect 60094 173360 60150 173369
rect 60094 173295 60150 173304
rect 3148 160064 3200 160070
rect 3148 160006 3200 160012
rect 3160 159225 3188 160006
rect 3146 159216 3202 159225
rect 3146 159151 3202 159160
rect 60002 159080 60058 159089
rect 60002 159015 60058 159024
rect 3240 143540 3292 143546
rect 3240 143482 3292 143488
rect 3252 142361 3280 143482
rect 3238 142352 3294 142361
rect 3238 142287 3294 142296
rect 60016 126954 60044 159015
rect 60108 143546 60136 173295
rect 60200 160070 60228 187575
rect 523696 165578 523724 191927
rect 523788 180810 523816 205255
rect 580172 195968 580224 195974
rect 580172 195910 580224 195916
rect 580184 195537 580212 195910
rect 580170 195528 580226 195537
rect 580170 195463 580226 195472
rect 523776 180804 523828 180810
rect 523776 180746 523828 180752
rect 580172 180804 580224 180810
rect 580172 180746 580224 180752
rect 580184 179897 580212 180746
rect 580170 179888 580226 179897
rect 580170 179823 580226 179832
rect 523866 178664 523922 178673
rect 523866 178599 523922 178608
rect 523684 165572 523736 165578
rect 523684 165514 523736 165520
rect 523774 165336 523830 165345
rect 523774 165271 523830 165280
rect 60188 160064 60240 160070
rect 60188 160006 60240 160012
rect 523682 152008 523738 152017
rect 523682 151943 523738 151952
rect 60186 144800 60242 144809
rect 60186 144735 60242 144744
rect 60096 143540 60148 143546
rect 60096 143482 60148 143488
rect 60094 130520 60150 130529
rect 60094 130455 60150 130464
rect 3240 126948 3292 126954
rect 3240 126890 3292 126896
rect 60004 126948 60056 126954
rect 60004 126890 60056 126896
rect 3252 125633 3280 126890
rect 3238 125624 3294 125633
rect 3238 125559 3294 125568
rect 60002 116240 60058 116249
rect 60002 116175 60058 116184
rect 3424 108996 3476 109002
rect 3424 108938 3476 108944
rect 3436 108905 3464 108938
rect 3422 108896 3478 108905
rect 3422 108831 3478 108840
rect 3332 92472 3384 92478
rect 3332 92414 3384 92420
rect 3344 92177 3372 92414
rect 3330 92168 3386 92177
rect 3330 92103 3386 92112
rect 60016 75886 60044 116175
rect 60108 92478 60136 130455
rect 60200 109002 60228 144735
rect 523696 118658 523724 151943
rect 523788 133890 523816 165271
rect 523880 149054 523908 178599
rect 580172 165572 580224 165578
rect 580172 165514 580224 165520
rect 580184 164257 580212 165514
rect 580170 164248 580226 164257
rect 580170 164183 580226 164192
rect 523868 149048 523920 149054
rect 523868 148990 523920 148996
rect 580172 149048 580224 149054
rect 580172 148990 580224 148996
rect 580184 148617 580212 148990
rect 580170 148608 580226 148617
rect 580170 148543 580226 148552
rect 523866 138680 523922 138689
rect 523866 138615 523922 138624
rect 523776 133884 523828 133890
rect 523776 133826 523828 133832
rect 523774 125352 523830 125361
rect 523774 125287 523830 125296
rect 523684 118652 523736 118658
rect 523684 118594 523736 118600
rect 523682 112024 523738 112033
rect 523682 111959 523738 111968
rect 60188 108996 60240 109002
rect 60188 108938 60240 108944
rect 60278 101960 60334 101969
rect 60278 101895 60334 101904
rect 60096 92472 60148 92478
rect 60096 92414 60148 92420
rect 60186 87680 60242 87689
rect 60186 87615 60242 87624
rect 3424 75880 3476 75886
rect 3424 75822 3476 75828
rect 60004 75880 60056 75886
rect 60004 75822 60056 75828
rect 3436 75313 3464 75822
rect 3422 75304 3478 75313
rect 3422 75239 3478 75248
rect 60094 73400 60150 73409
rect 60094 73335 60150 73344
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 60002 59120 60058 59129
rect 60002 59055 60058 59064
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 57888 49292 57940 49298
rect 57888 49234 57940 49240
rect 50988 49224 51040 49230
rect 50988 49166 51040 49172
rect 13084 49156 13136 49162
rect 13084 49098 13136 49104
rect 8944 49088 8996 49094
rect 8944 49030 8996 49036
rect 3424 42764 3476 42770
rect 3424 42706 3476 42712
rect 3436 41857 3464 42706
rect 3422 41848 3478 41857
rect 3422 41783 3478 41792
rect 3424 26240 3476 26246
rect 3424 26182 3476 26188
rect 3436 25129 3464 26182
rect 3422 25120 3478 25129
rect 3422 25055 3478 25064
rect 4068 10328 4120 10334
rect 4068 10270 4120 10276
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3436 8401 3464 9590
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 1676 7608 1728 7614
rect 1676 7550 1728 7556
rect 572 6180 624 6186
rect 572 6122 624 6128
rect 584 480 612 6122
rect 1688 480 1716 7550
rect 4080 3534 4108 10270
rect 8956 3806 8984 49030
rect 10324 47592 10376 47598
rect 10324 47534 10376 47540
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 5264 3800 5316 3806
rect 5264 3742 5316 3748
rect 8944 3800 8996 3806
rect 8944 3742 8996 3748
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 2884 480 2912 3470
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 480 4108 3334
rect 5276 480 5304 3742
rect 9048 3534 9076 11698
rect 10336 3670 10364 47534
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 3470
rect 10048 3256 10100 3262
rect 10048 3198 10100 3204
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8864 480 8892 2926
rect 10060 480 10088 3198
rect 10428 2990 10456 18566
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 11256 480 11284 3538
rect 12452 480 12480 4762
rect 13096 3262 13124 49098
rect 17224 49020 17276 49026
rect 17224 48962 17276 48968
rect 14464 36576 14516 36582
rect 14464 36518 14516 36524
rect 14476 3534 14504 36518
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 13084 3256 13136 3262
rect 13084 3198 13136 3204
rect 13648 480 13676 3470
rect 14844 480 14872 3538
rect 17236 3194 17264 48962
rect 22008 46232 22060 46238
rect 22008 46174 22060 46180
rect 19984 35216 20036 35222
rect 19984 35158 20036 35164
rect 17316 4888 17368 4894
rect 17316 4830 17368 4836
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16040 480 16068 3130
rect 17328 2530 17356 4830
rect 19996 3398 20024 35158
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 18328 3392 18380 3398
rect 19984 3392 20036 3398
rect 18328 3334 18380 3340
rect 19522 3360 19578 3369
rect 17236 2502 17356 2530
rect 17236 480 17264 2502
rect 18340 480 18368 3334
rect 19984 3334 20036 3340
rect 19522 3295 19578 3304
rect 19536 480 19564 3295
rect 20732 480 20760 3606
rect 22020 3482 22048 46174
rect 27528 44872 27580 44878
rect 27528 44814 27580 44820
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23400 3482 23428 22714
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 21928 3454 22048 3482
rect 23124 3454 23428 3482
rect 21928 480 21956 3454
rect 23124 480 23152 3454
rect 24320 480 24348 3674
rect 25502 3496 25558 3505
rect 25502 3431 25558 3440
rect 25516 480 25544 3431
rect 27540 3398 27568 44814
rect 34428 43444 34480 43450
rect 34428 43386 34480 43392
rect 28908 33788 28960 33794
rect 28908 33730 28960 33736
rect 28920 3398 28948 33730
rect 31668 32428 31720 32434
rect 31668 32370 31720 32376
rect 30288 13116 30340 13122
rect 30288 13058 30340 13064
rect 29092 3800 29144 3806
rect 29092 3742 29144 3748
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 26712 480 26740 3334
rect 27908 480 27936 3334
rect 29104 480 29132 3742
rect 30300 480 30328 13058
rect 31680 3482 31708 32370
rect 32680 3868 32732 3874
rect 32680 3810 32732 3816
rect 31496 3454 31708 3482
rect 31496 480 31524 3454
rect 32692 480 32720 3810
rect 34440 3398 34468 43386
rect 42708 42084 42760 42090
rect 42708 42026 42760 42032
rect 35808 31068 35860 31074
rect 35808 31010 35860 31016
rect 35820 3398 35848 31010
rect 38568 29640 38620 29646
rect 38568 29582 38620 29588
rect 38476 14476 38528 14482
rect 38476 14418 38528 14424
rect 36176 4004 36228 4010
rect 36176 3946 36228 3952
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 33888 480 33916 3334
rect 34992 480 35020 3334
rect 36188 480 36216 3946
rect 38488 3398 38516 14418
rect 37372 3392 37424 3398
rect 37372 3334 37424 3340
rect 38476 3392 38528 3398
rect 38476 3334 38528 3340
rect 37384 480 37412 3334
rect 38580 480 38608 29582
rect 41328 15904 41380 15910
rect 41328 15846 41380 15852
rect 39764 3936 39816 3942
rect 39764 3878 39816 3884
rect 39776 480 39804 3878
rect 41340 3482 41368 15846
rect 40972 3454 41368 3482
rect 40972 480 41000 3454
rect 42720 3398 42748 42026
rect 49608 40724 49660 40730
rect 49608 40666 49660 40672
rect 45468 17264 45520 17270
rect 45468 17206 45520 17212
rect 43352 4072 43404 4078
rect 43352 4014 43404 4020
rect 42156 3392 42208 3398
rect 42156 3334 42208 3340
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 42168 480 42196 3334
rect 43364 480 43392 4014
rect 45480 3330 45508 17206
rect 48136 4956 48188 4962
rect 48136 4898 48188 4904
rect 45744 4140 45796 4146
rect 45744 4082 45796 4088
rect 44548 3324 44600 3330
rect 44548 3266 44600 3272
rect 45468 3324 45520 3330
rect 45468 3266 45520 3272
rect 44560 480 44588 3266
rect 45756 480 45784 4082
rect 46940 3324 46992 3330
rect 46940 3266 46992 3272
rect 46952 480 46980 3266
rect 48148 480 48176 4898
rect 49620 3482 49648 40666
rect 49344 3454 49648 3482
rect 49344 480 49372 3454
rect 51000 3398 51028 49166
rect 53748 39364 53800 39370
rect 53748 39306 53800 39312
rect 51632 5024 51684 5030
rect 51632 4966 51684 4972
rect 50528 3392 50580 3398
rect 50528 3334 50580 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 50540 480 50568 3334
rect 51644 480 51672 4966
rect 53760 3398 53788 39306
rect 56416 37936 56468 37942
rect 56416 37878 56468 37884
rect 55220 5160 55272 5166
rect 55220 5102 55272 5108
rect 52828 3392 52880 3398
rect 52828 3334 52880 3340
rect 53748 3392 53800 3398
rect 53748 3334 53800 3340
rect 52840 480 52868 3334
rect 54024 3324 54076 3330
rect 54024 3266 54076 3272
rect 54036 480 54064 3266
rect 55232 480 55260 5102
rect 56428 480 56456 37878
rect 57900 3482 57928 49234
rect 60016 9654 60044 59055
rect 60108 26246 60136 73335
rect 60200 42770 60228 87615
rect 60292 59362 60320 101895
rect 523696 71738 523724 111959
rect 523788 86970 523816 125287
rect 523880 102134 523908 138615
rect 580172 133884 580224 133890
rect 580172 133826 580224 133832
rect 580184 132977 580212 133826
rect 580170 132968 580226 132977
rect 580170 132903 580226 132912
rect 580172 118652 580224 118658
rect 580172 118594 580224 118600
rect 580184 117337 580212 118594
rect 580170 117328 580226 117337
rect 580170 117263 580226 117272
rect 523868 102128 523920 102134
rect 523868 102070 523920 102076
rect 580172 102128 580224 102134
rect 580172 102070 580224 102076
rect 580184 101697 580212 102070
rect 580170 101688 580226 101697
rect 580170 101623 580226 101632
rect 523958 98696 524014 98705
rect 523958 98631 524014 98640
rect 523776 86964 523828 86970
rect 523776 86906 523828 86912
rect 523866 85368 523922 85377
rect 523866 85303 523922 85312
rect 523774 72040 523830 72049
rect 523774 71975 523830 71984
rect 523684 71732 523736 71738
rect 523684 71674 523736 71680
rect 60280 59356 60332 59362
rect 60280 59298 60332 59304
rect 523682 58712 523738 58721
rect 523682 58647 523738 58656
rect 75012 52142 75578 52170
rect 150912 52142 151662 52170
rect 168760 52142 169510 52170
rect 189368 52142 190118 52170
rect 197924 52142 198582 52170
rect 296194 52142 296668 52170
rect 62500 48346 62528 52020
rect 63144 52006 63434 52034
rect 63512 52006 64354 52034
rect 61384 48340 61436 48346
rect 61384 48282 61436 48288
rect 62488 48340 62540 48346
rect 62488 48282 62540 48288
rect 60188 42764 60240 42770
rect 60188 42706 60240 42712
rect 60096 26240 60148 26246
rect 60096 26182 60148 26188
rect 60648 21412 60700 21418
rect 60648 21354 60700 21360
rect 60004 9648 60056 9654
rect 60004 9590 60056 9596
rect 58808 5092 58860 5098
rect 58808 5034 58860 5040
rect 57624 3454 57928 3482
rect 57624 480 57652 3454
rect 58820 480 58848 5034
rect 60660 3466 60688 21354
rect 61396 6186 61424 48282
rect 63144 41410 63172 52006
rect 62396 41404 62448 41410
rect 62396 41346 62448 41352
rect 63132 41404 63184 41410
rect 63132 41346 63184 41352
rect 62408 31770 62436 41346
rect 62224 31742 62436 31770
rect 62224 31634 62252 31742
rect 62224 31606 62344 31634
rect 62316 28966 62344 31606
rect 62304 28960 62356 28966
rect 62304 28902 62356 28908
rect 62488 19372 62540 19378
rect 62488 19314 62540 19320
rect 62500 7614 62528 19314
rect 63512 10334 63540 52006
rect 64788 49360 64840 49366
rect 64788 49302 64840 49308
rect 64696 19984 64748 19990
rect 64696 19926 64748 19932
rect 63500 10328 63552 10334
rect 63500 10270 63552 10276
rect 62488 7608 62540 7614
rect 62488 7550 62540 7556
rect 61384 6180 61436 6186
rect 61384 6122 61436 6128
rect 62396 6180 62448 6186
rect 62396 6122 62448 6128
rect 60004 3460 60056 3466
rect 60004 3402 60056 3408
rect 60648 3460 60700 3466
rect 60648 3402 60700 3408
rect 60016 480 60044 3402
rect 61200 3256 61252 3262
rect 61200 3198 61252 3204
rect 61212 480 61240 3198
rect 62408 480 62436 6122
rect 64708 3602 64736 19926
rect 63592 3596 63644 3602
rect 63592 3538 63644 3544
rect 64696 3596 64748 3602
rect 64696 3538 64748 3544
rect 63604 480 63632 3538
rect 64800 480 64828 49302
rect 65260 47598 65288 52020
rect 66180 49094 66208 52020
rect 66364 52006 67206 52034
rect 67652 52006 68126 52034
rect 69046 52006 69152 52034
rect 66168 49088 66220 49094
rect 66168 49030 66220 49036
rect 65248 47592 65300 47598
rect 65248 47534 65300 47540
rect 65984 7608 66036 7614
rect 65984 7550 66036 7556
rect 65996 480 66024 7550
rect 66364 3194 66392 52006
rect 67548 24132 67600 24138
rect 67548 24074 67600 24080
rect 66352 3188 66404 3194
rect 66352 3130 66404 3136
rect 67560 626 67588 24074
rect 67652 11762 67680 52006
rect 69124 18630 69152 52006
rect 69952 49162 69980 52020
rect 70504 52006 70886 52034
rect 71792 52006 71898 52034
rect 72068 52006 72818 52034
rect 73172 52006 73738 52034
rect 69940 49156 69992 49162
rect 69940 49098 69992 49104
rect 70308 47592 70360 47598
rect 70308 47534 70360 47540
rect 69112 18624 69164 18630
rect 69112 18566 69164 18572
rect 67640 11756 67692 11762
rect 67640 11698 67692 11704
rect 70320 3534 70348 47534
rect 70504 3602 70532 52006
rect 71688 18624 71740 18630
rect 71688 18566 71740 18572
rect 71700 3670 71728 18566
rect 71792 4826 71820 52006
rect 72068 36582 72096 52006
rect 72056 36576 72108 36582
rect 72056 36518 72108 36524
rect 71780 4820 71832 4826
rect 71780 4762 71832 4768
rect 73068 4820 73120 4826
rect 73068 4762 73120 4768
rect 70676 3664 70728 3670
rect 70676 3606 70728 3612
rect 71688 3664 71740 3670
rect 71688 3606 71740 3612
rect 70492 3596 70544 3602
rect 70492 3538 70544 3544
rect 69480 3528 69532 3534
rect 69480 3470 69532 3476
rect 70308 3528 70360 3534
rect 70308 3470 70360 3476
rect 68284 3460 68336 3466
rect 68284 3402 68336 3408
rect 67192 598 67588 626
rect 67192 480 67220 598
rect 68296 480 68324 3402
rect 69492 480 69520 3470
rect 70688 480 70716 3606
rect 71872 3188 71924 3194
rect 71872 3130 71924 3136
rect 71884 480 71912 3130
rect 73080 480 73108 4762
rect 73172 3126 73200 52006
rect 74644 49026 74672 52020
rect 75012 51218 75040 52142
rect 74920 51190 75040 51218
rect 75932 52006 76590 52034
rect 74632 49020 74684 49026
rect 74632 48962 74684 48968
rect 74920 38690 74948 51190
rect 74724 38684 74776 38690
rect 74724 38626 74776 38632
rect 74908 38684 74960 38690
rect 74908 38626 74960 38632
rect 74448 25560 74500 25566
rect 74448 25502 74500 25508
rect 73160 3120 73212 3126
rect 73160 3062 73212 3068
rect 74460 610 74488 25502
rect 74736 22370 74764 38626
rect 75932 35222 75960 52006
rect 77392 46232 77444 46238
rect 77392 46174 77444 46180
rect 75920 35216 75972 35222
rect 75920 35158 75972 35164
rect 74724 22364 74776 22370
rect 74724 22306 74776 22312
rect 74724 19372 74776 19378
rect 74724 19314 74776 19320
rect 74736 4894 74764 19314
rect 76656 8968 76708 8974
rect 76656 8910 76708 8916
rect 74724 4888 74776 4894
rect 74724 4830 74776 4836
rect 75460 3596 75512 3602
rect 75460 3538 75512 3544
rect 74264 604 74316 610
rect 74264 546 74316 552
rect 74448 604 74500 610
rect 74448 546 74500 552
rect 74276 480 74304 546
rect 75472 480 75500 3538
rect 76668 480 76696 8910
rect 77404 3670 77432 46174
rect 77392 3664 77444 3670
rect 77392 3606 77444 3612
rect 77496 3369 77524 52020
rect 78048 52006 78430 52034
rect 78968 52006 79350 52034
rect 78048 46238 78076 52006
rect 78036 46232 78088 46238
rect 78036 46174 78088 46180
rect 78968 46170 78996 52006
rect 79968 49020 80020 49026
rect 79968 48962 80020 48968
rect 79324 48816 79376 48822
rect 79324 48758 79376 48764
rect 78956 46164 79008 46170
rect 78956 46106 79008 46112
rect 78588 26920 78640 26926
rect 78588 26862 78640 26868
rect 78600 3670 78628 26862
rect 79336 22778 79364 48758
rect 79324 22772 79376 22778
rect 79324 22714 79376 22720
rect 77852 3664 77904 3670
rect 77852 3606 77904 3612
rect 78588 3664 78640 3670
rect 78588 3606 78640 3612
rect 77482 3360 77538 3369
rect 77482 3295 77538 3304
rect 77864 480 77892 3606
rect 79980 882 80008 48962
rect 80256 48822 80284 52020
rect 80992 52006 81282 52034
rect 81544 52006 82202 52034
rect 82924 52006 83122 52034
rect 83752 52006 84042 52034
rect 84212 52006 84962 52034
rect 85592 52006 85974 52034
rect 86512 52006 86894 52034
rect 86972 52006 87814 52034
rect 88444 52006 88734 52034
rect 89272 52006 89654 52034
rect 89732 52006 90666 52034
rect 91112 52006 91586 52034
rect 92506 52006 92612 52034
rect 80244 48816 80296 48822
rect 80244 48758 80296 48764
rect 80992 46050 81020 52006
rect 80256 46022 81020 46050
rect 80256 27674 80284 46022
rect 80152 27668 80204 27674
rect 80152 27610 80204 27616
rect 80244 27668 80296 27674
rect 80244 27610 80296 27616
rect 80164 19281 80192 27610
rect 80150 19272 80206 19281
rect 80150 19207 80206 19216
rect 80426 19272 80482 19281
rect 80426 19207 80482 19216
rect 80440 12442 80468 19207
rect 80060 12436 80112 12442
rect 80060 12378 80112 12384
rect 80428 12436 80480 12442
rect 80428 12378 80480 12384
rect 80072 9602 80100 12378
rect 80244 10328 80296 10334
rect 80244 10270 80296 10276
rect 80072 9574 80192 9602
rect 80164 3738 80192 9574
rect 80152 3732 80204 3738
rect 80152 3674 80204 3680
rect 79048 876 79100 882
rect 79048 818 79100 824
rect 79968 876 80020 882
rect 79968 818 80020 824
rect 79060 480 79088 818
rect 80256 480 80284 10270
rect 81544 3505 81572 52006
rect 82924 44878 82952 52006
rect 82912 44872 82964 44878
rect 82912 44814 82964 44820
rect 83752 38690 83780 52006
rect 82820 38684 82872 38690
rect 82820 38626 82872 38632
rect 83740 38684 83792 38690
rect 83740 38626 83792 38632
rect 82832 33794 82860 38626
rect 82820 33788 82872 33794
rect 82820 33730 82872 33736
rect 82728 28280 82780 28286
rect 82728 28222 82780 28228
rect 81530 3496 81586 3505
rect 81530 3431 81586 3440
rect 82634 3360 82690 3369
rect 82634 3295 82690 3304
rect 81440 3120 81492 3126
rect 81440 3062 81492 3068
rect 81452 480 81480 3062
rect 82648 480 82676 3295
rect 82740 3126 82768 28222
rect 84108 11756 84160 11762
rect 84108 11698 84160 11704
rect 82728 3120 82780 3126
rect 82728 3062 82780 3068
rect 84120 610 84148 11698
rect 84212 3806 84240 52006
rect 85488 29708 85540 29714
rect 85488 29650 85540 29656
rect 85500 3874 85528 29650
rect 85592 13122 85620 52006
rect 86512 43518 86540 52006
rect 86500 43512 86552 43518
rect 86500 43454 86552 43460
rect 85764 38684 85816 38690
rect 85764 38626 85816 38632
rect 85776 32434 85804 38626
rect 85764 32428 85816 32434
rect 85764 32370 85816 32376
rect 85580 13116 85632 13122
rect 85580 13058 85632 13064
rect 84936 3868 84988 3874
rect 84936 3810 84988 3816
rect 85488 3868 85540 3874
rect 85488 3810 85540 3816
rect 84200 3800 84252 3806
rect 84200 3742 84252 3748
rect 83832 604 83884 610
rect 83832 546 83884 552
rect 84108 604 84160 610
rect 84108 546 84160 552
rect 83844 480 83872 546
rect 84948 480 84976 3810
rect 86972 3806 87000 52006
rect 88248 46232 88300 46238
rect 88248 46174 88300 46180
rect 86960 3800 87012 3806
rect 86960 3742 87012 3748
rect 86130 3496 86186 3505
rect 86130 3431 86186 3440
rect 86144 480 86172 3431
rect 88260 2922 88288 46174
rect 88444 43450 88472 52006
rect 88432 43444 88484 43450
rect 88432 43386 88484 43392
rect 89272 42922 89300 52006
rect 88352 42894 89300 42922
rect 88352 31074 88380 42894
rect 88340 31068 88392 31074
rect 88340 31010 88392 31016
rect 89628 31068 89680 31074
rect 89628 31010 89680 31016
rect 89640 3874 89668 31010
rect 89732 4010 89760 52006
rect 91008 22772 91060 22778
rect 91008 22714 91060 22720
rect 89720 4004 89772 4010
rect 89720 3946 89772 3952
rect 88524 3868 88576 3874
rect 88524 3810 88576 3816
rect 89628 3868 89680 3874
rect 89628 3810 89680 3816
rect 87328 2916 87380 2922
rect 87328 2858 87380 2864
rect 88248 2916 88300 2922
rect 88248 2858 88300 2864
rect 87340 480 87368 2858
rect 88536 480 88564 3810
rect 89720 3596 89772 3602
rect 89720 3538 89772 3544
rect 89732 480 89760 3538
rect 91020 592 91048 22714
rect 91112 14482 91140 52006
rect 92480 48816 92532 48822
rect 92480 48758 92532 48764
rect 92388 44872 92440 44878
rect 92388 44814 92440 44820
rect 91100 14476 91152 14482
rect 91100 14418 91152 14424
rect 92400 626 92428 44814
rect 92492 3942 92520 48758
rect 92584 29646 92612 52006
rect 93136 52006 93426 52034
rect 93872 52006 94346 52034
rect 93136 48822 93164 52006
rect 93124 48816 93176 48822
rect 93124 48758 93176 48764
rect 92572 29640 92624 29646
rect 92572 29582 92624 29588
rect 93872 15910 93900 52006
rect 95240 48816 95292 48822
rect 95240 48758 95292 48764
rect 93860 15904 93912 15910
rect 93860 15846 93912 15852
rect 95148 13116 95200 13122
rect 95148 13058 95200 13064
rect 92480 3936 92532 3942
rect 92480 3878 92532 3884
rect 93308 3664 93360 3670
rect 93308 3606 93360 3612
rect 92216 598 92428 626
rect 92216 592 92244 598
rect 90928 564 91048 592
rect 92124 564 92244 592
rect 90928 480 90956 564
rect 92124 480 92152 564
rect 93320 480 93348 3606
rect 95160 2922 95188 13058
rect 95252 3874 95280 48758
rect 95344 42090 95372 52020
rect 95896 52006 96278 52034
rect 96632 52006 97198 52034
rect 98012 52006 98118 52034
rect 98288 52006 99038 52034
rect 99392 52006 100050 52034
rect 100864 52006 100970 52034
rect 95896 48822 95924 52006
rect 95884 48816 95936 48822
rect 95884 48758 95936 48764
rect 95332 42084 95384 42090
rect 95332 42026 95384 42032
rect 96528 32428 96580 32434
rect 96528 32370 96580 32376
rect 95240 3868 95292 3874
rect 95240 3810 95292 3816
rect 96540 3398 96568 32370
rect 96632 17270 96660 52006
rect 96620 17264 96672 17270
rect 96620 17206 96672 17212
rect 98012 4146 98040 52006
rect 98288 35970 98316 52006
rect 98092 35964 98144 35970
rect 98092 35906 98144 35912
rect 98276 35964 98328 35970
rect 98276 35906 98328 35912
rect 98104 26194 98132 35906
rect 98104 26166 98316 26194
rect 98288 16658 98316 26166
rect 98092 16652 98144 16658
rect 98092 16594 98144 16600
rect 98276 16652 98328 16658
rect 98276 16594 98328 16600
rect 98104 6882 98132 16594
rect 99288 14476 99340 14482
rect 99288 14418 99340 14424
rect 98104 6854 98316 6882
rect 98000 4140 98052 4146
rect 98000 4082 98052 4088
rect 96896 3800 96948 3806
rect 96896 3742 96948 3748
rect 95700 3392 95752 3398
rect 95700 3334 95752 3340
rect 96528 3392 96580 3398
rect 96528 3334 96580 3340
rect 94504 2916 94556 2922
rect 94504 2858 94556 2864
rect 95148 2916 95200 2922
rect 95148 2858 95200 2864
rect 94516 480 94544 2858
rect 95712 480 95740 3334
rect 96908 480 96936 3742
rect 98288 3738 98316 6854
rect 99196 3868 99248 3874
rect 99196 3810 99248 3816
rect 98276 3732 98328 3738
rect 98276 3674 98328 3680
rect 98092 3392 98144 3398
rect 98092 3334 98144 3340
rect 98104 480 98132 3334
rect 99208 1986 99236 3810
rect 99300 3398 99328 14418
rect 99392 4962 99420 52006
rect 100864 40730 100892 52006
rect 101876 49230 101904 52020
rect 102152 52006 102810 52034
rect 103624 52006 103730 52034
rect 104360 52006 104742 52034
rect 104912 52006 105662 52034
rect 106384 52006 106582 52034
rect 101864 49224 101916 49230
rect 101864 49166 101916 49172
rect 100852 40724 100904 40730
rect 100852 40666 100904 40672
rect 102048 15904 102100 15910
rect 102048 15846 102100 15852
rect 99380 4956 99432 4962
rect 99380 4898 99432 4904
rect 100484 3732 100536 3738
rect 100484 3674 100536 3680
rect 99288 3392 99340 3398
rect 99288 3334 99340 3340
rect 99208 1958 99328 1986
rect 99300 480 99328 1958
rect 100496 480 100524 3674
rect 102060 3398 102088 15846
rect 102152 5030 102180 52006
rect 103428 49088 103480 49094
rect 103428 49030 103480 49036
rect 102140 5024 102192 5030
rect 102140 4966 102192 4972
rect 103440 3398 103468 49030
rect 103520 48816 103572 48822
rect 103520 48758 103572 48764
rect 101588 3392 101640 3398
rect 101588 3334 101640 3340
rect 102048 3392 102100 3398
rect 102048 3334 102100 3340
rect 102784 3392 102836 3398
rect 102784 3334 102836 3340
rect 103428 3392 103480 3398
rect 103428 3334 103480 3340
rect 101600 480 101628 3334
rect 102796 480 102824 3334
rect 103532 3330 103560 48758
rect 103624 39370 103652 52006
rect 104360 48822 104388 52006
rect 104348 48816 104400 48822
rect 104348 48758 104400 48764
rect 103612 39364 103664 39370
rect 103612 39306 103664 39312
rect 104912 5166 104940 52006
rect 106188 42084 106240 42090
rect 106188 42026 106240 42032
rect 104900 5160 104952 5166
rect 104900 5102 104952 5108
rect 103980 3936 104032 3942
rect 103980 3878 104032 3884
rect 103520 3324 103572 3330
rect 103520 3266 103572 3272
rect 103992 480 104020 3878
rect 106200 3398 106228 42026
rect 106384 37942 106412 52006
rect 107488 49298 107516 52020
rect 107672 52006 108514 52034
rect 107476 49292 107528 49298
rect 107476 49234 107528 49240
rect 107568 49156 107620 49162
rect 107568 49098 107620 49104
rect 106372 37936 106424 37942
rect 106372 37878 106424 37884
rect 106372 4140 106424 4146
rect 106372 4082 106424 4088
rect 105176 3392 105228 3398
rect 105176 3334 105228 3340
rect 106188 3392 106240 3398
rect 106188 3334 106240 3340
rect 105188 480 105216 3334
rect 106384 480 106412 4082
rect 107580 480 107608 49098
rect 107672 5098 107700 52006
rect 109420 48822 109448 52020
rect 110064 52006 110354 52034
rect 110432 52006 111274 52034
rect 108304 48816 108356 48822
rect 108304 48758 108356 48764
rect 109408 48816 109460 48822
rect 109408 48758 109460 48764
rect 108316 21418 108344 48758
rect 110064 38865 110092 52006
rect 110050 38856 110106 38865
rect 110050 38791 110106 38800
rect 109314 38720 109370 38729
rect 109370 38678 109448 38706
rect 109314 38655 109370 38664
rect 109420 38622 109448 38678
rect 109408 38616 109460 38622
rect 109408 38558 109460 38564
rect 109500 29028 109552 29034
rect 109500 28970 109552 28976
rect 109512 22250 109540 28970
rect 109420 22222 109540 22250
rect 108304 21412 108356 21418
rect 108304 21354 108356 21360
rect 108948 21412 109000 21418
rect 108948 21354 109000 21360
rect 107660 5092 107712 5098
rect 107660 5034 107712 5040
rect 108960 626 108988 21354
rect 109420 19378 109448 22222
rect 109316 19372 109368 19378
rect 109316 19314 109368 19320
rect 109408 19372 109460 19378
rect 109408 19314 109460 19320
rect 109328 12458 109356 19314
rect 109328 12430 109448 12458
rect 109420 3262 109448 12430
rect 110432 6186 110460 52006
rect 112180 48346 112208 52020
rect 113192 49366 113220 52020
rect 113284 52006 114126 52034
rect 114572 52006 115046 52034
rect 115966 52006 116164 52034
rect 113180 49360 113232 49366
rect 113180 49302 113232 49308
rect 111064 48340 111116 48346
rect 111064 48282 111116 48288
rect 112168 48340 112220 48346
rect 112168 48282 112220 48288
rect 111076 19990 111104 48282
rect 111064 19984 111116 19990
rect 111064 19926 111116 19932
rect 113284 7614 113312 52006
rect 114572 24138 114600 52006
rect 115848 49224 115900 49230
rect 115848 49166 115900 49172
rect 114560 24132 114612 24138
rect 114560 24074 114612 24080
rect 113272 7608 113324 7614
rect 113272 7550 113324 7556
rect 110420 6180 110472 6186
rect 110420 6122 110472 6128
rect 112352 6180 112404 6186
rect 112352 6122 112404 6128
rect 109960 4072 110012 4078
rect 109960 4014 110012 4020
rect 109408 3256 109460 3262
rect 109408 3198 109460 3204
rect 108776 598 108988 626
rect 108776 480 108804 598
rect 109972 480 110000 4014
rect 111156 4004 111208 4010
rect 111156 3946 111208 3952
rect 111168 480 111196 3946
rect 112364 480 112392 6122
rect 113548 3392 113600 3398
rect 113548 3334 113600 3340
rect 113560 480 113588 3334
rect 115860 3262 115888 49166
rect 115940 7608 115992 7614
rect 115940 7550 115992 7556
rect 114744 3256 114796 3262
rect 114744 3198 114796 3204
rect 115848 3256 115900 3262
rect 115848 3198 115900 3204
rect 114756 480 114784 3198
rect 115952 480 115980 7550
rect 116136 3466 116164 52006
rect 116872 47598 116900 52020
rect 117332 52006 117898 52034
rect 118818 52006 118924 52034
rect 116860 47592 116912 47598
rect 116860 47534 116912 47540
rect 117332 18630 117360 52006
rect 118792 46300 118844 46306
rect 118792 46242 118844 46248
rect 117320 18624 117372 18630
rect 117320 18566 117372 18572
rect 118804 4826 118832 46242
rect 118792 4820 118844 4826
rect 118792 4762 118844 4768
rect 116124 3460 116176 3466
rect 116124 3402 116176 3408
rect 118240 3460 118292 3466
rect 118240 3402 118292 3408
rect 117136 3324 117188 3330
rect 117136 3266 117188 3272
rect 117148 480 117176 3266
rect 118252 480 118280 3402
rect 118896 3126 118924 52006
rect 119448 52006 119738 52034
rect 120092 52006 120658 52034
rect 119448 46306 119476 52006
rect 119436 46300 119488 46306
rect 119436 46242 119488 46248
rect 120092 25566 120120 52006
rect 120724 48340 120776 48346
rect 120724 48282 120776 48288
rect 120080 25560 120132 25566
rect 120080 25502 120132 25508
rect 119436 9036 119488 9042
rect 119436 8978 119488 8984
rect 118884 3120 118936 3126
rect 118884 3062 118936 3068
rect 119448 480 119476 8978
rect 120736 8974 120764 48282
rect 120724 8968 120776 8974
rect 120724 8910 120776 8916
rect 120632 3256 120684 3262
rect 120632 3198 120684 3204
rect 120644 480 120672 3198
rect 121564 3194 121592 52020
rect 122576 48346 122604 52020
rect 122852 52006 123510 52034
rect 122748 49292 122800 49298
rect 122748 49234 122800 49240
rect 122564 48340 122616 48346
rect 122564 48282 122616 48288
rect 122760 3602 122788 49234
rect 122852 26926 122880 52006
rect 124416 49026 124444 52020
rect 124876 52006 125350 52034
rect 125612 52006 126270 52034
rect 127084 52006 127282 52034
rect 124404 49020 124456 49026
rect 124404 48962 124456 48968
rect 124876 46050 124904 52006
rect 125508 49020 125560 49026
rect 125508 48962 125560 48968
rect 124232 46022 124904 46050
rect 124232 41410 124260 46022
rect 124220 41404 124272 41410
rect 124220 41346 124272 41352
rect 124404 41404 124456 41410
rect 124404 41346 124456 41352
rect 124416 38622 124444 41346
rect 124404 38616 124456 38622
rect 124404 38558 124456 38564
rect 124312 29028 124364 29034
rect 124312 28970 124364 28976
rect 122840 26920 122892 26926
rect 122840 26862 122892 26868
rect 124128 26920 124180 26926
rect 124128 26862 124180 26868
rect 124140 3602 124168 26862
rect 124324 22166 124352 28970
rect 124312 22160 124364 22166
rect 124312 22102 124364 22108
rect 124312 22024 124364 22030
rect 124312 21966 124364 21972
rect 124324 12458 124352 21966
rect 124324 12430 124444 12458
rect 124416 10334 124444 12430
rect 124404 10328 124456 10334
rect 124404 10270 124456 10276
rect 125520 3602 125548 48962
rect 125612 28286 125640 52006
rect 126244 48340 126296 48346
rect 126244 48282 126296 48288
rect 125600 28280 125652 28286
rect 125600 28222 125652 28228
rect 126256 11762 126284 48282
rect 126244 11756 126296 11762
rect 126244 11698 126296 11704
rect 126612 4820 126664 4826
rect 126612 4762 126664 4768
rect 121828 3596 121880 3602
rect 121828 3538 121880 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 123024 3596 123076 3602
rect 123024 3538 123076 3544
rect 124128 3596 124180 3602
rect 124128 3538 124180 3544
rect 124220 3596 124272 3602
rect 124220 3538 124272 3544
rect 125508 3596 125560 3602
rect 125508 3538 125560 3544
rect 121552 3188 121604 3194
rect 121552 3130 121604 3136
rect 121840 480 121868 3538
rect 123036 480 123064 3538
rect 124232 480 124260 3538
rect 125416 3528 125468 3534
rect 125416 3470 125468 3476
rect 125428 480 125456 3470
rect 126624 480 126652 4762
rect 127084 3369 127112 52006
rect 128188 48346 128216 52020
rect 128372 52006 129122 52034
rect 129936 52006 130042 52034
rect 128176 48340 128228 48346
rect 128176 48282 128228 48288
rect 128372 29714 128400 52006
rect 129648 43444 129700 43450
rect 129648 43386 129700 43392
rect 128360 29708 128412 29714
rect 128360 29650 128412 29656
rect 128268 17264 128320 17270
rect 128268 17206 128320 17212
rect 128280 3534 128308 17206
rect 129660 3534 129688 43386
rect 127808 3528 127860 3534
rect 127808 3470 127860 3476
rect 128268 3528 128320 3534
rect 128268 3470 128320 3476
rect 129004 3528 129056 3534
rect 129004 3470 129056 3476
rect 129648 3528 129700 3534
rect 129936 3505 129964 52006
rect 130948 46238 130976 52020
rect 131132 52006 131974 52034
rect 132512 52006 132894 52034
rect 133432 52006 133814 52034
rect 133892 52006 134734 52034
rect 135272 52006 135654 52034
rect 130936 46232 130988 46238
rect 130936 46174 130988 46180
rect 131132 31074 131160 52006
rect 132408 46232 132460 46238
rect 132408 46174 132460 46180
rect 131120 31068 131172 31074
rect 131120 31010 131172 31016
rect 130200 6248 130252 6254
rect 130200 6190 130252 6196
rect 129648 3470 129700 3476
rect 129922 3496 129978 3505
rect 127070 3360 127126 3369
rect 127070 3295 127126 3304
rect 127820 480 127848 3470
rect 129016 480 129044 3470
rect 129922 3431 129978 3440
rect 130212 480 130240 6190
rect 132420 3602 132448 46174
rect 131396 3596 131448 3602
rect 131396 3538 131448 3544
rect 132408 3596 132460 3602
rect 132408 3538 132460 3544
rect 131408 480 131436 3538
rect 132512 3194 132540 52006
rect 133432 38690 133460 52006
rect 133892 44878 133920 52006
rect 133880 44872 133932 44878
rect 133880 44814 133932 44820
rect 132868 38684 132920 38690
rect 132868 38626 132920 38632
rect 133420 38684 133472 38690
rect 133420 38626 133472 38632
rect 132880 22778 132908 38626
rect 132868 22772 132920 22778
rect 132868 22714 132920 22720
rect 133788 22772 133840 22778
rect 133788 22714 133840 22720
rect 133696 7676 133748 7682
rect 133696 7618 133748 7624
rect 132592 3596 132644 3602
rect 132592 3538 132644 3544
rect 132500 3188 132552 3194
rect 132500 3130 132552 3136
rect 132604 480 132632 3538
rect 133708 1578 133736 7618
rect 133800 3602 133828 22714
rect 135168 18624 135220 18630
rect 135168 18566 135220 18572
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 133708 1550 133828 1578
rect 133800 480 133828 1550
rect 135180 626 135208 18566
rect 135272 3670 135300 52006
rect 136548 24132 136600 24138
rect 136548 24074 136600 24080
rect 135260 3664 135312 3670
rect 135260 3606 135312 3612
rect 136560 3602 136588 24074
rect 136652 13122 136680 52020
rect 136744 52006 137586 52034
rect 138032 52006 138506 52034
rect 139426 52006 139532 52034
rect 136744 32434 136772 52006
rect 136732 32428 136784 32434
rect 136732 32370 136784 32376
rect 136640 13116 136692 13122
rect 136640 13058 136692 13064
rect 137284 8968 137336 8974
rect 137284 8910 137336 8916
rect 136088 3596 136140 3602
rect 136088 3538 136140 3544
rect 136548 3596 136600 3602
rect 136548 3538 136600 3544
rect 134904 598 135208 626
rect 134904 480 134932 598
rect 136100 480 136128 3538
rect 137296 480 137324 8910
rect 138032 3806 138060 52006
rect 139400 48816 139452 48822
rect 139400 48758 139452 48764
rect 139308 44872 139360 44878
rect 139308 44814 139360 44820
rect 138020 3800 138072 3806
rect 138020 3742 138072 3748
rect 139320 3058 139348 44814
rect 139412 3874 139440 48758
rect 139504 14482 139532 52006
rect 140056 52006 140346 52034
rect 140792 52006 141358 52034
rect 140056 48822 140084 52006
rect 140044 48816 140096 48822
rect 140044 48758 140096 48764
rect 140688 25560 140740 25566
rect 140688 25502 140740 25508
rect 139492 14476 139544 14482
rect 139492 14418 139544 14424
rect 139400 3868 139452 3874
rect 139400 3810 139452 3816
rect 140700 3602 140728 25502
rect 140792 3738 140820 52006
rect 142068 19984 142120 19990
rect 142068 19926 142120 19932
rect 141976 10328 142028 10334
rect 141976 10270 142028 10276
rect 140780 3732 140832 3738
rect 140780 3674 140832 3680
rect 141988 3602 142016 10270
rect 139676 3596 139728 3602
rect 139676 3538 139728 3544
rect 140688 3596 140740 3602
rect 140688 3538 140740 3544
rect 140872 3596 140924 3602
rect 140872 3538 140924 3544
rect 141976 3596 142028 3602
rect 141976 3538 142028 3544
rect 138480 3052 138532 3058
rect 138480 2994 138532 3000
rect 139308 3052 139360 3058
rect 139308 2994 139360 3000
rect 138492 480 138520 2994
rect 139688 480 139716 3538
rect 140884 480 140912 3538
rect 142080 480 142108 19926
rect 142264 15910 142292 52020
rect 143184 49094 143212 52020
rect 143552 52006 144118 52034
rect 143172 49088 143224 49094
rect 143172 49030 143224 49036
rect 142252 15904 142304 15910
rect 142252 15846 142304 15852
rect 143552 3670 143580 52006
rect 144920 48816 144972 48822
rect 144920 48758 144972 48764
rect 144828 11756 144880 11762
rect 144828 11698 144880 11704
rect 143540 3664 143592 3670
rect 143540 3606 143592 3612
rect 143264 3596 143316 3602
rect 143264 3538 143316 3544
rect 143276 480 143304 3538
rect 144840 626 144868 11698
rect 144932 4146 144960 48758
rect 145024 42090 145052 52020
rect 145760 52006 146050 52034
rect 145760 48822 145788 52006
rect 146956 49162 146984 52020
rect 147772 51060 147824 51066
rect 147772 51002 147824 51008
rect 146944 49156 146996 49162
rect 146944 49098 146996 49104
rect 145748 48816 145800 48822
rect 145748 48758 145800 48764
rect 146944 48816 146996 48822
rect 146944 48758 146996 48764
rect 145012 42084 145064 42090
rect 145012 42026 145064 42032
rect 146208 21480 146260 21486
rect 146208 21422 146260 21428
rect 144920 4140 144972 4146
rect 144920 4082 144972 4088
rect 146220 3602 146248 21422
rect 146956 21418 146984 48758
rect 147784 31770 147812 51002
rect 147876 48822 147904 52020
rect 148060 52006 148810 52034
rect 149072 52006 149730 52034
rect 150544 52006 150742 52034
rect 148060 51066 148088 52006
rect 148048 51060 148100 51066
rect 148048 51002 148100 51008
rect 147864 48816 147916 48822
rect 147864 48758 147916 48764
rect 147784 31742 147904 31770
rect 146944 21412 146996 21418
rect 146944 21354 146996 21360
rect 147876 19310 147904 31742
rect 147864 19304 147916 19310
rect 147864 19246 147916 19252
rect 148968 13116 149020 13122
rect 148968 13058 149020 13064
rect 147772 9716 147824 9722
rect 147772 9658 147824 9664
rect 147784 4078 147812 9658
rect 147772 4072 147824 4078
rect 147772 4014 147824 4020
rect 146852 3732 146904 3738
rect 146852 3674 146904 3680
rect 145656 3596 145708 3602
rect 145656 3538 145708 3544
rect 146208 3596 146260 3602
rect 146208 3538 146260 3544
rect 144472 598 144868 626
rect 144472 480 144500 598
rect 145668 480 145696 3538
rect 146864 480 146892 3674
rect 148980 3534 149008 13058
rect 149072 4010 149100 52006
rect 150544 6186 150572 52006
rect 150912 26314 150940 52142
rect 152568 49230 152596 52020
rect 153304 52006 153502 52034
rect 154224 52006 154514 52034
rect 154684 52006 155434 52034
rect 156064 52006 156354 52034
rect 156984 52006 157274 52034
rect 152556 49224 152608 49230
rect 152556 49166 152608 49172
rect 153200 46300 153252 46306
rect 153200 46242 153252 46248
rect 150808 26308 150860 26314
rect 150808 26250 150860 26256
rect 150900 26308 150952 26314
rect 150900 26250 150952 26256
rect 150820 26194 150848 26250
rect 150636 26166 150848 26194
rect 150636 22166 150664 26166
rect 150624 22160 150676 22166
rect 150624 22102 150676 22108
rect 151728 14476 151780 14482
rect 151728 14418 151780 14424
rect 150808 9716 150860 9722
rect 150808 9658 150860 9664
rect 150532 6180 150584 6186
rect 150532 6122 150584 6128
rect 149060 4004 149112 4010
rect 149060 3946 149112 3952
rect 150440 3936 150492 3942
rect 150440 3878 150492 3884
rect 149244 3664 149296 3670
rect 149244 3606 149296 3612
rect 148048 3528 148100 3534
rect 148048 3470 148100 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 148060 480 148088 3470
rect 149256 480 149284 3606
rect 150452 480 150480 3878
rect 150820 3398 150848 9658
rect 150808 3392 150860 3398
rect 150808 3334 150860 3340
rect 151740 610 151768 14418
rect 152740 3392 152792 3398
rect 152740 3334 152792 3340
rect 151544 604 151596 610
rect 151544 546 151596 552
rect 151728 604 151780 610
rect 151728 546 151780 552
rect 151556 480 151584 546
rect 152752 480 152780 3334
rect 153212 3330 153240 46242
rect 153304 7614 153332 52006
rect 154224 46306 154252 52006
rect 154212 46300 154264 46306
rect 154212 46242 154264 46248
rect 153292 7608 153344 7614
rect 153292 7550 153344 7556
rect 153936 3868 153988 3874
rect 153936 3810 153988 3816
rect 153200 3324 153252 3330
rect 153200 3266 153252 3272
rect 153948 480 153976 3810
rect 154684 3806 154712 52006
rect 155868 47592 155920 47598
rect 155868 47534 155920 47540
rect 155880 4146 155908 47534
rect 155960 46300 156012 46306
rect 155960 46242 156012 46248
rect 155132 4140 155184 4146
rect 155132 4082 155184 4088
rect 155868 4140 155920 4146
rect 155868 4082 155920 4088
rect 154672 3800 154724 3806
rect 154672 3742 154724 3748
rect 155144 480 155172 4082
rect 155972 3262 156000 46242
rect 156064 9042 156092 52006
rect 156984 46306 157012 52006
rect 158180 49298 158208 52020
rect 158732 52006 159206 52034
rect 158168 49292 158220 49298
rect 158168 49234 158220 49240
rect 158628 49088 158680 49094
rect 158628 49030 158680 49036
rect 156972 46300 157024 46306
rect 156972 46242 157024 46248
rect 156052 9036 156104 9042
rect 156052 8978 156104 8984
rect 156328 4004 156380 4010
rect 156328 3946 156380 3952
rect 155960 3256 156012 3262
rect 155960 3198 156012 3204
rect 156340 480 156368 3946
rect 158640 3466 158668 49030
rect 158732 26926 158760 52006
rect 160008 49156 160060 49162
rect 160008 49098 160060 49104
rect 158720 26920 158772 26926
rect 158720 26862 158772 26868
rect 159916 15904 159968 15910
rect 159916 15846 159968 15852
rect 159928 4146 159956 15846
rect 158720 4140 158772 4146
rect 158720 4082 158772 4088
rect 159916 4140 159968 4146
rect 159916 4082 159968 4088
rect 157524 3460 157576 3466
rect 157524 3402 157576 3408
rect 158628 3460 158680 3466
rect 158628 3402 158680 3408
rect 157536 480 157564 3402
rect 158732 480 158760 4082
rect 160020 4026 160048 49098
rect 160112 49026 160140 52020
rect 160296 52006 161046 52034
rect 161492 52006 161966 52034
rect 160100 49020 160152 49026
rect 160100 48962 160152 48968
rect 159928 3998 160048 4026
rect 159928 480 159956 3998
rect 160296 3534 160324 52006
rect 161492 4826 161520 52006
rect 162872 48822 162900 52020
rect 162964 52006 163898 52034
rect 164252 52006 164818 52034
rect 162124 48816 162176 48822
rect 162124 48758 162176 48764
rect 162860 48816 162912 48822
rect 162860 48758 162912 48764
rect 162136 17270 162164 48758
rect 162964 43450 162992 52006
rect 162952 43444 163004 43450
rect 162952 43386 163004 43392
rect 162124 17264 162176 17270
rect 162124 17206 162176 17212
rect 164148 17264 164200 17270
rect 164148 17206 164200 17212
rect 161480 4820 161532 4826
rect 161480 4762 161532 4768
rect 162308 4820 162360 4826
rect 162308 4762 162360 4768
rect 160284 3528 160336 3534
rect 160284 3470 160336 3476
rect 161112 3460 161164 3466
rect 161112 3402 161164 3408
rect 161124 480 161152 3402
rect 162320 480 162348 4762
rect 164160 4146 164188 17206
rect 164252 6254 164280 52006
rect 165528 49020 165580 49026
rect 165528 48962 165580 48968
rect 164240 6248 164292 6254
rect 164240 6190 164292 6196
rect 163504 4140 163556 4146
rect 163504 4082 163556 4088
rect 164148 4140 164200 4146
rect 164148 4082 164200 4088
rect 163516 480 163544 4082
rect 165540 3126 165568 48962
rect 165724 46238 165752 52020
rect 165908 52006 166658 52034
rect 167012 52006 167578 52034
rect 168392 52006 168590 52034
rect 165712 46232 165764 46238
rect 165712 46174 165764 46180
rect 165908 46050 165936 52006
rect 165632 46022 165936 46050
rect 165632 22778 165660 46022
rect 165620 22772 165672 22778
rect 165620 22714 165672 22720
rect 167012 7682 167040 52006
rect 167644 48340 167696 48346
rect 167644 48282 167696 48288
rect 167656 8974 167684 48282
rect 168392 18630 168420 52006
rect 168760 48278 168788 52142
rect 170416 48346 170444 52020
rect 171244 52006 171350 52034
rect 171888 52006 172270 52034
rect 172532 52006 173282 52034
rect 174004 52006 174202 52034
rect 174832 52006 175122 52034
rect 175292 52006 176042 52034
rect 176764 52006 176962 52034
rect 177592 52006 177974 52034
rect 178052 52006 178894 52034
rect 179524 52006 179814 52034
rect 180352 52006 180734 52034
rect 180812 52006 181654 52034
rect 182192 52006 182666 52034
rect 170404 48340 170456 48346
rect 170404 48282 170456 48288
rect 168748 48272 168800 48278
rect 168748 48214 168800 48220
rect 171244 44878 171272 52006
rect 171232 44872 171284 44878
rect 171232 44814 171284 44820
rect 171888 44554 171916 52006
rect 172428 49224 172480 49230
rect 172428 49166 172480 49172
rect 171152 44526 171916 44554
rect 168840 38684 168892 38690
rect 168840 38626 168892 38632
rect 168852 24138 168880 38626
rect 171152 25566 171180 44526
rect 171140 25560 171192 25566
rect 171140 25502 171192 25508
rect 168840 24132 168892 24138
rect 168840 24074 168892 24080
rect 168380 18624 168432 18630
rect 168380 18566 168432 18572
rect 167644 8968 167696 8974
rect 167644 8910 167696 8916
rect 167000 7676 167052 7682
rect 167000 7618 167052 7624
rect 169392 7608 169444 7614
rect 169392 7550 169444 7556
rect 165896 6180 165948 6186
rect 165896 6122 165948 6128
rect 164700 3120 164752 3126
rect 164700 3062 164752 3068
rect 165528 3120 165580 3126
rect 165528 3062 165580 3068
rect 164712 480 164740 3062
rect 165908 480 165936 6122
rect 167092 4072 167144 4078
rect 167092 4014 167144 4020
rect 167104 480 167132 4014
rect 168196 3528 168248 3534
rect 168196 3470 168248 3476
rect 168208 480 168236 3470
rect 169404 480 169432 7550
rect 170588 4140 170640 4146
rect 170588 4082 170640 4088
rect 170600 480 170628 4082
rect 172440 3602 172468 49166
rect 172532 10334 172560 52006
rect 173900 46232 173952 46238
rect 173900 46174 173952 46180
rect 172520 10328 172572 10334
rect 172520 10270 172572 10276
rect 172980 8968 173032 8974
rect 172980 8910 173032 8916
rect 171784 3596 171836 3602
rect 171784 3538 171836 3544
rect 172428 3596 172480 3602
rect 172428 3538 172480 3544
rect 171796 480 171824 3538
rect 172992 480 173020 8910
rect 173912 3670 173940 46174
rect 174004 19990 174032 52006
rect 174832 46238 174860 52006
rect 174820 46232 174872 46238
rect 174820 46174 174872 46180
rect 173992 19984 174044 19990
rect 173992 19926 174044 19932
rect 175292 11762 175320 52006
rect 176660 46912 176712 46918
rect 176660 46854 176712 46860
rect 175280 11756 175332 11762
rect 175280 11698 175332 11704
rect 176568 10328 176620 10334
rect 176568 10270 176620 10276
rect 173900 3664 173952 3670
rect 173900 3606 173952 3612
rect 175372 3392 175424 3398
rect 175372 3334 175424 3340
rect 174176 3324 174228 3330
rect 174176 3266 174228 3272
rect 174188 480 174216 3266
rect 175384 480 175412 3334
rect 176580 480 176608 10270
rect 176672 3738 176700 46854
rect 176764 21486 176792 52006
rect 177592 46918 177620 52006
rect 177580 46912 177632 46918
rect 177580 46854 177632 46860
rect 176752 21480 176804 21486
rect 176752 21422 176804 21428
rect 178052 13122 178080 52006
rect 179328 49292 179380 49298
rect 179328 49234 179380 49240
rect 178040 13116 178092 13122
rect 178040 13058 178092 13064
rect 176660 3732 176712 3738
rect 176660 3674 176712 3680
rect 177764 3596 177816 3602
rect 177764 3538 177816 3544
rect 177776 480 177804 3538
rect 179340 3482 179368 49234
rect 179420 48816 179472 48822
rect 179420 48758 179472 48764
rect 179432 3942 179460 48758
rect 179420 3936 179472 3942
rect 179420 3878 179472 3884
rect 178972 3454 179368 3482
rect 178972 480 179000 3454
rect 179524 3262 179552 52006
rect 180352 48822 180380 52006
rect 180340 48816 180392 48822
rect 180340 48758 180392 48764
rect 180812 14482 180840 52006
rect 180800 14476 180852 14482
rect 180800 14418 180852 14424
rect 180708 11756 180760 11762
rect 180708 11698 180760 11704
rect 180720 3670 180748 11698
rect 182192 3806 182220 52006
rect 183572 3874 183600 52020
rect 184492 47598 184520 52020
rect 184952 52006 185426 52034
rect 184480 47592 184532 47598
rect 184480 47534 184532 47540
rect 183744 4888 183796 4894
rect 183744 4830 183796 4836
rect 183560 3868 183612 3874
rect 183560 3810 183612 3816
rect 182180 3800 182232 3806
rect 182180 3742 182232 3748
rect 182548 3800 182600 3806
rect 182548 3742 182600 3748
rect 180156 3664 180208 3670
rect 180156 3606 180208 3612
rect 180708 3664 180760 3670
rect 180708 3606 180760 3612
rect 181352 3664 181404 3670
rect 181352 3606 181404 3612
rect 179512 3256 179564 3262
rect 179512 3198 179564 3204
rect 180168 480 180196 3606
rect 181364 480 181392 3606
rect 182560 480 182588 3742
rect 183756 480 183784 4830
rect 184952 4010 184980 52006
rect 186228 49360 186280 49366
rect 186228 49302 186280 49308
rect 184940 4004 184992 4010
rect 184940 3946 184992 3952
rect 184848 3732 184900 3738
rect 184848 3674 184900 3680
rect 184860 480 184888 3674
rect 186240 626 186268 49302
rect 186332 49094 186360 52020
rect 186424 52006 187358 52034
rect 186320 49088 186372 49094
rect 186320 49030 186372 49036
rect 186424 15910 186452 52006
rect 188264 49162 188292 52020
rect 189092 52006 189198 52034
rect 188252 49156 188304 49162
rect 188252 49098 188304 49104
rect 186412 15904 186464 15910
rect 186412 15846 186464 15852
rect 187608 13116 187660 13122
rect 187608 13058 187660 13064
rect 186056 598 186268 626
rect 187620 610 187648 13058
rect 188436 3868 188488 3874
rect 188436 3810 188488 3816
rect 187240 604 187292 610
rect 186056 480 186084 598
rect 187240 546 187292 552
rect 187608 604 187660 610
rect 187608 546 187660 552
rect 187252 480 187280 546
rect 188448 480 188476 3810
rect 189092 3466 189120 52006
rect 189368 12458 189396 52142
rect 190472 52006 191038 52034
rect 190472 17270 190500 52006
rect 192036 49026 192064 52020
rect 192680 52006 192970 52034
rect 193232 52006 193890 52034
rect 194612 52006 194810 52034
rect 195440 52006 195730 52034
rect 195992 52006 196742 52034
rect 192024 49020 192076 49026
rect 192024 48962 192076 48968
rect 192680 46050 192708 52006
rect 192036 46022 192708 46050
rect 192036 22114 192064 46022
rect 191944 22086 192064 22114
rect 190460 17264 190512 17270
rect 190460 17206 190512 17212
rect 189184 12430 189396 12458
rect 189184 4826 189212 12430
rect 191944 6186 191972 22086
rect 191932 6180 191984 6186
rect 191932 6122 191984 6128
rect 189172 4820 189224 4826
rect 189172 4762 189224 4768
rect 193232 4078 193260 52006
rect 193220 4072 193272 4078
rect 193220 4014 193272 4020
rect 192024 3936 192076 3942
rect 192024 3878 192076 3884
rect 189080 3460 189132 3466
rect 189080 3402 189132 3408
rect 189632 3460 189684 3466
rect 189632 3402 189684 3408
rect 189644 480 189672 3402
rect 190826 3360 190882 3369
rect 190826 3295 190882 3304
rect 190840 480 190868 3295
rect 192036 480 192064 3878
rect 194612 3534 194640 52006
rect 195440 41478 195468 52006
rect 194784 41472 194836 41478
rect 194784 41414 194836 41420
rect 195428 41472 195480 41478
rect 195428 41414 195480 41420
rect 194796 22114 194824 41414
rect 194704 22086 194824 22114
rect 194704 7614 194732 22086
rect 194692 7608 194744 7614
rect 194692 7550 194744 7556
rect 195992 4146 196020 52006
rect 197648 49230 197676 52020
rect 197924 51218 197952 52142
rect 197832 51190 197952 51218
rect 198752 52006 199502 52034
rect 200132 52006 200514 52034
rect 201144 52006 201434 52034
rect 201512 52006 202354 52034
rect 197636 49224 197688 49230
rect 197636 49166 197688 49172
rect 197832 41562 197860 51190
rect 197556 41534 197860 41562
rect 197556 41426 197584 41534
rect 197464 41398 197584 41426
rect 197464 38622 197492 41398
rect 197452 38616 197504 38622
rect 197452 38558 197504 38564
rect 197452 31612 197504 31618
rect 197452 31554 197504 31560
rect 197464 8974 197492 31554
rect 197452 8968 197504 8974
rect 197452 8910 197504 8916
rect 195980 4140 196032 4146
rect 195980 4082 196032 4088
rect 196808 4072 196860 4078
rect 196808 4014 196860 4020
rect 195612 4004 195664 4010
rect 195612 3946 195664 3952
rect 194600 3528 194652 3534
rect 194414 3496 194470 3505
rect 194600 3470 194652 3476
rect 194414 3431 194470 3440
rect 193220 3256 193272 3262
rect 193220 3198 193272 3204
rect 193232 480 193260 3198
rect 194428 480 194456 3431
rect 195624 480 195652 3946
rect 196820 480 196848 4014
rect 198004 3528 198056 3534
rect 198004 3470 198056 3476
rect 198016 480 198044 3470
rect 198752 3330 198780 52006
rect 200132 3398 200160 52006
rect 201144 42090 201172 52006
rect 201132 42084 201184 42090
rect 201132 42026 201184 42032
rect 200488 31612 200540 31618
rect 200488 31554 200540 31560
rect 200500 24206 200528 31554
rect 200304 24200 200356 24206
rect 200304 24142 200356 24148
rect 200488 24200 200540 24206
rect 200488 24142 200540 24148
rect 200316 12458 200344 24142
rect 200316 12430 200436 12458
rect 200408 10334 200436 12430
rect 200396 10328 200448 10334
rect 200396 10270 200448 10276
rect 201512 3602 201540 52006
rect 203260 49298 203288 52020
rect 203904 52006 204194 52034
rect 204272 52006 205206 52034
rect 205652 52006 206126 52034
rect 203248 49292 203300 49298
rect 203248 49234 203300 49240
rect 202788 49020 202840 49026
rect 202788 48962 202840 48968
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 200120 3392 200172 3398
rect 200120 3334 200172 3340
rect 200396 3392 200448 3398
rect 200396 3334 200448 3340
rect 198740 3324 198792 3330
rect 198740 3266 198792 3272
rect 199200 3324 199252 3330
rect 199200 3266 199252 3272
rect 199212 480 199240 3266
rect 200408 480 200436 3334
rect 201500 3188 201552 3194
rect 201500 3130 201552 3136
rect 201512 480 201540 3130
rect 202800 626 202828 48962
rect 203904 38865 203932 52006
rect 203890 38856 203946 38865
rect 203890 38791 203946 38800
rect 203154 38720 203210 38729
rect 203210 38678 203288 38706
rect 203154 38655 203210 38664
rect 203260 38622 203288 38678
rect 203248 38616 203300 38622
rect 203248 38558 203300 38564
rect 203156 29028 203208 29034
rect 203156 28970 203208 28976
rect 203168 22114 203196 28970
rect 202984 22098 203196 22114
rect 202972 22092 203208 22098
rect 203024 22086 203156 22092
rect 202972 22034 203024 22040
rect 203156 22034 203208 22040
rect 203168 19310 203196 22034
rect 203156 19304 203208 19310
rect 203156 19246 203208 19252
rect 203892 3732 203944 3738
rect 203892 3674 203944 3680
rect 202708 598 202828 626
rect 202708 480 202736 598
rect 203904 480 203932 3674
rect 204272 3670 204300 52006
rect 204904 48748 204956 48754
rect 204904 48690 204956 48696
rect 204916 4894 204944 48690
rect 204904 4888 204956 4894
rect 204904 4830 204956 4836
rect 205652 3806 205680 52006
rect 206928 49156 206980 49162
rect 206928 49098 206980 49104
rect 205640 3800 205692 3806
rect 205640 3742 205692 3748
rect 204260 3664 204312 3670
rect 204260 3606 204312 3612
rect 206940 3602 206968 49098
rect 207032 48754 207060 52020
rect 207124 52006 207966 52034
rect 207020 48748 207072 48754
rect 207020 48690 207072 48696
rect 207124 4146 207152 52006
rect 208872 49366 208900 52020
rect 209884 49706 209912 52020
rect 209976 52006 210818 52034
rect 211172 52006 211738 52034
rect 209044 49700 209096 49706
rect 209044 49642 209096 49648
rect 209872 49700 209924 49706
rect 209872 49642 209924 49648
rect 208860 49360 208912 49366
rect 208860 49302 208912 49308
rect 208308 49224 208360 49230
rect 208308 49166 208360 49172
rect 207112 4140 207164 4146
rect 207112 4082 207164 4088
rect 208320 3602 208348 49166
rect 209056 13122 209084 49642
rect 209044 13116 209096 13122
rect 209044 13058 209096 13064
rect 209976 3874 210004 52006
rect 209964 3868 210016 3874
rect 209964 3810 210016 3816
rect 211068 3800 211120 3806
rect 211068 3742 211120 3748
rect 208676 3732 208728 3738
rect 208676 3674 208728 3680
rect 206284 3596 206336 3602
rect 206284 3538 206336 3544
rect 206928 3596 206980 3602
rect 206928 3538 206980 3544
rect 207480 3596 207532 3602
rect 207480 3538 207532 3544
rect 208308 3596 208360 3602
rect 208308 3538 208360 3544
rect 205088 3120 205140 3126
rect 205088 3062 205140 3068
rect 205100 480 205128 3062
rect 206296 480 206324 3538
rect 207492 480 207520 3538
rect 208688 480 208716 3674
rect 209872 3188 209924 3194
rect 209872 3130 209924 3136
rect 209884 480 209912 3130
rect 211080 480 211108 3742
rect 211172 3466 211200 52006
rect 212540 48816 212592 48822
rect 212540 48758 212592 48764
rect 212552 3942 212580 48758
rect 212540 3936 212592 3942
rect 212540 3878 212592 3884
rect 211160 3460 211212 3466
rect 211160 3402 211212 3408
rect 212264 3460 212316 3466
rect 212264 3402 212316 3408
rect 212276 480 212304 3402
rect 212644 3369 212672 52020
rect 213288 52006 213578 52034
rect 214024 52006 214590 52034
rect 215404 52006 215510 52034
rect 216048 52006 216430 52034
rect 216692 52006 217350 52034
rect 218164 52006 218270 52034
rect 218348 52006 219282 52034
rect 219544 52006 220202 52034
rect 220924 52006 221122 52034
rect 213288 48822 213316 52006
rect 213828 49088 213880 49094
rect 213828 49030 213880 49036
rect 213276 48816 213328 48822
rect 213276 48758 213328 48764
rect 212630 3360 212686 3369
rect 212630 3295 212686 3304
rect 213840 626 213868 49030
rect 214024 3262 214052 52006
rect 215208 49292 215260 49298
rect 215208 49234 215260 49240
rect 215220 3534 215248 49234
rect 215300 48816 215352 48822
rect 215300 48758 215352 48764
rect 215312 4010 215340 48758
rect 215300 4004 215352 4010
rect 215300 3946 215352 3952
rect 214656 3528 214708 3534
rect 214656 3470 214708 3476
rect 215208 3528 215260 3534
rect 215404 3505 215432 52006
rect 216048 48822 216076 52006
rect 216036 48816 216088 48822
rect 216036 48758 216088 48764
rect 216692 4078 216720 52006
rect 217968 49360 218020 49366
rect 217968 49302 218020 49308
rect 216680 4072 216732 4078
rect 216680 4014 216732 4020
rect 215852 3868 215904 3874
rect 215852 3810 215904 3816
rect 215208 3470 215260 3476
rect 215390 3496 215446 3505
rect 214012 3256 214064 3262
rect 214012 3198 214064 3204
rect 213472 598 213868 626
rect 213472 480 213500 598
rect 214668 480 214696 3470
rect 215390 3431 215446 3440
rect 215864 480 215892 3810
rect 217980 3534 218008 49302
rect 218164 3942 218192 52006
rect 218244 4072 218296 4078
rect 218244 4014 218296 4020
rect 218152 3936 218204 3942
rect 218152 3878 218204 3884
rect 217048 3528 217100 3534
rect 217048 3470 217100 3476
rect 217968 3528 218020 3534
rect 218256 3482 218284 4014
rect 217968 3470 218020 3476
rect 217060 480 217088 3470
rect 218164 3454 218284 3482
rect 218164 480 218192 3454
rect 218348 3330 218376 52006
rect 219348 49496 219400 49502
rect 219348 49438 219400 49444
rect 219360 4078 219388 49438
rect 219348 4072 219400 4078
rect 219348 4014 219400 4020
rect 219348 3528 219400 3534
rect 219348 3470 219400 3476
rect 218336 3324 218388 3330
rect 218336 3266 218388 3272
rect 219360 480 219388 3470
rect 219544 3398 219572 52006
rect 220728 49428 220780 49434
rect 220728 49370 220780 49376
rect 219532 3392 219584 3398
rect 219532 3334 219584 3340
rect 220740 610 220768 49370
rect 220924 3942 220952 52006
rect 222028 49026 222056 52020
rect 222212 52006 222962 52034
rect 223776 52006 223974 52034
rect 222016 49020 222068 49026
rect 222016 48962 222068 48968
rect 222108 49020 222160 49026
rect 222108 48962 222160 48968
rect 220912 3936 220964 3942
rect 220912 3878 220964 3884
rect 222120 626 222148 48962
rect 222212 3602 222240 52006
rect 223776 3738 223804 52006
rect 224880 49162 224908 52020
rect 225800 49230 225828 52020
rect 226444 52006 226734 52034
rect 227272 52006 227654 52034
rect 227732 52006 228666 52034
rect 229112 52006 229586 52034
rect 225788 49224 225840 49230
rect 225788 49166 225840 49172
rect 224868 49156 224920 49162
rect 224868 49098 224920 49104
rect 226248 49156 226300 49162
rect 226248 49098 226300 49104
rect 224132 3936 224184 3942
rect 224132 3878 224184 3884
rect 223764 3732 223816 3738
rect 223764 3674 223816 3680
rect 222936 3664 222988 3670
rect 222936 3606 222988 3612
rect 222200 3596 222252 3602
rect 222200 3538 222252 3544
rect 220544 604 220596 610
rect 220544 546 220596 552
rect 220728 604 220780 610
rect 220728 546 220780 552
rect 221752 598 222148 626
rect 220556 480 220584 546
rect 221752 480 221780 598
rect 222948 480 222976 3606
rect 224144 480 224172 3878
rect 226260 3602 226288 49098
rect 226340 48816 226392 48822
rect 226340 48758 226392 48764
rect 225328 3596 225380 3602
rect 225328 3538 225380 3544
rect 226248 3596 226300 3602
rect 226248 3538 226300 3544
rect 225340 480 225368 3538
rect 226352 3194 226380 48758
rect 226444 3806 226472 52006
rect 227272 48822 227300 52006
rect 227260 48816 227312 48822
rect 227260 48758 227312 48764
rect 227732 4010 227760 52006
rect 229008 49224 229060 49230
rect 229008 49166 229060 49172
rect 227720 4004 227772 4010
rect 227720 3946 227772 3952
rect 226432 3800 226484 3806
rect 226432 3742 226484 3748
rect 228916 3800 228968 3806
rect 228916 3742 228968 3748
rect 226524 3732 226576 3738
rect 226524 3674 226576 3680
rect 226340 3188 226392 3194
rect 226340 3130 226392 3136
rect 226536 480 226564 3674
rect 227720 3392 227772 3398
rect 227720 3334 227772 3340
rect 227732 480 227760 3334
rect 228928 480 228956 3742
rect 229020 3398 229048 49166
rect 229112 3466 229140 52006
rect 230492 49094 230520 52020
rect 231412 49298 231440 52020
rect 231872 52006 232346 52034
rect 231400 49292 231452 49298
rect 231400 49234 231452 49240
rect 230480 49088 230532 49094
rect 230480 49030 230532 49036
rect 231768 49088 231820 49094
rect 231768 49030 231820 49036
rect 231780 3534 231808 49030
rect 231872 3874 231900 52006
rect 232504 49700 232556 49706
rect 232504 49642 232556 49648
rect 231860 3868 231912 3874
rect 231860 3810 231912 3816
rect 232516 3806 232544 49642
rect 233344 49366 233372 52020
rect 234264 49502 234292 52020
rect 234632 52006 235198 52034
rect 234252 49496 234304 49502
rect 234252 49438 234304 49444
rect 233332 49360 233384 49366
rect 233332 49302 233384 49308
rect 234528 49360 234580 49366
rect 234528 49302 234580 49308
rect 233148 49292 233200 49298
rect 233148 49234 233200 49240
rect 232504 3800 232556 3806
rect 232504 3742 232556 3748
rect 233160 3534 233188 49234
rect 234540 3534 234568 49302
rect 234632 3602 234660 52006
rect 236104 49434 236132 52020
rect 236092 49428 236144 49434
rect 236092 49370 236144 49376
rect 237024 49026 237052 52020
rect 237392 52006 238050 52034
rect 238864 52006 238970 52034
rect 237196 49564 237248 49570
rect 237196 49506 237248 49512
rect 237012 49020 237064 49026
rect 237012 48962 237064 48968
rect 237208 3602 237236 49506
rect 237288 49428 237340 49434
rect 237288 49370 237340 49376
rect 234620 3596 234672 3602
rect 234620 3538 234672 3544
rect 236000 3596 236052 3602
rect 236000 3538 236052 3544
rect 237196 3596 237248 3602
rect 237196 3538 237248 3544
rect 231308 3528 231360 3534
rect 231308 3470 231360 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233700 3528 233752 3534
rect 233700 3470 233752 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234804 3528 234856 3534
rect 234804 3470 234856 3476
rect 229100 3460 229152 3466
rect 229100 3402 229152 3408
rect 230112 3460 230164 3466
rect 230112 3402 230164 3408
rect 229008 3392 229060 3398
rect 229008 3334 229060 3340
rect 230124 480 230152 3402
rect 231320 480 231348 3470
rect 232516 480 232544 3470
rect 233712 480 233740 3470
rect 234816 480 234844 3470
rect 236012 480 236040 3538
rect 237300 3482 237328 49370
rect 237392 3738 237420 52006
rect 238668 49496 238720 49502
rect 238668 49438 238720 49444
rect 237380 3732 237432 3738
rect 237380 3674 237432 3680
rect 237208 3454 237328 3482
rect 237208 480 237236 3454
rect 238680 610 238708 49438
rect 238864 3942 238892 52006
rect 239876 49162 239904 52020
rect 240152 52006 240810 52034
rect 239864 49156 239916 49162
rect 239864 49098 239916 49104
rect 240048 49020 240100 49026
rect 240048 48962 240100 48968
rect 238852 3936 238904 3942
rect 238852 3878 238904 3884
rect 240060 3534 240088 48962
rect 240152 4010 240180 52006
rect 241428 49632 241480 49638
rect 241428 49574 241480 49580
rect 240140 4004 240192 4010
rect 240140 3946 240192 3952
rect 241440 3534 241468 49574
rect 241716 49230 241744 52020
rect 242728 49706 242756 52020
rect 243004 52006 243662 52034
rect 242716 49700 242768 49706
rect 242716 49642 242768 49648
rect 241704 49224 241756 49230
rect 241704 49166 241756 49172
rect 242808 49224 242860 49230
rect 242808 49166 242860 49172
rect 242820 3534 242848 49166
rect 239588 3528 239640 3534
rect 239588 3470 239640 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 241980 3528 242032 3534
rect 241980 3470 242032 3476
rect 242808 3528 242860 3534
rect 242808 3470 242860 3476
rect 238392 604 238444 610
rect 238392 546 238444 552
rect 238668 604 238720 610
rect 238668 546 238720 552
rect 238404 480 238432 546
rect 239600 480 239628 3470
rect 240796 480 240824 3470
rect 241992 480 242020 3470
rect 243004 3466 243032 52006
rect 244188 49156 244240 49162
rect 244188 49098 244240 49104
rect 244200 3534 244228 49098
rect 244568 49094 244596 52020
rect 245488 49298 245516 52020
rect 245568 49700 245620 49706
rect 245568 49642 245620 49648
rect 245476 49292 245528 49298
rect 245476 49234 245528 49240
rect 245580 49178 245608 49642
rect 246500 49366 246528 52020
rect 247144 52006 247434 52034
rect 248064 52006 248354 52034
rect 246488 49360 246540 49366
rect 246488 49302 246540 49308
rect 246948 49292 247000 49298
rect 246948 49234 247000 49240
rect 245488 49150 245608 49178
rect 244556 49088 244608 49094
rect 244556 49030 244608 49036
rect 245488 3534 245516 49150
rect 245568 49088 245620 49094
rect 245568 49030 245620 49036
rect 243176 3528 243228 3534
rect 243176 3470 243228 3476
rect 244188 3528 244240 3534
rect 244188 3470 244240 3476
rect 244372 3528 244424 3534
rect 244372 3470 244424 3476
rect 245476 3528 245528 3534
rect 245476 3470 245528 3476
rect 242992 3460 243044 3466
rect 242992 3402 243044 3408
rect 243188 480 243216 3470
rect 244384 480 244412 3470
rect 245580 480 245608 49030
rect 246960 3346 246988 49234
rect 247144 3670 247172 52006
rect 248064 49570 248092 52006
rect 248052 49564 248104 49570
rect 248052 49506 248104 49512
rect 248328 49564 248380 49570
rect 248328 49506 248380 49512
rect 247132 3664 247184 3670
rect 247132 3606 247184 3612
rect 248340 3346 248368 49506
rect 249260 49434 249288 52020
rect 250180 49502 250208 52020
rect 250168 49496 250220 49502
rect 250168 49438 250220 49444
rect 249248 49428 249300 49434
rect 249248 49370 249300 49376
rect 249708 49428 249760 49434
rect 249708 49370 249760 49376
rect 249720 3534 249748 49370
rect 251088 49360 251140 49366
rect 251088 49302 251140 49308
rect 251100 3534 251128 49302
rect 251192 49026 251220 52020
rect 252112 49638 252140 52020
rect 252100 49632 252152 49638
rect 252100 49574 252152 49580
rect 253032 49230 253060 52020
rect 253020 49224 253072 49230
rect 253020 49166 253072 49172
rect 253848 49224 253900 49230
rect 253848 49166 253900 49172
rect 251180 49020 251232 49026
rect 251180 48962 251232 48968
rect 252468 49020 252520 49026
rect 252468 48962 252520 48968
rect 252480 3534 252508 48962
rect 253860 3534 253888 49166
rect 253952 49162 253980 52020
rect 254872 49706 254900 52020
rect 254860 49700 254912 49706
rect 254860 49642 254912 49648
rect 255228 49496 255280 49502
rect 255228 49438 255280 49444
rect 253940 49156 253992 49162
rect 253940 49098 253992 49104
rect 249156 3528 249208 3534
rect 249156 3470 249208 3476
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 250352 3528 250404 3534
rect 250352 3470 250404 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 251456 3528 251508 3534
rect 251456 3470 251508 3476
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 252652 3528 252704 3534
rect 252652 3470 252704 3476
rect 253848 3528 253900 3534
rect 255240 3482 255268 49438
rect 255884 49094 255912 52020
rect 256804 49298 256832 52020
rect 257344 49632 257396 49638
rect 257344 49574 257396 49580
rect 256792 49292 256844 49298
rect 256792 49234 256844 49240
rect 255872 49088 255924 49094
rect 255872 49030 255924 49036
rect 256608 49088 256660 49094
rect 256608 49030 256660 49036
rect 256620 3482 256648 49030
rect 253848 3470 253900 3476
rect 246776 3318 246988 3346
rect 247972 3318 248368 3346
rect 246776 480 246804 3318
rect 247972 480 248000 3318
rect 249168 480 249196 3470
rect 250364 480 250392 3470
rect 251468 480 251496 3470
rect 252664 480 252692 3470
rect 255056 3454 255268 3482
rect 256252 3454 256648 3482
rect 253848 3324 253900 3330
rect 253848 3266 253900 3272
rect 253860 480 253888 3266
rect 255056 480 255084 3454
rect 256252 480 256280 3454
rect 257356 3330 257384 49574
rect 257724 49570 257752 52020
rect 257712 49564 257764 49570
rect 257712 49506 257764 49512
rect 258644 49434 258672 52020
rect 258632 49428 258684 49434
rect 258632 49370 258684 49376
rect 259564 49366 259592 52020
rect 259552 49360 259604 49366
rect 259552 49302 259604 49308
rect 257988 49156 258040 49162
rect 257988 49098 258040 49104
rect 258000 3534 258028 49098
rect 260576 49026 260604 52020
rect 261496 49230 261524 52020
rect 262128 49700 262180 49706
rect 262128 49642 262180 49648
rect 261484 49224 261536 49230
rect 261484 49166 261536 49172
rect 260564 49020 260616 49026
rect 260564 48962 260616 48968
rect 259368 48816 259420 48822
rect 259368 48758 259420 48764
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 257344 3324 257396 3330
rect 257344 3266 257396 3272
rect 257448 480 257476 3470
rect 259380 3126 259408 48758
rect 261484 48408 261536 48414
rect 261484 48350 261536 48356
rect 261496 3534 261524 48350
rect 259828 3528 259880 3534
rect 259828 3470 259880 3476
rect 261484 3528 261536 3534
rect 261484 3470 261536 3476
rect 258632 3120 258684 3126
rect 258632 3062 258684 3068
rect 259368 3120 259420 3126
rect 259368 3062 259420 3068
rect 258644 480 258672 3062
rect 259840 480 259868 3470
rect 262140 3262 262168 49642
rect 262416 49638 262444 52020
rect 262404 49632 262456 49638
rect 262404 49574 262456 49580
rect 263336 49502 263364 52020
rect 263416 49632 263468 49638
rect 263416 49574 263468 49580
rect 263324 49496 263376 49502
rect 263324 49438 263376 49444
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 261024 3256 261076 3262
rect 261024 3198 261076 3204
rect 262128 3256 262180 3262
rect 262128 3198 262180 3204
rect 261036 480 261064 3198
rect 262232 480 262260 3470
rect 263428 480 263456 49574
rect 264256 49094 264284 52020
rect 265268 49162 265296 52020
rect 265256 49156 265308 49162
rect 265256 49098 265308 49104
rect 264244 49088 264296 49094
rect 264244 49030 264296 49036
rect 264888 49088 264940 49094
rect 264888 49030 264940 49036
rect 263508 48544 263560 48550
rect 263508 48486 263560 48492
rect 263520 3534 263548 48486
rect 263508 3528 263560 3534
rect 264900 3482 264928 49030
rect 266188 48822 266216 52020
rect 266268 49292 266320 49298
rect 266268 49234 266320 49240
rect 266176 48816 266228 48822
rect 266176 48758 266228 48764
rect 266280 3534 266308 49234
rect 267108 48414 267136 52020
rect 268028 49706 268056 52020
rect 268016 49700 268068 49706
rect 268016 49642 268068 49648
rect 267648 49156 267700 49162
rect 267648 49098 267700 49104
rect 267096 48408 267148 48414
rect 267096 48350 267148 48356
rect 263508 3470 263560 3476
rect 264624 3454 264928 3482
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 264624 480 264652 3454
rect 265820 480 265848 3470
rect 267660 3466 267688 49098
rect 268948 48550 268976 52020
rect 269960 49638 269988 52020
rect 269948 49632 270000 49638
rect 269948 49574 270000 49580
rect 270880 49094 270908 52020
rect 271800 49298 271828 52020
rect 271788 49292 271840 49298
rect 271788 49234 271840 49240
rect 272720 49162 272748 52020
rect 272708 49156 272760 49162
rect 272708 49098 272760 49104
rect 270868 49088 270920 49094
rect 270868 49030 270920 49036
rect 273168 49088 273220 49094
rect 273168 49030 273220 49036
rect 271788 48884 271840 48890
rect 271788 48826 271840 48832
rect 269028 48748 269080 48754
rect 269028 48690 269080 48696
rect 268936 48544 268988 48550
rect 268936 48486 268988 48492
rect 269040 3534 269068 48690
rect 270408 48612 270460 48618
rect 270408 48554 270460 48560
rect 268108 3528 268160 3534
rect 268108 3470 268160 3476
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267648 3460 267700 3466
rect 267648 3402 267700 3408
rect 267016 480 267044 3402
rect 268120 480 268148 3470
rect 270420 3058 270448 48554
rect 270500 3528 270552 3534
rect 271800 3482 271828 48826
rect 272524 48816 272576 48822
rect 272524 48758 272576 48764
rect 272536 3534 272564 48758
rect 270500 3470 270552 3476
rect 269304 3052 269356 3058
rect 269304 2994 269356 3000
rect 270408 3052 270460 3058
rect 270408 2994 270460 3000
rect 269316 480 269344 2994
rect 270512 480 270540 3470
rect 271708 3454 271828 3482
rect 272524 3528 272576 3534
rect 273180 3482 273208 49030
rect 273640 48754 273668 52020
rect 274548 49632 274600 49638
rect 274548 49574 274600 49580
rect 273628 48748 273680 48754
rect 273628 48690 273680 48696
rect 274560 3534 274588 49574
rect 274652 48618 274680 52020
rect 275572 48822 275600 52020
rect 275928 49700 275980 49706
rect 275928 49642 275980 49648
rect 275560 48816 275612 48822
rect 275560 48758 275612 48764
rect 274640 48612 274692 48618
rect 274640 48554 274692 48560
rect 275940 3534 275968 49642
rect 276492 48890 276520 52020
rect 277308 49156 277360 49162
rect 277308 49098 277360 49104
rect 276480 48884 276532 48890
rect 276480 48826 276532 48832
rect 277320 3534 277348 49098
rect 277412 49094 277440 52020
rect 278332 49638 278360 52020
rect 279344 49706 279372 52020
rect 279332 49700 279384 49706
rect 279332 49642 279384 49648
rect 278320 49632 278372 49638
rect 278320 49574 278372 49580
rect 280264 49162 280292 52020
rect 280448 52006 281198 52034
rect 280252 49156 280304 49162
rect 280252 49098 280304 49104
rect 277400 49088 277452 49094
rect 277400 49030 277452 49036
rect 280448 48770 280476 52006
rect 280068 48748 280120 48754
rect 280068 48690 280120 48696
rect 280264 48742 280476 48770
rect 281448 48816 281500 48822
rect 281448 48758 281500 48764
rect 279976 48612 280028 48618
rect 279976 48554 280028 48560
rect 279884 4956 279936 4962
rect 279884 4898 279936 4904
rect 279896 4146 279924 4898
rect 279988 4842 280016 48554
rect 280080 4962 280108 48690
rect 280068 4956 280120 4962
rect 280068 4898 280120 4904
rect 279988 4814 280108 4842
rect 278872 4140 278924 4146
rect 278872 4082 278924 4088
rect 279884 4140 279936 4146
rect 279884 4082 279936 4088
rect 272524 3470 272576 3476
rect 272904 3454 273208 3482
rect 274088 3528 274140 3534
rect 274088 3470 274140 3476
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 275284 3528 275336 3534
rect 275284 3470 275336 3476
rect 275928 3528 275980 3534
rect 275928 3470 275980 3476
rect 276480 3528 276532 3534
rect 276480 3470 276532 3476
rect 277308 3528 277360 3534
rect 277308 3470 277360 3476
rect 271708 480 271736 3454
rect 272904 480 272932 3454
rect 274100 480 274128 3470
rect 275296 480 275324 3470
rect 276492 480 276520 3470
rect 277676 3460 277728 3466
rect 277676 3402 277728 3408
rect 277688 480 277716 3402
rect 278884 480 278912 4082
rect 280080 480 280108 4814
rect 280264 3466 280292 48742
rect 281460 4842 281488 48758
rect 282104 48754 282132 52020
rect 282092 48748 282144 48754
rect 282092 48690 282144 48696
rect 283024 48618 283052 52020
rect 284036 48822 284064 52020
rect 284312 52006 284970 52034
rect 284024 48816 284076 48822
rect 284024 48758 284076 48764
rect 283012 48612 283064 48618
rect 283012 48554 283064 48560
rect 284208 48340 284260 48346
rect 284208 48282 284260 48288
rect 281276 4814 281488 4842
rect 280252 3460 280304 3466
rect 280252 3402 280304 3408
rect 281276 480 281304 4814
rect 282460 3188 282512 3194
rect 282460 3130 282512 3136
rect 282472 480 282500 3130
rect 284220 3126 284248 48282
rect 284312 3194 284340 52006
rect 285876 48346 285904 52020
rect 286060 52006 286810 52034
rect 285864 48340 285916 48346
rect 285864 48282 285916 48288
rect 286060 46050 286088 52006
rect 287716 48346 287744 52020
rect 288452 52006 288742 52034
rect 288452 48362 288480 52006
rect 286968 48340 287020 48346
rect 286968 48282 287020 48288
rect 287704 48340 287756 48346
rect 287704 48282 287756 48288
rect 288176 48334 288480 48362
rect 289648 48346 289676 52020
rect 289924 52006 290582 52034
rect 289636 48340 289688 48346
rect 285784 46022 286088 46050
rect 285784 4010 285812 46022
rect 284760 4004 284812 4010
rect 284760 3946 284812 3952
rect 285772 4004 285824 4010
rect 285772 3946 285824 3952
rect 284300 3188 284352 3194
rect 284300 3130 284352 3136
rect 283656 3120 283708 3126
rect 283656 3062 283708 3068
rect 284208 3120 284260 3126
rect 284208 3062 284260 3068
rect 283668 480 283696 3062
rect 284772 480 284800 3946
rect 286980 3670 287008 48282
rect 288176 36582 288204 48334
rect 289636 48282 289688 48288
rect 288256 48272 288308 48278
rect 288256 48214 288308 48220
rect 288164 36576 288216 36582
rect 288164 36518 288216 36524
rect 287152 4140 287204 4146
rect 287152 4082 287204 4088
rect 285956 3664 286008 3670
rect 285956 3606 286008 3612
rect 286968 3664 287020 3670
rect 286968 3606 287020 3612
rect 285968 480 285996 3606
rect 287164 480 287192 4082
rect 288268 4026 288296 48214
rect 288348 36576 288400 36582
rect 288348 36518 288400 36524
rect 288360 4146 288388 36518
rect 289924 4146 289952 52006
rect 291488 48346 291516 52020
rect 291672 52006 292514 52034
rect 292592 52006 293434 52034
rect 293972 52006 294354 52034
rect 290924 48340 290976 48346
rect 290924 48282 290976 48288
rect 291476 48340 291528 48346
rect 291476 48282 291528 48288
rect 290936 42106 290964 48282
rect 291672 45234 291700 52006
rect 290844 42078 290964 42106
rect 291396 45206 291700 45234
rect 290844 37194 290872 42078
rect 291396 38622 291424 45206
rect 291384 38616 291436 38622
rect 291384 38558 291436 38564
rect 290832 37188 290884 37194
rect 290832 37130 290884 37136
rect 291476 29028 291528 29034
rect 291476 28970 291528 28976
rect 291016 27668 291068 27674
rect 291016 27610 291068 27616
rect 291028 27554 291056 27610
rect 291028 27526 291148 27554
rect 291120 18630 291148 27526
rect 291488 22114 291516 28970
rect 291304 22098 291516 22114
rect 291292 22092 291528 22098
rect 291344 22086 291476 22092
rect 291292 22034 291344 22040
rect 291476 22034 291528 22040
rect 290648 18624 290700 18630
rect 290648 18566 290700 18572
rect 291108 18624 291160 18630
rect 291108 18566 291160 18572
rect 288348 4140 288400 4146
rect 288348 4082 288400 4088
rect 289544 4140 289596 4146
rect 289544 4082 289596 4088
rect 289912 4140 289964 4146
rect 289912 4082 289964 4088
rect 288268 3998 288388 4026
rect 288360 480 288388 3998
rect 289556 480 289584 4082
rect 290660 2666 290688 18566
rect 291488 12050 291516 22034
rect 291488 12022 291608 12050
rect 291580 11778 291608 12022
rect 291488 11750 291608 11778
rect 291488 4146 291516 11750
rect 292592 4146 292620 52006
rect 293972 46918 294000 52006
rect 293960 46912 294012 46918
rect 293960 46854 294012 46860
rect 293960 37324 294012 37330
rect 293960 37266 294012 37272
rect 293972 27606 294000 37266
rect 293960 27600 294012 27606
rect 293960 27542 294012 27548
rect 293960 18012 294012 18018
rect 293960 17954 294012 17960
rect 293972 14634 294000 17954
rect 293972 14606 294368 14634
rect 291476 4140 291528 4146
rect 291476 4082 291528 4088
rect 291936 4140 291988 4146
rect 291936 4082 291988 4088
rect 292580 4140 292632 4146
rect 292580 4082 292632 4088
rect 293132 4140 293184 4146
rect 293132 4082 293184 4088
rect 290660 2638 290780 2666
rect 290752 480 290780 2638
rect 291948 480 291976 4082
rect 293144 480 293172 4082
rect 294340 480 294368 14606
rect 295260 4026 295288 52020
rect 296640 48822 296668 52142
rect 296824 52006 297206 52034
rect 296628 48816 296680 48822
rect 296628 48758 296680 48764
rect 296720 4412 296772 4418
rect 296720 4354 296772 4360
rect 295260 3998 295564 4026
rect 295536 480 295564 3998
rect 296732 480 296760 4354
rect 296824 4146 296852 52006
rect 296904 48816 296956 48822
rect 296904 48758 296956 48764
rect 296916 41410 296944 48758
rect 296904 41404 296956 41410
rect 296904 41346 296956 41352
rect 297088 41404 297140 41410
rect 297088 41346 297140 41352
rect 297100 29034 297128 41346
rect 296996 29028 297048 29034
rect 296996 28970 297048 28976
rect 297088 29028 297140 29034
rect 297088 28970 297140 28976
rect 297008 27606 297036 28970
rect 296996 27600 297048 27606
rect 296996 27542 297048 27548
rect 297088 27600 297140 27606
rect 297088 27542 297140 27548
rect 297100 4418 297128 27542
rect 297088 4412 297140 4418
rect 297088 4354 297140 4360
rect 298112 4146 298140 52020
rect 299046 52006 299428 52034
rect 299400 4146 299428 52006
rect 299952 48822 299980 52020
rect 299940 48816 299992 48822
rect 299940 48758 299992 48764
rect 300872 48346 300900 52020
rect 301898 52006 302096 52034
rect 302818 52006 303568 52034
rect 301044 48816 301096 48822
rect 301044 48758 301096 48764
rect 300860 48340 300912 48346
rect 300860 48282 300912 48288
rect 301056 14498 301084 48758
rect 300964 14470 301084 14498
rect 300964 12306 300992 14470
rect 300952 12300 301004 12306
rect 300952 12242 301004 12248
rect 301412 12300 301464 12306
rect 301412 12242 301464 12248
rect 296812 4140 296864 4146
rect 296812 4082 296864 4088
rect 297916 4140 297968 4146
rect 297916 4082 297968 4088
rect 298100 4140 298152 4146
rect 298100 4082 298152 4088
rect 299112 4140 299164 4146
rect 299112 4082 299164 4088
rect 299388 4140 299440 4146
rect 299388 4082 299440 4088
rect 300308 4140 300360 4146
rect 300308 4082 300360 4088
rect 297928 480 297956 4082
rect 299124 480 299152 4082
rect 300320 480 300348 4082
rect 301424 480 301452 12242
rect 302068 3602 302096 52006
rect 302148 48340 302200 48346
rect 302148 48282 302200 48288
rect 302056 3596 302108 3602
rect 302056 3538 302108 3544
rect 302160 3534 302188 48282
rect 302148 3528 302200 3534
rect 302148 3470 302200 3476
rect 302608 3528 302660 3534
rect 302608 3470 302660 3476
rect 302620 480 302648 3470
rect 303540 3466 303568 52006
rect 303724 48482 303752 52020
rect 304658 52006 304856 52034
rect 305578 52006 306328 52034
rect 303712 48476 303764 48482
rect 303712 48418 303764 48424
rect 304828 4078 304856 52006
rect 304908 48476 304960 48482
rect 304908 48418 304960 48424
rect 304816 4072 304868 4078
rect 304816 4014 304868 4020
rect 303804 3596 303856 3602
rect 303804 3538 303856 3544
rect 303528 3460 303580 3466
rect 303528 3402 303580 3408
rect 303816 480 303844 3538
rect 304920 3534 304948 48418
rect 306300 4146 306328 52006
rect 306576 48686 306604 52020
rect 307510 52006 307708 52034
rect 308430 52006 309088 52034
rect 306564 48680 306616 48686
rect 306564 48622 306616 48628
rect 306288 4140 306340 4146
rect 306288 4082 306340 4088
rect 307392 4072 307444 4078
rect 307392 4014 307444 4020
rect 304908 3528 304960 3534
rect 304908 3470 304960 3476
rect 306196 3528 306248 3534
rect 306196 3470 306248 3476
rect 305000 3460 305052 3466
rect 305000 3402 305052 3408
rect 305012 480 305040 3402
rect 306208 480 306236 3470
rect 307404 480 307432 4014
rect 307680 3466 307708 52006
rect 308588 4140 308640 4146
rect 308588 4082 308640 4088
rect 307668 3460 307720 3466
rect 307668 3402 307720 3408
rect 308600 480 308628 4082
rect 309060 3602 309088 52006
rect 309336 48822 309364 52020
rect 310270 52006 310376 52034
rect 309324 48816 309376 48822
rect 309324 48758 309376 48764
rect 309324 48680 309376 48686
rect 309324 48622 309376 48628
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 309336 1442 309364 48622
rect 310348 3398 310376 52006
rect 311268 48822 311296 52020
rect 310428 48816 310480 48822
rect 310428 48758 310480 48764
rect 311256 48816 311308 48822
rect 311256 48758 311308 48764
rect 310440 3534 310468 48758
rect 312188 48754 312216 52020
rect 312544 48816 312596 48822
rect 312544 48758 312596 48764
rect 312176 48748 312228 48754
rect 312176 48690 312228 48696
rect 312176 3596 312228 3602
rect 312176 3538 312228 3544
rect 310428 3528 310480 3534
rect 310428 3470 310480 3476
rect 310980 3460 311032 3466
rect 310980 3402 311032 3408
rect 310336 3392 310388 3398
rect 310336 3334 310388 3340
rect 309336 1414 309732 1442
rect 309704 626 309732 1414
rect 309704 598 309824 626
rect 309796 480 309824 598
rect 310992 480 311020 3402
rect 312188 480 312216 3538
rect 312556 3262 312584 48758
rect 313108 3738 313136 52020
rect 314028 48822 314056 52020
rect 314016 48816 314068 48822
rect 314016 48758 314068 48764
rect 314948 48754 314976 52020
rect 315868 52006 315974 52034
rect 316894 52006 317368 52034
rect 315304 48816 315356 48822
rect 315304 48758 315356 48764
rect 313188 48748 313240 48754
rect 313188 48690 313240 48696
rect 314936 48748 314988 48754
rect 314936 48690 314988 48696
rect 313096 3732 313148 3738
rect 313096 3674 313148 3680
rect 313200 3466 313228 48690
rect 315316 3806 315344 48758
rect 315304 3800 315356 3806
rect 315304 3742 315356 3748
rect 313372 3528 313424 3534
rect 313372 3470 313424 3476
rect 313188 3460 313240 3466
rect 313188 3402 313240 3408
rect 312544 3256 312596 3262
rect 312544 3198 312596 3204
rect 313384 480 313412 3470
rect 315868 3466 315896 52006
rect 315948 48748 316000 48754
rect 315948 48690 316000 48696
rect 315960 3670 315988 48690
rect 315948 3664 316000 3670
rect 315948 3606 316000 3612
rect 316960 3528 317012 3534
rect 316960 3470 317012 3476
rect 315856 3460 315908 3466
rect 315856 3402 315908 3408
rect 314568 3392 314620 3398
rect 314568 3334 314620 3340
rect 314580 480 314608 3334
rect 315764 3256 315816 3262
rect 315764 3198 315816 3204
rect 315776 480 315804 3198
rect 316972 480 317000 3470
rect 317340 3262 317368 52006
rect 317800 48822 317828 52020
rect 317788 48816 317840 48822
rect 317788 48758 317840 48764
rect 318064 3732 318116 3738
rect 318064 3674 318116 3680
rect 317328 3256 317380 3262
rect 317328 3198 317380 3204
rect 318076 480 318104 3674
rect 318720 3534 318748 52020
rect 319654 52006 320128 52034
rect 320100 4010 320128 52006
rect 320652 48618 320680 52020
rect 321572 48822 321600 52020
rect 322506 52006 322888 52034
rect 320824 48816 320876 48822
rect 320824 48758 320876 48764
rect 321560 48816 321612 48822
rect 321560 48758 321612 48764
rect 322756 48816 322808 48822
rect 322756 48758 322808 48764
rect 320640 48612 320692 48618
rect 320640 48554 320692 48560
rect 320088 4004 320140 4010
rect 320088 3946 320140 3952
rect 319260 3800 319312 3806
rect 319260 3742 319312 3748
rect 318708 3528 318760 3534
rect 318708 3470 318760 3476
rect 319272 480 319300 3742
rect 320456 3664 320508 3670
rect 320456 3606 320508 3612
rect 320468 480 320496 3606
rect 320836 3330 320864 48758
rect 321468 48612 321520 48618
rect 321468 48554 321520 48560
rect 320824 3324 320876 3330
rect 320824 3266 320876 3272
rect 321480 3058 321508 48554
rect 322768 3602 322796 48758
rect 322756 3596 322808 3602
rect 322756 3538 322808 3544
rect 322860 3466 322888 52006
rect 323412 48618 323440 52020
rect 324332 49706 324360 52020
rect 325358 52006 325648 52034
rect 324320 49700 324372 49706
rect 324320 49642 324372 49648
rect 323400 48612 323452 48618
rect 323400 48554 323452 48560
rect 324228 48612 324280 48618
rect 324228 48554 324280 48560
rect 324240 3670 324268 48554
rect 325620 3738 325648 52006
rect 326264 48822 326292 52020
rect 326344 49700 326396 49706
rect 326344 49642 326396 49648
rect 326252 48816 326304 48822
rect 326252 48758 326304 48764
rect 325608 3732 325660 3738
rect 325608 3674 325660 3680
rect 324228 3664 324280 3670
rect 324228 3606 324280 3612
rect 326356 3534 326384 49642
rect 327184 48822 327212 52020
rect 328118 52006 328316 52034
rect 326988 48816 327040 48822
rect 326988 48758 327040 48764
rect 327172 48816 327224 48822
rect 327172 48758 327224 48764
rect 326436 4004 326488 4010
rect 326436 3946 326488 3952
rect 325240 3528 325292 3534
rect 325240 3470 325292 3476
rect 326344 3528 326396 3534
rect 326344 3470 326396 3476
rect 321652 3460 321704 3466
rect 321652 3402 321704 3408
rect 322848 3460 322900 3466
rect 322848 3402 322900 3408
rect 321468 3052 321520 3058
rect 321468 2994 321520 3000
rect 321664 480 321692 3402
rect 324044 3324 324096 3330
rect 324044 3266 324096 3272
rect 322848 3256 322900 3262
rect 322848 3198 322900 3204
rect 322860 480 322888 3198
rect 324056 480 324084 3266
rect 325252 480 325280 3470
rect 326448 480 326476 3946
rect 327000 2922 327028 48758
rect 328288 3398 328316 52006
rect 329024 48822 329052 52020
rect 330036 48822 330064 52020
rect 330970 52006 331076 52034
rect 331890 52006 332548 52034
rect 328368 48816 328420 48822
rect 328368 48758 328420 48764
rect 329012 48816 329064 48822
rect 329012 48758 329064 48764
rect 329748 48816 329800 48822
rect 329748 48758 329800 48764
rect 330024 48816 330076 48822
rect 330024 48758 330076 48764
rect 328380 3874 328408 48758
rect 328368 3868 328420 3874
rect 328368 3810 328420 3816
rect 329760 3602 329788 48758
rect 328828 3596 328880 3602
rect 328828 3538 328880 3544
rect 329748 3596 329800 3602
rect 329748 3538 329800 3544
rect 328276 3392 328328 3398
rect 328276 3334 328328 3340
rect 327632 3052 327684 3058
rect 327632 2994 327684 3000
rect 326988 2916 327040 2922
rect 326988 2858 327040 2864
rect 327644 480 327672 2994
rect 328840 480 328868 3538
rect 330024 3460 330076 3466
rect 330024 3402 330076 3408
rect 330036 480 330064 3402
rect 331048 3330 331076 52006
rect 331128 48816 331180 48822
rect 331128 48758 331180 48764
rect 331140 4078 331168 48758
rect 331128 4072 331180 4078
rect 331128 4014 331180 4020
rect 332520 4010 332548 52006
rect 332796 48822 332824 52020
rect 333730 52006 333836 52034
rect 334742 52006 335308 52034
rect 332784 48816 332836 48822
rect 332784 48758 332836 48764
rect 332508 4004 332560 4010
rect 332508 3946 332560 3952
rect 333808 3738 333836 52006
rect 333888 48816 333940 48822
rect 333888 48758 333940 48764
rect 333612 3732 333664 3738
rect 333612 3674 333664 3680
rect 333796 3732 333848 3738
rect 333796 3674 333848 3680
rect 331220 3664 331272 3670
rect 331220 3606 331272 3612
rect 331036 3324 331088 3330
rect 331036 3266 331088 3272
rect 331232 480 331260 3606
rect 332416 3528 332468 3534
rect 332416 3470 332468 3476
rect 332428 480 332456 3470
rect 333624 480 333652 3674
rect 333900 3398 333928 48758
rect 335280 3942 335308 52006
rect 335648 48822 335676 52020
rect 335636 48816 335688 48822
rect 335636 48758 335688 48764
rect 335268 3936 335320 3942
rect 335268 3878 335320 3884
rect 335912 3868 335964 3874
rect 335912 3810 335964 3816
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 334716 2916 334768 2922
rect 334716 2858 334768 2864
rect 334728 480 334756 2858
rect 335924 480 335952 3810
rect 336568 3670 336596 52020
rect 337502 52006 338068 52034
rect 336648 48816 336700 48822
rect 336648 48758 336700 48764
rect 336660 3874 336688 48758
rect 338040 4146 338068 52006
rect 338500 48822 338528 52020
rect 339328 52006 339434 52034
rect 340354 52006 340828 52034
rect 338488 48816 338540 48822
rect 338488 48758 338540 48764
rect 338028 4140 338080 4146
rect 338028 4082 338080 4088
rect 336648 3868 336700 3874
rect 336648 3810 336700 3816
rect 336556 3664 336608 3670
rect 336556 3606 336608 3612
rect 339328 3602 339356 52006
rect 339408 48816 339460 48822
rect 339408 48758 339460 48764
rect 339420 3806 339448 48758
rect 339500 4072 339552 4078
rect 339500 4014 339552 4020
rect 339408 3800 339460 3806
rect 339408 3742 339460 3748
rect 338304 3596 338356 3602
rect 338304 3538 338356 3544
rect 339316 3596 339368 3602
rect 339316 3538 339368 3544
rect 337108 3528 337160 3534
rect 337108 3470 337160 3476
rect 337120 480 337148 3470
rect 338316 480 338344 3538
rect 339512 480 339540 4014
rect 340696 3460 340748 3466
rect 340696 3402 340748 3408
rect 340708 480 340736 3402
rect 340800 3330 340828 52006
rect 341260 48822 341288 52020
rect 342088 52006 342194 52034
rect 343206 52006 343588 52034
rect 341248 48816 341300 48822
rect 341248 48758 341300 48764
rect 341892 4004 341944 4010
rect 341892 3946 341944 3952
rect 340788 3324 340840 3330
rect 340788 3266 340840 3272
rect 341904 480 341932 3946
rect 342088 3466 342116 52006
rect 342168 48816 342220 48822
rect 342168 48758 342220 48764
rect 342180 4078 342208 48758
rect 342168 4072 342220 4078
rect 342168 4014 342220 4020
rect 343560 3534 343588 52006
rect 344112 48822 344140 52020
rect 345032 48822 345060 52020
rect 345966 52006 346348 52034
rect 344100 48816 344152 48822
rect 344100 48758 344152 48764
rect 344928 48816 344980 48822
rect 344928 48758 344980 48764
rect 345020 48816 345072 48822
rect 345020 48758 345072 48764
rect 346216 48816 346268 48822
rect 346216 48758 346268 48764
rect 344284 3732 344336 3738
rect 344284 3674 344336 3680
rect 343548 3528 343600 3534
rect 343548 3470 343600 3476
rect 342076 3460 342128 3466
rect 342076 3402 342128 3408
rect 343088 3392 343140 3398
rect 343088 3334 343140 3340
rect 343100 480 343128 3334
rect 344296 480 344324 3674
rect 344940 3262 344968 48758
rect 345480 3936 345532 3942
rect 345480 3878 345532 3884
rect 344928 3256 344980 3262
rect 344928 3198 344980 3204
rect 345492 480 345520 3878
rect 346228 3398 346256 48758
rect 346320 4010 346348 52006
rect 346872 48550 346900 52020
rect 347884 48822 347912 52020
rect 348818 52006 349108 52034
rect 349738 52006 350488 52034
rect 347872 48816 347924 48822
rect 347872 48758 347924 48764
rect 348976 48816 349028 48822
rect 348976 48758 349028 48764
rect 346860 48544 346912 48550
rect 346860 48486 346912 48492
rect 347688 48544 347740 48550
rect 347688 48486 347740 48492
rect 346308 4004 346360 4010
rect 346308 3946 346360 3952
rect 347700 3942 347728 48486
rect 348884 4140 348936 4146
rect 348884 4082 348936 4088
rect 347688 3936 347740 3942
rect 347688 3878 347740 3884
rect 346676 3868 346728 3874
rect 346676 3810 346728 3816
rect 346216 3392 346268 3398
rect 346216 3334 346268 3340
rect 346688 480 346716 3810
rect 347872 3664 347924 3670
rect 347872 3606 347924 3612
rect 348896 3618 348924 4082
rect 348988 3738 349016 48758
rect 349080 3874 349108 52006
rect 350460 4146 350488 52006
rect 350644 49026 350672 52020
rect 351578 52006 351868 52034
rect 352590 52006 353248 52034
rect 350632 49020 350684 49026
rect 350632 48962 350684 48968
rect 350448 4140 350500 4146
rect 350448 4082 350500 4088
rect 349068 3868 349120 3874
rect 349068 3810 349120 3816
rect 351840 3806 351868 52006
rect 350264 3800 350316 3806
rect 350264 3742 350316 3748
rect 351828 3800 351880 3806
rect 351828 3742 351880 3748
rect 348976 3732 349028 3738
rect 348976 3674 349028 3680
rect 347884 480 347912 3606
rect 348896 3590 349108 3618
rect 349080 480 349108 3590
rect 350276 480 350304 3742
rect 351368 3596 351420 3602
rect 351368 3538 351420 3544
rect 351380 480 351408 3538
rect 353220 3330 353248 52006
rect 353496 48822 353524 52020
rect 354430 52006 354628 52034
rect 355350 52006 356008 52034
rect 353484 48816 353536 48822
rect 353484 48758 353536 48764
rect 354496 48816 354548 48822
rect 354496 48758 354548 48764
rect 353760 4072 353812 4078
rect 353760 4014 353812 4020
rect 352564 3324 352616 3330
rect 352564 3266 352616 3272
rect 353208 3324 353260 3330
rect 353208 3266 353260 3272
rect 352576 480 352604 3266
rect 353772 480 353800 4014
rect 354508 3602 354536 48758
rect 354600 4078 354628 52006
rect 354588 4072 354640 4078
rect 354588 4014 354640 4020
rect 355980 3670 356008 52006
rect 356256 48822 356284 52020
rect 357282 52006 357388 52034
rect 358202 52006 358768 52034
rect 356244 48816 356296 48822
rect 356244 48758 356296 48764
rect 357256 48816 357308 48822
rect 357256 48758 357308 48764
rect 357268 4826 357296 48758
rect 357256 4820 357308 4826
rect 357256 4762 357308 4768
rect 355968 3664 356020 3670
rect 355968 3606 356020 3612
rect 354496 3596 354548 3602
rect 354496 3538 354548 3544
rect 357360 3534 357388 52006
rect 356152 3528 356204 3534
rect 356152 3470 356204 3476
rect 357348 3528 357400 3534
rect 357348 3470 357400 3476
rect 354956 3460 355008 3466
rect 354956 3402 355008 3408
rect 354968 480 354996 3402
rect 356164 480 356192 3470
rect 358740 3398 358768 52006
rect 359108 48822 359136 52020
rect 360042 52006 360148 52034
rect 360962 52006 361528 52034
rect 359096 48816 359148 48822
rect 359096 48758 359148 48764
rect 360016 48816 360068 48822
rect 360016 48758 360068 48764
rect 360028 6186 360056 48758
rect 360016 6180 360068 6186
rect 360016 6122 360068 6128
rect 359740 4004 359792 4010
rect 359740 3946 359792 3952
rect 358544 3392 358596 3398
rect 358544 3334 358596 3340
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 357360 480 357388 3198
rect 358556 480 358584 3334
rect 359752 480 359780 3946
rect 360120 3466 360148 52006
rect 361500 4010 361528 52006
rect 361960 48822 361988 52020
rect 361948 48816 362000 48822
rect 361948 48758 362000 48764
rect 362776 48816 362828 48822
rect 362776 48758 362828 48764
rect 362788 7614 362816 48758
rect 362776 7608 362828 7614
rect 362776 7550 362828 7556
rect 361488 4004 361540 4010
rect 361488 3946 361540 3952
rect 360936 3936 360988 3942
rect 360936 3878 360988 3884
rect 360108 3460 360160 3466
rect 360108 3402 360160 3408
rect 360948 480 360976 3878
rect 362880 3738 362908 52020
rect 363814 52006 364288 52034
rect 364260 3942 364288 52006
rect 364720 48550 364748 52020
rect 364708 48544 364760 48550
rect 364708 48486 364760 48492
rect 364524 4140 364576 4146
rect 364524 4082 364576 4088
rect 364248 3936 364300 3942
rect 364248 3878 364300 3884
rect 363328 3868 363380 3874
rect 363328 3810 363380 3816
rect 362132 3732 362184 3738
rect 362132 3674 362184 3680
rect 362868 3732 362920 3738
rect 362868 3674 362920 3680
rect 362144 480 362172 3674
rect 363340 480 363368 3810
rect 364536 480 364564 4082
rect 365640 3874 365668 52020
rect 366666 52006 367048 52034
rect 365812 49020 365864 49026
rect 365812 48962 365864 48968
rect 365628 3868 365680 3874
rect 365628 3810 365680 3816
rect 365824 626 365852 48962
rect 367020 4146 367048 52006
rect 367572 48822 367600 52020
rect 368492 48822 368520 52020
rect 369426 52006 369808 52034
rect 367560 48816 367612 48822
rect 367560 48758 367612 48764
rect 368388 48816 368440 48822
rect 368388 48758 368440 48764
rect 368480 48816 368532 48822
rect 368480 48758 368532 48764
rect 369676 48816 369728 48822
rect 369676 48758 369728 48764
rect 368400 22778 368428 48758
rect 368388 22772 368440 22778
rect 368388 22714 368440 22720
rect 367008 4140 367060 4146
rect 367008 4082 367060 4088
rect 369688 3806 369716 48758
rect 366916 3800 366968 3806
rect 366916 3742 366968 3748
rect 369676 3800 369728 3806
rect 369676 3742 369728 3748
rect 365732 598 365852 626
rect 365732 480 365760 598
rect 366928 480 366956 3742
rect 369780 3602 369808 52006
rect 370332 48822 370360 52020
rect 371344 48822 371372 52020
rect 372278 52006 372568 52034
rect 370320 48816 370372 48822
rect 370320 48758 370372 48764
rect 371148 48816 371200 48822
rect 371148 48758 371200 48764
rect 371332 48816 371384 48822
rect 371332 48758 371384 48764
rect 372436 48816 372488 48822
rect 372436 48758 372488 48764
rect 371160 8974 371188 48758
rect 371148 8968 371200 8974
rect 371148 8910 371200 8916
rect 370412 4072 370464 4078
rect 370412 4014 370464 4020
rect 369216 3596 369268 3602
rect 369216 3538 369268 3544
rect 369768 3596 369820 3602
rect 369768 3538 369820 3544
rect 368020 3324 368072 3330
rect 368020 3266 368072 3272
rect 368032 480 368060 3266
rect 369228 480 369256 3538
rect 370424 480 370452 4014
rect 371608 3664 371660 3670
rect 371608 3606 371660 3612
rect 371620 480 371648 3606
rect 372448 3194 372476 48758
rect 372540 4078 372568 52006
rect 373184 49026 373212 52020
rect 373172 49020 373224 49026
rect 373172 48962 373224 48968
rect 374104 48822 374132 52020
rect 375038 52006 375236 52034
rect 376050 52006 376708 52034
rect 374092 48816 374144 48822
rect 374092 48758 374144 48764
rect 373264 48544 373316 48550
rect 373264 48486 373316 48492
rect 373276 4894 373304 48486
rect 373264 4888 373316 4894
rect 373264 4830 373316 4836
rect 372804 4820 372856 4826
rect 372804 4762 372856 4768
rect 372528 4072 372580 4078
rect 372528 4014 372580 4020
rect 372436 3188 372488 3194
rect 372436 3130 372488 3136
rect 372816 480 372844 4762
rect 375208 3534 375236 52006
rect 375288 48816 375340 48822
rect 375288 48758 375340 48764
rect 374000 3528 374052 3534
rect 374000 3470 374052 3476
rect 375196 3528 375248 3534
rect 375196 3470 375248 3476
rect 374012 480 374040 3470
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 375208 480 375236 3334
rect 375300 3262 375328 48758
rect 376680 6186 376708 52006
rect 376956 48822 376984 52020
rect 377890 52006 377996 52034
rect 376944 48816 376996 48822
rect 376944 48758 376996 48764
rect 376392 6180 376444 6186
rect 376392 6122 376444 6128
rect 376668 6180 376720 6186
rect 376668 6122 376720 6128
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 376404 480 376432 6122
rect 377968 3670 377996 52006
rect 378048 48816 378100 48822
rect 378048 48758 378100 48764
rect 377956 3664 378008 3670
rect 377956 3606 378008 3612
rect 377588 3460 377640 3466
rect 377588 3402 377640 3408
rect 377600 480 377628 3402
rect 378060 3398 378088 48758
rect 378796 48754 378824 52020
rect 379716 48822 379744 52020
rect 379704 48816 379756 48822
rect 379704 48758 379756 48764
rect 378784 48748 378836 48754
rect 378784 48690 378836 48696
rect 379980 7608 380032 7614
rect 379980 7550 380032 7556
rect 378784 4004 378836 4010
rect 378784 3946 378836 3952
rect 378048 3392 378100 3398
rect 378048 3334 378100 3340
rect 378796 480 378824 3946
rect 379992 480 380020 7550
rect 380728 3466 380756 52020
rect 381662 52006 382228 52034
rect 380808 48816 380860 48822
rect 380808 48758 380860 48764
rect 380716 3460 380768 3466
rect 380716 3402 380768 3408
rect 380820 3330 380848 48758
rect 381544 48748 381596 48754
rect 381544 48690 381596 48696
rect 381556 4826 381584 48690
rect 382200 7682 382228 52006
rect 382568 48822 382596 52020
rect 383502 52006 383608 52034
rect 384514 52006 384988 52034
rect 382556 48816 382608 48822
rect 382556 48758 382608 48764
rect 383476 48816 383528 48822
rect 383476 48758 383528 48764
rect 382188 7676 382240 7682
rect 382188 7618 382240 7624
rect 383384 4888 383436 4894
rect 383384 4830 383436 4836
rect 381544 4820 381596 4826
rect 381544 4762 381596 4768
rect 382372 3936 382424 3942
rect 382372 3878 382424 3884
rect 381176 3732 381228 3738
rect 381176 3674 381228 3680
rect 380808 3324 380860 3330
rect 380808 3266 380860 3272
rect 381188 480 381216 3674
rect 382384 480 382412 3878
rect 383396 3618 383424 4830
rect 383488 4010 383516 48758
rect 383476 4004 383528 4010
rect 383476 3946 383528 3952
rect 383580 3738 383608 52006
rect 384960 10334 384988 52006
rect 385420 48822 385448 52020
rect 385408 48816 385460 48822
rect 385408 48758 385460 48764
rect 386236 48816 386288 48822
rect 386236 48758 386288 48764
rect 384948 10328 385000 10334
rect 384948 10270 385000 10276
rect 386248 4146 386276 48758
rect 385868 4140 385920 4146
rect 385868 4082 385920 4088
rect 386236 4140 386288 4146
rect 386236 4082 386288 4088
rect 384672 3868 384724 3874
rect 384672 3810 384724 3816
rect 383568 3732 383620 3738
rect 383568 3674 383620 3680
rect 383396 3590 383608 3618
rect 383580 480 383608 3590
rect 384684 480 384712 3810
rect 385880 480 385908 4082
rect 386340 3942 386368 52020
rect 387274 52006 387748 52034
rect 386420 22772 386472 22778
rect 386420 22714 386472 22720
rect 386328 3936 386380 3942
rect 386328 3878 386380 3884
rect 386432 610 386460 22714
rect 387720 11762 387748 52006
rect 388180 48822 388208 52020
rect 389192 48822 389220 52020
rect 388168 48816 388220 48822
rect 388168 48758 388220 48764
rect 389088 48816 389140 48822
rect 389088 48758 389140 48764
rect 389180 48816 389232 48822
rect 389180 48758 389232 48764
rect 387708 11756 387760 11762
rect 387708 11698 387760 11704
rect 389100 3874 389128 48758
rect 390112 48754 390140 52020
rect 391032 49094 391060 52020
rect 391020 49088 391072 49094
rect 391020 49030 391072 49036
rect 391204 49020 391256 49026
rect 391204 48962 391256 48968
rect 390468 48816 390520 48822
rect 390468 48758 390520 48764
rect 390100 48748 390152 48754
rect 390100 48690 390152 48696
rect 389088 3868 389140 3874
rect 389088 3810 389140 3816
rect 390480 3806 390508 48758
rect 390652 8968 390704 8974
rect 390652 8910 390704 8916
rect 388260 3800 388312 3806
rect 388260 3742 388312 3748
rect 390468 3800 390520 3806
rect 390468 3742 390520 3748
rect 386420 604 386472 610
rect 386420 546 386472 552
rect 387064 604 387116 610
rect 387064 546 387116 552
rect 387076 480 387104 546
rect 388272 480 388300 3742
rect 389456 3596 389508 3602
rect 389456 3538 389508 3544
rect 389468 480 389496 3538
rect 390664 480 390692 8910
rect 391216 4690 391244 48962
rect 391952 48822 391980 52020
rect 392872 49638 392900 52020
rect 393898 52006 394648 52034
rect 392860 49632 392912 49638
rect 392860 49574 392912 49580
rect 393964 49632 394016 49638
rect 393964 49574 394016 49580
rect 391940 48816 391992 48822
rect 391940 48758 391992 48764
rect 393228 48816 393280 48822
rect 393228 48758 393280 48764
rect 391296 48748 391348 48754
rect 391296 48690 391348 48696
rect 391308 8974 391336 48690
rect 391296 8968 391348 8974
rect 391296 8910 391348 8916
rect 391204 4684 391256 4690
rect 391204 4626 391256 4632
rect 393240 4078 393268 48758
rect 393976 4894 394004 49574
rect 394620 15910 394648 52006
rect 394804 48822 394832 52020
rect 395738 52006 395936 52034
rect 394792 48816 394844 48822
rect 394792 48758 394844 48764
rect 394608 15904 394660 15910
rect 394608 15846 394660 15852
rect 395908 13190 395936 52006
rect 395988 48816 396040 48822
rect 395988 48758 396040 48764
rect 395896 13184 395948 13190
rect 395896 13126 395948 13132
rect 393964 4888 394016 4894
rect 393964 4830 394016 4836
rect 394240 4684 394292 4690
rect 394240 4626 394292 4632
rect 393044 4072 393096 4078
rect 393044 4014 393096 4020
rect 393228 4072 393280 4078
rect 393228 4014 393280 4020
rect 391848 3188 391900 3194
rect 391848 3130 391900 3136
rect 391860 480 391888 3130
rect 393056 480 393084 4014
rect 394252 480 394280 4626
rect 396000 3602 396028 48758
rect 396644 48686 396672 52020
rect 397564 48822 397592 52020
rect 398590 52006 398696 52034
rect 399510 52006 400168 52034
rect 397552 48816 397604 48822
rect 397552 48758 397604 48764
rect 396632 48680 396684 48686
rect 396632 48622 396684 48628
rect 398668 6186 398696 52006
rect 398748 48816 398800 48822
rect 398748 48758 398800 48764
rect 397828 6180 397880 6186
rect 397828 6122 397880 6128
rect 398656 6180 398708 6186
rect 398656 6122 398708 6128
rect 395988 3596 396040 3602
rect 395988 3538 396040 3544
rect 396632 3528 396684 3534
rect 396632 3470 396684 3476
rect 395436 3256 395488 3262
rect 395436 3198 395488 3204
rect 395448 480 395476 3198
rect 396644 480 396672 3470
rect 397840 480 397868 6122
rect 398760 3534 398788 48758
rect 399484 48680 399536 48686
rect 399484 48622 399536 48628
rect 399496 17270 399524 48622
rect 400140 18630 400168 52006
rect 400416 48822 400444 52020
rect 400404 48816 400456 48822
rect 400404 48758 400456 48764
rect 401336 48754 401364 52020
rect 402270 52006 402928 52034
rect 401508 48816 401560 48822
rect 401508 48758 401560 48764
rect 401324 48748 401376 48754
rect 401324 48690 401376 48696
rect 400128 18624 400180 18630
rect 400128 18566 400180 18572
rect 399484 17264 399536 17270
rect 399484 17206 399536 17212
rect 401324 4820 401376 4826
rect 401324 4762 401376 4768
rect 400220 3664 400272 3670
rect 400220 3606 400272 3612
rect 398748 3528 398800 3534
rect 398748 3470 398800 3476
rect 399024 3392 399076 3398
rect 399024 3334 399076 3340
rect 399036 480 399064 3334
rect 400232 480 400260 3606
rect 401336 480 401364 4762
rect 401520 3670 401548 48758
rect 402244 48748 402296 48754
rect 402244 48690 402296 48696
rect 402256 7614 402284 48690
rect 402900 22778 402928 52006
rect 403268 48822 403296 52020
rect 403256 48816 403308 48822
rect 403256 48758 403308 48764
rect 402888 22772 402940 22778
rect 402888 22714 402940 22720
rect 404188 14550 404216 52020
rect 405122 52006 405688 52034
rect 404268 48816 404320 48822
rect 404268 48758 404320 48764
rect 404176 14544 404228 14550
rect 404176 14486 404228 14492
rect 402244 7608 402296 7614
rect 402244 7550 402296 7556
rect 401508 3664 401560 3670
rect 401508 3606 401560 3612
rect 404280 3466 404308 48758
rect 405660 19990 405688 52006
rect 406028 49026 406056 52020
rect 406962 52006 407068 52034
rect 406016 49020 406068 49026
rect 406016 48962 406068 48968
rect 405648 19984 405700 19990
rect 405648 19926 405700 19932
rect 404912 7676 404964 7682
rect 404912 7618 404964 7624
rect 403716 3460 403768 3466
rect 403716 3402 403768 3408
rect 404268 3460 404320 3466
rect 404268 3402 404320 3408
rect 402520 3324 402572 3330
rect 402520 3266 402572 3272
rect 402532 480 402560 3266
rect 403728 480 403756 3402
rect 404924 480 404952 7618
rect 407040 4826 407068 52006
rect 407960 48754 407988 52020
rect 408880 48822 408908 52020
rect 409708 52006 409814 52034
rect 410734 52006 411208 52034
rect 408868 48816 408920 48822
rect 408868 48758 408920 48764
rect 407948 48748 408000 48754
rect 407948 48690 408000 48696
rect 409708 10334 409736 52006
rect 409788 48816 409840 48822
rect 409788 48758 409840 48764
rect 408592 10328 408644 10334
rect 408592 10270 408644 10276
rect 409696 10328 409748 10334
rect 409696 10270 409748 10276
rect 407028 4820 407080 4826
rect 407028 4762 407080 4768
rect 406108 4004 406160 4010
rect 406108 3946 406160 3952
rect 406120 480 406148 3946
rect 407304 3732 407356 3738
rect 407304 3674 407356 3680
rect 407316 480 407344 3674
rect 408604 3482 408632 10270
rect 409696 4140 409748 4146
rect 409696 4082 409748 4088
rect 408512 3454 408632 3482
rect 408512 480 408540 3454
rect 409708 480 409736 4082
rect 409800 4010 409828 48758
rect 410524 48748 410576 48754
rect 410524 48690 410576 48696
rect 410536 21418 410564 48690
rect 411180 24138 411208 52006
rect 411640 48822 411668 52020
rect 412652 48822 412680 52020
rect 413586 52006 413876 52034
rect 411628 48816 411680 48822
rect 411628 48758 411680 48764
rect 412548 48816 412600 48822
rect 412548 48758 412600 48764
rect 412640 48816 412692 48822
rect 412640 48758 412692 48764
rect 411168 24132 411220 24138
rect 411168 24074 411220 24080
rect 410524 21412 410576 21418
rect 410524 21354 410576 21360
rect 411260 11756 411312 11762
rect 411260 11698 411312 11704
rect 409788 4004 409840 4010
rect 409788 3946 409840 3952
rect 410892 3936 410944 3942
rect 410892 3878 410944 3884
rect 410904 480 410932 3878
rect 411272 3346 411300 11698
rect 412560 3942 412588 48758
rect 413848 25566 413876 52006
rect 414492 48822 414520 52020
rect 415412 48822 415440 52020
rect 416346 52006 416636 52034
rect 413928 48816 413980 48822
rect 413928 48758 413980 48764
rect 414480 48816 414532 48822
rect 414480 48758 414532 48764
rect 415308 48816 415360 48822
rect 415308 48758 415360 48764
rect 415400 48816 415452 48822
rect 415400 48758 415452 48764
rect 413836 25560 413888 25566
rect 413836 25502 413888 25508
rect 413940 11762 413968 48758
rect 413928 11756 413980 11762
rect 413928 11698 413980 11704
rect 412548 3936 412600 3942
rect 412548 3878 412600 3884
rect 415320 3874 415348 48758
rect 416608 26926 416636 52006
rect 416872 49088 416924 49094
rect 416872 49030 416924 49036
rect 416688 48816 416740 48822
rect 416688 48758 416740 48764
rect 416596 26920 416648 26926
rect 416596 26862 416648 26868
rect 416700 8974 416728 48758
rect 415676 8968 415728 8974
rect 415676 8910 415728 8916
rect 416688 8968 416740 8974
rect 416688 8910 416740 8916
rect 413284 3868 413336 3874
rect 413284 3810 413336 3816
rect 415308 3868 415360 3874
rect 415308 3810 415360 3816
rect 411272 3318 412128 3346
rect 412100 480 412128 3318
rect 413296 480 413324 3810
rect 414480 3800 414532 3806
rect 414480 3742 414532 3748
rect 414492 480 414520 3742
rect 415688 480 415716 8910
rect 416884 480 416912 49030
rect 417344 48482 417372 52020
rect 418264 48550 418292 52020
rect 419184 49366 419212 52020
rect 419172 49360 419224 49366
rect 419172 49302 419224 49308
rect 420104 48822 420132 52020
rect 421024 48822 421052 52020
rect 422050 52006 422156 52034
rect 422970 52006 423628 52034
rect 420092 48816 420144 48822
rect 420092 48758 420144 48764
rect 420828 48816 420880 48822
rect 420828 48758 420880 48764
rect 421012 48816 421064 48822
rect 421012 48758 421064 48764
rect 418252 48544 418304 48550
rect 418252 48486 418304 48492
rect 420184 48544 420236 48550
rect 420184 48486 420236 48492
rect 417332 48476 417384 48482
rect 417332 48418 417384 48424
rect 418068 48476 418120 48482
rect 418068 48418 418120 48424
rect 417976 4072 418028 4078
rect 417976 4014 418028 4020
rect 417988 480 418016 4014
rect 418080 3738 418108 48418
rect 420196 15910 420224 48486
rect 419540 15904 419592 15910
rect 419540 15846 419592 15852
rect 420184 15904 420236 15910
rect 420184 15846 420236 15852
rect 419172 4888 419224 4894
rect 419172 4830 419224 4836
rect 418068 3732 418120 3738
rect 418068 3674 418120 3680
rect 419184 480 419212 4830
rect 419552 3482 419580 15846
rect 419552 3454 420408 3482
rect 420380 480 420408 3454
rect 420840 3194 420868 48758
rect 422128 29646 422156 52006
rect 422944 49360 422996 49366
rect 422944 49302 422996 49308
rect 422208 48816 422260 48822
rect 422208 48758 422260 48764
rect 422116 29640 422168 29646
rect 422116 29582 422168 29588
rect 422220 13122 422248 48758
rect 422956 28286 422984 49302
rect 422944 28280 422996 28286
rect 422944 28222 422996 28228
rect 422300 13184 422352 13190
rect 422300 13126 422352 13132
rect 422208 13116 422260 13122
rect 422208 13058 422260 13064
rect 421564 3596 421616 3602
rect 421564 3538 421616 3544
rect 420828 3188 420880 3194
rect 420828 3130 420880 3136
rect 421576 480 421604 3538
rect 422312 3346 422340 13126
rect 423600 3806 423628 52006
rect 423876 48822 423904 52020
rect 424810 52006 425008 52034
rect 425730 52006 426388 52034
rect 423864 48816 423916 48822
rect 423864 48758 423916 48764
rect 424876 48816 424928 48822
rect 424876 48758 424928 48764
rect 424888 17338 424916 48758
rect 424876 17332 424928 17338
rect 424876 17274 424928 17280
rect 423680 17264 423732 17270
rect 423680 17206 423732 17212
rect 423588 3800 423640 3806
rect 423588 3742 423640 3748
rect 423692 3346 423720 17206
rect 424980 14482 425008 52006
rect 424968 14476 425020 14482
rect 424968 14418 425020 14424
rect 426256 6180 426308 6186
rect 426256 6122 426308 6128
rect 425152 3528 425204 3534
rect 425152 3470 425204 3476
rect 426268 3482 426296 6122
rect 426360 3602 426388 52006
rect 426728 49162 426756 52020
rect 427662 52006 427768 52034
rect 428582 52006 429148 52034
rect 426716 49156 426768 49162
rect 426716 49098 426768 49104
rect 427740 31074 427768 52006
rect 427728 31068 427780 31074
rect 427728 31010 427780 31016
rect 426440 18624 426492 18630
rect 426440 18566 426492 18572
rect 426348 3596 426400 3602
rect 426348 3538 426400 3544
rect 422312 3318 422800 3346
rect 423692 3318 423996 3346
rect 422772 480 422800 3318
rect 423968 480 423996 3318
rect 425164 480 425192 3470
rect 426268 3454 426388 3482
rect 426360 480 426388 3454
rect 426452 3346 426480 18566
rect 428740 3664 428792 3670
rect 428740 3606 428792 3612
rect 426452 3318 427584 3346
rect 427556 480 427584 3318
rect 428752 480 428780 3606
rect 429120 3262 429148 52006
rect 429488 48414 429516 52020
rect 430408 52006 430514 52034
rect 431434 52006 431908 52034
rect 429476 48408 429528 48414
rect 429476 48350 429528 48356
rect 430408 32434 430436 52006
rect 430488 48408 430540 48414
rect 430488 48350 430540 48356
rect 430396 32428 430448 32434
rect 430396 32370 430448 32376
rect 430500 18698 430528 48350
rect 430580 22772 430632 22778
rect 430580 22714 430632 22720
rect 430488 18692 430540 18698
rect 430488 18634 430540 18640
rect 429936 7608 429988 7614
rect 429936 7550 429988 7556
rect 429108 3256 429160 3262
rect 429108 3198 429160 3204
rect 429948 480 429976 7550
rect 430592 3346 430620 22714
rect 431880 3534 431908 52006
rect 432340 48822 432368 52020
rect 432328 48816 432380 48822
rect 432328 48758 432380 48764
rect 433260 33794 433288 52020
rect 434194 52006 434668 52034
rect 433984 48816 434036 48822
rect 433984 48758 434036 48764
rect 433248 33788 433300 33794
rect 433248 33730 433300 33736
rect 433996 19990 434024 48758
rect 433340 19984 433392 19990
rect 433340 19926 433392 19932
rect 433984 19984 434036 19990
rect 433984 19926 434036 19932
rect 431868 3528 431920 3534
rect 431868 3470 431920 3476
rect 433352 3466 433380 19926
rect 433432 14544 433484 14550
rect 433432 14486 433484 14492
rect 432328 3460 432380 3466
rect 432328 3402 432380 3408
rect 433340 3460 433392 3466
rect 433340 3402 433392 3408
rect 430592 3318 431172 3346
rect 431144 480 431172 3318
rect 432340 480 432368 3402
rect 433444 592 433472 14486
rect 434640 3670 434668 52006
rect 435192 49094 435220 52020
rect 435180 49088 435232 49094
rect 435180 49030 435232 49036
rect 434720 49020 434772 49026
rect 434720 48962 434772 48968
rect 434628 3664 434680 3670
rect 434628 3606 434680 3612
rect 434628 3460 434680 3466
rect 434628 3402 434680 3408
rect 433444 564 433564 592
rect 433536 480 433564 564
rect 434640 480 434668 3402
rect 434732 610 434760 48962
rect 436112 48822 436140 52020
rect 437046 52006 437428 52034
rect 436100 48816 436152 48822
rect 436100 48758 436152 48764
rect 437296 48816 437348 48822
rect 437296 48758 437348 48764
rect 437020 4820 437072 4826
rect 437020 4762 437072 4768
rect 434720 604 434772 610
rect 434720 546 434772 552
rect 435824 604 435876 610
rect 435824 546 435876 552
rect 435836 480 435864 546
rect 437032 480 437060 4762
rect 437308 3466 437336 48758
rect 437296 3460 437348 3466
rect 437296 3402 437348 3408
rect 437400 3398 437428 52006
rect 437952 48822 437980 52020
rect 438124 49156 438176 49162
rect 438124 49098 438176 49104
rect 437940 48816 437992 48822
rect 437940 48758 437992 48764
rect 438136 28966 438164 49098
rect 438872 48822 438900 52020
rect 439898 52006 440096 52034
rect 440818 52006 441568 52034
rect 438768 48816 438820 48822
rect 438768 48758 438820 48764
rect 438860 48816 438912 48822
rect 438860 48758 438912 48764
rect 438124 28960 438176 28966
rect 438124 28902 438176 28908
rect 438780 21486 438808 48758
rect 438768 21480 438820 21486
rect 438768 21422 438820 21428
rect 437480 21412 437532 21418
rect 437480 21354 437532 21360
rect 437388 3392 437440 3398
rect 437388 3334 437440 3340
rect 437492 610 437520 21354
rect 438308 19372 438360 19378
rect 438308 19314 438360 19320
rect 438320 4826 438348 19314
rect 438308 4820 438360 4826
rect 438308 4762 438360 4768
rect 440068 4078 440096 52006
rect 440148 48816 440200 48822
rect 440148 48758 440200 48764
rect 440056 4072 440108 4078
rect 440056 4014 440108 4020
rect 439412 4004 439464 4010
rect 439412 3946 439464 3952
rect 437480 604 437532 610
rect 437480 546 437532 552
rect 438216 604 438268 610
rect 438216 546 438268 552
rect 438228 480 438256 546
rect 439424 480 439452 3946
rect 440160 3330 440188 48758
rect 440240 10328 440292 10334
rect 440240 10270 440292 10276
rect 440148 3324 440200 3330
rect 440148 3266 440200 3272
rect 440252 626 440280 10270
rect 441540 6186 441568 52006
rect 441724 48822 441752 52020
rect 442658 52006 442948 52034
rect 441712 48816 441764 48822
rect 441712 48758 441764 48764
rect 442816 48816 442868 48822
rect 442816 48758 442868 48764
rect 441620 24132 441672 24138
rect 441620 24074 441672 24080
rect 441528 6180 441580 6186
rect 441528 6122 441580 6128
rect 440252 598 440556 626
rect 441632 610 441660 24074
rect 442828 4146 442856 48758
rect 442816 4140 442868 4146
rect 442816 4082 442868 4088
rect 442920 3505 442948 52006
rect 443564 48754 443592 52020
rect 444576 48822 444604 52020
rect 445510 52006 445708 52034
rect 446430 52006 447088 52034
rect 444564 48816 444616 48822
rect 444564 48758 444616 48764
rect 445576 48816 445628 48822
rect 445576 48758 445628 48764
rect 443552 48748 443604 48754
rect 443552 48690 443604 48696
rect 444380 25560 444432 25566
rect 444380 25502 444432 25508
rect 443092 11756 443144 11762
rect 443092 11698 443144 11704
rect 443000 3936 443052 3942
rect 443000 3878 443052 3884
rect 442906 3496 442962 3505
rect 442906 3431 442962 3440
rect 440528 592 440556 598
rect 441620 604 441672 610
rect 440528 564 440648 592
rect 440620 480 440648 564
rect 441620 546 441672 552
rect 441804 604 441856 610
rect 441804 546 441856 552
rect 441816 480 441844 546
rect 443012 480 443040 3878
rect 443104 610 443132 11698
rect 444392 610 444420 25502
rect 445588 22846 445616 48758
rect 445576 22840 445628 22846
rect 445576 22782 445628 22788
rect 445680 3942 445708 52006
rect 446404 48748 446456 48754
rect 446404 48690 446456 48696
rect 446416 6254 446444 48690
rect 447060 7682 447088 52006
rect 447336 47598 447364 52020
rect 448270 52006 448376 52034
rect 449282 52006 449848 52034
rect 447324 47592 447376 47598
rect 447324 47534 447376 47540
rect 447784 8968 447836 8974
rect 447784 8910 447836 8916
rect 447048 7676 447100 7682
rect 447048 7618 447100 7624
rect 446404 6248 446456 6254
rect 446404 6190 446456 6196
rect 445668 3936 445720 3942
rect 445668 3878 445720 3884
rect 446588 3868 446640 3874
rect 446588 3810 446640 3816
rect 443092 604 443144 610
rect 443092 546 443144 552
rect 444196 604 444248 610
rect 444196 546 444248 552
rect 444380 604 444432 610
rect 444380 546 444432 552
rect 445392 604 445444 610
rect 445392 546 445444 552
rect 444208 480 444236 546
rect 445404 480 445432 546
rect 446600 480 446628 3810
rect 447796 480 447824 8910
rect 448348 4010 448376 52006
rect 448520 26920 448572 26926
rect 448520 26862 448572 26868
rect 448336 4004 448388 4010
rect 448336 3946 448388 3952
rect 448532 610 448560 26862
rect 449820 9042 449848 52006
rect 450188 49706 450216 52020
rect 451122 52006 451228 52034
rect 452042 52006 452608 52034
rect 450176 49700 450228 49706
rect 450176 49642 450228 49648
rect 449808 9036 449860 9042
rect 449808 8978 449860 8984
rect 451200 3874 451228 52006
rect 451924 49700 451976 49706
rect 451924 49642 451976 49648
rect 451280 28280 451332 28286
rect 451280 28222 451332 28228
rect 451188 3868 451240 3874
rect 451188 3810 451240 3816
rect 451292 3738 451320 28222
rect 451936 24138 451964 49642
rect 451924 24132 451976 24138
rect 451924 24074 451976 24080
rect 451372 15904 451424 15910
rect 451372 15846 451424 15852
rect 450176 3732 450228 3738
rect 450176 3674 450228 3680
rect 451280 3732 451332 3738
rect 451280 3674 451332 3680
rect 448520 604 448572 610
rect 448520 546 448572 552
rect 448980 604 449032 610
rect 448980 546 449032 552
rect 448992 480 449020 546
rect 450188 480 450216 3674
rect 451384 3482 451412 15846
rect 452580 10334 452608 52006
rect 452948 48822 452976 52020
rect 452936 48816 452988 48822
rect 452936 48758 452988 48764
rect 453856 48816 453908 48822
rect 453856 48758 453908 48764
rect 453868 17270 453896 48758
rect 453856 17264 453908 17270
rect 453856 17206 453908 17212
rect 452568 10328 452620 10334
rect 452568 10270 452620 10276
rect 453960 3738 453988 52020
rect 454880 49026 454908 52020
rect 454868 49020 454920 49026
rect 454868 48962 454920 48968
rect 455800 46238 455828 52020
rect 455788 46232 455840 46238
rect 455788 46174 455840 46180
rect 455420 29640 455472 29646
rect 455420 29582 455472 29588
rect 454040 13116 454092 13122
rect 454040 13058 454092 13064
rect 452476 3732 452528 3738
rect 452476 3674 452528 3680
rect 453948 3732 454000 3738
rect 453948 3674 454000 3680
rect 451292 3454 451412 3482
rect 451292 480 451320 3454
rect 452488 480 452516 3674
rect 454052 3346 454080 13058
rect 455432 3346 455460 29582
rect 456720 3369 456748 52020
rect 457654 52006 458128 52034
rect 457444 49088 457496 49094
rect 457444 49030 457496 49036
rect 457456 4894 457484 49030
rect 458100 11762 458128 52006
rect 458652 48822 458680 52020
rect 459572 48822 459600 52020
rect 460506 52006 460796 52034
rect 458640 48816 458692 48822
rect 458640 48758 458692 48764
rect 459468 48816 459520 48822
rect 459468 48758 459520 48764
rect 459560 48816 459612 48822
rect 459560 48758 459612 48764
rect 459480 25566 459508 48758
rect 459468 25560 459520 25566
rect 459468 25502 459520 25508
rect 458180 17332 458232 17338
rect 458180 17274 458232 17280
rect 458088 11756 458140 11762
rect 458088 11698 458140 11704
rect 457444 4888 457496 4894
rect 457444 4830 457496 4836
rect 457260 3800 457312 3806
rect 457260 3742 457312 3748
rect 456706 3360 456762 3369
rect 454052 3318 454908 3346
rect 455432 3318 456104 3346
rect 453672 3188 453724 3194
rect 453672 3130 453724 3136
rect 453684 480 453712 3130
rect 454880 480 454908 3318
rect 456076 480 456104 3318
rect 456706 3295 456762 3304
rect 457272 480 457300 3742
rect 458192 3346 458220 17274
rect 459652 14476 459704 14482
rect 459652 14418 459704 14424
rect 458192 3318 458496 3346
rect 458468 480 458496 3318
rect 459664 480 459692 14418
rect 460768 13190 460796 52006
rect 460848 48816 460900 48822
rect 460848 48758 460900 48764
rect 460756 13184 460808 13190
rect 460756 13126 460808 13132
rect 460860 3806 460888 48758
rect 461412 48754 461440 52020
rect 462332 48822 462360 52020
rect 463358 52006 463556 52034
rect 462320 48816 462372 48822
rect 462320 48758 462372 48764
rect 461400 48748 461452 48754
rect 461400 48690 461452 48696
rect 462320 31068 462372 31074
rect 462320 31010 462372 31016
rect 462044 4820 462096 4826
rect 462044 4762 462096 4768
rect 460848 3800 460900 3806
rect 460848 3742 460900 3748
rect 460848 3596 460900 3602
rect 460848 3538 460900 3544
rect 460860 480 460888 3538
rect 462056 480 462084 4762
rect 462332 3346 462360 31010
rect 463528 14482 463556 52006
rect 464264 48822 464292 52020
rect 465184 49366 465212 52020
rect 466118 52006 466408 52034
rect 465172 49360 465224 49366
rect 465172 49302 465224 49308
rect 463608 48816 463660 48822
rect 463608 48758 463660 48764
rect 464252 48816 464304 48822
rect 464252 48758 464304 48764
rect 464988 48816 465040 48822
rect 464988 48758 465040 48764
rect 463516 14476 463568 14482
rect 463516 14418 463568 14424
rect 463620 3602 463648 48758
rect 464344 48748 464396 48754
rect 464344 48690 464396 48696
rect 464356 26926 464384 48690
rect 464344 26920 464396 26926
rect 464344 26862 464396 26868
rect 465000 18630 465028 48758
rect 465080 18692 465132 18698
rect 465080 18634 465132 18640
rect 464988 18624 465040 18630
rect 464988 18566 465040 18572
rect 463608 3596 463660 3602
rect 463608 3538 463660 3544
rect 465092 3346 465120 18634
rect 466380 7614 466408 52006
rect 467024 48822 467052 52020
rect 468036 48822 468064 52020
rect 467012 48816 467064 48822
rect 467012 48758 467064 48764
rect 467748 48816 467800 48822
rect 467748 48758 467800 48764
rect 468024 48816 468076 48822
rect 468024 48758 468076 48764
rect 466460 32428 466512 32434
rect 466460 32370 466512 32376
rect 466368 7608 466420 7614
rect 466368 7550 466420 7556
rect 466472 3346 466500 32370
rect 467760 8974 467788 48758
rect 468956 48754 468984 52020
rect 469890 52006 470548 52034
rect 469128 48816 469180 48822
rect 469128 48758 469180 48764
rect 468944 48748 468996 48754
rect 468944 48690 468996 48696
rect 467932 19984 467984 19990
rect 467932 19926 467984 19932
rect 467748 8968 467800 8974
rect 467748 8910 467800 8916
rect 467944 3534 467972 19926
rect 469140 5250 469168 48758
rect 469864 48748 469916 48754
rect 469864 48690 469916 48696
rect 469220 33788 469272 33794
rect 469220 33730 469272 33736
rect 469048 5222 469168 5250
rect 469048 3602 469076 5222
rect 469036 3596 469088 3602
rect 469036 3538 469088 3544
rect 467840 3528 467892 3534
rect 467840 3470 467892 3476
rect 467932 3528 467984 3534
rect 467932 3470 467984 3476
rect 469128 3528 469180 3534
rect 469128 3470 469180 3476
rect 467852 3346 467880 3470
rect 462332 3318 463280 3346
rect 465092 3318 465672 3346
rect 466472 3318 466868 3346
rect 467852 3318 467972 3346
rect 463252 480 463280 3318
rect 464436 3256 464488 3262
rect 464436 3198 464488 3204
rect 464448 480 464476 3198
rect 465644 480 465672 3318
rect 466840 480 466868 3318
rect 467944 480 467972 3318
rect 469140 480 469168 3470
rect 469232 3346 469260 33730
rect 469876 15910 469904 48690
rect 470520 28286 470548 52006
rect 470796 48822 470824 52020
rect 471730 52006 471836 52034
rect 470784 48816 470836 48822
rect 470784 48758 470836 48764
rect 470508 28280 470560 28286
rect 470508 28222 470560 28228
rect 469864 15904 469916 15910
rect 469864 15846 469916 15852
rect 471808 5370 471836 52006
rect 471888 48816 471940 48822
rect 471888 48758 471940 48764
rect 471796 5364 471848 5370
rect 471796 5306 471848 5312
rect 471900 3670 471928 48758
rect 472728 48754 472756 52020
rect 473648 48822 473676 52020
rect 473636 48816 473688 48822
rect 473636 48758 473688 48764
rect 472716 48748 472768 48754
rect 472716 48690 472768 48696
rect 474568 5302 474596 52020
rect 475502 52006 476068 52034
rect 474648 48816 474700 48822
rect 474648 48758 474700 48764
rect 474556 5296 474608 5302
rect 474556 5238 474608 5244
rect 472716 4820 472768 4826
rect 472716 4762 472768 4768
rect 471520 3664 471572 3670
rect 471520 3606 471572 3612
rect 471888 3664 471940 3670
rect 471888 3606 471940 3612
rect 469232 3318 470364 3346
rect 470336 480 470364 3318
rect 471532 480 471560 3606
rect 472728 480 472756 4762
rect 474660 3466 474688 48758
rect 475384 48748 475436 48754
rect 475384 48690 475436 48696
rect 475396 19990 475424 48690
rect 476040 21418 476068 52006
rect 476500 49298 476528 52020
rect 476488 49292 476540 49298
rect 476488 49234 476540 49240
rect 476120 21480 476172 21486
rect 476120 21422 476172 21428
rect 476028 21412 476080 21418
rect 476028 21354 476080 21360
rect 475384 19984 475436 19990
rect 475384 19926 475436 19932
rect 473912 3460 473964 3466
rect 473912 3402 473964 3408
rect 474648 3460 474700 3466
rect 474648 3402 474700 3408
rect 473924 480 473952 3402
rect 475108 3392 475160 3398
rect 475108 3334 475160 3340
rect 475120 480 475148 3334
rect 476132 626 476160 21422
rect 477420 5166 477448 52020
rect 478354 52006 478828 52034
rect 478800 31074 478828 52006
rect 479260 48822 479288 52020
rect 480088 52006 480194 52034
rect 481206 52006 481588 52034
rect 479248 48816 479300 48822
rect 479248 48758 479300 48764
rect 478788 31068 478840 31074
rect 478788 31010 478840 31016
rect 479892 6180 479944 6186
rect 479892 6122 479944 6128
rect 477408 5160 477460 5166
rect 477408 5102 477460 5108
rect 478696 4072 478748 4078
rect 478696 4014 478748 4020
rect 477500 3324 477552 3330
rect 477500 3266 477552 3272
rect 476132 598 476344 626
rect 476316 480 476344 598
rect 477512 480 477540 3266
rect 478708 480 478736 4014
rect 479904 480 479932 6122
rect 480088 5098 480116 52006
rect 480168 48816 480220 48822
rect 480168 48758 480220 48764
rect 480076 5092 480128 5098
rect 480076 5034 480128 5040
rect 480180 3262 480208 48758
rect 481560 22778 481588 52006
rect 482112 49230 482140 52020
rect 482100 49224 482152 49230
rect 482100 49166 482152 49172
rect 482284 49020 482336 49026
rect 482284 48962 482336 48968
rect 481548 22772 481600 22778
rect 481548 22714 481600 22720
rect 482296 6186 482324 48962
rect 483032 48822 483060 52020
rect 483966 52006 484256 52034
rect 483020 48816 483072 48822
rect 483020 48758 483072 48764
rect 484228 40730 484256 52006
rect 484872 48822 484900 52020
rect 484308 48816 484360 48822
rect 484308 48758 484360 48764
rect 484860 48816 484912 48822
rect 484860 48758 484912 48764
rect 485688 48816 485740 48822
rect 485688 48758 485740 48764
rect 484216 40724 484268 40730
rect 484216 40666 484268 40672
rect 483480 6248 483532 6254
rect 483480 6190 483532 6196
rect 482284 6180 482336 6186
rect 482284 6122 482336 6128
rect 481088 4140 481140 4146
rect 481088 4082 481140 4088
rect 480168 3256 480220 3262
rect 480168 3198 480220 3204
rect 481100 480 481128 4082
rect 482282 3496 482338 3505
rect 482282 3431 482338 3440
rect 482296 480 482324 3431
rect 483492 480 483520 6190
rect 484320 5234 484348 48758
rect 484400 22840 484452 22846
rect 484400 22782 484452 22788
rect 484308 5228 484360 5234
rect 484308 5170 484360 5176
rect 484412 3346 484440 22782
rect 484412 3318 484624 3346
rect 485700 3330 485728 48758
rect 485884 48550 485912 52020
rect 486818 52006 487016 52034
rect 485872 48544 485924 48550
rect 485872 48486 485924 48492
rect 486988 37942 487016 52006
rect 487724 49162 487752 52020
rect 488658 52006 489040 52034
rect 489578 52006 489776 52034
rect 490590 52006 491248 52034
rect 487712 49156 487764 49162
rect 487712 49098 487764 49104
rect 487068 48544 487120 48550
rect 487068 48486 487120 48492
rect 486976 37936 487028 37942
rect 486976 37878 487028 37884
rect 486976 7676 487028 7682
rect 486976 7618 487028 7624
rect 485780 3936 485832 3942
rect 485780 3878 485832 3884
rect 484596 480 484624 3318
rect 485688 3324 485740 3330
rect 485688 3266 485740 3272
rect 485792 480 485820 3878
rect 486988 480 487016 7618
rect 487080 4962 487108 48486
rect 489012 48346 489040 52006
rect 489000 48340 489052 48346
rect 489000 48282 489052 48288
rect 489644 48340 489696 48346
rect 489644 48282 489696 48288
rect 489656 48210 489684 48282
rect 489644 48204 489696 48210
rect 489644 48146 489696 48152
rect 487160 47592 487212 47598
rect 487160 47534 487212 47540
rect 487172 38622 487200 47534
rect 489748 41478 489776 52006
rect 489736 41472 489788 41478
rect 489736 41414 489788 41420
rect 489736 41336 489788 41342
rect 489736 41278 489788 41284
rect 487160 38616 487212 38622
rect 487160 38558 487212 38564
rect 489644 31748 489696 31754
rect 489644 31690 489696 31696
rect 487160 29028 487212 29034
rect 487160 28970 487212 28976
rect 487172 19310 487200 28970
rect 489656 26874 489684 31690
rect 489748 29646 489776 41278
rect 489828 38684 489880 38690
rect 489828 38626 489880 38632
rect 489840 31754 489868 38626
rect 489828 31748 489880 31754
rect 489828 31690 489880 31696
rect 489736 29640 489788 29646
rect 489736 29582 489788 29588
rect 489656 26846 489776 26874
rect 487160 19304 487212 19310
rect 487160 19246 487212 19252
rect 489748 12458 489776 26846
rect 489656 12430 489776 12458
rect 487160 9716 487212 9722
rect 487160 9658 487212 9664
rect 487068 4956 487120 4962
rect 487068 4898 487120 4904
rect 487172 2938 487200 9658
rect 489656 5030 489684 12430
rect 490564 9036 490616 9042
rect 490564 8978 490616 8984
rect 489644 5024 489696 5030
rect 489644 4966 489696 4972
rect 489368 4004 489420 4010
rect 489368 3946 489420 3952
rect 487080 2910 487200 2938
rect 487080 610 487108 2910
rect 487068 604 487120 610
rect 487068 546 487120 552
rect 488172 604 488224 610
rect 488172 546 488224 552
rect 488184 480 488212 546
rect 489380 480 489408 3946
rect 490576 480 490604 8978
rect 491220 3942 491248 52006
rect 491496 48550 491524 52020
rect 492430 52006 492536 52034
rect 491484 48544 491536 48550
rect 491484 48486 491536 48492
rect 492508 36582 492536 52006
rect 493336 49094 493364 52020
rect 493324 49088 493376 49094
rect 493324 49030 493376 49036
rect 492588 48544 492640 48550
rect 492588 48486 492640 48492
rect 492496 36576 492548 36582
rect 492496 36518 492548 36524
rect 491300 24132 491352 24138
rect 491300 24074 491352 24080
rect 491208 3936 491260 3942
rect 491208 3878 491260 3884
rect 491312 2938 491340 24074
rect 492600 4894 492628 48486
rect 494256 48346 494284 52020
rect 495268 49722 495296 52020
rect 496202 52006 496768 52034
rect 495176 49694 495296 49722
rect 495176 48346 495204 49694
rect 494244 48340 494296 48346
rect 494244 48282 494296 48288
rect 495072 48340 495124 48346
rect 495072 48282 495124 48288
rect 495164 48340 495216 48346
rect 495164 48282 495216 48288
rect 496084 48340 496136 48346
rect 496084 48282 496136 48288
rect 495084 48226 495112 48282
rect 494992 48198 495112 48226
rect 494992 41290 495020 48198
rect 494992 41262 495112 41290
rect 495084 31754 495112 41262
rect 495072 31748 495124 31754
rect 495072 31690 495124 31696
rect 495256 31748 495308 31754
rect 495256 31690 495308 31696
rect 495268 22166 495296 31690
rect 495256 22160 495308 22166
rect 495256 22102 495308 22108
rect 495256 22024 495308 22030
rect 495256 21966 495308 21972
rect 494060 17264 494112 17270
rect 494060 17206 494112 17212
rect 494072 7682 494100 17206
rect 495268 12458 495296 21966
rect 496096 17270 496124 48282
rect 496084 17264 496136 17270
rect 496084 17206 496136 17212
rect 495176 12430 495296 12458
rect 494152 10328 494204 10334
rect 494152 10270 494204 10276
rect 494060 7676 494112 7682
rect 494060 7618 494112 7624
rect 492588 4888 492640 4894
rect 492588 4830 492640 4836
rect 492956 3868 493008 3874
rect 492956 3810 493008 3816
rect 491220 2910 491340 2938
rect 491220 610 491248 2910
rect 491208 604 491260 610
rect 491208 546 491260 552
rect 491760 604 491812 610
rect 491760 546 491812 552
rect 491772 480 491800 546
rect 492968 480 492996 3810
rect 494164 480 494192 10270
rect 495176 4826 495204 12430
rect 495348 7676 495400 7682
rect 495348 7618 495400 7624
rect 495164 4820 495216 4826
rect 495164 4762 495216 4768
rect 495360 480 495388 7618
rect 496740 4146 496768 52006
rect 497108 47598 497136 52020
rect 497096 47592 497148 47598
rect 497096 47534 497148 47540
rect 498028 35222 498056 52020
rect 498948 49026 498976 52020
rect 498936 49020 498988 49026
rect 498936 48962 498988 48968
rect 499960 46238 499988 52020
rect 498200 46232 498252 46238
rect 498200 46174 498252 46180
rect 499948 46232 500000 46238
rect 499948 46174 500000 46180
rect 498016 35216 498068 35222
rect 498016 35158 498068 35164
rect 497740 6180 497792 6186
rect 497740 6122 497792 6128
rect 496728 4140 496780 4146
rect 496728 4082 496780 4088
rect 496544 3732 496596 3738
rect 496544 3674 496596 3680
rect 496556 480 496584 3674
rect 497752 480 497780 6122
rect 498212 3346 498240 46174
rect 500880 13122 500908 52020
rect 501814 52006 502288 52034
rect 500868 13116 500920 13122
rect 500868 13058 500920 13064
rect 500960 11756 501012 11762
rect 500960 11698 501012 11704
rect 500130 3360 500186 3369
rect 498212 3318 498976 3346
rect 498948 480 498976 3318
rect 500972 3346 501000 11698
rect 502260 4078 502288 52006
rect 502720 44878 502748 52020
rect 502708 44872 502760 44878
rect 502708 44814 502760 44820
rect 503640 25566 503668 52020
rect 504666 52006 505048 52034
rect 502432 25560 502484 25566
rect 502432 25502 502484 25508
rect 503628 25560 503680 25566
rect 503628 25502 503680 25508
rect 502248 4072 502300 4078
rect 502248 4014 502300 4020
rect 500972 3318 501276 3346
rect 500130 3295 500186 3304
rect 500144 480 500172 3295
rect 501248 480 501276 3318
rect 502444 480 502472 25502
rect 503720 13184 503772 13190
rect 503720 13126 503772 13132
rect 503628 3800 503680 3806
rect 503628 3742 503680 3748
rect 503640 480 503668 3742
rect 503732 3346 503760 13126
rect 505020 4010 505048 52006
rect 505572 48346 505600 52020
rect 506492 48822 506520 52020
rect 507426 52006 507808 52034
rect 506480 48816 506532 48822
rect 506480 48758 506532 48764
rect 507676 48816 507728 48822
rect 507676 48758 507728 48764
rect 505560 48340 505612 48346
rect 505560 48282 505612 48288
rect 506388 48340 506440 48346
rect 506388 48282 506440 48288
rect 505100 26920 505152 26926
rect 505100 26862 505152 26868
rect 505008 4004 505060 4010
rect 505008 3946 505060 3952
rect 505112 3346 505140 26862
rect 506400 6186 506428 48282
rect 507688 33794 507716 48758
rect 507676 33788 507728 33794
rect 507676 33730 507728 33736
rect 506388 6180 506440 6186
rect 506388 6122 506440 6128
rect 507780 3942 507808 52006
rect 508332 48346 508360 52020
rect 509344 48686 509372 52020
rect 510278 52006 510568 52034
rect 509332 48680 509384 48686
rect 509332 48622 509384 48628
rect 510436 48680 510488 48686
rect 510436 48622 510488 48628
rect 508320 48340 508372 48346
rect 508320 48282 508372 48288
rect 509148 48340 509200 48346
rect 509148 48282 509200 48288
rect 509160 43450 509188 48282
rect 509148 43444 509200 43450
rect 509148 43386 509200 43392
rect 509240 18624 509292 18630
rect 509240 18566 509292 18572
rect 507860 14476 507912 14482
rect 507860 14418 507912 14424
rect 507768 3936 507820 3942
rect 507768 3878 507820 3884
rect 507216 3596 507268 3602
rect 507216 3538 507268 3544
rect 503732 3318 504864 3346
rect 505112 3318 506060 3346
rect 504836 480 504864 3318
rect 506032 480 506060 3318
rect 507228 480 507256 3538
rect 507872 3346 507900 14418
rect 509252 3346 509280 18566
rect 510448 14482 510476 48622
rect 510436 14476 510488 14482
rect 510436 14418 510488 14424
rect 510540 3874 510568 52006
rect 510712 49360 510764 49366
rect 510712 49302 510764 49308
rect 510528 3868 510580 3874
rect 510528 3810 510580 3816
rect 510724 3482 510752 49302
rect 511184 48822 511212 52020
rect 511172 48816 511224 48822
rect 511172 48758 511224 48764
rect 511908 48816 511960 48822
rect 511908 48758 511960 48764
rect 511920 42090 511948 48758
rect 512104 48686 512132 52020
rect 513038 52006 513328 52034
rect 514050 52006 514708 52034
rect 512092 48680 512144 48686
rect 512092 48622 512144 48628
rect 513196 48680 513248 48686
rect 513196 48622 513248 48628
rect 511908 42084 511960 42090
rect 511908 42026 511960 42032
rect 513208 12034 513236 48622
rect 513196 12028 513248 12034
rect 513196 11970 513248 11976
rect 513300 11914 513328 52006
rect 513116 11886 513328 11914
rect 512000 7608 512052 7614
rect 512000 7550 512052 7556
rect 510724 3454 510844 3482
rect 507872 3318 508452 3346
rect 509252 3318 509648 3346
rect 508424 480 508452 3318
rect 509620 480 509648 3318
rect 510816 480 510844 3454
rect 512012 480 512040 7550
rect 513116 3602 513144 11886
rect 513288 11824 513340 11830
rect 513288 11766 513340 11772
rect 513196 8968 513248 8974
rect 513196 8910 513248 8916
rect 513104 3596 513156 3602
rect 513104 3538 513156 3544
rect 513208 480 513236 8910
rect 513300 3738 513328 11766
rect 514680 8974 514708 52006
rect 514956 48822 514984 52020
rect 515890 52006 515996 52034
rect 516810 52006 517468 52034
rect 514944 48816 514996 48822
rect 514944 48758 514996 48764
rect 514760 15904 514812 15910
rect 514760 15846 514812 15852
rect 514668 8968 514720 8974
rect 514668 8910 514720 8916
rect 513288 3732 513340 3738
rect 513288 3674 513340 3680
rect 514392 3528 514444 3534
rect 514392 3470 514444 3476
rect 514404 480 514432 3470
rect 514772 3346 514800 15846
rect 515968 3534 515996 52006
rect 516048 48816 516100 48822
rect 516048 48758 516100 48764
rect 516060 3806 516088 48758
rect 516140 28280 516192 28286
rect 516140 28222 516192 28228
rect 516048 3800 516100 3806
rect 516048 3742 516100 3748
rect 515956 3528 516008 3534
rect 515956 3470 516008 3476
rect 516152 3346 516180 28222
rect 517440 11762 517468 52006
rect 517716 48822 517744 52020
rect 517704 48816 517756 48822
rect 517704 48758 517756 48764
rect 517428 11756 517480 11762
rect 517428 11698 517480 11704
rect 517888 3664 517940 3670
rect 517888 3606 517940 3612
rect 514772 3318 515628 3346
rect 516152 3318 516824 3346
rect 515600 480 515628 3318
rect 516796 480 516824 3318
rect 517900 480 517928 3606
rect 518728 3369 518756 52020
rect 519662 52006 520228 52034
rect 518808 48816 518860 48822
rect 518808 48758 518860 48764
rect 518820 3670 518848 48758
rect 520200 10334 520228 52006
rect 520568 48822 520596 52020
rect 521502 52006 521608 52034
rect 520556 48816 520608 48822
rect 520556 48758 520608 48764
rect 521476 48816 521528 48822
rect 521476 48758 521528 48764
rect 520372 19984 520424 19990
rect 520372 19926 520424 19932
rect 520188 10328 520240 10334
rect 520188 10270 520240 10276
rect 519084 5364 519136 5370
rect 519084 5306 519136 5312
rect 518808 3664 518860 3670
rect 518808 3606 518860 3612
rect 518714 3360 518770 3369
rect 518714 3295 518770 3304
rect 519096 480 519124 5306
rect 520384 3482 520412 19926
rect 520292 3454 520412 3482
rect 521488 3482 521516 48758
rect 521580 3641 521608 52006
rect 523040 21412 523092 21418
rect 523040 21354 523092 21360
rect 522672 5296 522724 5302
rect 522672 5238 522724 5244
rect 521566 3632 521622 3641
rect 521566 3567 521622 3576
rect 521488 3466 521608 3482
rect 521384 3460 521436 3466
rect 520292 480 520320 3454
rect 521488 3460 521620 3466
rect 521488 3454 521568 3460
rect 521384 3402 521436 3408
rect 521568 3402 521620 3408
rect 521396 3346 521424 3402
rect 521396 3318 521516 3346
rect 521488 480 521516 3318
rect 522684 480 522712 5238
rect 523052 3346 523080 21354
rect 523696 8294 523724 58647
rect 523788 24818 523816 71975
rect 523880 40050 523908 85303
rect 523972 55214 524000 98631
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86057 580212 86906
rect 580170 86048 580226 86057
rect 580170 85983 580226 85992
rect 580172 71732 580224 71738
rect 580172 71674 580224 71680
rect 580184 70417 580212 71674
rect 580170 70408 580226 70417
rect 580170 70343 580226 70352
rect 523960 55208 524012 55214
rect 523960 55150 524012 55156
rect 580172 55208 580224 55214
rect 580172 55150 580224 55156
rect 580184 54777 580212 55150
rect 580170 54768 580226 54777
rect 580170 54703 580226 54712
rect 524420 49292 524472 49298
rect 524420 49234 524472 49240
rect 523868 40044 523920 40050
rect 523868 39986 523920 39992
rect 523776 24812 523828 24818
rect 523776 24754 523828 24760
rect 523684 8288 523736 8294
rect 523684 8230 523736 8236
rect 524432 3346 524460 49234
rect 531320 49224 531372 49230
rect 531320 49166 531372 49172
rect 527180 31068 527232 31074
rect 527180 31010 527232 31016
rect 526260 5160 526312 5166
rect 526260 5102 526312 5108
rect 523052 3318 523908 3346
rect 524432 3318 525104 3346
rect 523880 480 523908 3318
rect 525076 480 525104 3318
rect 526272 480 526300 5102
rect 527192 3346 527220 31010
rect 529940 22772 529992 22778
rect 529940 22714 529992 22720
rect 529848 5092 529900 5098
rect 529848 5034 529900 5040
rect 527192 3318 527496 3346
rect 527468 480 527496 3318
rect 528652 3256 528704 3262
rect 528652 3198 528704 3204
rect 528664 480 528692 3198
rect 529860 480 529888 5034
rect 529952 3482 529980 22714
rect 531332 3482 531360 49166
rect 538220 49156 538272 49162
rect 538220 49098 538272 49104
rect 534080 40724 534132 40730
rect 534080 40666 534132 40672
rect 533436 5228 533488 5234
rect 533436 5170 533488 5176
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 5170
rect 534092 3482 534120 40666
rect 536840 37936 536892 37942
rect 536840 37878 536892 37884
rect 534092 3454 534580 3482
rect 534552 480 534580 3454
rect 536852 3330 536880 37878
rect 536932 4956 536984 4962
rect 536932 4898 536984 4904
rect 535736 3324 535788 3330
rect 535736 3266 535788 3272
rect 536840 3324 536892 3330
rect 536840 3266 536892 3272
rect 535748 480 535776 3266
rect 536944 480 536972 4898
rect 538232 3482 538260 49098
rect 546500 49088 546552 49094
rect 546500 49030 546552 49036
rect 545120 36576 545172 36582
rect 545120 36518 545172 36524
rect 540980 29640 541032 29646
rect 540980 29582 541032 29588
rect 540520 5160 540572 5166
rect 540520 5102 540572 5108
rect 538232 3454 539364 3482
rect 538128 3324 538180 3330
rect 538128 3266 538180 3272
rect 538140 480 538168 3266
rect 539336 480 539364 3454
rect 540532 480 540560 5102
rect 540992 3482 541020 29582
rect 544108 4888 544160 4894
rect 544108 4830 544160 4836
rect 540992 3454 541756 3482
rect 541728 480 541756 3454
rect 542912 3392 542964 3398
rect 542912 3334 542964 3340
rect 542924 480 542952 3334
rect 544120 480 544148 4830
rect 545132 3482 545160 36518
rect 545132 3454 545344 3482
rect 545316 480 545344 3454
rect 546512 480 546540 49030
rect 553400 49020 553452 49026
rect 553400 48962 553452 48968
rect 550640 47592 550692 47598
rect 550640 47534 550692 47540
rect 547880 17264 547932 17270
rect 547880 17206 547932 17212
rect 547696 4820 547748 4826
rect 547696 4762 547748 4768
rect 547708 480 547736 4762
rect 547892 3482 547920 17206
rect 550088 4140 550140 4146
rect 550088 4082 550140 4088
rect 547892 3454 548932 3482
rect 548904 480 548932 3454
rect 550100 480 550128 4082
rect 550652 3482 550680 47534
rect 552020 35216 552072 35222
rect 552020 35158 552072 35164
rect 552032 3482 552060 35158
rect 553412 3482 553440 48962
rect 554780 46232 554832 46238
rect 554780 46174 554832 46180
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 553412 3454 553624 3482
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3454
rect 554792 480 554820 46174
rect 557540 44872 557592 44878
rect 557540 44814 557592 44820
rect 554872 13116 554924 13122
rect 554872 13058 554924 13064
rect 554884 3482 554912 13058
rect 557172 4072 557224 4078
rect 557172 4014 557224 4020
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 4014
rect 557552 3482 557580 44814
rect 564440 43444 564492 43450
rect 564440 43386 564492 43392
rect 563152 33788 563204 33794
rect 563152 33730 563204 33736
rect 558920 25560 558972 25566
rect 558920 25502 558972 25508
rect 558932 3482 558960 25502
rect 561956 6180 562008 6186
rect 561956 6122 562008 6128
rect 560760 4004 560812 4010
rect 560760 3946 560812 3952
rect 557552 3454 558408 3482
rect 558932 3454 559604 3482
rect 558380 480 558408 3454
rect 559576 480 559604 3454
rect 560772 480 560800 3946
rect 561968 480 561996 6122
rect 563164 480 563192 33730
rect 564348 3936 564400 3942
rect 564348 3878 564400 3884
rect 564360 480 564388 3878
rect 564452 3482 564480 43386
rect 568580 42084 568632 42090
rect 568580 42026 568632 42032
rect 565820 14476 565872 14482
rect 565820 14418 565872 14424
rect 565832 3482 565860 14418
rect 567844 3868 567896 3874
rect 567844 3810 567896 3816
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3810
rect 568592 3482 568620 42026
rect 580172 40044 580224 40050
rect 580172 39986 580224 39992
rect 580184 39137 580212 39986
rect 580170 39128 580226 39137
rect 580170 39063 580226 39072
rect 580172 24812 580224 24818
rect 580172 24754 580224 24760
rect 580184 23497 580212 24754
rect 580170 23488 580226 23497
rect 580170 23423 580226 23432
rect 574744 11756 574796 11762
rect 574744 11698 574796 11704
rect 572628 8968 572680 8974
rect 572628 8910 572680 8916
rect 570236 3732 570288 3738
rect 570236 3674 570288 3680
rect 568592 3454 569080 3482
rect 569052 480 569080 3454
rect 570248 480 570276 3674
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 571444 480 571472 3538
rect 572640 480 572668 8910
rect 573824 3800 573876 3806
rect 573824 3742 573876 3748
rect 573836 480 573864 3742
rect 574756 3534 574784 11698
rect 579620 10328 579672 10334
rect 579620 10270 579672 10276
rect 577412 3664 577464 3670
rect 577412 3606 577464 3612
rect 575020 3596 575072 3602
rect 575020 3538 575072 3544
rect 574744 3528 574796 3534
rect 574744 3470 574796 3476
rect 575032 480 575060 3538
rect 576216 3528 576268 3534
rect 576216 3470 576268 3476
rect 576228 480 576256 3470
rect 577424 480 577452 3606
rect 578606 3360 578662 3369
rect 578606 3295 578662 3304
rect 578620 480 578648 3295
rect 579632 610 579660 10270
rect 580172 8288 580224 8294
rect 580172 8230 580224 8236
rect 580184 7857 580212 8230
rect 580170 7848 580226 7857
rect 580170 7783 580226 7792
rect 582194 3632 582250 3641
rect 582194 3567 582250 3576
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 579620 604 579672 610
rect 579620 546 579672 552
rect 579804 604 579856 610
rect 579804 546 579856 552
rect 579816 480 579844 546
rect 581012 480 581040 3402
rect 582208 480 582236 3567
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 695408 3478 695464
rect 3514 678680 3570 678736
rect 3606 661952 3662 662008
rect 3422 628360 3478 628416
rect 580170 695952 580226 696008
rect 3698 645224 3754 645280
rect 3514 611632 3570 611688
rect 3422 578176 3478 578232
rect 580170 680348 580172 680368
rect 580172 680348 580224 680368
rect 580224 680348 580226 680368
rect 523682 645224 523738 645280
rect 59358 644680 59414 644736
rect 59358 630400 59414 630456
rect 59358 616120 59414 616176
rect 523130 605240 523186 605296
rect 59358 601840 59414 601896
rect 3606 594904 3662 594960
rect 3514 561312 3570 561368
rect 580170 680312 580226 680348
rect 580262 664672 580318 664728
rect 580170 633428 580172 633448
rect 580172 633428 580224 633448
rect 580224 633428 580226 633448
rect 580170 633392 580226 633428
rect 523774 631896 523830 631952
rect 580354 649032 580410 649088
rect 524326 618568 524382 618624
rect 580262 617752 580318 617808
rect 580170 602112 580226 602168
rect 523682 591912 523738 591968
rect 59358 587560 59414 587616
rect 59358 573280 59414 573336
rect 59358 559000 59414 559056
rect 580170 586508 580172 586528
rect 580172 586508 580224 586528
rect 580224 586508 580226 586528
rect 580170 586472 580226 586508
rect 524326 578584 524382 578640
rect 580262 570832 580318 570888
rect 523774 565256 523830 565312
rect 580170 555192 580226 555248
rect 523682 551928 523738 551984
rect 59358 544720 59414 544776
rect 3606 544584 3662 544640
rect 3422 527856 3478 527912
rect 523682 538600 523738 538656
rect 59358 530440 59414 530496
rect 59358 516160 59414 516216
rect 580170 539588 580172 539608
rect 580172 539588 580224 539608
rect 580224 539588 580226 539608
rect 580170 539552 580226 539588
rect 523774 525272 523830 525328
rect 580170 523912 580226 523968
rect 523682 511944 523738 512000
rect 3514 511128 3570 511184
rect 3422 494264 3478 494320
rect 59358 501880 59414 501936
rect 59358 487600 59414 487656
rect 580170 508272 580226 508328
rect 523774 498616 523830 498672
rect 580170 492668 580172 492688
rect 580172 492668 580224 492688
rect 580224 492668 580226 492688
rect 523682 485288 523738 485344
rect 3514 477536 3570 477592
rect 3422 460808 3478 460864
rect 59358 473320 59414 473376
rect 59358 459040 59414 459096
rect 580170 492632 580226 492668
rect 580170 476992 580226 477048
rect 523774 471960 523830 472016
rect 580170 461352 580226 461408
rect 523682 458632 523738 458688
rect 59358 444760 59414 444816
rect 3422 444080 3478 444136
rect 580170 445748 580172 445768
rect 580172 445748 580224 445768
rect 580224 445748 580226 445768
rect 580170 445712 580226 445748
rect 523774 445304 523830 445360
rect 523682 431976 523738 432032
rect 59358 430516 59360 430536
rect 59360 430516 59412 430536
rect 59412 430516 59414 430536
rect 59358 430480 59414 430516
rect 580170 430072 580226 430128
rect 3422 427216 3478 427272
rect 523682 418648 523738 418704
rect 59358 416200 59414 416256
rect 580170 414432 580226 414488
rect 3422 410488 3478 410544
rect 523682 405320 523738 405376
rect 59358 401920 59414 401976
rect 580170 398828 580172 398848
rect 580172 398828 580224 398848
rect 580224 398828 580226 398848
rect 3882 393760 3938 393816
rect 580170 398792 580226 398828
rect 523682 391992 523738 392048
rect 59358 387640 59414 387696
rect 580170 383152 580226 383208
rect 523130 378664 523186 378720
rect 3422 377032 3478 377088
rect 59358 373360 59414 373416
rect 580170 367512 580226 367568
rect 523314 365336 523370 365392
rect 3422 360304 3478 360360
rect 59358 359080 59414 359136
rect 524326 351872 524382 351928
rect 580170 351872 580226 351928
rect 59358 344664 59414 344720
rect 3422 343440 3478 343496
rect 523406 338544 523462 338600
rect 580170 336232 580226 336288
rect 59358 330384 59414 330440
rect 3330 326712 3386 326768
rect 523130 325216 523186 325272
rect 580170 320592 580226 320648
rect 60002 316104 60058 316160
rect 523682 311888 523738 311944
rect 3422 309984 3478 310040
rect 580170 304952 580226 305008
rect 60002 301824 60058 301880
rect 523682 298560 523738 298616
rect 3146 293256 3202 293312
rect 580170 289312 580226 289368
rect 60002 287544 60058 287600
rect 523682 285232 523738 285288
rect 3422 276392 3478 276448
rect 580170 273672 580226 273728
rect 60002 273264 60058 273320
rect 523682 271904 523738 271960
rect 3422 259664 3478 259720
rect 60002 258984 60058 259040
rect 523774 258576 523830 258632
rect 523682 245248 523738 245304
rect 60094 244704 60150 244760
rect 3422 242936 3478 242992
rect 60002 230424 60058 230480
rect 3422 226244 3424 226264
rect 3424 226244 3476 226264
rect 3476 226244 3478 226264
rect 3422 226208 3478 226244
rect 580170 258032 580226 258088
rect 580170 242392 580226 242448
rect 523774 231920 523830 231976
rect 523682 218592 523738 218648
rect 60094 216144 60150 216200
rect 3422 209344 3478 209400
rect 60002 201864 60058 201920
rect 3514 192616 3570 192672
rect 580170 226752 580226 226808
rect 580170 211112 580226 211168
rect 523774 205264 523830 205320
rect 523682 191936 523738 191992
rect 60186 187584 60242 187640
rect 3422 175888 3478 175944
rect 60094 173304 60150 173360
rect 3146 159160 3202 159216
rect 60002 159024 60058 159080
rect 3238 142296 3294 142352
rect 580170 195472 580226 195528
rect 580170 179832 580226 179888
rect 523866 178608 523922 178664
rect 523774 165280 523830 165336
rect 523682 151952 523738 152008
rect 60186 144744 60242 144800
rect 60094 130464 60150 130520
rect 3238 125568 3294 125624
rect 60002 116184 60058 116240
rect 3422 108840 3478 108896
rect 3330 92112 3386 92168
rect 580170 164192 580226 164248
rect 580170 148552 580226 148608
rect 523866 138624 523922 138680
rect 523774 125296 523830 125352
rect 523682 111968 523738 112024
rect 60278 101904 60334 101960
rect 60186 87624 60242 87680
rect 3422 75248 3478 75304
rect 60094 73344 60150 73400
rect 60002 59064 60058 59120
rect 3054 58520 3110 58576
rect 3422 41792 3478 41848
rect 3422 25064 3478 25120
rect 3422 8336 3478 8392
rect 19522 3304 19578 3360
rect 25502 3440 25558 3496
rect 580170 132912 580226 132968
rect 580170 117272 580226 117328
rect 580170 101632 580226 101688
rect 523958 98640 524014 98696
rect 523866 85312 523922 85368
rect 523774 71984 523830 72040
rect 523682 58656 523738 58712
rect 77482 3304 77538 3360
rect 80150 19216 80206 19272
rect 80426 19216 80482 19272
rect 81530 3440 81586 3496
rect 82634 3304 82690 3360
rect 86130 3440 86186 3496
rect 110050 38800 110106 38856
rect 109314 38664 109370 38720
rect 127070 3304 127126 3360
rect 129922 3440 129978 3496
rect 190826 3304 190882 3360
rect 194414 3440 194470 3496
rect 203890 38800 203946 38856
rect 203154 38664 203210 38720
rect 212630 3304 212686 3360
rect 215390 3440 215446 3496
rect 442906 3440 442962 3496
rect 456706 3304 456762 3360
rect 482282 3440 482338 3496
rect 500130 3304 500186 3360
rect 518714 3304 518770 3360
rect 521566 3576 521622 3632
rect 580170 85992 580226 86048
rect 580170 70352 580226 70408
rect 580170 54712 580226 54768
rect 580170 39072 580226 39128
rect 580170 23432 580226 23488
rect 578606 3304 578662 3360
rect 580170 7792 580226 7848
rect 582194 3576 582250 3632
<< metal3 >>
rect 580165 696010 580231 696013
rect 583520 696010 584960 696100
rect 580165 696008 584960 696010
rect 580165 695952 580170 696008
rect 580226 695952 584960 696008
rect 580165 695950 584960 695952
rect 580165 695947 580231 695950
rect 583520 695860 584960 695950
rect -960 695466 480 695556
rect 3417 695466 3483 695469
rect -960 695464 3483 695466
rect -960 695408 3422 695464
rect 3478 695408 3483 695464
rect -960 695406 3483 695408
rect -960 695316 480 695406
rect 3417 695403 3483 695406
rect 580165 680370 580231 680373
rect 583520 680370 584960 680460
rect 580165 680368 584960 680370
rect 580165 680312 580170 680368
rect 580226 680312 584960 680368
rect 580165 680310 584960 680312
rect 580165 680307 580231 680310
rect 583520 680220 584960 680310
rect -960 678738 480 678828
rect 3509 678738 3575 678741
rect -960 678736 3575 678738
rect -960 678680 3514 678736
rect 3570 678680 3575 678736
rect -960 678678 3575 678680
rect -960 678588 480 678678
rect 3509 678675 3575 678678
rect 580257 664730 580323 664733
rect 583520 664730 584960 664820
rect 580257 664728 584960 664730
rect 580257 664672 580262 664728
rect 580318 664672 584960 664728
rect 580257 664670 584960 664672
rect 580257 664667 580323 664670
rect 583520 664580 584960 664670
rect -960 662010 480 662100
rect 3601 662010 3667 662013
rect -960 662008 3667 662010
rect -960 661952 3606 662008
rect 3662 661952 3667 662008
rect -960 661950 3667 661952
rect -960 661860 480 661950
rect 3601 661947 3667 661950
rect 580349 649090 580415 649093
rect 583520 649090 584960 649180
rect 580349 649088 584960 649090
rect 580349 649032 580354 649088
rect 580410 649032 584960 649088
rect 580349 649030 584960 649032
rect 580349 649027 580415 649030
rect 583520 648940 584960 649030
rect -960 645282 480 645372
rect 3693 645282 3759 645285
rect 523677 645282 523743 645285
rect -960 645280 3759 645282
rect -960 645224 3698 645280
rect 3754 645224 3759 645280
rect -960 645222 3759 645224
rect 521916 645280 523743 645282
rect 521916 645224 523682 645280
rect 523738 645224 523743 645280
rect 521916 645222 523743 645224
rect -960 645132 480 645222
rect 3693 645219 3759 645222
rect 523677 645219 523743 645222
rect 59353 644738 59419 644741
rect 59353 644736 62100 644738
rect 59353 644680 59358 644736
rect 59414 644680 62100 644736
rect 59353 644678 62100 644680
rect 59353 644675 59419 644678
rect 580165 633450 580231 633453
rect 583520 633450 584960 633540
rect 580165 633448 584960 633450
rect 580165 633392 580170 633448
rect 580226 633392 584960 633448
rect 580165 633390 584960 633392
rect 580165 633387 580231 633390
rect 583520 633300 584960 633390
rect 523769 631954 523835 631957
rect 521916 631952 523835 631954
rect 521916 631896 523774 631952
rect 523830 631896 523835 631952
rect 521916 631894 523835 631896
rect 523769 631891 523835 631894
rect 59353 630458 59419 630461
rect 59353 630456 62100 630458
rect 59353 630400 59358 630456
rect 59414 630400 62100 630456
rect 59353 630398 62100 630400
rect 59353 630395 59419 630398
rect -960 628418 480 628508
rect 3417 628418 3483 628421
rect -960 628416 3483 628418
rect -960 628360 3422 628416
rect 3478 628360 3483 628416
rect -960 628358 3483 628360
rect -960 628268 480 628358
rect 3417 628355 3483 628358
rect 524321 618626 524387 618629
rect 521916 618624 524387 618626
rect 521916 618568 524326 618624
rect 524382 618568 524387 618624
rect 521916 618566 524387 618568
rect 524321 618563 524387 618566
rect 580257 617810 580323 617813
rect 583520 617810 584960 617900
rect 580257 617808 584960 617810
rect 580257 617752 580262 617808
rect 580318 617752 584960 617808
rect 580257 617750 584960 617752
rect 580257 617747 580323 617750
rect 583520 617660 584960 617750
rect 59353 616178 59419 616181
rect 59353 616176 62100 616178
rect 59353 616120 59358 616176
rect 59414 616120 62100 616176
rect 59353 616118 62100 616120
rect 59353 616115 59419 616118
rect -960 611690 480 611780
rect 3509 611690 3575 611693
rect -960 611688 3575 611690
rect -960 611632 3514 611688
rect 3570 611632 3575 611688
rect -960 611630 3575 611632
rect -960 611540 480 611630
rect 3509 611627 3575 611630
rect 523125 605298 523191 605301
rect 521916 605296 523191 605298
rect 521916 605240 523130 605296
rect 523186 605240 523191 605296
rect 521916 605238 523191 605240
rect 523125 605235 523191 605238
rect 580165 602170 580231 602173
rect 583520 602170 584960 602260
rect 580165 602168 584960 602170
rect 580165 602112 580170 602168
rect 580226 602112 584960 602168
rect 580165 602110 584960 602112
rect 580165 602107 580231 602110
rect 583520 602020 584960 602110
rect 59353 601898 59419 601901
rect 59353 601896 62100 601898
rect 59353 601840 59358 601896
rect 59414 601840 62100 601896
rect 59353 601838 62100 601840
rect 59353 601835 59419 601838
rect -960 594962 480 595052
rect 3601 594962 3667 594965
rect -960 594960 3667 594962
rect -960 594904 3606 594960
rect 3662 594904 3667 594960
rect -960 594902 3667 594904
rect -960 594812 480 594902
rect 3601 594899 3667 594902
rect 523677 591970 523743 591973
rect 521916 591968 523743 591970
rect 521916 591912 523682 591968
rect 523738 591912 523743 591968
rect 521916 591910 523743 591912
rect 523677 591907 523743 591910
rect 59353 587618 59419 587621
rect 59353 587616 62100 587618
rect 59353 587560 59358 587616
rect 59414 587560 62100 587616
rect 59353 587558 62100 587560
rect 59353 587555 59419 587558
rect 580165 586530 580231 586533
rect 583520 586530 584960 586620
rect 580165 586528 584960 586530
rect 580165 586472 580170 586528
rect 580226 586472 584960 586528
rect 580165 586470 584960 586472
rect 580165 586467 580231 586470
rect 583520 586380 584960 586470
rect 524321 578642 524387 578645
rect 521916 578640 524387 578642
rect 521916 578584 524326 578640
rect 524382 578584 524387 578640
rect 521916 578582 524387 578584
rect 524321 578579 524387 578582
rect -960 578234 480 578324
rect 3417 578234 3483 578237
rect -960 578232 3483 578234
rect -960 578176 3422 578232
rect 3478 578176 3483 578232
rect -960 578174 3483 578176
rect -960 578084 480 578174
rect 3417 578171 3483 578174
rect 59353 573338 59419 573341
rect 59353 573336 62100 573338
rect 59353 573280 59358 573336
rect 59414 573280 62100 573336
rect 59353 573278 62100 573280
rect 59353 573275 59419 573278
rect 580257 570890 580323 570893
rect 583520 570890 584960 570980
rect 580257 570888 584960 570890
rect 580257 570832 580262 570888
rect 580318 570832 584960 570888
rect 580257 570830 584960 570832
rect 580257 570827 580323 570830
rect 583520 570740 584960 570830
rect 523769 565314 523835 565317
rect 521916 565312 523835 565314
rect 521916 565256 523774 565312
rect 523830 565256 523835 565312
rect 521916 565254 523835 565256
rect 523769 565251 523835 565254
rect -960 561370 480 561460
rect 3509 561370 3575 561373
rect -960 561368 3575 561370
rect -960 561312 3514 561368
rect 3570 561312 3575 561368
rect -960 561310 3575 561312
rect -960 561220 480 561310
rect 3509 561307 3575 561310
rect 59353 559058 59419 559061
rect 59353 559056 62100 559058
rect 59353 559000 59358 559056
rect 59414 559000 62100 559056
rect 59353 558998 62100 559000
rect 59353 558995 59419 558998
rect 580165 555250 580231 555253
rect 583520 555250 584960 555340
rect 580165 555248 584960 555250
rect 580165 555192 580170 555248
rect 580226 555192 584960 555248
rect 580165 555190 584960 555192
rect 580165 555187 580231 555190
rect 583520 555100 584960 555190
rect 523677 551986 523743 551989
rect 521916 551984 523743 551986
rect 521916 551928 523682 551984
rect 523738 551928 523743 551984
rect 521916 551926 523743 551928
rect 523677 551923 523743 551926
rect 59353 544778 59419 544781
rect 59353 544776 62100 544778
rect -960 544642 480 544732
rect 59353 544720 59358 544776
rect 59414 544720 62100 544776
rect 59353 544718 62100 544720
rect 59353 544715 59419 544718
rect 3601 544642 3667 544645
rect -960 544640 3667 544642
rect -960 544584 3606 544640
rect 3662 544584 3667 544640
rect -960 544582 3667 544584
rect -960 544492 480 544582
rect 3601 544579 3667 544582
rect 580165 539610 580231 539613
rect 583520 539610 584960 539700
rect 580165 539608 584960 539610
rect 580165 539552 580170 539608
rect 580226 539552 584960 539608
rect 580165 539550 584960 539552
rect 580165 539547 580231 539550
rect 583520 539460 584960 539550
rect 523677 538658 523743 538661
rect 521916 538656 523743 538658
rect 521916 538600 523682 538656
rect 523738 538600 523743 538656
rect 521916 538598 523743 538600
rect 523677 538595 523743 538598
rect 59353 530498 59419 530501
rect 59353 530496 62100 530498
rect 59353 530440 59358 530496
rect 59414 530440 62100 530496
rect 59353 530438 62100 530440
rect 59353 530435 59419 530438
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 523769 525330 523835 525333
rect 521916 525328 523835 525330
rect 521916 525272 523774 525328
rect 523830 525272 523835 525328
rect 521916 525270 523835 525272
rect 523769 525267 523835 525270
rect 580165 523970 580231 523973
rect 583520 523970 584960 524060
rect 580165 523968 584960 523970
rect 580165 523912 580170 523968
rect 580226 523912 584960 523968
rect 580165 523910 584960 523912
rect 580165 523907 580231 523910
rect 583520 523820 584960 523910
rect 59353 516218 59419 516221
rect 59353 516216 62100 516218
rect 59353 516160 59358 516216
rect 59414 516160 62100 516216
rect 59353 516158 62100 516160
rect 59353 516155 59419 516158
rect 523677 512002 523743 512005
rect 521916 512000 523743 512002
rect 521916 511944 523682 512000
rect 523738 511944 523743 512000
rect 521916 511942 523743 511944
rect 523677 511939 523743 511942
rect -960 511186 480 511276
rect 3509 511186 3575 511189
rect -960 511184 3575 511186
rect -960 511128 3514 511184
rect 3570 511128 3575 511184
rect -960 511126 3575 511128
rect -960 511036 480 511126
rect 3509 511123 3575 511126
rect 580165 508330 580231 508333
rect 583520 508330 584960 508420
rect 580165 508328 584960 508330
rect 580165 508272 580170 508328
rect 580226 508272 584960 508328
rect 580165 508270 584960 508272
rect 580165 508267 580231 508270
rect 583520 508180 584960 508270
rect 59353 501938 59419 501941
rect 59353 501936 62100 501938
rect 59353 501880 59358 501936
rect 59414 501880 62100 501936
rect 59353 501878 62100 501880
rect 59353 501875 59419 501878
rect 523769 498674 523835 498677
rect 521916 498672 523835 498674
rect 521916 498616 523774 498672
rect 523830 498616 523835 498672
rect 521916 498614 523835 498616
rect 523769 498611 523835 498614
rect -960 494322 480 494412
rect 3417 494322 3483 494325
rect -960 494320 3483 494322
rect -960 494264 3422 494320
rect 3478 494264 3483 494320
rect -960 494262 3483 494264
rect -960 494172 480 494262
rect 3417 494259 3483 494262
rect 580165 492690 580231 492693
rect 583520 492690 584960 492780
rect 580165 492688 584960 492690
rect 580165 492632 580170 492688
rect 580226 492632 584960 492688
rect 580165 492630 584960 492632
rect 580165 492627 580231 492630
rect 583520 492540 584960 492630
rect 59353 487658 59419 487661
rect 59353 487656 62100 487658
rect 59353 487600 59358 487656
rect 59414 487600 62100 487656
rect 59353 487598 62100 487600
rect 59353 487595 59419 487598
rect 523677 485346 523743 485349
rect 521916 485344 523743 485346
rect 521916 485288 523682 485344
rect 523738 485288 523743 485344
rect 521916 485286 523743 485288
rect 523677 485283 523743 485286
rect -960 477594 480 477684
rect 3509 477594 3575 477597
rect -960 477592 3575 477594
rect -960 477536 3514 477592
rect 3570 477536 3575 477592
rect -960 477534 3575 477536
rect -960 477444 480 477534
rect 3509 477531 3575 477534
rect 580165 477050 580231 477053
rect 583520 477050 584960 477140
rect 580165 477048 584960 477050
rect 580165 476992 580170 477048
rect 580226 476992 584960 477048
rect 580165 476990 584960 476992
rect 580165 476987 580231 476990
rect 583520 476900 584960 476990
rect 59353 473378 59419 473381
rect 59353 473376 62100 473378
rect 59353 473320 59358 473376
rect 59414 473320 62100 473376
rect 59353 473318 62100 473320
rect 59353 473315 59419 473318
rect 523769 472018 523835 472021
rect 521916 472016 523835 472018
rect 521916 471960 523774 472016
rect 523830 471960 523835 472016
rect 521916 471958 523835 471960
rect 523769 471955 523835 471958
rect 580165 461410 580231 461413
rect 583520 461410 584960 461500
rect 580165 461408 584960 461410
rect 580165 461352 580170 461408
rect 580226 461352 584960 461408
rect 580165 461350 584960 461352
rect 580165 461347 580231 461350
rect 583520 461260 584960 461350
rect -960 460866 480 460956
rect 3417 460866 3483 460869
rect -960 460864 3483 460866
rect -960 460808 3422 460864
rect 3478 460808 3483 460864
rect -960 460806 3483 460808
rect -960 460716 480 460806
rect 3417 460803 3483 460806
rect 59353 459098 59419 459101
rect 59353 459096 62100 459098
rect 59353 459040 59358 459096
rect 59414 459040 62100 459096
rect 59353 459038 62100 459040
rect 59353 459035 59419 459038
rect 523677 458690 523743 458693
rect 521916 458688 523743 458690
rect 521916 458632 523682 458688
rect 523738 458632 523743 458688
rect 521916 458630 523743 458632
rect 523677 458627 523743 458630
rect 580165 445770 580231 445773
rect 583520 445770 584960 445860
rect 580165 445768 584960 445770
rect 580165 445712 580170 445768
rect 580226 445712 584960 445768
rect 580165 445710 584960 445712
rect 580165 445707 580231 445710
rect 583520 445620 584960 445710
rect 523769 445362 523835 445365
rect 521916 445360 523835 445362
rect 521916 445304 523774 445360
rect 523830 445304 523835 445360
rect 521916 445302 523835 445304
rect 523769 445299 523835 445302
rect 59353 444818 59419 444821
rect 59353 444816 62100 444818
rect 59353 444760 59358 444816
rect 59414 444760 62100 444816
rect 59353 444758 62100 444760
rect 59353 444755 59419 444758
rect -960 444138 480 444228
rect 3417 444138 3483 444141
rect -960 444136 3483 444138
rect -960 444080 3422 444136
rect 3478 444080 3483 444136
rect -960 444078 3483 444080
rect -960 443988 480 444078
rect 3417 444075 3483 444078
rect 523677 432034 523743 432037
rect 521916 432032 523743 432034
rect 521916 431976 523682 432032
rect 523738 431976 523743 432032
rect 521916 431974 523743 431976
rect 523677 431971 523743 431974
rect 59353 430538 59419 430541
rect 59353 430536 62100 430538
rect 59353 430480 59358 430536
rect 59414 430480 62100 430536
rect 59353 430478 62100 430480
rect 59353 430475 59419 430478
rect 580165 430130 580231 430133
rect 583520 430130 584960 430220
rect 580165 430128 584960 430130
rect 580165 430072 580170 430128
rect 580226 430072 584960 430128
rect 580165 430070 584960 430072
rect 580165 430067 580231 430070
rect 583520 429980 584960 430070
rect -960 427274 480 427364
rect 3417 427274 3483 427277
rect -960 427272 3483 427274
rect -960 427216 3422 427272
rect 3478 427216 3483 427272
rect -960 427214 3483 427216
rect -960 427124 480 427214
rect 3417 427211 3483 427214
rect 523677 418706 523743 418709
rect 521916 418704 523743 418706
rect 521916 418648 523682 418704
rect 523738 418648 523743 418704
rect 521916 418646 523743 418648
rect 523677 418643 523743 418646
rect 59353 416258 59419 416261
rect 59353 416256 62100 416258
rect 59353 416200 59358 416256
rect 59414 416200 62100 416256
rect 59353 416198 62100 416200
rect 59353 416195 59419 416198
rect 580165 414490 580231 414493
rect 583520 414490 584960 414580
rect 580165 414488 584960 414490
rect 580165 414432 580170 414488
rect 580226 414432 584960 414488
rect 580165 414430 584960 414432
rect 580165 414427 580231 414430
rect 583520 414340 584960 414430
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 523677 405378 523743 405381
rect 521916 405376 523743 405378
rect 521916 405320 523682 405376
rect 523738 405320 523743 405376
rect 521916 405318 523743 405320
rect 523677 405315 523743 405318
rect 59353 401978 59419 401981
rect 59353 401976 62100 401978
rect 59353 401920 59358 401976
rect 59414 401920 62100 401976
rect 59353 401918 62100 401920
rect 59353 401915 59419 401918
rect 580165 398850 580231 398853
rect 583520 398850 584960 398940
rect 580165 398848 584960 398850
rect 580165 398792 580170 398848
rect 580226 398792 584960 398848
rect 580165 398790 584960 398792
rect 580165 398787 580231 398790
rect 583520 398700 584960 398790
rect -960 393818 480 393908
rect 3877 393818 3943 393821
rect -960 393816 3943 393818
rect -960 393760 3882 393816
rect 3938 393760 3943 393816
rect -960 393758 3943 393760
rect -960 393668 480 393758
rect 3877 393755 3943 393758
rect 523677 392050 523743 392053
rect 521916 392048 523743 392050
rect 521916 391992 523682 392048
rect 523738 391992 523743 392048
rect 521916 391990 523743 391992
rect 523677 391987 523743 391990
rect 59353 387698 59419 387701
rect 59353 387696 62100 387698
rect 59353 387640 59358 387696
rect 59414 387640 62100 387696
rect 59353 387638 62100 387640
rect 59353 387635 59419 387638
rect 580165 383210 580231 383213
rect 583520 383210 584960 383300
rect 580165 383208 584960 383210
rect 580165 383152 580170 383208
rect 580226 383152 584960 383208
rect 580165 383150 584960 383152
rect 580165 383147 580231 383150
rect 583520 383060 584960 383150
rect 523125 378722 523191 378725
rect 521916 378720 523191 378722
rect 521916 378664 523130 378720
rect 523186 378664 523191 378720
rect 521916 378662 523191 378664
rect 523125 378659 523191 378662
rect -960 377090 480 377180
rect 3417 377090 3483 377093
rect -960 377088 3483 377090
rect -960 377032 3422 377088
rect 3478 377032 3483 377088
rect -960 377030 3483 377032
rect -960 376940 480 377030
rect 3417 377027 3483 377030
rect 59353 373418 59419 373421
rect 59353 373416 62100 373418
rect 59353 373360 59358 373416
rect 59414 373360 62100 373416
rect 59353 373358 62100 373360
rect 59353 373355 59419 373358
rect 580165 367570 580231 367573
rect 583520 367570 584960 367660
rect 580165 367568 584960 367570
rect 580165 367512 580170 367568
rect 580226 367512 584960 367568
rect 580165 367510 584960 367512
rect 580165 367507 580231 367510
rect 583520 367420 584960 367510
rect 523309 365394 523375 365397
rect 521916 365392 523375 365394
rect 521916 365336 523314 365392
rect 523370 365336 523375 365392
rect 521916 365334 523375 365336
rect 523309 365331 523375 365334
rect -960 360362 480 360452
rect 3417 360362 3483 360365
rect -960 360360 3483 360362
rect -960 360304 3422 360360
rect 3478 360304 3483 360360
rect -960 360302 3483 360304
rect -960 360212 480 360302
rect 3417 360299 3483 360302
rect 59353 359138 59419 359141
rect 59353 359136 62100 359138
rect 59353 359080 59358 359136
rect 59414 359080 62100 359136
rect 59353 359078 62100 359080
rect 59353 359075 59419 359078
rect 524321 351930 524387 351933
rect 521916 351928 524387 351930
rect 521916 351872 524326 351928
rect 524382 351872 524387 351928
rect 521916 351870 524387 351872
rect 524321 351867 524387 351870
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 59353 344722 59419 344725
rect 59353 344720 62100 344722
rect 59353 344664 59358 344720
rect 59414 344664 62100 344720
rect 59353 344662 62100 344664
rect 59353 344659 59419 344662
rect -960 343498 480 343588
rect 3417 343498 3483 343501
rect -960 343496 3483 343498
rect -960 343440 3422 343496
rect 3478 343440 3483 343496
rect -960 343438 3483 343440
rect -960 343348 480 343438
rect 3417 343435 3483 343438
rect 523401 338602 523467 338605
rect 521916 338600 523467 338602
rect 521916 338544 523406 338600
rect 523462 338544 523467 338600
rect 521916 338542 523467 338544
rect 523401 338539 523467 338542
rect 580165 336290 580231 336293
rect 583520 336290 584960 336380
rect 580165 336288 584960 336290
rect 580165 336232 580170 336288
rect 580226 336232 584960 336288
rect 580165 336230 584960 336232
rect 580165 336227 580231 336230
rect 583520 336140 584960 336230
rect 59353 330442 59419 330445
rect 59353 330440 62100 330442
rect 59353 330384 59358 330440
rect 59414 330384 62100 330440
rect 59353 330382 62100 330384
rect 59353 330379 59419 330382
rect -960 326770 480 326860
rect 3325 326770 3391 326773
rect -960 326768 3391 326770
rect -960 326712 3330 326768
rect 3386 326712 3391 326768
rect -960 326710 3391 326712
rect -960 326620 480 326710
rect 3325 326707 3391 326710
rect 523125 325274 523191 325277
rect 521916 325272 523191 325274
rect 521916 325216 523130 325272
rect 523186 325216 523191 325272
rect 521916 325214 523191 325216
rect 523125 325211 523191 325214
rect 580165 320650 580231 320653
rect 583520 320650 584960 320740
rect 580165 320648 584960 320650
rect 580165 320592 580170 320648
rect 580226 320592 584960 320648
rect 580165 320590 584960 320592
rect 580165 320587 580231 320590
rect 583520 320500 584960 320590
rect 59997 316162 60063 316165
rect 59997 316160 62100 316162
rect 59997 316104 60002 316160
rect 60058 316104 62100 316160
rect 59997 316102 62100 316104
rect 59997 316099 60063 316102
rect 523677 311946 523743 311949
rect 521916 311944 523743 311946
rect 521916 311888 523682 311944
rect 523738 311888 523743 311944
rect 521916 311886 523743 311888
rect 523677 311883 523743 311886
rect -960 310042 480 310132
rect 3417 310042 3483 310045
rect -960 310040 3483 310042
rect -960 309984 3422 310040
rect 3478 309984 3483 310040
rect -960 309982 3483 309984
rect -960 309892 480 309982
rect 3417 309979 3483 309982
rect 580165 305010 580231 305013
rect 583520 305010 584960 305100
rect 580165 305008 584960 305010
rect 580165 304952 580170 305008
rect 580226 304952 584960 305008
rect 580165 304950 584960 304952
rect 580165 304947 580231 304950
rect 583520 304860 584960 304950
rect 59997 301882 60063 301885
rect 59997 301880 62100 301882
rect 59997 301824 60002 301880
rect 60058 301824 62100 301880
rect 59997 301822 62100 301824
rect 59997 301819 60063 301822
rect 523677 298618 523743 298621
rect 521916 298616 523743 298618
rect 521916 298560 523682 298616
rect 523738 298560 523743 298616
rect 521916 298558 523743 298560
rect 523677 298555 523743 298558
rect -960 293314 480 293404
rect 3141 293314 3207 293317
rect -960 293312 3207 293314
rect -960 293256 3146 293312
rect 3202 293256 3207 293312
rect -960 293254 3207 293256
rect -960 293164 480 293254
rect 3141 293251 3207 293254
rect 580165 289370 580231 289373
rect 583520 289370 584960 289460
rect 580165 289368 584960 289370
rect 580165 289312 580170 289368
rect 580226 289312 584960 289368
rect 580165 289310 584960 289312
rect 580165 289307 580231 289310
rect 583520 289220 584960 289310
rect 59997 287602 60063 287605
rect 59997 287600 62100 287602
rect 59997 287544 60002 287600
rect 60058 287544 62100 287600
rect 59997 287542 62100 287544
rect 59997 287539 60063 287542
rect 523677 285290 523743 285293
rect 521916 285288 523743 285290
rect 521916 285232 523682 285288
rect 523738 285232 523743 285288
rect 521916 285230 523743 285232
rect 523677 285227 523743 285230
rect -960 276450 480 276540
rect 3417 276450 3483 276453
rect -960 276448 3483 276450
rect -960 276392 3422 276448
rect 3478 276392 3483 276448
rect -960 276390 3483 276392
rect -960 276300 480 276390
rect 3417 276387 3483 276390
rect 580165 273730 580231 273733
rect 583520 273730 584960 273820
rect 580165 273728 584960 273730
rect 580165 273672 580170 273728
rect 580226 273672 584960 273728
rect 580165 273670 584960 273672
rect 580165 273667 580231 273670
rect 583520 273580 584960 273670
rect 59997 273322 60063 273325
rect 59997 273320 62100 273322
rect 59997 273264 60002 273320
rect 60058 273264 62100 273320
rect 59997 273262 62100 273264
rect 59997 273259 60063 273262
rect 523677 271962 523743 271965
rect 521916 271960 523743 271962
rect 521916 271904 523682 271960
rect 523738 271904 523743 271960
rect 521916 271902 523743 271904
rect 523677 271899 523743 271902
rect -960 259722 480 259812
rect 3417 259722 3483 259725
rect -960 259720 3483 259722
rect -960 259664 3422 259720
rect 3478 259664 3483 259720
rect -960 259662 3483 259664
rect -960 259572 480 259662
rect 3417 259659 3483 259662
rect 59997 259042 60063 259045
rect 59997 259040 62100 259042
rect 59997 258984 60002 259040
rect 60058 258984 62100 259040
rect 59997 258982 62100 258984
rect 59997 258979 60063 258982
rect 523769 258634 523835 258637
rect 521916 258632 523835 258634
rect 521916 258576 523774 258632
rect 523830 258576 523835 258632
rect 521916 258574 523835 258576
rect 523769 258571 523835 258574
rect 580165 258090 580231 258093
rect 583520 258090 584960 258180
rect 580165 258088 584960 258090
rect 580165 258032 580170 258088
rect 580226 258032 584960 258088
rect 580165 258030 584960 258032
rect 580165 258027 580231 258030
rect 583520 257940 584960 258030
rect 523677 245306 523743 245309
rect 521916 245304 523743 245306
rect 521916 245248 523682 245304
rect 523738 245248 523743 245304
rect 521916 245246 523743 245248
rect 523677 245243 523743 245246
rect 60089 244762 60155 244765
rect 60089 244760 62100 244762
rect 60089 244704 60094 244760
rect 60150 244704 62100 244760
rect 60089 244702 62100 244704
rect 60089 244699 60155 244702
rect -960 242994 480 243084
rect 3417 242994 3483 242997
rect -960 242992 3483 242994
rect -960 242936 3422 242992
rect 3478 242936 3483 242992
rect -960 242934 3483 242936
rect -960 242844 480 242934
rect 3417 242931 3483 242934
rect 580165 242450 580231 242453
rect 583520 242450 584960 242540
rect 580165 242448 584960 242450
rect 580165 242392 580170 242448
rect 580226 242392 584960 242448
rect 580165 242390 584960 242392
rect 580165 242387 580231 242390
rect 583520 242300 584960 242390
rect 523769 231978 523835 231981
rect 521916 231976 523835 231978
rect 521916 231920 523774 231976
rect 523830 231920 523835 231976
rect 521916 231918 523835 231920
rect 523769 231915 523835 231918
rect 59997 230482 60063 230485
rect 59997 230480 62100 230482
rect 59997 230424 60002 230480
rect 60058 230424 62100 230480
rect 59997 230422 62100 230424
rect 59997 230419 60063 230422
rect 580165 226810 580231 226813
rect 583520 226810 584960 226900
rect 580165 226808 584960 226810
rect 580165 226752 580170 226808
rect 580226 226752 584960 226808
rect 580165 226750 584960 226752
rect 580165 226747 580231 226750
rect 583520 226660 584960 226750
rect -960 226266 480 226356
rect 3417 226266 3483 226269
rect -960 226264 3483 226266
rect -960 226208 3422 226264
rect 3478 226208 3483 226264
rect -960 226206 3483 226208
rect -960 226116 480 226206
rect 3417 226203 3483 226206
rect 523677 218650 523743 218653
rect 521916 218648 523743 218650
rect 521916 218592 523682 218648
rect 523738 218592 523743 218648
rect 521916 218590 523743 218592
rect 523677 218587 523743 218590
rect 60089 216202 60155 216205
rect 60089 216200 62100 216202
rect 60089 216144 60094 216200
rect 60150 216144 62100 216200
rect 60089 216142 62100 216144
rect 60089 216139 60155 216142
rect 580165 211170 580231 211173
rect 583520 211170 584960 211260
rect 580165 211168 584960 211170
rect 580165 211112 580170 211168
rect 580226 211112 584960 211168
rect 580165 211110 584960 211112
rect 580165 211107 580231 211110
rect 583520 211020 584960 211110
rect -960 209402 480 209492
rect 3417 209402 3483 209405
rect -960 209400 3483 209402
rect -960 209344 3422 209400
rect 3478 209344 3483 209400
rect -960 209342 3483 209344
rect -960 209252 480 209342
rect 3417 209339 3483 209342
rect 523769 205322 523835 205325
rect 521916 205320 523835 205322
rect 521916 205264 523774 205320
rect 523830 205264 523835 205320
rect 521916 205262 523835 205264
rect 523769 205259 523835 205262
rect 59997 201922 60063 201925
rect 59997 201920 62100 201922
rect 59997 201864 60002 201920
rect 60058 201864 62100 201920
rect 59997 201862 62100 201864
rect 59997 201859 60063 201862
rect 580165 195530 580231 195533
rect 583520 195530 584960 195620
rect 580165 195528 584960 195530
rect 580165 195472 580170 195528
rect 580226 195472 584960 195528
rect 580165 195470 584960 195472
rect 580165 195467 580231 195470
rect 583520 195380 584960 195470
rect -960 192674 480 192764
rect 3509 192674 3575 192677
rect -960 192672 3575 192674
rect -960 192616 3514 192672
rect 3570 192616 3575 192672
rect -960 192614 3575 192616
rect -960 192524 480 192614
rect 3509 192611 3575 192614
rect 523677 191994 523743 191997
rect 521916 191992 523743 191994
rect 521916 191936 523682 191992
rect 523738 191936 523743 191992
rect 521916 191934 523743 191936
rect 523677 191931 523743 191934
rect 60181 187642 60247 187645
rect 60181 187640 62100 187642
rect 60181 187584 60186 187640
rect 60242 187584 62100 187640
rect 60181 187582 62100 187584
rect 60181 187579 60247 187582
rect 580165 179890 580231 179893
rect 583520 179890 584960 179980
rect 580165 179888 584960 179890
rect 580165 179832 580170 179888
rect 580226 179832 584960 179888
rect 580165 179830 584960 179832
rect 580165 179827 580231 179830
rect 583520 179740 584960 179830
rect 523861 178666 523927 178669
rect 521916 178664 523927 178666
rect 521916 178608 523866 178664
rect 523922 178608 523927 178664
rect 521916 178606 523927 178608
rect 523861 178603 523927 178606
rect -960 175946 480 176036
rect 3417 175946 3483 175949
rect -960 175944 3483 175946
rect -960 175888 3422 175944
rect 3478 175888 3483 175944
rect -960 175886 3483 175888
rect -960 175796 480 175886
rect 3417 175883 3483 175886
rect 60089 173362 60155 173365
rect 60089 173360 62100 173362
rect 60089 173304 60094 173360
rect 60150 173304 62100 173360
rect 60089 173302 62100 173304
rect 60089 173299 60155 173302
rect 523769 165338 523835 165341
rect 521916 165336 523835 165338
rect 521916 165280 523774 165336
rect 523830 165280 523835 165336
rect 521916 165278 523835 165280
rect 523769 165275 523835 165278
rect 580165 164250 580231 164253
rect 583520 164250 584960 164340
rect 580165 164248 584960 164250
rect 580165 164192 580170 164248
rect 580226 164192 584960 164248
rect 580165 164190 584960 164192
rect 580165 164187 580231 164190
rect 583520 164100 584960 164190
rect -960 159218 480 159308
rect 3141 159218 3207 159221
rect -960 159216 3207 159218
rect -960 159160 3146 159216
rect 3202 159160 3207 159216
rect -960 159158 3207 159160
rect -960 159068 480 159158
rect 3141 159155 3207 159158
rect 59997 159082 60063 159085
rect 59997 159080 62100 159082
rect 59997 159024 60002 159080
rect 60058 159024 62100 159080
rect 59997 159022 62100 159024
rect 59997 159019 60063 159022
rect 523677 152010 523743 152013
rect 521916 152008 523743 152010
rect 521916 151952 523682 152008
rect 523738 151952 523743 152008
rect 521916 151950 523743 151952
rect 523677 151947 523743 151950
rect 580165 148610 580231 148613
rect 583520 148610 584960 148700
rect 580165 148608 584960 148610
rect 580165 148552 580170 148608
rect 580226 148552 584960 148608
rect 580165 148550 584960 148552
rect 580165 148547 580231 148550
rect 583520 148460 584960 148550
rect 60181 144802 60247 144805
rect 60181 144800 62100 144802
rect 60181 144744 60186 144800
rect 60242 144744 62100 144800
rect 60181 144742 62100 144744
rect 60181 144739 60247 144742
rect -960 142354 480 142444
rect 3233 142354 3299 142357
rect -960 142352 3299 142354
rect -960 142296 3238 142352
rect 3294 142296 3299 142352
rect -960 142294 3299 142296
rect -960 142204 480 142294
rect 3233 142291 3299 142294
rect 523861 138682 523927 138685
rect 521916 138680 523927 138682
rect 521916 138624 523866 138680
rect 523922 138624 523927 138680
rect 521916 138622 523927 138624
rect 523861 138619 523927 138622
rect 580165 132970 580231 132973
rect 583520 132970 584960 133060
rect 580165 132968 584960 132970
rect 580165 132912 580170 132968
rect 580226 132912 584960 132968
rect 580165 132910 584960 132912
rect 580165 132907 580231 132910
rect 583520 132820 584960 132910
rect 60089 130522 60155 130525
rect 60089 130520 62100 130522
rect 60089 130464 60094 130520
rect 60150 130464 62100 130520
rect 60089 130462 62100 130464
rect 60089 130459 60155 130462
rect -960 125626 480 125716
rect 3233 125626 3299 125629
rect -960 125624 3299 125626
rect -960 125568 3238 125624
rect 3294 125568 3299 125624
rect -960 125566 3299 125568
rect -960 125476 480 125566
rect 3233 125563 3299 125566
rect 523769 125354 523835 125357
rect 521916 125352 523835 125354
rect 521916 125296 523774 125352
rect 523830 125296 523835 125352
rect 521916 125294 523835 125296
rect 523769 125291 523835 125294
rect 580165 117330 580231 117333
rect 583520 117330 584960 117420
rect 580165 117328 584960 117330
rect 580165 117272 580170 117328
rect 580226 117272 584960 117328
rect 580165 117270 584960 117272
rect 580165 117267 580231 117270
rect 583520 117180 584960 117270
rect 59997 116242 60063 116245
rect 59997 116240 62100 116242
rect 59997 116184 60002 116240
rect 60058 116184 62100 116240
rect 59997 116182 62100 116184
rect 59997 116179 60063 116182
rect 523677 112026 523743 112029
rect 521916 112024 523743 112026
rect 521916 111968 523682 112024
rect 523738 111968 523743 112024
rect 521916 111966 523743 111968
rect 523677 111963 523743 111966
rect -960 108898 480 108988
rect 3417 108898 3483 108901
rect -960 108896 3483 108898
rect -960 108840 3422 108896
rect 3478 108840 3483 108896
rect -960 108838 3483 108840
rect -960 108748 480 108838
rect 3417 108835 3483 108838
rect 60273 101962 60339 101965
rect 60273 101960 62100 101962
rect 60273 101904 60278 101960
rect 60334 101904 62100 101960
rect 60273 101902 62100 101904
rect 60273 101899 60339 101902
rect 580165 101690 580231 101693
rect 583520 101690 584960 101780
rect 580165 101688 584960 101690
rect 580165 101632 580170 101688
rect 580226 101632 584960 101688
rect 580165 101630 584960 101632
rect 580165 101627 580231 101630
rect 583520 101540 584960 101630
rect 523953 98698 524019 98701
rect 521916 98696 524019 98698
rect 521916 98640 523958 98696
rect 524014 98640 524019 98696
rect 521916 98638 524019 98640
rect 523953 98635 524019 98638
rect -960 92170 480 92260
rect 3325 92170 3391 92173
rect -960 92168 3391 92170
rect -960 92112 3330 92168
rect 3386 92112 3391 92168
rect -960 92110 3391 92112
rect -960 92020 480 92110
rect 3325 92107 3391 92110
rect 60181 87682 60247 87685
rect 60181 87680 62100 87682
rect 60181 87624 60186 87680
rect 60242 87624 62100 87680
rect 60181 87622 62100 87624
rect 60181 87619 60247 87622
rect 580165 86050 580231 86053
rect 583520 86050 584960 86140
rect 580165 86048 584960 86050
rect 580165 85992 580170 86048
rect 580226 85992 584960 86048
rect 580165 85990 584960 85992
rect 580165 85987 580231 85990
rect 583520 85900 584960 85990
rect 523861 85370 523927 85373
rect 521916 85368 523927 85370
rect 521916 85312 523866 85368
rect 523922 85312 523927 85368
rect 521916 85310 523927 85312
rect 523861 85307 523927 85310
rect -960 75306 480 75396
rect 3417 75306 3483 75309
rect -960 75304 3483 75306
rect -960 75248 3422 75304
rect 3478 75248 3483 75304
rect -960 75246 3483 75248
rect -960 75156 480 75246
rect 3417 75243 3483 75246
rect 60089 73402 60155 73405
rect 60089 73400 62100 73402
rect 60089 73344 60094 73400
rect 60150 73344 62100 73400
rect 60089 73342 62100 73344
rect 60089 73339 60155 73342
rect 523769 72042 523835 72045
rect 521916 72040 523835 72042
rect 521916 71984 523774 72040
rect 523830 71984 523835 72040
rect 521916 71982 523835 71984
rect 523769 71979 523835 71982
rect 580165 70410 580231 70413
rect 583520 70410 584960 70500
rect 580165 70408 584960 70410
rect 580165 70352 580170 70408
rect 580226 70352 584960 70408
rect 580165 70350 584960 70352
rect 580165 70347 580231 70350
rect 583520 70260 584960 70350
rect 59997 59122 60063 59125
rect 59997 59120 62100 59122
rect 59997 59064 60002 59120
rect 60058 59064 62100 59120
rect 59997 59062 62100 59064
rect 59997 59059 60063 59062
rect 523677 58714 523743 58717
rect 521916 58712 523743 58714
rect -960 58578 480 58668
rect 521916 58656 523682 58712
rect 523738 58656 523743 58712
rect 521916 58654 523743 58656
rect 523677 58651 523743 58654
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 54770 580231 54773
rect 583520 54770 584960 54860
rect 580165 54768 584960 54770
rect 580165 54712 580170 54768
rect 580226 54712 584960 54768
rect 580165 54710 584960 54712
rect 580165 54707 580231 54710
rect 583520 54620 584960 54710
rect -960 41850 480 41940
rect 3417 41850 3483 41853
rect -960 41848 3483 41850
rect -960 41792 3422 41848
rect 3478 41792 3483 41848
rect -960 41790 3483 41792
rect -960 41700 480 41790
rect 3417 41787 3483 41790
rect 580165 39130 580231 39133
rect 583520 39130 584960 39220
rect 580165 39128 584960 39130
rect 580165 39072 580170 39128
rect 580226 39072 584960 39128
rect 580165 39070 584960 39072
rect 580165 39067 580231 39070
rect 583520 38980 584960 39070
rect 110045 38858 110111 38861
rect 203885 38858 203951 38861
rect 109174 38856 110111 38858
rect 109174 38800 110050 38856
rect 110106 38800 110111 38856
rect 109174 38798 110111 38800
rect 109174 38722 109234 38798
rect 110045 38795 110111 38798
rect 203014 38856 203951 38858
rect 203014 38800 203890 38856
rect 203946 38800 203951 38856
rect 203014 38798 203951 38800
rect 109309 38722 109375 38725
rect 109174 38720 109375 38722
rect 109174 38664 109314 38720
rect 109370 38664 109375 38720
rect 109174 38662 109375 38664
rect 203014 38722 203074 38798
rect 203885 38795 203951 38798
rect 203149 38722 203215 38725
rect 203014 38720 203215 38722
rect 203014 38664 203154 38720
rect 203210 38664 203215 38720
rect 203014 38662 203215 38664
rect 109309 38659 109375 38662
rect 203149 38659 203215 38662
rect -960 25122 480 25212
rect 3417 25122 3483 25125
rect -960 25120 3483 25122
rect -960 25064 3422 25120
rect 3478 25064 3483 25120
rect -960 25062 3483 25064
rect -960 24972 480 25062
rect 3417 25059 3483 25062
rect 580165 23490 580231 23493
rect 583520 23490 584960 23580
rect 580165 23488 584960 23490
rect 580165 23432 580170 23488
rect 580226 23432 584960 23488
rect 580165 23430 584960 23432
rect 580165 23427 580231 23430
rect 583520 23340 584960 23430
rect 80145 19274 80211 19277
rect 80421 19274 80487 19277
rect 80145 19272 80487 19274
rect 80145 19216 80150 19272
rect 80206 19216 80426 19272
rect 80482 19216 80487 19272
rect 80145 19214 80487 19216
rect 80145 19211 80211 19214
rect 80421 19211 80487 19214
rect -960 8394 480 8484
rect 3417 8394 3483 8397
rect -960 8392 3483 8394
rect -960 8336 3422 8392
rect 3478 8336 3483 8392
rect -960 8334 3483 8336
rect -960 8244 480 8334
rect 3417 8331 3483 8334
rect 580165 7850 580231 7853
rect 583520 7850 584960 7940
rect 580165 7848 584960 7850
rect 580165 7792 580170 7848
rect 580226 7792 584960 7848
rect 580165 7790 584960 7792
rect 580165 7787 580231 7790
rect 583520 7700 584960 7790
rect 521561 3634 521627 3637
rect 582189 3634 582255 3637
rect 521561 3632 582255 3634
rect 521561 3576 521566 3632
rect 521622 3576 582194 3632
rect 582250 3576 582255 3632
rect 521561 3574 582255 3576
rect 521561 3571 521627 3574
rect 582189 3571 582255 3574
rect 25497 3498 25563 3501
rect 81525 3498 81591 3501
rect 25497 3496 81591 3498
rect 25497 3440 25502 3496
rect 25558 3440 81530 3496
rect 81586 3440 81591 3496
rect 25497 3438 81591 3440
rect 25497 3435 25563 3438
rect 81525 3435 81591 3438
rect 86125 3498 86191 3501
rect 129917 3498 129983 3501
rect 86125 3496 129983 3498
rect 86125 3440 86130 3496
rect 86186 3440 129922 3496
rect 129978 3440 129983 3496
rect 86125 3438 129983 3440
rect 86125 3435 86191 3438
rect 129917 3435 129983 3438
rect 194409 3498 194475 3501
rect 215385 3498 215451 3501
rect 194409 3496 215451 3498
rect 194409 3440 194414 3496
rect 194470 3440 215390 3496
rect 215446 3440 215451 3496
rect 194409 3438 215451 3440
rect 194409 3435 194475 3438
rect 215385 3435 215451 3438
rect 442901 3498 442967 3501
rect 482277 3498 482343 3501
rect 442901 3496 482343 3498
rect 442901 3440 442906 3496
rect 442962 3440 482282 3496
rect 482338 3440 482343 3496
rect 442901 3438 482343 3440
rect 442901 3435 442967 3438
rect 482277 3435 482343 3438
rect 19517 3362 19583 3365
rect 77477 3362 77543 3365
rect 19517 3360 77543 3362
rect 19517 3304 19522 3360
rect 19578 3304 77482 3360
rect 77538 3304 77543 3360
rect 19517 3302 77543 3304
rect 19517 3299 19583 3302
rect 77477 3299 77543 3302
rect 82629 3362 82695 3365
rect 127065 3362 127131 3365
rect 82629 3360 127131 3362
rect 82629 3304 82634 3360
rect 82690 3304 127070 3360
rect 127126 3304 127131 3360
rect 82629 3302 127131 3304
rect 82629 3299 82695 3302
rect 127065 3299 127131 3302
rect 190821 3362 190887 3365
rect 212625 3362 212691 3365
rect 190821 3360 212691 3362
rect 190821 3304 190826 3360
rect 190882 3304 212630 3360
rect 212686 3304 212691 3360
rect 190821 3302 212691 3304
rect 190821 3299 190887 3302
rect 212625 3299 212691 3302
rect 456701 3362 456767 3365
rect 500125 3362 500191 3365
rect 456701 3360 500191 3362
rect 456701 3304 456706 3360
rect 456762 3304 500130 3360
rect 500186 3304 500191 3360
rect 456701 3302 500191 3304
rect 456701 3299 456767 3302
rect 500125 3299 500191 3302
rect 518709 3362 518775 3365
rect 578601 3362 578667 3365
rect 518709 3360 578667 3362
rect 518709 3304 518714 3360
rect 518770 3304 578606 3360
rect 578662 3304 578667 3360
rect 518709 3302 578667 3304
rect 518709 3299 518775 3302
rect 578601 3299 578667 3302
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 652000 62604 675098
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 652000 66204 678698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 652000 73404 685898
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 652000 77004 653498
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 652000 80604 657098
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 652000 84204 660698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 652000 91404 667898
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 652000 95004 671498
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 652000 98604 675098
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 652000 102204 678698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 652000 109404 685898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 652000 113004 653498
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 652000 116604 657098
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 652000 120204 660698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 652000 127404 667898
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 652000 131004 671498
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 652000 134604 675098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 652000 138204 678698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 652000 145404 685898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 652000 149004 653498
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 652000 152604 657098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 652000 156204 660698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 652000 163404 667898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 652000 167004 671498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 652000 170604 675098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 652000 174204 678698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 652000 181404 685898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 652000 185004 653498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 652000 188604 657098
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 652000 192204 660698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 652000 199404 667898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 652000 203004 671498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 652000 206604 675098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 652000 210204 678698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 652000 217404 685898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 652000 221004 653498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 652000 224604 657098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 652000 228204 660698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 652000 235404 667898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 652000 239004 671498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 652000 242604 675098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 652000 246204 678698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 652000 253404 685898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 652000 257004 653498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 652000 260604 657098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 652000 264204 660698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 652000 271404 667898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 652000 275004 671498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 652000 278604 675098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 652000 282204 678698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 652000 289404 685898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 652000 293004 653498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 652000 296604 657098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 652000 300204 660698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 652000 307404 667898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 652000 311004 671498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 652000 314604 675098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 652000 318204 678698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 652000 325404 685898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 652000 329004 653498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 652000 332604 657098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 652000 336204 660698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 652000 343404 667898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 652000 347004 671498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 652000 350604 675098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 652000 354204 678698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 652000 361404 685898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 652000 365004 653498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 652000 368604 657098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 652000 372204 660698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 652000 379404 667898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 652000 383004 671498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 652000 386604 675098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 652000 390204 678698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 652000 397404 685898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 652000 401004 653498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 652000 404604 657098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 652000 408204 660698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 652000 415404 667898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 652000 419004 671498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 652000 422604 675098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 652000 426204 678698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 652000 433404 685898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 652000 437004 653498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 652000 440604 657098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 652000 444204 660698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 652000 451404 667898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 652000 455004 671498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 652000 458604 675098
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 652000 462204 678698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 652000 469404 685898
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 652000 473004 653498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 652000 476604 657098
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 652000 480204 660698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 652000 487404 667898
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 652000 491004 671498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 652000 494604 675098
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 652000 498204 678698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 652000 505404 685898
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 652000 509004 653498
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 652000 512604 657098
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 652000 516204 660698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 27654 62604 52000
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 31254 66204 52000
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 38454 73404 52000
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 42054 77004 52000
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 45654 80604 52000
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 49254 84204 52000
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 20454 91404 52000
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 24054 95004 52000
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 27654 98604 52000
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 31254 102204 52000
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 38454 109404 52000
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 42054 113004 52000
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 45654 116604 52000
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 49254 120204 52000
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 20454 127404 52000
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 24054 131004 52000
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 27654 134604 52000
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 31254 138204 52000
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 38454 145404 52000
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 42054 149004 52000
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 45654 152604 52000
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 49254 156204 52000
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 20454 163404 52000
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 24054 167004 52000
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 27654 170604 52000
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 31254 174204 52000
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 38454 181404 52000
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 42054 185004 52000
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 45654 188604 52000
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 49254 192204 52000
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 20454 199404 52000
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 24054 203004 52000
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 27654 206604 52000
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 31254 210204 52000
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 38454 217404 52000
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 42054 221004 52000
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 45654 224604 52000
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 49254 228204 52000
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 20454 235404 52000
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 24054 239004 52000
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 27654 242604 52000
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 31254 246204 52000
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 38454 253404 52000
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 42054 257004 52000
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 45654 260604 52000
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 49254 264204 52000
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 20454 271404 52000
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 24054 275004 52000
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 27654 278604 52000
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 31254 282204 52000
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 38454 289404 52000
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 42054 293004 52000
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 45654 296604 52000
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 49254 300204 52000
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 20454 307404 52000
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 24054 311004 52000
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 27654 314604 52000
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 31254 318204 52000
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 38454 325404 52000
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 42054 329004 52000
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 45654 332604 52000
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 49254 336204 52000
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 20454 343404 52000
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 24054 347004 52000
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 27654 350604 52000
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 31254 354204 52000
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 38454 361404 52000
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 42054 365004 52000
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 45654 368604 52000
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 49254 372204 52000
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 20454 379404 52000
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 24054 383004 52000
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 27654 386604 52000
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 31254 390204 52000
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 38454 397404 52000
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 42054 401004 52000
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 45654 404604 52000
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 49254 408204 52000
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 20454 415404 52000
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 24054 419004 52000
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 27654 422604 52000
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 31254 426204 52000
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 38454 433404 52000
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 42054 437004 52000
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 45654 440604 52000
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 49254 444204 52000
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 20454 451404 52000
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 24054 455004 52000
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 27654 458604 52000
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 31254 462204 52000
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 38454 469404 52000
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 42054 473004 52000
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 45654 476604 52000
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 49254 480204 52000
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 20454 487404 52000
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 24054 491004 52000
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 27654 494604 52000
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 31254 498204 52000
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 38454 505404 52000
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 42054 509004 52000
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 45654 512604 52000
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 49254 516204 52000
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use ghazi_top_dffram_csv  mprj
timestamp 1607490450
transform 1 0 62000 0 1 52000
box 0 0 460000 600000
<< labels >>
rlabel metal3 s 583520 7700 584960 7940 6 io_in[0]
port 0 nsew default input
rlabel metal3 s 583520 476900 584960 477140 6 io_in[10]
port 1 nsew default input
rlabel metal3 s 583520 523820 584960 524060 6 io_in[11]
port 2 nsew default input
rlabel metal3 s 583520 570740 584960 570980 6 io_in[12]
port 3 nsew default input
rlabel metal3 s 583520 617660 584960 617900 6 io_in[13]
port 4 nsew default input
rlabel metal3 s 583520 664580 584960 664820 6 io_in[14]
port 5 nsew default input
rlabel metal2 s 573058 703520 573170 704960 6 io_in[15]
port 6 nsew default input
rlabel metal2 s 508198 703520 508310 704960 6 io_in[16]
port 7 nsew default input
rlabel metal2 s 443338 703520 443450 704960 6 io_in[17]
port 8 nsew default input
rlabel metal2 s 378386 703520 378498 704960 6 io_in[18]
port 9 nsew default input
rlabel metal2 s 313526 703520 313638 704960 6 io_in[19]
port 10 nsew default input
rlabel metal3 s 583520 54620 584960 54860 6 io_in[1]
port 11 nsew default input
rlabel metal2 s 248666 703520 248778 704960 6 io_in[20]
port 12 nsew default input
rlabel metal2 s 183714 703520 183826 704960 6 io_in[21]
port 13 nsew default input
rlabel metal2 s 118854 703520 118966 704960 6 io_in[22]
port 14 nsew default input
rlabel metal2 s 53994 703520 54106 704960 6 io_in[23]
port 15 nsew default input
rlabel metal3 s -960 695316 480 695556 4 io_in[24]
port 16 nsew default input
rlabel metal3 s -960 645132 480 645372 4 io_in[25]
port 17 nsew default input
rlabel metal3 s -960 594812 480 595052 4 io_in[26]
port 18 nsew default input
rlabel metal3 s -960 544492 480 544732 4 io_in[27]
port 19 nsew default input
rlabel metal3 s -960 494172 480 494412 4 io_in[28]
port 20 nsew default input
rlabel metal3 s -960 443988 480 444228 4 io_in[29]
port 21 nsew default input
rlabel metal3 s 583520 101540 584960 101780 6 io_in[2]
port 22 nsew default input
rlabel metal3 s -960 393668 480 393908 4 io_in[30]
port 23 nsew default input
rlabel metal3 s -960 343348 480 343588 4 io_in[31]
port 24 nsew default input
rlabel metal3 s -960 293164 480 293404 4 io_in[32]
port 25 nsew default input
rlabel metal3 s -960 242844 480 243084 4 io_in[33]
port 26 nsew default input
rlabel metal3 s -960 192524 480 192764 4 io_in[34]
port 27 nsew default input
rlabel metal3 s -960 142204 480 142444 4 io_in[35]
port 28 nsew default input
rlabel metal3 s -960 92020 480 92260 4 io_in[36]
port 29 nsew default input
rlabel metal3 s -960 41700 480 41940 4 io_in[37]
port 30 nsew default input
rlabel metal3 s 583520 148460 584960 148700 6 io_in[3]
port 31 nsew default input
rlabel metal3 s 583520 195380 584960 195620 6 io_in[4]
port 32 nsew default input
rlabel metal3 s 583520 242300 584960 242540 6 io_in[5]
port 33 nsew default input
rlabel metal3 s 583520 289220 584960 289460 6 io_in[6]
port 34 nsew default input
rlabel metal3 s 583520 336140 584960 336380 6 io_in[7]
port 35 nsew default input
rlabel metal3 s 583520 383060 584960 383300 6 io_in[8]
port 36 nsew default input
rlabel metal3 s 583520 429980 584960 430220 6 io_in[9]
port 37 nsew default input
rlabel metal3 s 583520 38980 584960 39220 6 io_oeb[0]
port 38 nsew default tristate
rlabel metal3 s 583520 508180 584960 508420 6 io_oeb[10]
port 39 nsew default tristate
rlabel metal3 s 583520 555100 584960 555340 6 io_oeb[11]
port 40 nsew default tristate
rlabel metal3 s 583520 602020 584960 602260 6 io_oeb[12]
port 41 nsew default tristate
rlabel metal3 s 583520 648940 584960 649180 6 io_oeb[13]
port 42 nsew default tristate
rlabel metal3 s 583520 695860 584960 696100 6 io_oeb[14]
port 43 nsew default tristate
rlabel metal2 s 529818 703520 529930 704960 6 io_oeb[15]
port 44 nsew default tristate
rlabel metal2 s 464958 703520 465070 704960 6 io_oeb[16]
port 45 nsew default tristate
rlabel metal2 s 400098 703520 400210 704960 6 io_oeb[17]
port 46 nsew default tristate
rlabel metal2 s 335146 703520 335258 704960 6 io_oeb[18]
port 47 nsew default tristate
rlabel metal2 s 270286 703520 270398 704960 6 io_oeb[19]
port 48 nsew default tristate
rlabel metal3 s 583520 85900 584960 86140 6 io_oeb[1]
port 49 nsew default tristate
rlabel metal2 s 205426 703520 205538 704960 6 io_oeb[20]
port 50 nsew default tristate
rlabel metal2 s 140474 703520 140586 704960 6 io_oeb[21]
port 51 nsew default tristate
rlabel metal2 s 75614 703520 75726 704960 6 io_oeb[22]
port 52 nsew default tristate
rlabel metal2 s 10754 703520 10866 704960 6 io_oeb[23]
port 53 nsew default tristate
rlabel metal3 s -960 661860 480 662100 4 io_oeb[24]
port 54 nsew default tristate
rlabel metal3 s -960 611540 480 611780 4 io_oeb[25]
port 55 nsew default tristate
rlabel metal3 s -960 561220 480 561460 4 io_oeb[26]
port 56 nsew default tristate
rlabel metal3 s -960 511036 480 511276 4 io_oeb[27]
port 57 nsew default tristate
rlabel metal3 s -960 460716 480 460956 4 io_oeb[28]
port 58 nsew default tristate
rlabel metal3 s -960 410396 480 410636 4 io_oeb[29]
port 59 nsew default tristate
rlabel metal3 s 583520 132820 584960 133060 6 io_oeb[2]
port 60 nsew default tristate
rlabel metal3 s -960 360212 480 360452 4 io_oeb[30]
port 61 nsew default tristate
rlabel metal3 s -960 309892 480 310132 4 io_oeb[31]
port 62 nsew default tristate
rlabel metal3 s -960 259572 480 259812 4 io_oeb[32]
port 63 nsew default tristate
rlabel metal3 s -960 209252 480 209492 4 io_oeb[33]
port 64 nsew default tristate
rlabel metal3 s -960 159068 480 159308 4 io_oeb[34]
port 65 nsew default tristate
rlabel metal3 s -960 108748 480 108988 4 io_oeb[35]
port 66 nsew default tristate
rlabel metal3 s -960 58428 480 58668 4 io_oeb[36]
port 67 nsew default tristate
rlabel metal3 s -960 8244 480 8484 4 io_oeb[37]
port 68 nsew default tristate
rlabel metal3 s 583520 179740 584960 179980 6 io_oeb[3]
port 69 nsew default tristate
rlabel metal3 s 583520 226660 584960 226900 6 io_oeb[4]
port 70 nsew default tristate
rlabel metal3 s 583520 273580 584960 273820 6 io_oeb[5]
port 71 nsew default tristate
rlabel metal3 s 583520 320500 584960 320740 6 io_oeb[6]
port 72 nsew default tristate
rlabel metal3 s 583520 367420 584960 367660 6 io_oeb[7]
port 73 nsew default tristate
rlabel metal3 s 583520 414340 584960 414580 6 io_oeb[8]
port 74 nsew default tristate
rlabel metal3 s 583520 461260 584960 461500 6 io_oeb[9]
port 75 nsew default tristate
rlabel metal3 s 583520 23340 584960 23580 6 io_out[0]
port 76 nsew default tristate
rlabel metal3 s 583520 492540 584960 492780 6 io_out[10]
port 77 nsew default tristate
rlabel metal3 s 583520 539460 584960 539700 6 io_out[11]
port 78 nsew default tristate
rlabel metal3 s 583520 586380 584960 586620 6 io_out[12]
port 79 nsew default tristate
rlabel metal3 s 583520 633300 584960 633540 6 io_out[13]
port 80 nsew default tristate
rlabel metal3 s 583520 680220 584960 680460 6 io_out[14]
port 81 nsew default tristate
rlabel metal2 s 551438 703520 551550 704960 6 io_out[15]
port 82 nsew default tristate
rlabel metal2 s 486578 703520 486690 704960 6 io_out[16]
port 83 nsew default tristate
rlabel metal2 s 421718 703520 421830 704960 6 io_out[17]
port 84 nsew default tristate
rlabel metal2 s 356766 703520 356878 704960 6 io_out[18]
port 85 nsew default tristate
rlabel metal2 s 291906 703520 292018 704960 6 io_out[19]
port 86 nsew default tristate
rlabel metal3 s 583520 70260 584960 70500 6 io_out[1]
port 87 nsew default tristate
rlabel metal2 s 227046 703520 227158 704960 6 io_out[20]
port 88 nsew default tristate
rlabel metal2 s 162094 703520 162206 704960 6 io_out[21]
port 89 nsew default tristate
rlabel metal2 s 97234 703520 97346 704960 6 io_out[22]
port 90 nsew default tristate
rlabel metal2 s 32374 703520 32486 704960 6 io_out[23]
port 91 nsew default tristate
rlabel metal3 s -960 678588 480 678828 4 io_out[24]
port 92 nsew default tristate
rlabel metal3 s -960 628268 480 628508 4 io_out[25]
port 93 nsew default tristate
rlabel metal3 s -960 578084 480 578324 4 io_out[26]
port 94 nsew default tristate
rlabel metal3 s -960 527764 480 528004 4 io_out[27]
port 95 nsew default tristate
rlabel metal3 s -960 477444 480 477684 4 io_out[28]
port 96 nsew default tristate
rlabel metal3 s -960 427124 480 427364 4 io_out[29]
port 97 nsew default tristate
rlabel metal3 s 583520 117180 584960 117420 6 io_out[2]
port 98 nsew default tristate
rlabel metal3 s -960 376940 480 377180 4 io_out[30]
port 99 nsew default tristate
rlabel metal3 s -960 326620 480 326860 4 io_out[31]
port 100 nsew default tristate
rlabel metal3 s -960 276300 480 276540 4 io_out[32]
port 101 nsew default tristate
rlabel metal3 s -960 226116 480 226356 4 io_out[33]
port 102 nsew default tristate
rlabel metal3 s -960 175796 480 176036 4 io_out[34]
port 103 nsew default tristate
rlabel metal3 s -960 125476 480 125716 4 io_out[35]
port 104 nsew default tristate
rlabel metal3 s -960 75156 480 75396 4 io_out[36]
port 105 nsew default tristate
rlabel metal3 s -960 24972 480 25212 4 io_out[37]
port 106 nsew default tristate
rlabel metal3 s 583520 164100 584960 164340 6 io_out[3]
port 107 nsew default tristate
rlabel metal3 s 583520 211020 584960 211260 6 io_out[4]
port 108 nsew default tristate
rlabel metal3 s 583520 257940 584960 258180 6 io_out[5]
port 109 nsew default tristate
rlabel metal3 s 583520 304860 584960 305100 6 io_out[6]
port 110 nsew default tristate
rlabel metal3 s 583520 351780 584960 352020 6 io_out[7]
port 111 nsew default tristate
rlabel metal3 s 583520 398700 584960 398940 6 io_out[8]
port 112 nsew default tristate
rlabel metal3 s 583520 445620 584960 445860 6 io_out[9]
port 113 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 114 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 115 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 116 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 117 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 118 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 119 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 120 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 121 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 122 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 123 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 124 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 125 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 126 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 127 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 128 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 129 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 130 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 131 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 132 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 133 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 134 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 135 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 136 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 137 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 138 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 139 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 140 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 141 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 142 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 143 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 144 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 145 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 146 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 147 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 148 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 149 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 150 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 151 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 152 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 153 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 154 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 155 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 156 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 157 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 158 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 159 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 160 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 161 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 162 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 163 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 164 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 165 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 166 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 167 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 168 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 169 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 170 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 171 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 172 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 173 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 174 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 175 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 176 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 177 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 178 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 179 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 180 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 181 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 182 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 183 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 184 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 185 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 186 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 187 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 188 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 189 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 190 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 191 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 192 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 193 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 194 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 195 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 196 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 197 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 198 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 199 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 200 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 201 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 202 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 203 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 204 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 205 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 206 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 207 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 208 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 209 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 210 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 211 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 212 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 213 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 214 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 215 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 216 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 217 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 218 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 219 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 220 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 221 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 222 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 223 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 224 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 225 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 226 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 227 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 228 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 229 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 230 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 231 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 232 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 233 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 234 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 235 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 236 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 237 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 238 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 239 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 240 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 241 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 242 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 243 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 244 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 245 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 246 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 247 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 248 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 249 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 250 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 251 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 252 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 253 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 254 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 255 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 256 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 257 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 258 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 259 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 260 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 261 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 262 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 263 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 264 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 265 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 266 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 267 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 268 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 269 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 270 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 271 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 272 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 273 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 274 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 275 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 276 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 277 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 278 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 279 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 280 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 281 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 282 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 283 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 284 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 285 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 286 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 287 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 288 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 289 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 290 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 291 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 292 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 293 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 294 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 295 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 296 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 297 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 298 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 299 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 300 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 301 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 302 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 303 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 304 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 305 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 306 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 307 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 308 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 309 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 310 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 311 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 312 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 313 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 314 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 315 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 316 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 317 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 318 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 319 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 320 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 321 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 322 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 323 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 324 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 325 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 326 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 327 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 328 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 329 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 330 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 331 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 332 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 333 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 334 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 335 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 336 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 337 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 338 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 339 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 340 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 341 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 342 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 343 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 344 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 345 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 346 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 347 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 348 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 349 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 350 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 351 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 352 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 353 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 354 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 355 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 356 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 357 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 358 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 359 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 360 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 361 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 362 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 363 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 364 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 365 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 366 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 367 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 368 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 369 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 370 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 371 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 372 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 373 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 374 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 375 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 376 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 377 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 378 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 379 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 380 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 381 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 382 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 383 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 384 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 385 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 386 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 387 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 388 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 389 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 390 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 391 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 392 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 393 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 394 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 395 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 396 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 397 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 398 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 399 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 400 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 401 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 402 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 403 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 404 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 405 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 406 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 407 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 408 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 409 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 410 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 411 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 412 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 413 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 414 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 415 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 416 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 417 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 418 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 419 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 420 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 421 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 422 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 423 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 424 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 425 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 426 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 427 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 428 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 429 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 430 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 431 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 432 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 433 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 434 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 435 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 436 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 437 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 438 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 439 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 440 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 441 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 442 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 443 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 444 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 445 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 446 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 447 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 448 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 449 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 450 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 451 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 452 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 453 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 454 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 455 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 456 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 457 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 458 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 459 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 460 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 461 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 462 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 463 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 464 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 465 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 466 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 467 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 468 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 469 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 470 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 471 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 472 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 473 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 474 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 475 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 476 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 477 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 478 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 479 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 480 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 481 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 482 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 483 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 484 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 485 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 486 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 487 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 488 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 489 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 490 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 491 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 492 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 493 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 494 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 495 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 496 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 497 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 498 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 499 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 500 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 501 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 502 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 503 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 504 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 505 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 506 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 507 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 508 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 509 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 510 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 511 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 512 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 513 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 514 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 515 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 516 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 517 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 518 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 519 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 520 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 521 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 522 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 523 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 524 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 525 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 526 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 527 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 528 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 529 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 530 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 531 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 532 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 533 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 534 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 535 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 536 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 537 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 538 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 539 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 540 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 541 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 542 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 543 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 544 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 545 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 546 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 547 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 548 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 549 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 550 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 551 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 552 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 553 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 554 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 555 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 556 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 557 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 558 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 559 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 560 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 561 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 562 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 563 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 564 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 565 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 566 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 567 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 568 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 569 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 570 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 571 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 572 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 573 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 574 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 575 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 576 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 577 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 578 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 579 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 580 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 581 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 582 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 583 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 584 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 585 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 586 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 587 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 588 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 589 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 590 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 591 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 592 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 593 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 594 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 595 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 596 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 597 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 598 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 599 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 600 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 601 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 602 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 603 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 604 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 605 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 606 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 607 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 608 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 609 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 610 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 611 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 612 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
