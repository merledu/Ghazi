VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 89.660 2619.630 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2619.310 89.520 2899.310 89.660 ;
        RECT 2619.310 89.460 2619.630 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2619.340 89.460 2619.600 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2619.330 293.235 2619.610 293.605 ;
        RECT 2619.400 89.750 2619.540 293.235 ;
        RECT 2619.340 89.430 2619.600 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2619.330 293.280 2619.610 293.560 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2606.000 293.570 2610.000 293.960 ;
        RECT 2619.305 293.570 2619.635 293.585 ;
        RECT 2606.000 293.360 2619.635 293.570 ;
        RECT 2609.580 293.270 2619.635 293.360 ;
        RECT 2619.305 293.255 2619.635 293.270 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 2297.620 2621.930 2297.680 ;
        RECT 2901.290 2297.620 2901.610 2297.680 ;
        RECT 2621.610 2297.480 2901.610 2297.620 ;
        RECT 2621.610 2297.420 2621.930 2297.480 ;
        RECT 2901.290 2297.420 2901.610 2297.480 ;
      LAYER via ;
        RECT 2621.640 2297.420 2621.900 2297.680 ;
        RECT 2901.320 2297.420 2901.580 2297.680 ;
      LAYER met2 ;
        RECT 2901.310 2433.875 2901.590 2434.245 ;
        RECT 2901.380 2297.710 2901.520 2433.875 ;
        RECT 2621.640 2297.390 2621.900 2297.710 ;
        RECT 2901.320 2297.390 2901.580 2297.710 ;
        RECT 2621.700 2293.485 2621.840 2297.390 ;
        RECT 2621.630 2293.115 2621.910 2293.485 ;
      LAYER via2 ;
        RECT 2901.310 2433.920 2901.590 2434.200 ;
        RECT 2621.630 2293.160 2621.910 2293.440 ;
      LAYER met3 ;
        RECT 2901.285 2434.210 2901.615 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2901.285 2433.910 2924.800 2434.210 ;
        RECT 2901.285 2433.895 2901.615 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2606.000 2293.450 2610.000 2293.840 ;
        RECT 2621.605 2293.450 2621.935 2293.465 ;
        RECT 2606.000 2293.240 2621.935 2293.450 ;
        RECT 2609.580 2293.150 2621.935 2293.240 ;
        RECT 2621.605 2293.135 2621.935 2293.150 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2497.540 2618.710 2497.600 ;
        RECT 2901.290 2497.540 2901.610 2497.600 ;
        RECT 2618.390 2497.400 2901.610 2497.540 ;
        RECT 2618.390 2497.340 2618.710 2497.400 ;
        RECT 2901.290 2497.340 2901.610 2497.400 ;
      LAYER via ;
        RECT 2618.420 2497.340 2618.680 2497.600 ;
        RECT 2901.320 2497.340 2901.580 2497.600 ;
      LAYER met2 ;
        RECT 2901.310 2669.155 2901.590 2669.525 ;
        RECT 2901.380 2497.630 2901.520 2669.155 ;
        RECT 2618.420 2497.310 2618.680 2497.630 ;
        RECT 2901.320 2497.310 2901.580 2497.630 ;
        RECT 2618.480 2493.405 2618.620 2497.310 ;
        RECT 2618.410 2493.035 2618.690 2493.405 ;
      LAYER via2 ;
        RECT 2901.310 2669.200 2901.590 2669.480 ;
        RECT 2618.410 2493.080 2618.690 2493.360 ;
      LAYER met3 ;
        RECT 2901.285 2669.490 2901.615 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2901.285 2669.190 2924.800 2669.490 ;
        RECT 2901.285 2669.175 2901.615 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2606.000 2493.370 2610.000 2493.760 ;
        RECT 2618.385 2493.370 2618.715 2493.385 ;
        RECT 2606.000 2493.160 2618.715 2493.370 ;
        RECT 2609.580 2493.070 2618.715 2493.160 ;
        RECT 2618.385 2493.055 2618.715 2493.070 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2697.800 2618.710 2697.860 ;
        RECT 2901.290 2697.800 2901.610 2697.860 ;
        RECT 2618.390 2697.660 2901.610 2697.800 ;
        RECT 2618.390 2697.600 2618.710 2697.660 ;
        RECT 2901.290 2697.600 2901.610 2697.660 ;
      LAYER via ;
        RECT 2618.420 2697.600 2618.680 2697.860 ;
        RECT 2901.320 2697.600 2901.580 2697.860 ;
      LAYER met2 ;
        RECT 2901.310 2903.755 2901.590 2904.125 ;
        RECT 2901.380 2697.890 2901.520 2903.755 ;
        RECT 2618.420 2697.570 2618.680 2697.890 ;
        RECT 2901.320 2697.570 2901.580 2697.890 ;
        RECT 2618.480 2693.325 2618.620 2697.570 ;
        RECT 2618.410 2692.955 2618.690 2693.325 ;
      LAYER via2 ;
        RECT 2901.310 2903.800 2901.590 2904.080 ;
        RECT 2618.410 2693.000 2618.690 2693.280 ;
      LAYER met3 ;
        RECT 2901.285 2904.090 2901.615 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2901.285 2903.790 2924.800 2904.090 ;
        RECT 2901.285 2903.775 2901.615 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2606.000 2693.290 2610.000 2693.680 ;
        RECT 2618.385 2693.290 2618.715 2693.305 ;
        RECT 2606.000 2693.080 2618.715 2693.290 ;
        RECT 2609.580 2692.990 2618.715 2693.080 ;
        RECT 2618.385 2692.975 2618.715 2692.990 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 2898.060 2621.930 2898.120 ;
        RECT 2901.750 2898.060 2902.070 2898.120 ;
        RECT 2621.610 2897.920 2902.070 2898.060 ;
        RECT 2621.610 2897.860 2621.930 2897.920 ;
        RECT 2901.750 2897.860 2902.070 2897.920 ;
      LAYER via ;
        RECT 2621.640 2897.860 2621.900 2898.120 ;
        RECT 2901.780 2897.860 2902.040 2898.120 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 2901.840 2898.150 2901.980 3138.355 ;
        RECT 2621.640 2897.830 2621.900 2898.150 ;
        RECT 2901.780 2897.830 2902.040 2898.150 ;
        RECT 2621.700 2893.245 2621.840 2897.830 ;
        RECT 2621.630 2892.875 2621.910 2893.245 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
        RECT 2621.630 2892.920 2621.910 2893.200 ;
      LAYER met3 ;
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2606.000 2893.210 2610.000 2893.600 ;
        RECT 2621.605 2893.210 2621.935 2893.225 ;
        RECT 2606.000 2893.000 2621.935 2893.210 ;
        RECT 2609.580 2892.910 2621.935 2893.000 ;
        RECT 2621.605 2892.895 2621.935 2892.910 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 3097.980 2621.930 3098.040 ;
        RECT 2901.290 3097.980 2901.610 3098.040 ;
        RECT 2621.610 3097.840 2901.610 3097.980 ;
        RECT 2621.610 3097.780 2621.930 3097.840 ;
        RECT 2901.290 3097.780 2901.610 3097.840 ;
      LAYER via ;
        RECT 2621.640 3097.780 2621.900 3098.040 ;
        RECT 2901.320 3097.780 2901.580 3098.040 ;
      LAYER met2 ;
        RECT 2901.310 3372.955 2901.590 3373.325 ;
        RECT 2901.380 3098.070 2901.520 3372.955 ;
        RECT 2621.640 3097.750 2621.900 3098.070 ;
        RECT 2901.320 3097.750 2901.580 3098.070 ;
        RECT 2621.700 3093.165 2621.840 3097.750 ;
        RECT 2621.630 3092.795 2621.910 3093.165 ;
      LAYER via2 ;
        RECT 2901.310 3373.000 2901.590 3373.280 ;
        RECT 2621.630 3092.840 2621.910 3093.120 ;
      LAYER met3 ;
        RECT 2901.285 3373.290 2901.615 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2901.285 3372.990 2924.800 3373.290 ;
        RECT 2901.285 3372.975 2901.615 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2606.000 3093.130 2610.000 3093.520 ;
        RECT 2621.605 3093.130 2621.935 3093.145 ;
        RECT 2606.000 3092.920 2621.935 3093.130 ;
        RECT 2609.580 3092.830 2621.935 3092.920 ;
        RECT 2621.605 3092.815 2621.935 3092.830 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 3502.240 2573.630 3502.300 ;
        RECT 2798.250 3502.240 2798.570 3502.300 ;
        RECT 2573.310 3502.100 2798.570 3502.240 ;
        RECT 2573.310 3502.040 2573.630 3502.100 ;
        RECT 2798.250 3502.040 2798.570 3502.100 ;
        RECT 2566.870 3276.480 2567.190 3276.540 ;
        RECT 2573.310 3276.480 2573.630 3276.540 ;
        RECT 2566.870 3276.340 2573.630 3276.480 ;
        RECT 2566.870 3276.280 2567.190 3276.340 ;
        RECT 2573.310 3276.280 2573.630 3276.340 ;
      LAYER via ;
        RECT 2573.340 3502.040 2573.600 3502.300 ;
        RECT 2798.280 3502.040 2798.540 3502.300 ;
        RECT 2566.900 3276.280 2567.160 3276.540 ;
        RECT 2573.340 3276.280 2573.600 3276.540 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3502.330 2798.480 3517.600 ;
        RECT 2573.340 3502.010 2573.600 3502.330 ;
        RECT 2798.280 3502.010 2798.540 3502.330 ;
        RECT 2573.400 3276.570 2573.540 3502.010 ;
        RECT 2566.900 3276.250 2567.160 3276.570 ;
        RECT 2573.340 3276.250 2573.600 3276.570 ;
        RECT 2566.960 3260.000 2567.100 3276.250 ;
        RECT 2566.850 3256.000 2567.130 3260.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2318.010 3502.240 2318.330 3502.300 ;
        RECT 2473.950 3502.240 2474.270 3502.300 ;
        RECT 2318.010 3502.100 2474.270 3502.240 ;
        RECT 2318.010 3502.040 2318.330 3502.100 ;
        RECT 2473.950 3502.040 2474.270 3502.100 ;
        RECT 2311.570 3277.500 2311.890 3277.560 ;
        RECT 2318.010 3277.500 2318.330 3277.560 ;
        RECT 2311.570 3277.360 2318.330 3277.500 ;
        RECT 2311.570 3277.300 2311.890 3277.360 ;
        RECT 2318.010 3277.300 2318.330 3277.360 ;
      LAYER via ;
        RECT 2318.040 3502.040 2318.300 3502.300 ;
        RECT 2473.980 3502.040 2474.240 3502.300 ;
        RECT 2311.600 3277.300 2311.860 3277.560 ;
        RECT 2318.040 3277.300 2318.300 3277.560 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3502.330 2474.180 3517.600 ;
        RECT 2318.040 3502.010 2318.300 3502.330 ;
        RECT 2473.980 3502.010 2474.240 3502.330 ;
        RECT 2318.100 3277.590 2318.240 3502.010 ;
        RECT 2311.600 3277.270 2311.860 3277.590 ;
        RECT 2318.040 3277.270 2318.300 3277.590 ;
        RECT 2311.660 3260.000 2311.800 3277.270 ;
        RECT 2311.550 3256.000 2311.830 3260.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 3502.240 2056.130 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 2055.810 3502.100 2149.510 3502.240 ;
        RECT 2055.810 3502.040 2056.130 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
      LAYER via ;
        RECT 2055.840 3502.040 2056.100 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 2055.840 3502.010 2056.100 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 2055.900 3260.000 2056.040 3502.010 ;
        RECT 2055.790 3256.000 2056.070 3260.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.510 3498.500 1800.830 3498.560 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1800.510 3498.360 1825.210 3498.500 ;
        RECT 1800.510 3498.300 1800.830 3498.360 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
      LAYER via ;
        RECT 1800.540 3498.300 1800.800 3498.560 ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1800.540 3498.270 1800.800 3498.590 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1800.600 3260.000 1800.740 3498.270 ;
        RECT 1800.490 3256.000 1800.770 3260.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 3270.700 1504.130 3270.760 ;
        RECT 1544.750 3270.700 1545.070 3270.760 ;
        RECT 1503.810 3270.560 1545.070 3270.700 ;
        RECT 1503.810 3270.500 1504.130 3270.560 ;
        RECT 1544.750 3270.500 1545.070 3270.560 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 3270.500 1504.100 3270.760 ;
        RECT 1544.780 3270.500 1545.040 3270.760 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3270.790 1504.040 3498.270 ;
        RECT 1503.840 3270.470 1504.100 3270.790 ;
        RECT 1544.780 3270.470 1545.040 3270.790 ;
        RECT 1544.840 3260.000 1544.980 3270.470 ;
        RECT 1544.730 3256.000 1545.010 3260.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 324.260 2619.630 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2619.310 324.120 2899.310 324.260 ;
        RECT 2619.310 324.060 2619.630 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2619.340 324.060 2619.600 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2619.330 493.155 2619.610 493.525 ;
        RECT 2619.400 324.350 2619.540 493.155 ;
        RECT 2619.340 324.030 2619.600 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2619.330 493.200 2619.610 493.480 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2606.000 493.490 2610.000 493.880 ;
        RECT 2619.305 493.490 2619.635 493.505 ;
        RECT 2606.000 493.280 2619.635 493.490 ;
        RECT 2609.580 493.190 2619.635 493.280 ;
        RECT 2619.305 493.175 2619.635 493.190 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3274.100 1179.830 3274.160 ;
        RECT 1289.450 3274.100 1289.770 3274.160 ;
        RECT 1179.510 3273.960 1289.770 3274.100 ;
        RECT 1179.510 3273.900 1179.830 3273.960 ;
        RECT 1289.450 3273.900 1289.770 3273.960 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3273.900 1179.800 3274.160 ;
        RECT 1289.480 3273.900 1289.740 3274.160 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3274.190 1179.740 3498.270 ;
        RECT 1179.540 3273.870 1179.800 3274.190 ;
        RECT 1289.480 3273.870 1289.740 3274.190 ;
        RECT 1289.540 3260.000 1289.680 3273.870 ;
        RECT 1289.430 3256.000 1289.710 3260.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 855.210 3501.220 855.530 3501.280 ;
        RECT 851.530 3501.080 855.530 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 855.210 3501.020 855.530 3501.080 ;
        RECT 855.210 3274.440 855.530 3274.500 ;
        RECT 1033.690 3274.440 1034.010 3274.500 ;
        RECT 855.210 3274.300 1034.010 3274.440 ;
        RECT 855.210 3274.240 855.530 3274.300 ;
        RECT 1033.690 3274.240 1034.010 3274.300 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 855.240 3501.020 855.500 3501.280 ;
        RECT 855.240 3274.240 855.500 3274.500 ;
        RECT 1033.720 3274.240 1033.980 3274.500 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 855.240 3500.990 855.500 3501.310 ;
        RECT 855.300 3274.530 855.440 3500.990 ;
        RECT 855.240 3274.210 855.500 3274.530 ;
        RECT 1033.720 3274.210 1033.980 3274.530 ;
        RECT 1033.780 3260.000 1033.920 3274.210 ;
        RECT 1033.670 3256.000 1033.950 3260.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 3274.780 531.230 3274.840 ;
        RECT 777.930 3274.780 778.250 3274.840 ;
        RECT 530.910 3274.640 778.250 3274.780 ;
        RECT 530.910 3274.580 531.230 3274.640 ;
        RECT 777.930 3274.580 778.250 3274.640 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 3274.580 531.200 3274.840 ;
        RECT 777.960 3274.580 778.220 3274.840 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 3274.870 531.140 3498.270 ;
        RECT 530.940 3274.550 531.200 3274.870 ;
        RECT 777.960 3274.550 778.220 3274.870 ;
        RECT 778.020 3260.000 778.160 3274.550 ;
        RECT 777.910 3256.000 778.190 3260.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 3274.780 206.930 3274.840 ;
        RECT 522.630 3274.780 522.950 3274.840 ;
        RECT 206.610 3274.640 522.950 3274.780 ;
        RECT 206.610 3274.580 206.930 3274.640 ;
        RECT 522.630 3274.580 522.950 3274.640 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 3274.580 206.900 3274.840 ;
        RECT 522.660 3274.580 522.920 3274.840 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 3274.870 206.840 3501.670 ;
        RECT 206.640 3274.550 206.900 3274.870 ;
        RECT 522.660 3274.550 522.920 3274.870 ;
        RECT 522.720 3260.000 522.860 3274.550 ;
        RECT 522.610 3256.000 522.890 3260.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3229.220 17.870 3229.280 ;
        RECT 296.770 3229.220 297.090 3229.280 ;
        RECT 17.550 3229.080 297.090 3229.220 ;
        RECT 17.550 3229.020 17.870 3229.080 ;
        RECT 296.770 3229.020 297.090 3229.080 ;
      LAYER via ;
        RECT 17.580 3229.020 17.840 3229.280 ;
        RECT 296.800 3229.020 297.060 3229.280 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3229.310 17.780 3411.035 ;
        RECT 17.580 3228.990 17.840 3229.310 ;
        RECT 296.800 3228.990 297.060 3229.310 ;
        RECT 296.860 3223.725 297.000 3228.990 ;
        RECT 296.790 3223.355 297.070 3223.725 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
        RECT 296.790 3223.400 297.070 3223.680 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
        RECT 296.765 3223.690 297.095 3223.705 ;
        RECT 310.000 3223.690 314.000 3224.080 ;
        RECT 296.765 3223.480 314.000 3223.690 ;
        RECT 296.765 3223.390 310.500 3223.480 ;
        RECT 296.765 3223.375 297.095 3223.390 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3015.360 17.870 3015.420 ;
        RECT 296.770 3015.360 297.090 3015.420 ;
        RECT 17.550 3015.220 297.090 3015.360 ;
        RECT 17.550 3015.160 17.870 3015.220 ;
        RECT 296.770 3015.160 297.090 3015.220 ;
      LAYER via ;
        RECT 17.580 3015.160 17.840 3015.420 ;
        RECT 296.800 3015.160 297.060 3015.420 ;
      LAYER met2 ;
        RECT 17.570 3124.075 17.850 3124.445 ;
        RECT 17.640 3015.450 17.780 3124.075 ;
        RECT 17.580 3015.130 17.840 3015.450 ;
        RECT 296.800 3015.130 297.060 3015.450 ;
        RECT 296.860 3009.525 297.000 3015.130 ;
        RECT 296.790 3009.155 297.070 3009.525 ;
      LAYER via2 ;
        RECT 17.570 3124.120 17.850 3124.400 ;
        RECT 296.790 3009.200 297.070 3009.480 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.545 3124.410 17.875 3124.425 ;
        RECT -4.800 3124.110 17.875 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.545 3124.095 17.875 3124.110 ;
        RECT 296.765 3009.490 297.095 3009.505 ;
        RECT 310.000 3009.490 314.000 3009.880 ;
        RECT 296.765 3009.280 314.000 3009.490 ;
        RECT 296.765 3009.190 310.500 3009.280 ;
        RECT 296.765 3009.175 297.095 3009.190 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2801.160 17.410 2801.220 ;
        RECT 296.770 2801.160 297.090 2801.220 ;
        RECT 17.090 2801.020 297.090 2801.160 ;
        RECT 17.090 2800.960 17.410 2801.020 ;
        RECT 296.770 2800.960 297.090 2801.020 ;
      LAYER via ;
        RECT 17.120 2800.960 17.380 2801.220 ;
        RECT 296.800 2800.960 297.060 2801.220 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2801.250 17.320 2836.435 ;
        RECT 17.120 2800.930 17.380 2801.250 ;
        RECT 296.800 2800.930 297.060 2801.250 ;
        RECT 296.860 2795.325 297.000 2800.930 ;
        RECT 296.790 2794.955 297.070 2795.325 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
        RECT 296.790 2795.000 297.070 2795.280 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
        RECT 296.765 2795.290 297.095 2795.305 ;
        RECT 310.000 2795.290 314.000 2795.680 ;
        RECT 296.765 2795.080 314.000 2795.290 ;
        RECT 296.765 2794.990 310.500 2795.080 ;
        RECT 296.765 2794.975 297.095 2794.990 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 2552.960 16.030 2553.020 ;
        RECT 296.770 2552.960 297.090 2553.020 ;
        RECT 15.710 2552.820 297.090 2552.960 ;
        RECT 15.710 2552.760 16.030 2552.820 ;
        RECT 296.770 2552.760 297.090 2552.820 ;
      LAYER via ;
        RECT 15.740 2552.760 16.000 2553.020 ;
        RECT 296.800 2552.760 297.060 2553.020 ;
      LAYER met2 ;
        RECT 296.790 2580.755 297.070 2581.125 ;
        RECT 296.860 2553.050 297.000 2580.755 ;
        RECT 15.740 2552.730 16.000 2553.050 ;
        RECT 296.800 2552.730 297.060 2553.050 ;
        RECT 15.800 2549.845 15.940 2552.730 ;
        RECT 15.730 2549.475 16.010 2549.845 ;
      LAYER via2 ;
        RECT 296.790 2580.800 297.070 2581.080 ;
        RECT 15.730 2549.520 16.010 2549.800 ;
      LAYER met3 ;
        RECT 296.765 2581.090 297.095 2581.105 ;
        RECT 310.000 2581.090 314.000 2581.480 ;
        RECT 296.765 2580.880 314.000 2581.090 ;
        RECT 296.765 2580.790 310.500 2580.880 ;
        RECT 296.765 2580.775 297.095 2580.790 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 15.705 2549.810 16.035 2549.825 ;
        RECT -4.800 2549.510 16.035 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 15.705 2549.495 16.035 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2262.940 17.410 2263.000 ;
        RECT 299.990 2262.940 300.310 2263.000 ;
        RECT 17.090 2262.800 300.310 2262.940 ;
        RECT 17.090 2262.740 17.410 2262.800 ;
        RECT 299.990 2262.740 300.310 2262.800 ;
      LAYER via ;
        RECT 17.120 2262.740 17.380 2263.000 ;
        RECT 300.020 2262.740 300.280 2263.000 ;
      LAYER met2 ;
        RECT 300.010 2366.555 300.290 2366.925 ;
        RECT 300.080 2263.030 300.220 2366.555 ;
        RECT 17.120 2262.710 17.380 2263.030 ;
        RECT 300.020 2262.710 300.280 2263.030 ;
        RECT 17.180 2262.205 17.320 2262.710 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
      LAYER via2 ;
        RECT 300.010 2366.600 300.290 2366.880 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
        RECT 299.985 2366.890 300.315 2366.905 ;
        RECT 310.000 2366.890 314.000 2367.280 ;
        RECT 299.985 2366.680 314.000 2366.890 ;
        RECT 299.985 2366.590 310.500 2366.680 ;
        RECT 299.985 2366.575 300.315 2366.590 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 300.450 1980.060 300.770 1980.120 ;
        RECT 15.710 1979.920 300.770 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 300.450 1979.860 300.770 1979.920 ;
      LAYER via ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 300.480 1979.860 300.740 1980.120 ;
      LAYER met2 ;
        RECT 300.470 2152.355 300.750 2152.725 ;
        RECT 300.540 1980.150 300.680 2152.355 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 300.480 1979.830 300.740 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 300.470 2152.400 300.750 2152.680 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT 300.445 2152.690 300.775 2152.705 ;
        RECT 310.000 2152.690 314.000 2153.080 ;
        RECT 300.445 2152.480 314.000 2152.690 ;
        RECT 300.445 2152.390 310.500 2152.480 ;
        RECT 300.445 2152.375 300.775 2152.390 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 558.860 2619.630 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2619.310 558.720 2899.310 558.860 ;
        RECT 2619.310 558.660 2619.630 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2619.340 558.660 2619.600 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2619.330 693.075 2619.610 693.445 ;
        RECT 2619.400 558.950 2619.540 693.075 ;
        RECT 2619.340 558.630 2619.600 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2619.330 693.120 2619.610 693.400 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2606.000 693.410 2610.000 693.800 ;
        RECT 2619.305 693.410 2619.635 693.425 ;
        RECT 2606.000 693.200 2619.635 693.410 ;
        RECT 2609.580 693.110 2619.635 693.200 ;
        RECT 2619.305 693.095 2619.635 693.110 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 300.450 1690.380 300.770 1690.440 ;
        RECT 17.090 1690.240 300.770 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 300.450 1690.180 300.770 1690.240 ;
      LAYER via ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 300.480 1690.180 300.740 1690.440 ;
      LAYER met2 ;
        RECT 300.470 1938.155 300.750 1938.525 ;
        RECT 300.540 1690.470 300.680 1938.155 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 300.480 1690.150 300.740 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 300.470 1938.200 300.750 1938.480 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT 300.445 1938.490 300.775 1938.505 ;
        RECT 310.000 1938.490 314.000 1938.880 ;
        RECT 300.445 1938.280 314.000 1938.490 ;
        RECT 300.445 1938.190 310.500 1938.280 ;
        RECT 300.445 1938.175 300.775 1938.190 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1476.520 17.410 1476.580 ;
        RECT 301.830 1476.520 302.150 1476.580 ;
        RECT 17.090 1476.380 302.150 1476.520 ;
        RECT 17.090 1476.320 17.410 1476.380 ;
        RECT 301.830 1476.320 302.150 1476.380 ;
      LAYER via ;
        RECT 17.120 1476.320 17.380 1476.580 ;
        RECT 301.860 1476.320 302.120 1476.580 ;
      LAYER met2 ;
        RECT 301.850 1723.275 302.130 1723.645 ;
        RECT 301.920 1476.610 302.060 1723.275 ;
        RECT 17.120 1476.290 17.380 1476.610 ;
        RECT 301.860 1476.290 302.120 1476.610 ;
        RECT 17.180 1472.045 17.320 1476.290 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 301.850 1723.320 302.130 1723.600 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT 301.825 1723.610 302.155 1723.625 ;
        RECT 310.000 1723.610 314.000 1724.000 ;
        RECT 301.825 1723.400 314.000 1723.610 ;
        RECT 301.825 1723.310 310.500 1723.400 ;
        RECT 301.825 1723.295 302.155 1723.310 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1262.660 17.410 1262.720 ;
        RECT 302.290 1262.660 302.610 1262.720 ;
        RECT 17.090 1262.520 302.610 1262.660 ;
        RECT 17.090 1262.460 17.410 1262.520 ;
        RECT 302.290 1262.460 302.610 1262.520 ;
      LAYER via ;
        RECT 17.120 1262.460 17.380 1262.720 ;
        RECT 302.320 1262.460 302.580 1262.720 ;
      LAYER met2 ;
        RECT 302.310 1509.075 302.590 1509.445 ;
        RECT 302.380 1262.750 302.520 1509.075 ;
        RECT 17.120 1262.430 17.380 1262.750 ;
        RECT 302.320 1262.430 302.580 1262.750 ;
        RECT 17.180 1256.485 17.320 1262.430 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
      LAYER via2 ;
        RECT 302.310 1509.120 302.590 1509.400 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
      LAYER met3 ;
        RECT 302.285 1509.410 302.615 1509.425 ;
        RECT 310.000 1509.410 314.000 1509.800 ;
        RECT 302.285 1509.200 314.000 1509.410 ;
        RECT 302.285 1509.110 310.500 1509.200 ;
        RECT 302.285 1509.095 302.615 1509.110 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 300.450 1041.660 300.770 1041.720 ;
        RECT 17.090 1041.520 300.770 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 300.450 1041.460 300.770 1041.520 ;
      LAYER via ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 300.480 1041.460 300.740 1041.720 ;
      LAYER met2 ;
        RECT 300.470 1294.875 300.750 1295.245 ;
        RECT 300.540 1041.750 300.680 1294.875 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 300.480 1041.430 300.740 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 300.470 1294.920 300.750 1295.200 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT 300.445 1295.210 300.775 1295.225 ;
        RECT 310.000 1295.210 314.000 1295.600 ;
        RECT 300.445 1295.000 314.000 1295.210 ;
        RECT 300.445 1294.910 310.500 1295.000 ;
        RECT 300.445 1294.895 300.775 1294.910 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 300.910 827.800 301.230 827.860 ;
        RECT 17.550 827.660 301.230 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 300.910 827.600 301.230 827.660 ;
      LAYER via ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 300.940 827.600 301.200 827.860 ;
      LAYER met2 ;
        RECT 300.930 1080.675 301.210 1081.045 ;
        RECT 301.000 827.890 301.140 1080.675 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 300.940 827.570 301.200 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 300.930 1080.720 301.210 1081.000 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT 300.905 1081.010 301.235 1081.025 ;
        RECT 310.000 1081.010 314.000 1081.400 ;
        RECT 300.905 1080.800 314.000 1081.010 ;
        RECT 300.905 1080.710 310.500 1080.800 ;
        RECT 300.905 1080.695 301.235 1080.710 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 613.940 17.410 614.000 ;
        RECT 301.830 613.940 302.150 614.000 ;
        RECT 17.090 613.800 302.150 613.940 ;
        RECT 17.090 613.740 17.410 613.800 ;
        RECT 301.830 613.740 302.150 613.800 ;
      LAYER via ;
        RECT 17.120 613.740 17.380 614.000 ;
        RECT 301.860 613.740 302.120 614.000 ;
      LAYER met2 ;
        RECT 301.850 866.475 302.130 866.845 ;
        RECT 301.920 614.030 302.060 866.475 ;
        RECT 17.120 613.710 17.380 614.030 ;
        RECT 301.860 613.710 302.120 614.030 ;
        RECT 17.180 610.485 17.320 613.710 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 301.850 866.520 302.130 866.800 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT 301.825 866.810 302.155 866.825 ;
        RECT 310.000 866.810 314.000 867.200 ;
        RECT 301.825 866.600 314.000 866.810 ;
        RECT 301.825 866.510 310.500 866.600 ;
        RECT 301.825 866.495 302.155 866.510 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 400.080 17.410 400.140 ;
        RECT 299.990 400.080 300.310 400.140 ;
        RECT 17.090 399.940 300.310 400.080 ;
        RECT 17.090 399.880 17.410 399.940 ;
        RECT 299.990 399.880 300.310 399.940 ;
      LAYER via ;
        RECT 17.120 399.880 17.380 400.140 ;
        RECT 300.020 399.880 300.280 400.140 ;
      LAYER met2 ;
        RECT 300.010 652.275 300.290 652.645 ;
        RECT 300.080 400.170 300.220 652.275 ;
        RECT 17.120 399.850 17.380 400.170 ;
        RECT 300.020 399.850 300.280 400.170 ;
        RECT 17.180 394.925 17.320 399.850 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 300.010 652.320 300.290 652.600 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT 299.985 652.610 300.315 652.625 ;
        RECT 310.000 652.610 314.000 653.000 ;
        RECT 299.985 652.400 314.000 652.610 ;
        RECT 299.985 652.310 310.500 652.400 ;
        RECT 299.985 652.295 300.315 652.310 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 300.910 179.420 301.230 179.480 ;
        RECT 17.090 179.280 301.230 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 300.910 179.220 301.230 179.280 ;
      LAYER via ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 300.940 179.220 301.200 179.480 ;
      LAYER met2 ;
        RECT 300.930 438.075 301.210 438.445 ;
        RECT 301.000 179.510 301.140 438.075 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 300.940 179.190 301.200 179.510 ;
      LAYER via2 ;
        RECT 300.930 438.120 301.210 438.400 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 300.905 438.410 301.235 438.425 ;
        RECT 310.000 438.410 314.000 438.800 ;
        RECT 300.905 438.200 314.000 438.410 ;
        RECT 300.905 438.110 310.500 438.200 ;
        RECT 300.905 438.095 301.235 438.110 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 793.460 2619.630 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2619.310 793.320 2899.310 793.460 ;
        RECT 2619.310 793.260 2619.630 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2619.340 793.260 2619.600 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2619.330 892.995 2619.610 893.365 ;
        RECT 2619.400 793.550 2619.540 892.995 ;
        RECT 2619.340 793.230 2619.600 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2619.330 893.040 2619.610 893.320 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2606.000 893.330 2610.000 893.720 ;
        RECT 2619.305 893.330 2619.635 893.345 ;
        RECT 2606.000 893.120 2619.635 893.330 ;
        RECT 2609.580 893.030 2619.635 893.120 ;
        RECT 2619.305 893.015 2619.635 893.030 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 1028.060 2619.630 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2619.310 1027.920 2899.310 1028.060 ;
        RECT 2619.310 1027.860 2619.630 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2619.340 1027.860 2619.600 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2619.330 1092.915 2619.610 1093.285 ;
        RECT 2619.400 1028.150 2619.540 1092.915 ;
        RECT 2619.340 1027.830 2619.600 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2619.330 1092.960 2619.610 1093.240 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2606.000 1093.250 2610.000 1093.640 ;
        RECT 2619.305 1093.250 2619.635 1093.265 ;
        RECT 2606.000 1093.040 2619.635 1093.250 ;
        RECT 2609.580 1092.950 2619.635 1093.040 ;
        RECT 2619.305 1092.935 2619.635 1092.950 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1262.660 2618.710 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 2618.390 1262.520 2899.310 1262.660 ;
        RECT 2618.390 1262.460 2618.710 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 2618.420 1262.460 2618.680 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 2618.410 1292.835 2618.690 1293.205 ;
        RECT 2618.480 1262.750 2618.620 1292.835 ;
        RECT 2618.420 1262.430 2618.680 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2618.410 1292.880 2618.690 1293.160 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2606.000 1293.170 2610.000 1293.560 ;
        RECT 2618.385 1293.170 2618.715 1293.185 ;
        RECT 2606.000 1292.960 2618.715 1293.170 ;
        RECT 2609.580 1292.870 2618.715 1292.960 ;
        RECT 2618.385 1292.855 2618.715 1292.870 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1493.860 2621.930 1493.920 ;
        RECT 2900.830 1493.860 2901.150 1493.920 ;
        RECT 2621.610 1493.720 2901.150 1493.860 ;
        RECT 2621.610 1493.660 2621.930 1493.720 ;
        RECT 2900.830 1493.660 2901.150 1493.720 ;
      LAYER via ;
        RECT 2621.640 1493.660 2621.900 1493.920 ;
        RECT 2900.860 1493.660 2901.120 1493.920 ;
      LAYER met2 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
        RECT 2900.920 1493.950 2901.060 1495.475 ;
        RECT 2621.640 1493.630 2621.900 1493.950 ;
        RECT 2900.860 1493.630 2901.120 1493.950 ;
        RECT 2621.700 1493.125 2621.840 1493.630 ;
        RECT 2621.630 1492.755 2621.910 1493.125 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
        RECT 2621.630 1492.800 2621.910 1493.080 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2606.000 1493.090 2610.000 1493.480 ;
        RECT 2621.605 1493.090 2621.935 1493.105 ;
        RECT 2606.000 1492.880 2621.935 1493.090 ;
        RECT 2609.580 1492.790 2621.935 1492.880 ;
        RECT 2621.605 1492.775 2621.935 1492.790 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1725.400 2619.170 1725.460 ;
        RECT 2900.830 1725.400 2901.150 1725.460 ;
        RECT 2618.850 1725.260 2901.150 1725.400 ;
        RECT 2618.850 1725.200 2619.170 1725.260 ;
        RECT 2900.830 1725.200 2901.150 1725.260 ;
      LAYER via ;
        RECT 2618.880 1725.200 2619.140 1725.460 ;
        RECT 2900.860 1725.200 2901.120 1725.460 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 2900.920 1725.490 2901.060 1730.075 ;
        RECT 2618.880 1725.170 2619.140 1725.490 ;
        RECT 2900.860 1725.170 2901.120 1725.490 ;
        RECT 2618.940 1693.045 2619.080 1725.170 ;
        RECT 2618.870 1692.675 2619.150 1693.045 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
        RECT 2618.870 1692.720 2619.150 1693.000 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2606.000 1693.010 2610.000 1693.400 ;
        RECT 2618.845 1693.010 2619.175 1693.025 ;
        RECT 2606.000 1692.800 2619.175 1693.010 ;
        RECT 2609.580 1692.710 2619.175 1692.800 ;
        RECT 2618.845 1692.695 2619.175 1692.710 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1960.000 2618.710 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 2618.390 1959.860 2901.150 1960.000 ;
        RECT 2618.390 1959.800 2618.710 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
      LAYER via ;
        RECT 2618.420 1959.800 2618.680 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 2618.420 1959.770 2618.680 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 2618.480 1893.645 2618.620 1959.770 ;
        RECT 2618.410 1893.275 2618.690 1893.645 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
        RECT 2618.410 1893.320 2618.690 1893.600 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2606.000 1893.610 2610.000 1894.000 ;
        RECT 2618.385 1893.610 2618.715 1893.625 ;
        RECT 2606.000 1893.400 2618.715 1893.610 ;
        RECT 2609.580 1893.310 2618.715 1893.400 ;
        RECT 2618.385 1893.295 2618.715 1893.310 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2194.600 2618.710 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2618.390 2194.460 2901.150 2194.600 ;
        RECT 2618.390 2194.400 2618.710 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
      LAYER via ;
        RECT 2618.420 2194.400 2618.680 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2618.420 2194.370 2618.680 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2618.480 2093.565 2618.620 2194.370 ;
        RECT 2618.410 2093.195 2618.690 2093.565 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2618.410 2093.240 2618.690 2093.520 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2606.000 2093.530 2610.000 2093.920 ;
        RECT 2618.385 2093.530 2618.715 2093.545 ;
        RECT 2606.000 2093.320 2618.715 2093.530 ;
        RECT 2609.580 2093.230 2618.715 2093.320 ;
        RECT 2618.385 2093.215 2618.715 2093.230 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 206.960 2618.710 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2618.390 206.820 2901.150 206.960 ;
        RECT 2618.390 206.760 2618.710 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2618.420 206.760 2618.680 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2618.410 426.515 2618.690 426.885 ;
        RECT 2618.480 207.050 2618.620 426.515 ;
        RECT 2618.420 206.730 2618.680 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2618.410 426.560 2618.690 426.840 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2606.000 426.850 2610.000 427.240 ;
        RECT 2618.385 426.850 2618.715 426.865 ;
        RECT 2606.000 426.640 2618.715 426.850 ;
        RECT 2609.580 426.550 2618.715 426.640 ;
        RECT 2618.385 426.535 2618.715 426.550 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2546.500 2619.170 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2618.850 2546.360 2901.150 2546.500 ;
        RECT 2618.850 2546.300 2619.170 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
      LAYER via ;
        RECT 2618.880 2546.300 2619.140 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2618.880 2546.270 2619.140 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2618.940 2426.765 2619.080 2546.270 ;
        RECT 2618.870 2426.395 2619.150 2426.765 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2618.870 2426.440 2619.150 2426.720 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2606.000 2426.730 2610.000 2427.120 ;
        RECT 2618.845 2426.730 2619.175 2426.745 ;
        RECT 2606.000 2426.520 2619.175 2426.730 ;
        RECT 2609.580 2426.430 2619.175 2426.520 ;
        RECT 2618.845 2426.415 2619.175 2426.430 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2781.100 2619.170 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2618.850 2780.960 2901.150 2781.100 ;
        RECT 2618.850 2780.900 2619.170 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 2618.880 2780.900 2619.140 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2618.880 2780.870 2619.140 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2618.940 2626.685 2619.080 2780.870 ;
        RECT 2618.870 2626.315 2619.150 2626.685 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2618.870 2626.360 2619.150 2626.640 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2606.000 2626.650 2610.000 2627.040 ;
        RECT 2618.845 2626.650 2619.175 2626.665 ;
        RECT 2606.000 2626.440 2619.175 2626.650 ;
        RECT 2609.580 2626.350 2619.175 2626.440 ;
        RECT 2618.845 2626.335 2619.175 2626.350 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.630 2829.040 2615.950 2829.100 ;
        RECT 2902.210 2829.040 2902.530 2829.100 ;
        RECT 2615.630 2828.900 2902.530 2829.040 ;
        RECT 2615.630 2828.840 2615.950 2828.900 ;
        RECT 2902.210 2828.840 2902.530 2828.900 ;
      LAYER via ;
        RECT 2615.660 2828.840 2615.920 2829.100 ;
        RECT 2902.240 2828.840 2902.500 2829.100 ;
      LAYER met2 ;
        RECT 2902.230 3020.715 2902.510 3021.085 ;
        RECT 2902.300 2829.130 2902.440 3020.715 ;
        RECT 2615.660 2828.810 2615.920 2829.130 ;
        RECT 2902.240 2828.810 2902.500 2829.130 ;
        RECT 2615.720 2826.605 2615.860 2828.810 ;
        RECT 2615.650 2826.235 2615.930 2826.605 ;
      LAYER via2 ;
        RECT 2902.230 3020.760 2902.510 3021.040 ;
        RECT 2615.650 2826.280 2615.930 2826.560 ;
      LAYER met3 ;
        RECT 2902.205 3021.050 2902.535 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2902.205 3020.750 2924.800 3021.050 ;
        RECT 2902.205 3020.735 2902.535 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2606.000 2826.570 2610.000 2826.960 ;
        RECT 2615.625 2826.570 2615.955 2826.585 ;
        RECT 2606.000 2826.360 2615.955 2826.570 ;
        RECT 2609.580 2826.270 2615.955 2826.360 ;
        RECT 2615.625 2826.255 2615.955 2826.270 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.630 3028.960 2615.950 3029.020 ;
        RECT 2902.210 3028.960 2902.530 3029.020 ;
        RECT 2615.630 3028.820 2902.530 3028.960 ;
        RECT 2615.630 3028.760 2615.950 3028.820 ;
        RECT 2902.210 3028.760 2902.530 3028.820 ;
      LAYER via ;
        RECT 2615.660 3028.760 2615.920 3029.020 ;
        RECT 2902.240 3028.760 2902.500 3029.020 ;
      LAYER met2 ;
        RECT 2902.230 3255.315 2902.510 3255.685 ;
        RECT 2902.300 3029.050 2902.440 3255.315 ;
        RECT 2615.660 3028.730 2615.920 3029.050 ;
        RECT 2902.240 3028.730 2902.500 3029.050 ;
        RECT 2615.720 3026.525 2615.860 3028.730 ;
        RECT 2615.650 3026.155 2615.930 3026.525 ;
      LAYER via2 ;
        RECT 2902.230 3255.360 2902.510 3255.640 ;
        RECT 2615.650 3026.200 2615.930 3026.480 ;
      LAYER met3 ;
        RECT 2902.205 3255.650 2902.535 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2902.205 3255.350 2924.800 3255.650 ;
        RECT 2902.205 3255.335 2902.535 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2606.000 3026.490 2610.000 3026.880 ;
        RECT 2615.625 3026.490 2615.955 3026.505 ;
        RECT 2606.000 3026.280 2615.955 3026.490 ;
        RECT 2609.580 3026.190 2615.955 3026.280 ;
        RECT 2615.625 3026.175 2615.955 3026.190 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3484.900 2619.170 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2618.850 3484.760 2901.150 3484.900 ;
        RECT 2618.850 3484.700 2619.170 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 2618.880 3484.700 2619.140 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2618.880 3484.670 2619.140 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2618.940 3226.445 2619.080 3484.670 ;
        RECT 2618.870 3226.075 2619.150 3226.445 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2618.870 3226.120 2619.150 3226.400 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2606.000 3226.410 2610.000 3226.800 ;
        RECT 2618.845 3226.410 2619.175 3226.425 ;
        RECT 2606.000 3226.200 2619.175 3226.410 ;
        RECT 2609.580 3226.110 2619.175 3226.200 ;
        RECT 2618.845 3226.095 2619.175 3226.110 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2400.810 3501.560 2401.130 3501.620 ;
        RECT 2635.870 3501.560 2636.190 3501.620 ;
        RECT 2400.810 3501.420 2636.190 3501.560 ;
        RECT 2400.810 3501.360 2401.130 3501.420 ;
        RECT 2635.870 3501.360 2636.190 3501.420 ;
        RECT 2396.670 3277.500 2396.990 3277.560 ;
        RECT 2400.810 3277.500 2401.130 3277.560 ;
        RECT 2396.670 3277.360 2401.130 3277.500 ;
        RECT 2396.670 3277.300 2396.990 3277.360 ;
        RECT 2400.810 3277.300 2401.130 3277.360 ;
      LAYER via ;
        RECT 2400.840 3501.360 2401.100 3501.620 ;
        RECT 2635.900 3501.360 2636.160 3501.620 ;
        RECT 2396.700 3277.300 2396.960 3277.560 ;
        RECT 2400.840 3277.300 2401.100 3277.560 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.650 2636.100 3517.600 ;
        RECT 2400.840 3501.330 2401.100 3501.650 ;
        RECT 2635.900 3501.330 2636.160 3501.650 ;
        RECT 2400.900 3277.590 2401.040 3501.330 ;
        RECT 2396.700 3277.270 2396.960 3277.590 ;
        RECT 2400.840 3277.270 2401.100 3277.590 ;
        RECT 2396.760 3260.000 2396.900 3277.270 ;
        RECT 2396.650 3256.000 2396.930 3260.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2145.510 3501.560 2145.830 3501.620 ;
        RECT 2311.570 3501.560 2311.890 3501.620 ;
        RECT 2145.510 3501.420 2311.890 3501.560 ;
        RECT 2145.510 3501.360 2145.830 3501.420 ;
        RECT 2311.570 3501.360 2311.890 3501.420 ;
        RECT 2140.910 3277.500 2141.230 3277.560 ;
        RECT 2145.510 3277.500 2145.830 3277.560 ;
        RECT 2140.910 3277.360 2145.830 3277.500 ;
        RECT 2140.910 3277.300 2141.230 3277.360 ;
        RECT 2145.510 3277.300 2145.830 3277.360 ;
      LAYER via ;
        RECT 2145.540 3501.360 2145.800 3501.620 ;
        RECT 2311.600 3501.360 2311.860 3501.620 ;
        RECT 2140.940 3277.300 2141.200 3277.560 ;
        RECT 2145.540 3277.300 2145.800 3277.560 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.650 2311.800 3517.600 ;
        RECT 2145.540 3501.330 2145.800 3501.650 ;
        RECT 2311.600 3501.330 2311.860 3501.650 ;
        RECT 2145.600 3277.590 2145.740 3501.330 ;
        RECT 2140.940 3277.270 2141.200 3277.590 ;
        RECT 2145.540 3277.270 2145.800 3277.590 ;
        RECT 2141.000 3260.000 2141.140 3277.270 ;
        RECT 2140.890 3256.000 2141.170 3260.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1890.210 3501.560 1890.530 3501.620 ;
        RECT 1987.270 3501.560 1987.590 3501.620 ;
        RECT 1890.210 3501.420 1987.590 3501.560 ;
        RECT 1890.210 3501.360 1890.530 3501.420 ;
        RECT 1987.270 3501.360 1987.590 3501.420 ;
        RECT 1885.610 3277.500 1885.930 3277.560 ;
        RECT 1890.210 3277.500 1890.530 3277.560 ;
        RECT 1885.610 3277.360 1890.530 3277.500 ;
        RECT 1885.610 3277.300 1885.930 3277.360 ;
        RECT 1890.210 3277.300 1890.530 3277.360 ;
      LAYER via ;
        RECT 1890.240 3501.360 1890.500 3501.620 ;
        RECT 1987.300 3501.360 1987.560 3501.620 ;
        RECT 1885.640 3277.300 1885.900 3277.560 ;
        RECT 1890.240 3277.300 1890.500 3277.560 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3501.650 1987.500 3517.600 ;
        RECT 1890.240 3501.330 1890.500 3501.650 ;
        RECT 1987.300 3501.330 1987.560 3501.650 ;
        RECT 1890.300 3277.590 1890.440 3501.330 ;
        RECT 1885.640 3277.270 1885.900 3277.590 ;
        RECT 1890.240 3277.270 1890.500 3277.590 ;
        RECT 1885.700 3260.000 1885.840 3277.270 ;
        RECT 1885.590 3256.000 1885.870 3260.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1634.910 3498.500 1635.230 3498.560 ;
        RECT 1662.510 3498.500 1662.830 3498.560 ;
        RECT 1634.910 3498.360 1662.830 3498.500 ;
        RECT 1634.910 3498.300 1635.230 3498.360 ;
        RECT 1662.510 3498.300 1662.830 3498.360 ;
        RECT 1629.850 3275.800 1630.170 3275.860 ;
        RECT 1634.910 3275.800 1635.230 3275.860 ;
        RECT 1629.850 3275.660 1635.230 3275.800 ;
        RECT 1629.850 3275.600 1630.170 3275.660 ;
        RECT 1634.910 3275.600 1635.230 3275.660 ;
      LAYER via ;
        RECT 1634.940 3498.300 1635.200 3498.560 ;
        RECT 1662.540 3498.300 1662.800 3498.560 ;
        RECT 1629.880 3275.600 1630.140 3275.860 ;
        RECT 1634.940 3275.600 1635.200 3275.860 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3498.590 1662.740 3517.600 ;
        RECT 1634.940 3498.270 1635.200 3498.590 ;
        RECT 1662.540 3498.270 1662.800 3498.590 ;
        RECT 1635.000 3275.890 1635.140 3498.270 ;
        RECT 1629.880 3275.570 1630.140 3275.890 ;
        RECT 1634.940 3275.570 1635.200 3275.890 ;
        RECT 1629.940 3260.000 1630.080 3275.570 ;
        RECT 1629.830 3256.000 1630.110 3260.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3274.100 1338.530 3274.160 ;
        RECT 1374.550 3274.100 1374.870 3274.160 ;
        RECT 1338.210 3273.960 1374.870 3274.100 ;
        RECT 1338.210 3273.900 1338.530 3273.960 ;
        RECT 1374.550 3273.900 1374.870 3273.960 ;
      LAYER via ;
        RECT 1338.240 3273.900 1338.500 3274.160 ;
        RECT 1374.580 3273.900 1374.840 3274.160 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3274.190 1338.440 3517.600 ;
        RECT 1338.240 3273.870 1338.500 3274.190 ;
        RECT 1374.580 3273.870 1374.840 3274.190 ;
        RECT 1374.640 3260.000 1374.780 3273.870 ;
        RECT 1374.530 3256.000 1374.810 3260.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 441.560 2618.710 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2618.390 441.420 2901.150 441.560 ;
        RECT 2618.390 441.360 2618.710 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2618.420 441.360 2618.680 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2618.410 626.435 2618.690 626.805 ;
        RECT 2618.480 441.650 2618.620 626.435 ;
        RECT 2618.420 441.330 2618.680 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2618.410 626.480 2618.690 626.760 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2606.000 626.770 2610.000 627.160 ;
        RECT 2618.385 626.770 2618.715 626.785 ;
        RECT 2606.000 626.560 2618.715 626.770 ;
        RECT 2609.580 626.470 2618.715 626.560 ;
        RECT 2618.385 626.455 2618.715 626.470 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3274.100 1014.230 3274.160 ;
        RECT 1118.790 3274.100 1119.110 3274.160 ;
        RECT 1013.910 3273.960 1119.110 3274.100 ;
        RECT 1013.910 3273.900 1014.230 3273.960 ;
        RECT 1118.790 3273.900 1119.110 3273.960 ;
      LAYER via ;
        RECT 1013.940 3273.900 1014.200 3274.160 ;
        RECT 1118.820 3273.900 1119.080 3274.160 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3274.190 1014.140 3517.600 ;
        RECT 1013.940 3273.870 1014.200 3274.190 ;
        RECT 1118.820 3273.870 1119.080 3274.190 ;
        RECT 1118.880 3260.000 1119.020 3273.870 ;
        RECT 1118.770 3256.000 1119.050 3260.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 689.225 3429.325 689.395 3477.435 ;
      LAYER mcon ;
        RECT 689.225 3477.265 689.395 3477.435 ;
      LAYER met1 ;
        RECT 688.690 3491.360 689.010 3491.420 ;
        RECT 689.610 3491.360 689.930 3491.420 ;
        RECT 688.690 3491.220 689.930 3491.360 ;
        RECT 688.690 3491.160 689.010 3491.220 ;
        RECT 689.610 3491.160 689.930 3491.220 ;
        RECT 689.165 3477.420 689.455 3477.465 ;
        RECT 689.610 3477.420 689.930 3477.480 ;
        RECT 689.165 3477.280 689.930 3477.420 ;
        RECT 689.165 3477.235 689.455 3477.280 ;
        RECT 689.610 3477.220 689.930 3477.280 ;
        RECT 689.150 3429.480 689.470 3429.540 ;
        RECT 688.955 3429.340 689.470 3429.480 ;
        RECT 689.150 3429.280 689.470 3429.340 ;
        RECT 689.150 3395.140 689.470 3395.200 ;
        RECT 688.780 3395.000 689.470 3395.140 ;
        RECT 688.780 3394.860 688.920 3395.000 ;
        RECT 689.150 3394.940 689.470 3395.000 ;
        RECT 688.690 3394.600 689.010 3394.860 ;
        RECT 688.690 3367.600 689.010 3367.660 ;
        RECT 689.610 3367.600 689.930 3367.660 ;
        RECT 688.690 3367.460 689.930 3367.600 ;
        RECT 688.690 3367.400 689.010 3367.460 ;
        RECT 689.610 3367.400 689.930 3367.460 ;
        RECT 688.690 3274.100 689.010 3274.160 ;
        RECT 863.490 3274.100 863.810 3274.160 ;
        RECT 688.690 3273.960 863.810 3274.100 ;
        RECT 688.690 3273.900 689.010 3273.960 ;
        RECT 863.490 3273.900 863.810 3273.960 ;
      LAYER via ;
        RECT 688.720 3491.160 688.980 3491.420 ;
        RECT 689.640 3491.160 689.900 3491.420 ;
        RECT 689.640 3477.220 689.900 3477.480 ;
        RECT 689.180 3429.280 689.440 3429.540 ;
        RECT 689.180 3394.940 689.440 3395.200 ;
        RECT 688.720 3394.600 688.980 3394.860 ;
        RECT 688.720 3367.400 688.980 3367.660 ;
        RECT 689.640 3367.400 689.900 3367.660 ;
        RECT 688.720 3273.900 688.980 3274.160 ;
        RECT 863.520 3273.900 863.780 3274.160 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.780 3517.230 689.380 3517.370 ;
        RECT 688.780 3491.450 688.920 3517.230 ;
        RECT 688.720 3491.130 688.980 3491.450 ;
        RECT 689.640 3491.130 689.900 3491.450 ;
        RECT 689.700 3477.510 689.840 3491.130 ;
        RECT 689.640 3477.190 689.900 3477.510 ;
        RECT 689.180 3429.250 689.440 3429.570 ;
        RECT 689.240 3395.230 689.380 3429.250 ;
        RECT 689.180 3394.910 689.440 3395.230 ;
        RECT 688.720 3394.570 688.980 3394.890 ;
        RECT 688.780 3367.690 688.920 3394.570 ;
        RECT 688.720 3367.370 688.980 3367.690 ;
        RECT 689.640 3367.370 689.900 3367.690 ;
        RECT 689.700 3318.810 689.840 3367.370 ;
        RECT 688.780 3318.670 689.840 3318.810 ;
        RECT 688.780 3274.190 688.920 3318.670 ;
        RECT 688.720 3273.870 688.980 3274.190 ;
        RECT 863.520 3273.870 863.780 3274.190 ;
        RECT 863.580 3260.000 863.720 3273.870 ;
        RECT 863.470 3256.000 863.750 3260.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 362.625 3416.065 362.795 3463.835 ;
        RECT 363.545 3394.305 363.715 3415.555 ;
        RECT 364.005 3284.485 364.175 3332.595 ;
      LAYER mcon ;
        RECT 362.625 3463.665 362.795 3463.835 ;
        RECT 363.545 3415.385 363.715 3415.555 ;
        RECT 364.005 3332.425 364.175 3332.595 ;
      LAYER met1 ;
        RECT 362.565 3463.820 362.855 3463.865 ;
        RECT 363.470 3463.820 363.790 3463.880 ;
        RECT 362.565 3463.680 363.790 3463.820 ;
        RECT 362.565 3463.635 362.855 3463.680 ;
        RECT 363.470 3463.620 363.790 3463.680 ;
        RECT 362.550 3416.220 362.870 3416.280 ;
        RECT 362.355 3416.080 362.870 3416.220 ;
        RECT 362.550 3416.020 362.870 3416.080 ;
        RECT 362.550 3415.540 362.870 3415.600 ;
        RECT 363.485 3415.540 363.775 3415.585 ;
        RECT 362.550 3415.400 363.775 3415.540 ;
        RECT 362.550 3415.340 362.870 3415.400 ;
        RECT 363.485 3415.355 363.775 3415.400 ;
        RECT 363.470 3394.460 363.790 3394.520 ;
        RECT 363.275 3394.320 363.790 3394.460 ;
        RECT 363.470 3394.260 363.790 3394.320 ;
        RECT 363.470 3346.520 363.790 3346.580 ;
        RECT 364.390 3346.520 364.710 3346.580 ;
        RECT 363.470 3346.380 364.710 3346.520 ;
        RECT 363.470 3346.320 363.790 3346.380 ;
        RECT 364.390 3346.320 364.710 3346.380 ;
        RECT 363.945 3332.580 364.235 3332.625 ;
        RECT 364.390 3332.580 364.710 3332.640 ;
        RECT 363.945 3332.440 364.710 3332.580 ;
        RECT 363.945 3332.395 364.235 3332.440 ;
        RECT 364.390 3332.380 364.710 3332.440 ;
        RECT 363.930 3284.640 364.250 3284.700 ;
        RECT 363.735 3284.500 364.250 3284.640 ;
        RECT 363.930 3284.440 364.250 3284.500 ;
        RECT 363.930 3274.100 364.250 3274.160 ;
        RECT 607.730 3274.100 608.050 3274.160 ;
        RECT 363.930 3273.960 608.050 3274.100 ;
        RECT 363.930 3273.900 364.250 3273.960 ;
        RECT 607.730 3273.900 608.050 3273.960 ;
      LAYER via ;
        RECT 363.500 3463.620 363.760 3463.880 ;
        RECT 362.580 3416.020 362.840 3416.280 ;
        RECT 362.580 3415.340 362.840 3415.600 ;
        RECT 363.500 3394.260 363.760 3394.520 ;
        RECT 363.500 3346.320 363.760 3346.580 ;
        RECT 364.420 3346.320 364.680 3346.580 ;
        RECT 364.420 3332.380 364.680 3332.640 ;
        RECT 363.960 3284.440 364.220 3284.700 ;
        RECT 363.960 3273.900 364.220 3274.160 ;
        RECT 607.760 3273.900 608.020 3274.160 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3463.910 363.700 3491.390 ;
        RECT 363.500 3463.590 363.760 3463.910 ;
        RECT 362.580 3415.990 362.840 3416.310 ;
        RECT 362.640 3415.630 362.780 3415.990 ;
        RECT 362.580 3415.310 362.840 3415.630 ;
        RECT 363.500 3394.230 363.760 3394.550 ;
        RECT 363.560 3346.610 363.700 3394.230 ;
        RECT 363.500 3346.290 363.760 3346.610 ;
        RECT 364.420 3346.290 364.680 3346.610 ;
        RECT 364.480 3332.670 364.620 3346.290 ;
        RECT 364.420 3332.350 364.680 3332.670 ;
        RECT 363.960 3284.410 364.220 3284.730 ;
        RECT 364.020 3274.190 364.160 3284.410 ;
        RECT 363.960 3273.870 364.220 3274.190 ;
        RECT 607.760 3273.870 608.020 3274.190 ;
        RECT 607.820 3260.000 607.960 3273.870 ;
        RECT 607.710 3256.000 607.990 3260.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3274.100 40.410 3274.160 ;
        RECT 352.430 3274.100 352.750 3274.160 ;
        RECT 40.090 3273.960 352.750 3274.100 ;
        RECT 40.090 3273.900 40.410 3273.960 ;
        RECT 352.430 3273.900 352.750 3273.960 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3273.900 40.380 3274.160 ;
        RECT 352.460 3273.900 352.720 3274.160 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3274.190 40.320 3318.670 ;
        RECT 40.120 3273.870 40.380 3274.190 ;
        RECT 352.460 3273.870 352.720 3274.190 ;
        RECT 352.520 3260.000 352.660 3273.870 ;
        RECT 352.410 3256.000 352.690 3260.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 3084.040 18.330 3084.100 ;
        RECT 296.770 3084.040 297.090 3084.100 ;
        RECT 18.010 3083.900 297.090 3084.040 ;
        RECT 18.010 3083.840 18.330 3083.900 ;
        RECT 296.770 3083.840 297.090 3083.900 ;
      LAYER via ;
        RECT 18.040 3083.840 18.300 3084.100 ;
        RECT 296.800 3083.840 297.060 3084.100 ;
      LAYER met2 ;
        RECT 18.030 3267.555 18.310 3267.925 ;
        RECT 18.100 3084.130 18.240 3267.555 ;
        RECT 18.040 3083.810 18.300 3084.130 ;
        RECT 296.800 3083.810 297.060 3084.130 ;
        RECT 296.860 3080.925 297.000 3083.810 ;
        RECT 296.790 3080.555 297.070 3080.925 ;
      LAYER via2 ;
        RECT 18.030 3267.600 18.310 3267.880 ;
        RECT 296.790 3080.600 297.070 3080.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 18.005 3267.890 18.335 3267.905 ;
        RECT -4.800 3267.590 18.335 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 18.005 3267.575 18.335 3267.590 ;
        RECT 296.765 3080.890 297.095 3080.905 ;
        RECT 310.000 3080.890 314.000 3081.280 ;
        RECT 296.765 3080.680 314.000 3080.890 ;
        RECT 296.765 3080.590 310.500 3080.680 ;
        RECT 296.765 3080.575 297.095 3080.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2870.180 17.870 2870.240 ;
        RECT 296.770 2870.180 297.090 2870.240 ;
        RECT 17.550 2870.040 297.090 2870.180 ;
        RECT 17.550 2869.980 17.870 2870.040 ;
        RECT 296.770 2869.980 297.090 2870.040 ;
      LAYER via ;
        RECT 17.580 2869.980 17.840 2870.240 ;
        RECT 296.800 2869.980 297.060 2870.240 ;
      LAYER met2 ;
        RECT 17.570 2979.915 17.850 2980.285 ;
        RECT 17.640 2870.270 17.780 2979.915 ;
        RECT 17.580 2869.950 17.840 2870.270 ;
        RECT 296.800 2869.950 297.060 2870.270 ;
        RECT 296.860 2866.725 297.000 2869.950 ;
        RECT 296.790 2866.355 297.070 2866.725 ;
      LAYER via2 ;
        RECT 17.570 2979.960 17.850 2980.240 ;
        RECT 296.790 2866.400 297.070 2866.680 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 17.545 2980.250 17.875 2980.265 ;
        RECT -4.800 2979.950 17.875 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 17.545 2979.935 17.875 2979.950 ;
        RECT 296.765 2866.690 297.095 2866.705 ;
        RECT 310.000 2866.690 314.000 2867.080 ;
        RECT 296.765 2866.480 314.000 2866.690 ;
        RECT 296.765 2866.390 310.500 2866.480 ;
        RECT 296.765 2866.375 297.095 2866.390 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2656.320 17.410 2656.380 ;
        RECT 296.770 2656.320 297.090 2656.380 ;
        RECT 17.090 2656.180 297.090 2656.320 ;
        RECT 17.090 2656.120 17.410 2656.180 ;
        RECT 296.770 2656.120 297.090 2656.180 ;
      LAYER via ;
        RECT 17.120 2656.120 17.380 2656.380 ;
        RECT 296.800 2656.120 297.060 2656.380 ;
      LAYER met2 ;
        RECT 17.110 2692.955 17.390 2693.325 ;
        RECT 17.180 2656.410 17.320 2692.955 ;
        RECT 17.120 2656.090 17.380 2656.410 ;
        RECT 296.800 2656.090 297.060 2656.410 ;
        RECT 296.860 2652.525 297.000 2656.090 ;
        RECT 296.790 2652.155 297.070 2652.525 ;
      LAYER via2 ;
        RECT 17.110 2693.000 17.390 2693.280 ;
        RECT 296.790 2652.200 297.070 2652.480 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.085 2693.290 17.415 2693.305 ;
        RECT -4.800 2692.990 17.415 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.085 2692.975 17.415 2692.990 ;
        RECT 296.765 2652.490 297.095 2652.505 ;
        RECT 310.000 2652.490 314.000 2652.880 ;
        RECT 296.765 2652.280 314.000 2652.490 ;
        RECT 296.765 2652.190 310.500 2652.280 ;
        RECT 296.765 2652.175 297.095 2652.190 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2408.120 17.870 2408.180 ;
        RECT 296.770 2408.120 297.090 2408.180 ;
        RECT 17.550 2407.980 297.090 2408.120 ;
        RECT 17.550 2407.920 17.870 2407.980 ;
        RECT 296.770 2407.920 297.090 2407.980 ;
      LAYER via ;
        RECT 17.580 2407.920 17.840 2408.180 ;
        RECT 296.800 2407.920 297.060 2408.180 ;
      LAYER met2 ;
        RECT 296.790 2437.955 297.070 2438.325 ;
        RECT 296.860 2408.210 297.000 2437.955 ;
        RECT 17.580 2407.890 17.840 2408.210 ;
        RECT 296.800 2407.890 297.060 2408.210 ;
        RECT 17.640 2405.685 17.780 2407.890 ;
        RECT 17.570 2405.315 17.850 2405.685 ;
      LAYER via2 ;
        RECT 296.790 2438.000 297.070 2438.280 ;
        RECT 17.570 2405.360 17.850 2405.640 ;
      LAYER met3 ;
        RECT 296.765 2438.290 297.095 2438.305 ;
        RECT 310.000 2438.290 314.000 2438.680 ;
        RECT 296.765 2438.080 314.000 2438.290 ;
        RECT 296.765 2437.990 310.500 2438.080 ;
        RECT 296.765 2437.975 297.095 2437.990 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 17.545 2405.650 17.875 2405.665 ;
        RECT -4.800 2405.350 17.875 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 17.545 2405.335 17.875 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2125.240 16.490 2125.300 ;
        RECT 299.990 2125.240 300.310 2125.300 ;
        RECT 16.170 2125.100 300.310 2125.240 ;
        RECT 16.170 2125.040 16.490 2125.100 ;
        RECT 299.990 2125.040 300.310 2125.100 ;
      LAYER via ;
        RECT 16.200 2125.040 16.460 2125.300 ;
        RECT 300.020 2125.040 300.280 2125.300 ;
      LAYER met2 ;
        RECT 300.010 2223.755 300.290 2224.125 ;
        RECT 300.080 2125.330 300.220 2223.755 ;
        RECT 16.200 2125.010 16.460 2125.330 ;
        RECT 300.020 2125.010 300.280 2125.330 ;
        RECT 16.260 2118.725 16.400 2125.010 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
      LAYER via2 ;
        RECT 300.010 2223.800 300.290 2224.080 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
      LAYER met3 ;
        RECT 299.985 2224.090 300.315 2224.105 ;
        RECT 310.000 2224.090 314.000 2224.480 ;
        RECT 299.985 2223.880 314.000 2224.090 ;
        RECT 299.985 2223.790 310.500 2223.880 ;
        RECT 299.985 2223.775 300.315 2223.790 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 299.990 1835.220 300.310 1835.280 ;
        RECT 15.710 1835.080 300.310 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 299.990 1835.020 300.310 1835.080 ;
      LAYER via ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 300.020 1835.020 300.280 1835.280 ;
      LAYER met2 ;
        RECT 300.010 2009.555 300.290 2009.925 ;
        RECT 300.080 1835.310 300.220 2009.555 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 300.020 1834.990 300.280 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 300.010 2009.600 300.290 2009.880 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT 299.985 2009.890 300.315 2009.905 ;
        RECT 310.000 2009.890 314.000 2010.280 ;
        RECT 299.985 2009.680 314.000 2009.890 ;
        RECT 299.985 2009.590 310.500 2009.680 ;
        RECT 299.985 2009.575 300.315 2009.590 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 676.160 2618.710 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2618.390 676.020 2901.150 676.160 ;
        RECT 2618.390 675.960 2618.710 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2618.420 675.960 2618.680 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2618.410 826.355 2618.690 826.725 ;
        RECT 2618.480 676.250 2618.620 826.355 ;
        RECT 2618.420 675.930 2618.680 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2618.410 826.400 2618.690 826.680 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2606.000 826.690 2610.000 827.080 ;
        RECT 2618.385 826.690 2618.715 826.705 ;
        RECT 2606.000 826.480 2618.715 826.690 ;
        RECT 2609.580 826.390 2618.715 826.480 ;
        RECT 2618.385 826.375 2618.715 826.390 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 299.990 1545.540 300.310 1545.600 ;
        RECT 16.630 1545.400 300.310 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 299.990 1545.340 300.310 1545.400 ;
      LAYER via ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 300.020 1545.340 300.280 1545.600 ;
      LAYER met2 ;
        RECT 300.010 1795.355 300.290 1795.725 ;
        RECT 300.080 1545.630 300.220 1795.355 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 300.020 1545.310 300.280 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 300.010 1795.400 300.290 1795.680 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 299.985 1795.690 300.315 1795.705 ;
        RECT 310.000 1795.690 314.000 1796.080 ;
        RECT 299.985 1795.480 314.000 1795.690 ;
        RECT 299.985 1795.390 310.500 1795.480 ;
        RECT 299.985 1795.375 300.315 1795.390 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1331.680 16.030 1331.740 ;
        RECT 301.370 1331.680 301.690 1331.740 ;
        RECT 15.710 1331.540 301.690 1331.680 ;
        RECT 15.710 1331.480 16.030 1331.540 ;
        RECT 301.370 1331.480 301.690 1331.540 ;
      LAYER via ;
        RECT 15.740 1331.480 16.000 1331.740 ;
        RECT 301.400 1331.480 301.660 1331.740 ;
      LAYER met2 ;
        RECT 301.390 1580.475 301.670 1580.845 ;
        RECT 301.460 1331.770 301.600 1580.475 ;
        RECT 15.740 1331.450 16.000 1331.770 ;
        RECT 301.400 1331.450 301.660 1331.770 ;
        RECT 15.800 1328.565 15.940 1331.450 ;
        RECT 15.730 1328.195 16.010 1328.565 ;
      LAYER via2 ;
        RECT 301.390 1580.520 301.670 1580.800 ;
        RECT 15.730 1328.240 16.010 1328.520 ;
      LAYER met3 ;
        RECT 301.365 1580.810 301.695 1580.825 ;
        RECT 310.000 1580.810 314.000 1581.200 ;
        RECT 301.365 1580.600 314.000 1580.810 ;
        RECT 301.365 1580.510 310.500 1580.600 ;
        RECT 301.365 1580.495 301.695 1580.510 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 15.705 1328.530 16.035 1328.545 ;
        RECT -4.800 1328.230 16.035 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 15.705 1328.215 16.035 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 300.910 1117.820 301.230 1117.880 ;
        RECT 15.710 1117.680 301.230 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 300.910 1117.620 301.230 1117.680 ;
      LAYER via ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 300.940 1117.620 301.200 1117.880 ;
      LAYER met2 ;
        RECT 300.930 1366.275 301.210 1366.645 ;
        RECT 301.000 1117.910 301.140 1366.275 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 300.940 1117.590 301.200 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 300.930 1366.320 301.210 1366.600 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 300.905 1366.610 301.235 1366.625 ;
        RECT 310.000 1366.610 314.000 1367.000 ;
        RECT 300.905 1366.400 314.000 1366.610 ;
        RECT 300.905 1366.310 310.500 1366.400 ;
        RECT 300.905 1366.295 301.235 1366.310 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 301.830 903.960 302.150 904.020 ;
        RECT 16.170 903.820 302.150 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 301.830 903.760 302.150 903.820 ;
      LAYER via ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 301.860 903.760 302.120 904.020 ;
      LAYER met2 ;
        RECT 301.850 1152.075 302.130 1152.445 ;
        RECT 301.920 904.050 302.060 1152.075 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 301.860 903.730 302.120 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 301.850 1152.120 302.130 1152.400 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 301.825 1152.410 302.155 1152.425 ;
        RECT 310.000 1152.410 314.000 1152.800 ;
        RECT 301.825 1152.200 314.000 1152.410 ;
        RECT 301.825 1152.110 310.500 1152.200 ;
        RECT 301.825 1152.095 302.155 1152.110 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 299.990 682.960 300.310 683.020 ;
        RECT 16.170 682.820 300.310 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 299.990 682.760 300.310 682.820 ;
      LAYER via ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 300.020 682.760 300.280 683.020 ;
      LAYER met2 ;
        RECT 300.010 937.875 300.290 938.245 ;
        RECT 300.080 683.050 300.220 937.875 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 300.020 682.730 300.280 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 300.010 937.920 300.290 938.200 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 299.985 938.210 300.315 938.225 ;
        RECT 310.000 938.210 314.000 938.600 ;
        RECT 299.985 938.000 314.000 938.210 ;
        RECT 299.985 937.910 310.500 938.000 ;
        RECT 299.985 937.895 300.315 937.910 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 300.910 469.100 301.230 469.160 ;
        RECT 17.090 468.960 301.230 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 300.910 468.900 301.230 468.960 ;
      LAYER via ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 300.940 468.900 301.200 469.160 ;
      LAYER met2 ;
        RECT 300.930 723.675 301.210 724.045 ;
        RECT 301.000 469.190 301.140 723.675 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 300.940 468.870 301.200 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 300.930 723.720 301.210 724.000 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 300.905 724.010 301.235 724.025 ;
        RECT 310.000 724.010 314.000 724.400 ;
        RECT 300.905 723.800 314.000 724.010 ;
        RECT 300.905 723.710 310.500 723.800 ;
        RECT 300.905 723.695 301.235 723.710 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 301.370 255.240 301.690 255.300 ;
        RECT 17.090 255.100 301.690 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 301.370 255.040 301.690 255.100 ;
      LAYER via ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 301.400 255.040 301.660 255.300 ;
      LAYER met2 ;
        RECT 301.390 509.475 301.670 509.845 ;
        RECT 301.460 255.330 301.600 509.475 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 301.400 255.010 301.660 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 301.390 509.520 301.670 509.800 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 301.365 509.810 301.695 509.825 ;
        RECT 310.000 509.810 314.000 510.200 ;
        RECT 301.365 509.600 314.000 509.810 ;
        RECT 301.365 509.510 310.500 509.600 ;
        RECT 301.365 509.495 301.695 509.510 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 300.450 41.380 300.770 41.440 ;
        RECT 17.090 41.240 300.770 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 300.450 41.180 300.770 41.240 ;
      LAYER via ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 300.480 41.180 300.740 41.440 ;
      LAYER met2 ;
        RECT 300.470 295.275 300.750 295.645 ;
        RECT 300.540 41.470 300.680 295.275 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 300.480 41.150 300.740 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 300.470 295.320 300.750 295.600 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 300.445 295.610 300.775 295.625 ;
        RECT 310.000 295.610 314.000 296.000 ;
        RECT 300.445 295.400 314.000 295.610 ;
        RECT 300.445 295.310 310.500 295.400 ;
        RECT 300.445 295.295 300.775 295.310 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 910.760 2618.710 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2618.390 910.620 2901.150 910.760 ;
        RECT 2618.390 910.560 2618.710 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2618.420 910.560 2618.680 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2618.410 1026.275 2618.690 1026.645 ;
        RECT 2618.480 910.850 2618.620 1026.275 ;
        RECT 2618.420 910.530 2618.680 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2618.410 1026.320 2618.690 1026.600 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2606.000 1026.610 2610.000 1027.000 ;
        RECT 2618.385 1026.610 2618.715 1026.625 ;
        RECT 2606.000 1026.400 2618.715 1026.610 ;
        RECT 2609.580 1026.310 2618.715 1026.400 ;
        RECT 2618.385 1026.295 2618.715 1026.310 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1145.360 2618.710 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2618.390 1145.220 2901.150 1145.360 ;
        RECT 2618.390 1145.160 2618.710 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2618.420 1145.160 2618.680 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2618.410 1226.195 2618.690 1226.565 ;
        RECT 2618.480 1145.450 2618.620 1226.195 ;
        RECT 2618.420 1145.130 2618.680 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2618.410 1226.240 2618.690 1226.520 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2606.000 1226.530 2610.000 1226.920 ;
        RECT 2618.385 1226.530 2618.715 1226.545 ;
        RECT 2606.000 1226.320 2618.715 1226.530 ;
        RECT 2609.580 1226.230 2618.715 1226.320 ;
        RECT 2618.385 1226.215 2618.715 1226.230 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1379.960 2618.710 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2618.390 1379.820 2901.150 1379.960 ;
        RECT 2618.390 1379.760 2618.710 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 2618.420 1379.760 2618.680 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 2618.410 1426.115 2618.690 1426.485 ;
        RECT 2618.480 1380.050 2618.620 1426.115 ;
        RECT 2618.420 1379.730 2618.680 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2618.410 1426.160 2618.690 1426.440 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2606.000 1426.450 2610.000 1426.840 ;
        RECT 2618.385 1426.450 2618.715 1426.465 ;
        RECT 2606.000 1426.240 2618.715 1426.450 ;
        RECT 2609.580 1426.150 2618.715 1426.240 ;
        RECT 2618.385 1426.135 2618.715 1426.150 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1614.560 2621.930 1614.620 ;
        RECT 2900.830 1614.560 2901.150 1614.620 ;
        RECT 2621.610 1614.420 2901.150 1614.560 ;
        RECT 2621.610 1614.360 2621.930 1614.420 ;
        RECT 2900.830 1614.360 2901.150 1614.420 ;
      LAYER via ;
        RECT 2621.640 1614.360 2621.900 1614.620 ;
        RECT 2900.860 1614.360 2901.120 1614.620 ;
      LAYER met2 ;
        RECT 2621.630 1626.035 2621.910 1626.405 ;
        RECT 2621.700 1614.650 2621.840 1626.035 ;
        RECT 2621.640 1614.330 2621.900 1614.650 ;
        RECT 2900.860 1614.330 2901.120 1614.650 ;
        RECT 2900.920 1613.485 2901.060 1614.330 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2621.630 1626.080 2621.910 1626.360 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2606.000 1626.370 2610.000 1626.760 ;
        RECT 2621.605 1626.370 2621.935 1626.385 ;
        RECT 2606.000 1626.160 2621.935 1626.370 ;
        RECT 2609.580 1626.070 2621.935 1626.160 ;
        RECT 2621.605 1626.055 2621.935 1626.070 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2621.150 1842.700 2621.470 1842.760 ;
        RECT 2900.830 1842.700 2901.150 1842.760 ;
        RECT 2621.150 1842.560 2901.150 1842.700 ;
        RECT 2621.150 1842.500 2621.470 1842.560 ;
        RECT 2900.830 1842.500 2901.150 1842.560 ;
      LAYER via ;
        RECT 2621.180 1842.500 2621.440 1842.760 ;
        RECT 2900.860 1842.500 2901.120 1842.760 ;
      LAYER met2 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
        RECT 2900.920 1842.790 2901.060 1847.715 ;
        RECT 2621.180 1842.470 2621.440 1842.790 ;
        RECT 2900.860 1842.470 2901.120 1842.790 ;
        RECT 2621.240 1827.005 2621.380 1842.470 ;
        RECT 2621.170 1826.635 2621.450 1827.005 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
        RECT 2621.170 1826.680 2621.450 1826.960 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2606.000 1826.970 2610.000 1827.360 ;
        RECT 2621.145 1826.970 2621.475 1826.985 ;
        RECT 2606.000 1826.760 2621.475 1826.970 ;
        RECT 2609.580 1826.670 2621.475 1826.760 ;
        RECT 2621.145 1826.655 2621.475 1826.670 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2077.300 2618.710 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 2618.390 2077.160 2901.150 2077.300 ;
        RECT 2618.390 2077.100 2618.710 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
      LAYER via ;
        RECT 2618.420 2077.100 2618.680 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 2618.420 2077.070 2618.680 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 2618.480 2026.925 2618.620 2077.070 ;
        RECT 2618.410 2026.555 2618.690 2026.925 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
        RECT 2618.410 2026.600 2618.690 2026.880 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2606.000 2026.890 2610.000 2027.280 ;
        RECT 2618.385 2026.890 2618.715 2026.905 ;
        RECT 2606.000 2026.680 2618.715 2026.890 ;
        RECT 2609.580 2026.590 2618.715 2026.680 ;
        RECT 2618.385 2026.575 2618.715 2026.590 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2311.900 2618.710 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2618.390 2311.760 2901.150 2311.900 ;
        RECT 2618.390 2311.700 2618.710 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
      LAYER via ;
        RECT 2618.420 2311.700 2618.680 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2618.420 2311.670 2618.680 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2618.480 2226.845 2618.620 2311.670 ;
        RECT 2618.410 2226.475 2618.690 2226.845 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2618.410 2226.520 2618.690 2226.800 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2606.000 2226.810 2610.000 2227.200 ;
        RECT 2618.385 2226.810 2618.715 2226.825 ;
        RECT 2606.000 2226.600 2618.715 2226.810 ;
        RECT 2609.580 2226.510 2618.715 2226.600 ;
        RECT 2618.385 2226.495 2618.715 2226.510 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 151.540 2619.170 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2618.850 151.400 2901.150 151.540 ;
        RECT 2618.850 151.340 2619.170 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2618.880 151.340 2619.140 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2618.870 359.875 2619.150 360.245 ;
        RECT 2618.940 151.630 2619.080 359.875 ;
        RECT 2618.880 151.310 2619.140 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2618.870 359.920 2619.150 360.200 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2606.000 360.210 2610.000 360.600 ;
        RECT 2618.845 360.210 2619.175 360.225 ;
        RECT 2606.000 360.000 2619.175 360.210 ;
        RECT 2609.580 359.910 2619.175 360.000 ;
        RECT 2618.845 359.895 2619.175 359.910 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2491.080 2618.710 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 2618.390 2490.940 2901.150 2491.080 ;
        RECT 2618.390 2490.880 2618.710 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
      LAYER via ;
        RECT 2618.420 2490.880 2618.680 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 2618.420 2490.850 2618.680 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 2618.480 2360.125 2618.620 2490.850 ;
        RECT 2618.410 2359.755 2618.690 2360.125 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 2618.410 2359.800 2618.690 2360.080 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2606.000 2360.090 2610.000 2360.480 ;
        RECT 2618.385 2360.090 2618.715 2360.105 ;
        RECT 2606.000 2359.880 2618.715 2360.090 ;
        RECT 2609.580 2359.790 2618.715 2359.880 ;
        RECT 2618.385 2359.775 2618.715 2359.790 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2617.470 2725.680 2617.790 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2617.470 2725.540 2901.150 2725.680 ;
        RECT 2617.470 2725.480 2617.790 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 2617.500 2725.480 2617.760 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2617.500 2725.450 2617.760 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 2617.560 2691.170 2617.700 2725.450 ;
        RECT 2617.560 2691.030 2618.620 2691.170 ;
        RECT 2618.480 2560.045 2618.620 2691.030 ;
        RECT 2618.410 2559.675 2618.690 2560.045 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 2618.410 2559.720 2618.690 2560.000 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2606.000 2560.010 2610.000 2560.400 ;
        RECT 2618.385 2560.010 2618.715 2560.025 ;
        RECT 2606.000 2559.800 2618.715 2560.010 ;
        RECT 2609.580 2559.710 2618.715 2559.800 ;
        RECT 2618.385 2559.695 2618.715 2559.710 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2960.280 2618.710 2960.340 ;
        RECT 2898.990 2960.280 2899.310 2960.340 ;
        RECT 2618.390 2960.140 2899.310 2960.280 ;
        RECT 2618.390 2960.080 2618.710 2960.140 ;
        RECT 2898.990 2960.080 2899.310 2960.140 ;
      LAYER via ;
        RECT 2618.420 2960.080 2618.680 2960.340 ;
        RECT 2899.020 2960.080 2899.280 2960.340 ;
      LAYER met2 ;
        RECT 2899.010 2962.235 2899.290 2962.605 ;
        RECT 2899.080 2960.370 2899.220 2962.235 ;
        RECT 2618.420 2960.050 2618.680 2960.370 ;
        RECT 2899.020 2960.050 2899.280 2960.370 ;
        RECT 2618.480 2759.965 2618.620 2960.050 ;
        RECT 2618.410 2759.595 2618.690 2759.965 ;
      LAYER via2 ;
        RECT 2899.010 2962.280 2899.290 2962.560 ;
        RECT 2618.410 2759.640 2618.690 2759.920 ;
      LAYER met3 ;
        RECT 2898.985 2962.570 2899.315 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2898.985 2962.270 2924.800 2962.570 ;
        RECT 2898.985 2962.255 2899.315 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2606.000 2759.930 2610.000 2760.320 ;
        RECT 2618.385 2759.930 2618.715 2759.945 ;
        RECT 2606.000 2759.720 2618.715 2759.930 ;
        RECT 2609.580 2759.630 2618.715 2759.720 ;
        RECT 2618.385 2759.615 2618.715 2759.630 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3194.880 2619.170 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2618.850 3194.740 2901.150 3194.880 ;
        RECT 2618.850 3194.680 2619.170 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 2618.880 3194.680 2619.140 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2618.880 3194.650 2619.140 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 2618.940 2959.885 2619.080 3194.650 ;
        RECT 2618.870 2959.515 2619.150 2959.885 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 2618.870 2959.560 2619.150 2959.840 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2606.000 2959.850 2610.000 2960.240 ;
        RECT 2618.845 2959.850 2619.175 2959.865 ;
        RECT 2606.000 2959.640 2619.175 2959.850 ;
        RECT 2609.580 2959.550 2619.175 2959.640 ;
        RECT 2618.845 2959.535 2619.175 2959.550 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 3429.480 2618.710 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2618.390 3429.340 2901.150 3429.480 ;
        RECT 2618.390 3429.280 2618.710 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 2618.420 3429.280 2618.680 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 2618.420 3429.250 2618.680 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 2618.480 3159.805 2618.620 3429.250 ;
        RECT 2618.410 3159.435 2618.690 3159.805 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 2618.410 3159.480 2618.690 3159.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2606.000 3159.770 2610.000 3160.160 ;
        RECT 2618.385 3159.770 2618.715 3159.785 ;
        RECT 2606.000 3159.560 2618.715 3159.770 ;
        RECT 2609.580 3159.470 2618.715 3159.560 ;
        RECT 2618.385 3159.455 2618.715 3159.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2483.610 3501.900 2483.930 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 2483.610 3501.760 2717.610 3501.900 ;
        RECT 2483.610 3501.700 2483.930 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 2483.640 3501.700 2483.900 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 2483.640 3501.670 2483.900 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 2481.750 3259.650 2482.030 3260.000 ;
        RECT 2483.700 3259.650 2483.840 3501.670 ;
        RECT 2481.750 3259.510 2483.840 3259.650 ;
        RECT 2481.750 3256.000 2482.030 3259.510 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2228.310 3501.900 2228.630 3501.960 ;
        RECT 2392.530 3501.900 2392.850 3501.960 ;
        RECT 2228.310 3501.760 2392.850 3501.900 ;
        RECT 2228.310 3501.700 2228.630 3501.760 ;
        RECT 2392.530 3501.700 2392.850 3501.760 ;
      LAYER via ;
        RECT 2228.340 3501.700 2228.600 3501.960 ;
        RECT 2392.560 3501.700 2392.820 3501.960 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.990 2392.760 3517.600 ;
        RECT 2228.340 3501.670 2228.600 3501.990 ;
        RECT 2392.560 3501.670 2392.820 3501.990 ;
        RECT 2226.450 3259.650 2226.730 3260.000 ;
        RECT 2228.400 3259.650 2228.540 3501.670 ;
        RECT 2226.450 3259.510 2228.540 3259.650 ;
        RECT 2226.450 3256.000 2226.730 3259.510 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 3501.900 1973.330 3501.960 ;
        RECT 2068.230 3501.900 2068.550 3501.960 ;
        RECT 1973.010 3501.760 2068.550 3501.900 ;
        RECT 1973.010 3501.700 1973.330 3501.760 ;
        RECT 2068.230 3501.700 2068.550 3501.760 ;
      LAYER via ;
        RECT 1973.040 3501.700 1973.300 3501.960 ;
        RECT 2068.260 3501.700 2068.520 3501.960 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.990 2068.460 3517.600 ;
        RECT 1973.040 3501.670 1973.300 3501.990 ;
        RECT 2068.260 3501.670 2068.520 3501.990 ;
        RECT 1970.690 3258.970 1970.970 3260.000 ;
        RECT 1973.100 3258.970 1973.240 3501.670 ;
        RECT 1970.690 3258.830 1973.240 3258.970 ;
        RECT 1970.690 3256.000 1970.970 3258.830 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1717.710 3501.560 1718.030 3501.620 ;
        RECT 1743.930 3501.560 1744.250 3501.620 ;
        RECT 1717.710 3501.420 1744.250 3501.560 ;
        RECT 1717.710 3501.360 1718.030 3501.420 ;
        RECT 1743.930 3501.360 1744.250 3501.420 ;
      LAYER via ;
        RECT 1717.740 3501.360 1718.000 3501.620 ;
        RECT 1743.960 3501.360 1744.220 3501.620 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3501.650 1744.160 3517.600 ;
        RECT 1717.740 3501.330 1718.000 3501.650 ;
        RECT 1743.960 3501.330 1744.220 3501.650 ;
        RECT 1714.930 3258.970 1715.210 3260.000 ;
        RECT 1717.800 3258.970 1717.940 3501.330 ;
        RECT 1714.930 3258.830 1717.940 3258.970 ;
        RECT 1714.930 3256.000 1715.210 3258.830 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1420.165 3381.045 1420.335 3429.155 ;
      LAYER mcon ;
        RECT 1420.165 3428.985 1420.335 3429.155 ;
      LAYER met1 ;
        RECT 1419.170 3477.760 1419.490 3477.820 ;
        RECT 1419.630 3477.760 1419.950 3477.820 ;
        RECT 1419.170 3477.620 1419.950 3477.760 ;
        RECT 1419.170 3477.560 1419.490 3477.620 ;
        RECT 1419.630 3477.560 1419.950 3477.620 ;
        RECT 1419.630 3443.080 1419.950 3443.140 ;
        RECT 1420.550 3443.080 1420.870 3443.140 ;
        RECT 1419.630 3442.940 1420.870 3443.080 ;
        RECT 1419.630 3442.880 1419.950 3442.940 ;
        RECT 1420.550 3442.880 1420.870 3442.940 ;
        RECT 1420.105 3429.140 1420.395 3429.185 ;
        RECT 1420.550 3429.140 1420.870 3429.200 ;
        RECT 1420.105 3429.000 1420.870 3429.140 ;
        RECT 1420.105 3428.955 1420.395 3429.000 ;
        RECT 1420.550 3428.940 1420.870 3429.000 ;
        RECT 1420.090 3381.200 1420.410 3381.260 ;
        RECT 1419.895 3381.060 1420.410 3381.200 ;
        RECT 1420.090 3381.000 1420.410 3381.060 ;
        RECT 1420.090 3367.600 1420.410 3367.660 ;
        RECT 1421.010 3367.600 1421.330 3367.660 ;
        RECT 1420.090 3367.460 1421.330 3367.600 ;
        RECT 1420.090 3367.400 1420.410 3367.460 ;
        RECT 1421.010 3367.400 1421.330 3367.460 ;
        RECT 1420.090 3274.100 1420.410 3274.160 ;
        RECT 1459.650 3274.100 1459.970 3274.160 ;
        RECT 1420.090 3273.960 1459.970 3274.100 ;
        RECT 1420.090 3273.900 1420.410 3273.960 ;
        RECT 1459.650 3273.900 1459.970 3273.960 ;
      LAYER via ;
        RECT 1419.200 3477.560 1419.460 3477.820 ;
        RECT 1419.660 3477.560 1419.920 3477.820 ;
        RECT 1419.660 3442.880 1419.920 3443.140 ;
        RECT 1420.580 3442.880 1420.840 3443.140 ;
        RECT 1420.580 3428.940 1420.840 3429.200 ;
        RECT 1420.120 3381.000 1420.380 3381.260 ;
        RECT 1420.120 3367.400 1420.380 3367.660 ;
        RECT 1421.040 3367.400 1421.300 3367.660 ;
        RECT 1420.120 3273.900 1420.380 3274.160 ;
        RECT 1459.680 3273.900 1459.940 3274.160 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3477.850 1419.400 3517.600 ;
        RECT 1419.200 3477.530 1419.460 3477.850 ;
        RECT 1419.660 3477.530 1419.920 3477.850 ;
        RECT 1419.720 3443.170 1419.860 3477.530 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3274.190 1420.320 3318.670 ;
        RECT 1420.120 3273.870 1420.380 3274.190 ;
        RECT 1459.680 3273.870 1459.940 3274.190 ;
        RECT 1459.740 3260.000 1459.880 3273.870 ;
        RECT 1459.630 3256.000 1459.910 3260.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 386.140 2619.170 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2618.850 386.000 2901.150 386.140 ;
        RECT 2618.850 385.940 2619.170 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2618.880 385.940 2619.140 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2618.870 559.795 2619.150 560.165 ;
        RECT 2618.940 386.230 2619.080 559.795 ;
        RECT 2618.880 385.910 2619.140 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2618.870 559.840 2619.150 560.120 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 2606.000 560.130 2610.000 560.520 ;
        RECT 2618.845 560.130 2619.175 560.145 ;
        RECT 2606.000 559.920 2619.175 560.130 ;
        RECT 2609.580 559.830 2619.175 559.920 ;
        RECT 2618.845 559.815 2619.175 559.830 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1095.405 3284.485 1095.575 3332.595 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1095.405 3332.425 1095.575 3332.595 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1095.330 3395.140 1095.650 3395.200 ;
        RECT 1094.960 3395.000 1095.650 3395.140 ;
        RECT 1094.960 3394.860 1095.100 3395.000 ;
        RECT 1095.330 3394.940 1095.650 3395.000 ;
        RECT 1094.870 3394.600 1095.190 3394.860 ;
        RECT 1094.870 3346.520 1095.190 3346.580 ;
        RECT 1095.790 3346.520 1096.110 3346.580 ;
        RECT 1094.870 3346.380 1096.110 3346.520 ;
        RECT 1094.870 3346.320 1095.190 3346.380 ;
        RECT 1095.790 3346.320 1096.110 3346.380 ;
        RECT 1095.345 3332.580 1095.635 3332.625 ;
        RECT 1095.790 3332.580 1096.110 3332.640 ;
        RECT 1095.345 3332.440 1096.110 3332.580 ;
        RECT 1095.345 3332.395 1095.635 3332.440 ;
        RECT 1095.790 3332.380 1096.110 3332.440 ;
        RECT 1095.330 3284.640 1095.650 3284.700 ;
        RECT 1095.135 3284.500 1095.650 3284.640 ;
        RECT 1095.330 3284.440 1095.650 3284.500 ;
        RECT 1095.330 3274.440 1095.650 3274.500 ;
        RECT 1203.890 3274.440 1204.210 3274.500 ;
        RECT 1095.330 3274.300 1204.210 3274.440 ;
        RECT 1095.330 3274.240 1095.650 3274.300 ;
        RECT 1203.890 3274.240 1204.210 3274.300 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1095.360 3394.940 1095.620 3395.200 ;
        RECT 1094.900 3394.600 1095.160 3394.860 ;
        RECT 1094.900 3346.320 1095.160 3346.580 ;
        RECT 1095.820 3346.320 1096.080 3346.580 ;
        RECT 1095.820 3332.380 1096.080 3332.640 ;
        RECT 1095.360 3284.440 1095.620 3284.700 ;
        RECT 1095.360 3274.240 1095.620 3274.500 ;
        RECT 1203.920 3274.240 1204.180 3274.500 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3395.230 1095.560 3429.250 ;
        RECT 1095.360 3394.910 1095.620 3395.230 ;
        RECT 1094.900 3394.570 1095.160 3394.890 ;
        RECT 1094.960 3346.610 1095.100 3394.570 ;
        RECT 1094.900 3346.290 1095.160 3346.610 ;
        RECT 1095.820 3346.290 1096.080 3346.610 ;
        RECT 1095.880 3332.670 1096.020 3346.290 ;
        RECT 1095.820 3332.350 1096.080 3332.670 ;
        RECT 1095.360 3284.410 1095.620 3284.730 ;
        RECT 1095.420 3274.530 1095.560 3284.410 ;
        RECT 1095.360 3274.210 1095.620 3274.530 ;
        RECT 1203.920 3274.210 1204.180 3274.530 ;
        RECT 1203.980 3260.000 1204.120 3274.210 ;
        RECT 1203.870 3256.000 1204.150 3260.000 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3275.120 771.810 3275.180 ;
        RECT 948.590 3275.120 948.910 3275.180 ;
        RECT 771.490 3274.980 948.910 3275.120 ;
        RECT 771.490 3274.920 771.810 3274.980 ;
        RECT 948.590 3274.920 948.910 3274.980 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3274.920 771.780 3275.180 ;
        RECT 948.620 3274.920 948.880 3275.180 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3275.210 771.720 3318.670 ;
        RECT 771.520 3274.890 771.780 3275.210 ;
        RECT 948.620 3274.890 948.880 3275.210 ;
        RECT 948.680 3260.000 948.820 3274.890 ;
        RECT 948.570 3256.000 948.850 3260.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 3274.440 448.430 3274.500 ;
        RECT 692.830 3274.440 693.150 3274.500 ;
        RECT 448.110 3274.300 693.150 3274.440 ;
        RECT 448.110 3274.240 448.430 3274.300 ;
        RECT 692.830 3274.240 693.150 3274.300 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 3274.240 448.400 3274.500 ;
        RECT 692.860 3274.240 693.120 3274.500 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 3274.530 448.340 3498.270 ;
        RECT 448.140 3274.210 448.400 3274.530 ;
        RECT 692.860 3274.210 693.120 3274.530 ;
        RECT 692.920 3260.000 693.060 3274.210 ;
        RECT 692.810 3256.000 693.090 3260.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 3274.440 124.130 3274.500 ;
        RECT 437.530 3274.440 437.850 3274.500 ;
        RECT 123.810 3274.300 437.850 3274.440 ;
        RECT 123.810 3274.240 124.130 3274.300 ;
        RECT 437.530 3274.240 437.850 3274.300 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 3274.240 124.100 3274.500 ;
        RECT 437.560 3274.240 437.820 3274.500 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 3274.530 124.040 3498.270 ;
        RECT 123.840 3274.210 124.100 3274.530 ;
        RECT 437.560 3274.210 437.820 3274.530 ;
        RECT 437.620 3260.000 437.760 3274.210 ;
        RECT 437.510 3256.000 437.790 3260.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3153.060 17.410 3153.120 ;
        RECT 296.770 3153.060 297.090 3153.120 ;
        RECT 17.090 3152.920 297.090 3153.060 ;
        RECT 17.090 3152.860 17.410 3152.920 ;
        RECT 296.770 3152.860 297.090 3152.920 ;
      LAYER via ;
        RECT 17.120 3152.860 17.380 3153.120 ;
        RECT 296.800 3152.860 297.060 3153.120 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 3153.150 17.320 3339.635 ;
        RECT 17.120 3152.830 17.380 3153.150 ;
        RECT 296.800 3152.830 297.060 3153.150 ;
        RECT 296.860 3152.325 297.000 3152.830 ;
        RECT 296.790 3151.955 297.070 3152.325 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 296.790 3152.000 297.070 3152.280 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 296.765 3152.290 297.095 3152.305 ;
        RECT 310.000 3152.290 314.000 3152.680 ;
        RECT 296.765 3152.080 314.000 3152.290 ;
        RECT 296.765 3151.990 310.500 3152.080 ;
        RECT 296.765 3151.975 297.095 3151.990 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2939.200 17.410 2939.260 ;
        RECT 296.770 2939.200 297.090 2939.260 ;
        RECT 17.090 2939.060 297.090 2939.200 ;
        RECT 17.090 2939.000 17.410 2939.060 ;
        RECT 296.770 2939.000 297.090 2939.060 ;
      LAYER via ;
        RECT 17.120 2939.000 17.380 2939.260 ;
        RECT 296.800 2939.000 297.060 2939.260 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 2939.290 17.320 3051.995 ;
        RECT 17.120 2938.970 17.380 2939.290 ;
        RECT 296.800 2938.970 297.060 2939.290 ;
        RECT 296.860 2938.125 297.000 2938.970 ;
        RECT 296.790 2937.755 297.070 2938.125 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 296.790 2937.800 297.070 2938.080 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 296.765 2938.090 297.095 2938.105 ;
        RECT 310.000 2938.090 314.000 2938.480 ;
        RECT 296.765 2937.880 314.000 2938.090 ;
        RECT 296.765 2937.790 310.500 2937.880 ;
        RECT 296.765 2937.775 297.095 2937.790 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2725.340 17.410 2725.400 ;
        RECT 296.770 2725.340 297.090 2725.400 ;
        RECT 17.090 2725.200 297.090 2725.340 ;
        RECT 17.090 2725.140 17.410 2725.200 ;
        RECT 296.770 2725.140 297.090 2725.200 ;
      LAYER via ;
        RECT 17.120 2725.140 17.380 2725.400 ;
        RECT 296.800 2725.140 297.060 2725.400 ;
      LAYER met2 ;
        RECT 17.110 2765.035 17.390 2765.405 ;
        RECT 17.180 2725.430 17.320 2765.035 ;
        RECT 17.120 2725.110 17.380 2725.430 ;
        RECT 296.800 2725.110 297.060 2725.430 ;
        RECT 296.860 2723.925 297.000 2725.110 ;
        RECT 296.790 2723.555 297.070 2723.925 ;
      LAYER via2 ;
        RECT 17.110 2765.080 17.390 2765.360 ;
        RECT 296.790 2723.600 297.070 2723.880 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 17.085 2765.370 17.415 2765.385 ;
        RECT -4.800 2765.070 17.415 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 17.085 2765.055 17.415 2765.070 ;
        RECT 296.765 2723.890 297.095 2723.905 ;
        RECT 310.000 2723.890 314.000 2724.280 ;
        RECT 296.765 2723.680 314.000 2723.890 ;
        RECT 296.765 2723.590 310.500 2723.680 ;
        RECT 296.765 2723.575 297.095 2723.590 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2483.940 17.410 2484.000 ;
        RECT 299.990 2483.940 300.310 2484.000 ;
        RECT 17.090 2483.800 300.310 2483.940 ;
        RECT 17.090 2483.740 17.410 2483.800 ;
        RECT 299.990 2483.740 300.310 2483.800 ;
      LAYER via ;
        RECT 17.120 2483.740 17.380 2484.000 ;
        RECT 300.020 2483.740 300.280 2484.000 ;
      LAYER met2 ;
        RECT 300.010 2509.355 300.290 2509.725 ;
        RECT 300.080 2484.030 300.220 2509.355 ;
        RECT 17.120 2483.710 17.380 2484.030 ;
        RECT 300.020 2483.710 300.280 2484.030 ;
        RECT 17.180 2477.765 17.320 2483.710 ;
        RECT 17.110 2477.395 17.390 2477.765 ;
      LAYER via2 ;
        RECT 300.010 2509.400 300.290 2509.680 ;
        RECT 17.110 2477.440 17.390 2477.720 ;
      LAYER met3 ;
        RECT 299.985 2509.690 300.315 2509.705 ;
        RECT 310.000 2509.690 314.000 2510.080 ;
        RECT 299.985 2509.480 314.000 2509.690 ;
        RECT 299.985 2509.390 310.500 2509.480 ;
        RECT 299.985 2509.375 300.315 2509.390 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.085 2477.730 17.415 2477.745 ;
        RECT -4.800 2477.430 17.415 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.085 2477.415 17.415 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2194.260 16.030 2194.320 ;
        RECT 300.450 2194.260 300.770 2194.320 ;
        RECT 15.710 2194.120 300.770 2194.260 ;
        RECT 15.710 2194.060 16.030 2194.120 ;
        RECT 300.450 2194.060 300.770 2194.120 ;
      LAYER via ;
        RECT 15.740 2194.060 16.000 2194.320 ;
        RECT 300.480 2194.060 300.740 2194.320 ;
      LAYER met2 ;
        RECT 300.470 2295.155 300.750 2295.525 ;
        RECT 300.540 2194.350 300.680 2295.155 ;
        RECT 15.740 2194.030 16.000 2194.350 ;
        RECT 300.480 2194.030 300.740 2194.350 ;
        RECT 15.800 2190.125 15.940 2194.030 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
      LAYER via2 ;
        RECT 300.470 2295.200 300.750 2295.480 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
      LAYER met3 ;
        RECT 300.445 2295.490 300.775 2295.505 ;
        RECT 310.000 2295.490 314.000 2295.880 ;
        RECT 300.445 2295.280 314.000 2295.490 ;
        RECT 300.445 2295.190 310.500 2295.280 ;
        RECT 300.445 2295.175 300.775 2295.190 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.800 2189.790 16.035 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1904.240 16.490 1904.300 ;
        RECT 300.910 1904.240 301.230 1904.300 ;
        RECT 16.170 1904.100 301.230 1904.240 ;
        RECT 16.170 1904.040 16.490 1904.100 ;
        RECT 300.910 1904.040 301.230 1904.100 ;
      LAYER via ;
        RECT 16.200 1904.040 16.460 1904.300 ;
        RECT 300.940 1904.040 301.200 1904.300 ;
      LAYER met2 ;
        RECT 300.930 2080.955 301.210 2081.325 ;
        RECT 301.000 1904.330 301.140 2080.955 ;
        RECT 16.200 1904.010 16.460 1904.330 ;
        RECT 300.940 1904.010 301.200 1904.330 ;
        RECT 16.260 1903.165 16.400 1904.010 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
      LAYER via2 ;
        RECT 300.930 2081.000 301.210 2081.280 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT 300.905 2081.290 301.235 2081.305 ;
        RECT 310.000 2081.290 314.000 2081.680 ;
        RECT 300.905 2081.080 314.000 2081.290 ;
        RECT 300.905 2080.990 310.500 2081.080 ;
        RECT 300.905 2080.975 301.235 2080.990 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 620.740 2619.170 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2618.850 620.600 2901.150 620.740 ;
        RECT 2618.850 620.540 2619.170 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2618.880 620.540 2619.140 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2618.870 759.715 2619.150 760.085 ;
        RECT 2618.940 620.830 2619.080 759.715 ;
        RECT 2618.880 620.510 2619.140 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2618.870 759.760 2619.150 760.040 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2606.000 760.050 2610.000 760.440 ;
        RECT 2618.845 760.050 2619.175 760.065 ;
        RECT 2606.000 759.840 2619.175 760.050 ;
        RECT 2609.580 759.750 2619.175 759.840 ;
        RECT 2618.845 759.735 2619.175 759.750 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 300.910 1621.360 301.230 1621.420 ;
        RECT 16.170 1621.220 301.230 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 300.910 1621.160 301.230 1621.220 ;
      LAYER via ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 300.940 1621.160 301.200 1621.420 ;
      LAYER met2 ;
        RECT 300.930 1866.755 301.210 1867.125 ;
        RECT 301.000 1621.450 301.140 1866.755 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 300.940 1621.130 301.200 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 300.930 1866.800 301.210 1867.080 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT 300.905 1867.090 301.235 1867.105 ;
        RECT 310.000 1867.090 314.000 1867.480 ;
        RECT 300.905 1866.880 314.000 1867.090 ;
        RECT 300.905 1866.790 310.500 1866.880 ;
        RECT 300.905 1866.775 301.235 1866.790 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 300.450 1400.700 300.770 1400.760 ;
        RECT 17.090 1400.560 300.770 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 300.450 1400.500 300.770 1400.560 ;
      LAYER via ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 300.480 1400.500 300.740 1400.760 ;
      LAYER met2 ;
        RECT 300.470 1651.875 300.750 1652.245 ;
        RECT 300.540 1400.790 300.680 1651.875 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 300.480 1400.470 300.740 1400.790 ;
      LAYER via2 ;
        RECT 300.470 1651.920 300.750 1652.200 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 300.445 1652.210 300.775 1652.225 ;
        RECT 310.000 1652.210 314.000 1652.600 ;
        RECT 300.445 1652.000 314.000 1652.210 ;
        RECT 300.445 1651.910 310.500 1652.000 ;
        RECT 300.445 1651.895 300.775 1651.910 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 299.990 1186.840 300.310 1186.900 ;
        RECT 17.090 1186.700 300.310 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 299.990 1186.640 300.310 1186.700 ;
      LAYER via ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 300.020 1186.640 300.280 1186.900 ;
      LAYER met2 ;
        RECT 300.010 1437.675 300.290 1438.045 ;
        RECT 300.080 1186.930 300.220 1437.675 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 300.020 1186.610 300.280 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 300.010 1437.720 300.290 1438.000 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT 299.985 1438.010 300.315 1438.025 ;
        RECT 310.000 1438.010 314.000 1438.400 ;
        RECT 299.985 1437.800 314.000 1438.010 ;
        RECT 299.985 1437.710 310.500 1437.800 ;
        RECT 299.985 1437.695 300.315 1437.710 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 301.370 972.640 301.690 972.700 ;
        RECT 15.710 972.500 301.690 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 301.370 972.440 301.690 972.500 ;
      LAYER via ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 301.400 972.440 301.660 972.700 ;
      LAYER met2 ;
        RECT 301.390 1223.475 301.670 1223.845 ;
        RECT 301.460 972.730 301.600 1223.475 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 301.400 972.410 301.660 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 301.390 1223.520 301.670 1223.800 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT 301.365 1223.810 301.695 1223.825 ;
        RECT 310.000 1223.810 314.000 1224.200 ;
        RECT 301.365 1223.600 314.000 1223.810 ;
        RECT 301.365 1223.510 310.500 1223.600 ;
        RECT 301.365 1223.495 301.695 1223.510 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 300.450 758.780 300.770 758.840 ;
        RECT 15.710 758.640 300.770 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 300.450 758.580 300.770 758.640 ;
      LAYER via ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 300.480 758.580 300.740 758.840 ;
      LAYER met2 ;
        RECT 300.470 1009.275 300.750 1009.645 ;
        RECT 300.540 758.870 300.680 1009.275 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 300.480 758.550 300.740 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 300.470 1009.320 300.750 1009.600 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 300.445 1009.610 300.775 1009.625 ;
        RECT 310.000 1009.610 314.000 1010.000 ;
        RECT 300.445 1009.400 314.000 1009.610 ;
        RECT 300.445 1009.310 310.500 1009.400 ;
        RECT 300.445 1009.295 300.775 1009.310 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 301.370 544.920 301.690 544.980 ;
        RECT 16.170 544.780 301.690 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 301.370 544.720 301.690 544.780 ;
      LAYER via ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 301.400 544.720 301.660 544.980 ;
      LAYER met2 ;
        RECT 301.390 795.075 301.670 795.445 ;
        RECT 301.460 545.010 301.600 795.075 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 301.400 544.690 301.660 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 301.390 795.120 301.670 795.400 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 301.365 795.410 301.695 795.425 ;
        RECT 310.000 795.410 314.000 795.800 ;
        RECT 301.365 795.200 314.000 795.410 ;
        RECT 301.365 795.110 310.500 795.200 ;
        RECT 301.365 795.095 301.695 795.110 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 300.450 324.260 300.770 324.320 ;
        RECT 16.630 324.120 300.770 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 300.450 324.060 300.770 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 300.480 324.060 300.740 324.320 ;
      LAYER met2 ;
        RECT 300.470 580.875 300.750 581.245 ;
        RECT 300.540 324.350 300.680 580.875 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 300.480 324.030 300.740 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 300.470 580.920 300.750 581.200 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 300.445 581.210 300.775 581.225 ;
        RECT 310.000 581.210 314.000 581.600 ;
        RECT 300.445 581.000 314.000 581.210 ;
        RECT 300.445 580.910 310.500 581.000 ;
        RECT 300.445 580.895 300.775 580.910 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 299.990 110.400 300.310 110.460 ;
        RECT 15.710 110.260 300.310 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 299.990 110.200 300.310 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 300.020 110.200 300.280 110.460 ;
      LAYER met2 ;
        RECT 300.010 366.675 300.290 367.045 ;
        RECT 300.080 110.490 300.220 366.675 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 300.020 110.170 300.280 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 300.010 366.720 300.290 367.000 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 299.985 367.010 300.315 367.025 ;
        RECT 310.000 367.010 314.000 367.400 ;
        RECT 299.985 366.800 314.000 367.010 ;
        RECT 299.985 366.710 310.500 366.800 ;
        RECT 299.985 366.695 300.315 366.710 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 855.340 2619.170 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2618.850 855.200 2901.150 855.340 ;
        RECT 2618.850 855.140 2619.170 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2618.880 855.140 2619.140 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2618.870 959.635 2619.150 960.005 ;
        RECT 2618.940 855.430 2619.080 959.635 ;
        RECT 2618.880 855.110 2619.140 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2618.870 959.680 2619.150 959.960 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2606.000 959.970 2610.000 960.360 ;
        RECT 2618.845 959.970 2619.175 959.985 ;
        RECT 2606.000 959.760 2619.175 959.970 ;
        RECT 2609.580 959.670 2619.175 959.760 ;
        RECT 2618.845 959.655 2619.175 959.670 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1089.940 2619.170 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2618.850 1089.800 2901.150 1089.940 ;
        RECT 2618.850 1089.740 2619.170 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2618.880 1089.740 2619.140 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2618.870 1159.555 2619.150 1159.925 ;
        RECT 2618.940 1090.030 2619.080 1159.555 ;
        RECT 2618.880 1089.710 2619.140 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2618.870 1159.600 2619.150 1159.880 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2606.000 1159.890 2610.000 1160.280 ;
        RECT 2618.845 1159.890 2619.175 1159.905 ;
        RECT 2606.000 1159.680 2619.175 1159.890 ;
        RECT 2609.580 1159.590 2619.175 1159.680 ;
        RECT 2618.845 1159.575 2619.175 1159.590 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1324.540 2618.710 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2618.390 1324.400 2901.150 1324.540 ;
        RECT 2618.390 1324.340 2618.710 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 2618.420 1324.340 2618.680 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 2618.410 1359.475 2618.690 1359.845 ;
        RECT 2618.480 1324.630 2618.620 1359.475 ;
        RECT 2618.420 1324.310 2618.680 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2618.410 1359.520 2618.690 1359.800 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2606.000 1359.810 2610.000 1360.200 ;
        RECT 2618.385 1359.810 2618.715 1359.825 ;
        RECT 2606.000 1359.600 2618.715 1359.810 ;
        RECT 2609.580 1359.510 2618.715 1359.600 ;
        RECT 2618.385 1359.495 2618.715 1359.510 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1559.140 2621.930 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2621.610 1559.000 2901.150 1559.140 ;
        RECT 2621.610 1558.940 2621.930 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 2621.640 1558.940 2621.900 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 2621.630 1559.395 2621.910 1559.765 ;
        RECT 2621.700 1559.230 2621.840 1559.395 ;
        RECT 2621.640 1558.910 2621.900 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2621.630 1559.440 2621.910 1559.720 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2606.000 1559.730 2610.000 1560.120 ;
        RECT 2621.605 1559.730 2621.935 1559.745 ;
        RECT 2606.000 1559.520 2621.935 1559.730 ;
        RECT 2609.580 1559.430 2621.935 1559.520 ;
        RECT 2621.605 1559.415 2621.935 1559.430 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1787.280 2618.710 1787.340 ;
        RECT 2900.830 1787.280 2901.150 1787.340 ;
        RECT 2618.390 1787.140 2901.150 1787.280 ;
        RECT 2618.390 1787.080 2618.710 1787.140 ;
        RECT 2900.830 1787.080 2901.150 1787.140 ;
      LAYER via ;
        RECT 2618.420 1787.080 2618.680 1787.340 ;
        RECT 2900.860 1787.080 2901.120 1787.340 ;
      LAYER met2 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
        RECT 2900.920 1787.370 2901.060 1789.235 ;
        RECT 2618.420 1787.050 2618.680 1787.370 ;
        RECT 2900.860 1787.050 2901.120 1787.370 ;
        RECT 2618.480 1759.685 2618.620 1787.050 ;
        RECT 2618.410 1759.315 2618.690 1759.685 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
        RECT 2618.410 1759.360 2618.690 1759.640 ;
      LAYER met3 ;
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2606.000 1759.650 2610.000 1760.040 ;
        RECT 2618.385 1759.650 2618.715 1759.665 ;
        RECT 2606.000 1759.440 2618.715 1759.650 ;
        RECT 2609.580 1759.350 2618.715 1759.440 ;
        RECT 2618.385 1759.335 2618.715 1759.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2021.880 2619.170 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 2618.850 2021.740 2901.150 2021.880 ;
        RECT 2618.850 2021.680 2619.170 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 2618.880 2021.680 2619.140 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 2618.880 2021.650 2619.140 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 2618.940 1960.285 2619.080 2021.650 ;
        RECT 2618.870 1959.915 2619.150 1960.285 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
        RECT 2618.870 1959.960 2619.150 1960.240 ;
      LAYER met3 ;
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2606.000 1960.250 2610.000 1960.640 ;
        RECT 2618.845 1960.250 2619.175 1960.265 ;
        RECT 2606.000 1960.040 2619.175 1960.250 ;
        RECT 2609.580 1959.950 2619.175 1960.040 ;
        RECT 2618.845 1959.935 2619.175 1959.950 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2256.480 2619.170 2256.540 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 2618.850 2256.340 2901.150 2256.480 ;
        RECT 2618.850 2256.280 2619.170 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
      LAYER via ;
        RECT 2618.880 2256.280 2619.140 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 2618.880 2256.250 2619.140 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 2618.940 2160.205 2619.080 2256.250 ;
        RECT 2618.870 2159.835 2619.150 2160.205 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
        RECT 2618.870 2159.880 2619.150 2160.160 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2606.000 2160.170 2610.000 2160.560 ;
        RECT 2618.845 2160.170 2619.175 2160.185 ;
        RECT 2606.000 2159.960 2619.175 2160.170 ;
        RECT 2609.580 2159.870 2619.175 2159.960 ;
        RECT 2618.845 2159.855 2619.175 2159.870 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 324.370 243.680 324.690 243.740 ;
        RECT 330.810 243.680 331.130 243.740 ;
        RECT 324.370 243.540 331.130 243.680 ;
        RECT 324.370 243.480 324.690 243.540 ;
        RECT 330.810 243.480 331.130 243.540 ;
        RECT 330.810 24.040 331.130 24.100 ;
        RECT 633.030 24.040 633.350 24.100 ;
        RECT 330.810 23.900 633.350 24.040 ;
        RECT 330.810 23.840 331.130 23.900 ;
        RECT 633.030 23.840 633.350 23.900 ;
      LAYER via ;
        RECT 324.400 243.480 324.660 243.740 ;
        RECT 330.840 243.480 331.100 243.740 ;
        RECT 330.840 23.840 331.100 24.100 ;
        RECT 633.060 23.840 633.320 24.100 ;
      LAYER met2 ;
        RECT 324.350 260.000 324.630 264.000 ;
        RECT 324.460 243.770 324.600 260.000 ;
        RECT 324.400 243.450 324.660 243.770 ;
        RECT 330.840 243.450 331.100 243.770 ;
        RECT 330.900 24.130 331.040 243.450 ;
        RECT 330.840 23.810 331.100 24.130 ;
        RECT 633.060 23.810 633.320 24.130 ;
        RECT 633.120 2.400 633.260 23.810 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2111.930 244.020 2112.250 244.080 ;
        RECT 2117.910 244.020 2118.230 244.080 ;
        RECT 2111.930 243.880 2118.230 244.020 ;
        RECT 2111.930 243.820 2112.250 243.880 ;
        RECT 2117.910 243.820 2118.230 243.880 ;
        RECT 2117.910 38.320 2118.230 38.380 ;
        RECT 2417.370 38.320 2417.690 38.380 ;
        RECT 2117.910 38.180 2417.690 38.320 ;
        RECT 2117.910 38.120 2118.230 38.180 ;
        RECT 2417.370 38.120 2417.690 38.180 ;
      LAYER via ;
        RECT 2111.960 243.820 2112.220 244.080 ;
        RECT 2117.940 243.820 2118.200 244.080 ;
        RECT 2117.940 38.120 2118.200 38.380 ;
        RECT 2417.400 38.120 2417.660 38.380 ;
      LAYER met2 ;
        RECT 2111.910 260.000 2112.190 264.000 ;
        RECT 2112.020 244.110 2112.160 260.000 ;
        RECT 2111.960 243.790 2112.220 244.110 ;
        RECT 2117.940 243.790 2118.200 244.110 ;
        RECT 2118.000 38.410 2118.140 243.790 ;
        RECT 2117.940 38.090 2118.200 38.410 ;
        RECT 2417.400 38.090 2417.660 38.410 ;
        RECT 2417.460 2.400 2417.600 38.090 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2129.870 237.900 2130.190 237.960 ;
        RECT 2428.870 237.900 2429.190 237.960 ;
        RECT 2129.870 237.760 2429.190 237.900 ;
        RECT 2129.870 237.700 2130.190 237.760 ;
        RECT 2428.870 237.700 2429.190 237.760 ;
        RECT 2428.870 18.260 2429.190 18.320 ;
        RECT 2434.850 18.260 2435.170 18.320 ;
        RECT 2428.870 18.120 2435.170 18.260 ;
        RECT 2428.870 18.060 2429.190 18.120 ;
        RECT 2434.850 18.060 2435.170 18.120 ;
      LAYER via ;
        RECT 2129.900 237.700 2130.160 237.960 ;
        RECT 2428.900 237.700 2429.160 237.960 ;
        RECT 2428.900 18.060 2429.160 18.320 ;
        RECT 2434.880 18.060 2435.140 18.320 ;
      LAYER met2 ;
        RECT 2129.850 260.000 2130.130 264.000 ;
        RECT 2129.960 237.990 2130.100 260.000 ;
        RECT 2129.900 237.670 2130.160 237.990 ;
        RECT 2428.900 237.670 2429.160 237.990 ;
        RECT 2428.960 18.350 2429.100 237.670 ;
        RECT 2428.900 18.030 2429.160 18.350 ;
        RECT 2434.880 18.030 2435.140 18.350 ;
        RECT 2434.940 2.400 2435.080 18.030 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2147.810 244.020 2148.130 244.080 ;
        RECT 2152.410 244.020 2152.730 244.080 ;
        RECT 2147.810 243.880 2152.730 244.020 ;
        RECT 2147.810 243.820 2148.130 243.880 ;
        RECT 2152.410 243.820 2152.730 243.880 ;
        RECT 2152.410 30.840 2152.730 30.900 ;
        RECT 2452.790 30.840 2453.110 30.900 ;
        RECT 2152.410 30.700 2453.110 30.840 ;
        RECT 2152.410 30.640 2152.730 30.700 ;
        RECT 2452.790 30.640 2453.110 30.700 ;
      LAYER via ;
        RECT 2147.840 243.820 2148.100 244.080 ;
        RECT 2152.440 243.820 2152.700 244.080 ;
        RECT 2152.440 30.640 2152.700 30.900 ;
        RECT 2452.820 30.640 2453.080 30.900 ;
      LAYER met2 ;
        RECT 2147.790 260.000 2148.070 264.000 ;
        RECT 2147.900 244.110 2148.040 260.000 ;
        RECT 2147.840 243.790 2148.100 244.110 ;
        RECT 2152.440 243.790 2152.700 244.110 ;
        RECT 2152.500 30.930 2152.640 243.790 ;
        RECT 2152.440 30.610 2152.700 30.930 ;
        RECT 2452.820 30.610 2453.080 30.930 ;
        RECT 2452.880 2.400 2453.020 30.610 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2165.750 244.020 2166.070 244.080 ;
        RECT 2169.890 244.020 2170.210 244.080 ;
        RECT 2165.750 243.880 2170.210 244.020 ;
        RECT 2165.750 243.820 2166.070 243.880 ;
        RECT 2169.890 243.820 2170.210 243.880 ;
        RECT 2169.890 44.780 2170.210 44.840 ;
        RECT 2470.730 44.780 2471.050 44.840 ;
        RECT 2169.890 44.640 2471.050 44.780 ;
        RECT 2169.890 44.580 2170.210 44.640 ;
        RECT 2470.730 44.580 2471.050 44.640 ;
      LAYER via ;
        RECT 2165.780 243.820 2166.040 244.080 ;
        RECT 2169.920 243.820 2170.180 244.080 ;
        RECT 2169.920 44.580 2170.180 44.840 ;
        RECT 2470.760 44.580 2471.020 44.840 ;
      LAYER met2 ;
        RECT 2165.730 260.000 2166.010 264.000 ;
        RECT 2165.840 244.110 2165.980 260.000 ;
        RECT 2165.780 243.790 2166.040 244.110 ;
        RECT 2169.920 243.790 2170.180 244.110 ;
        RECT 2169.980 44.870 2170.120 243.790 ;
        RECT 2169.920 44.550 2170.180 44.870 ;
        RECT 2470.760 44.550 2471.020 44.870 ;
        RECT 2470.820 2.400 2470.960 44.550 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2183.690 243.680 2184.010 243.740 ;
        RECT 2190.590 243.680 2190.910 243.740 ;
        RECT 2183.690 243.540 2190.910 243.680 ;
        RECT 2183.690 243.480 2184.010 243.540 ;
        RECT 2190.590 243.480 2190.910 243.540 ;
        RECT 2190.590 51.920 2190.910 51.980 ;
        RECT 2484.070 51.920 2484.390 51.980 ;
        RECT 2190.590 51.780 2484.390 51.920 ;
        RECT 2190.590 51.720 2190.910 51.780 ;
        RECT 2484.070 51.720 2484.390 51.780 ;
      LAYER via ;
        RECT 2183.720 243.480 2183.980 243.740 ;
        RECT 2190.620 243.480 2190.880 243.740 ;
        RECT 2190.620 51.720 2190.880 51.980 ;
        RECT 2484.100 51.720 2484.360 51.980 ;
      LAYER met2 ;
        RECT 2183.670 260.000 2183.950 264.000 ;
        RECT 2183.780 243.770 2183.920 260.000 ;
        RECT 2183.720 243.450 2183.980 243.770 ;
        RECT 2190.620 243.450 2190.880 243.770 ;
        RECT 2190.680 52.010 2190.820 243.450 ;
        RECT 2190.620 51.690 2190.880 52.010 ;
        RECT 2484.100 51.690 2484.360 52.010 ;
        RECT 2484.160 17.410 2484.300 51.690 ;
        RECT 2484.160 17.270 2488.900 17.410 ;
        RECT 2488.760 2.400 2488.900 17.270 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2201.630 248.440 2201.950 248.500 ;
        RECT 2211.290 248.440 2211.610 248.500 ;
        RECT 2201.630 248.300 2211.610 248.440 ;
        RECT 2201.630 248.240 2201.950 248.300 ;
        RECT 2211.290 248.240 2211.610 248.300 ;
        RECT 2211.290 59.060 2211.610 59.120 ;
        RECT 2504.770 59.060 2505.090 59.120 ;
        RECT 2211.290 58.920 2505.090 59.060 ;
        RECT 2211.290 58.860 2211.610 58.920 ;
        RECT 2504.770 58.860 2505.090 58.920 ;
      LAYER via ;
        RECT 2201.660 248.240 2201.920 248.500 ;
        RECT 2211.320 248.240 2211.580 248.500 ;
        RECT 2211.320 58.860 2211.580 59.120 ;
        RECT 2504.800 58.860 2505.060 59.120 ;
      LAYER met2 ;
        RECT 2201.610 260.000 2201.890 264.000 ;
        RECT 2201.720 248.530 2201.860 260.000 ;
        RECT 2201.660 248.210 2201.920 248.530 ;
        RECT 2211.320 248.210 2211.580 248.530 ;
        RECT 2211.380 59.150 2211.520 248.210 ;
        RECT 2211.320 58.830 2211.580 59.150 ;
        RECT 2504.800 58.830 2505.060 59.150 ;
        RECT 2504.860 16.730 2505.000 58.830 ;
        RECT 2504.860 16.590 2506.380 16.730 ;
        RECT 2506.240 2.400 2506.380 16.590 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2219.570 231.440 2219.890 231.500 ;
        RECT 2518.570 231.440 2518.890 231.500 ;
        RECT 2219.570 231.300 2518.890 231.440 ;
        RECT 2219.570 231.240 2219.890 231.300 ;
        RECT 2518.570 231.240 2518.890 231.300 ;
      LAYER via ;
        RECT 2219.600 231.240 2219.860 231.500 ;
        RECT 2518.600 231.240 2518.860 231.500 ;
      LAYER met2 ;
        RECT 2219.550 260.000 2219.830 264.000 ;
        RECT 2219.660 231.530 2219.800 260.000 ;
        RECT 2219.600 231.210 2219.860 231.530 ;
        RECT 2518.600 231.210 2518.860 231.530 ;
        RECT 2518.660 16.730 2518.800 231.210 ;
        RECT 2518.660 16.590 2524.320 16.730 ;
        RECT 2524.180 2.400 2524.320 16.590 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2237.050 244.020 2237.370 244.080 ;
        RECT 2242.110 244.020 2242.430 244.080 ;
        RECT 2237.050 243.880 2242.430 244.020 ;
        RECT 2237.050 243.820 2237.370 243.880 ;
        RECT 2242.110 243.820 2242.430 243.880 ;
        RECT 2242.110 65.520 2242.430 65.580 ;
        RECT 2539.270 65.520 2539.590 65.580 ;
        RECT 2242.110 65.380 2539.590 65.520 ;
        RECT 2242.110 65.320 2242.430 65.380 ;
        RECT 2539.270 65.320 2539.590 65.380 ;
      LAYER via ;
        RECT 2237.080 243.820 2237.340 244.080 ;
        RECT 2242.140 243.820 2242.400 244.080 ;
        RECT 2242.140 65.320 2242.400 65.580 ;
        RECT 2539.300 65.320 2539.560 65.580 ;
      LAYER met2 ;
        RECT 2237.030 260.000 2237.310 264.000 ;
        RECT 2237.140 244.110 2237.280 260.000 ;
        RECT 2237.080 243.790 2237.340 244.110 ;
        RECT 2242.140 243.790 2242.400 244.110 ;
        RECT 2242.200 65.610 2242.340 243.790 ;
        RECT 2242.140 65.290 2242.400 65.610 ;
        RECT 2539.300 65.290 2539.560 65.610 ;
        RECT 2539.360 16.730 2539.500 65.290 ;
        RECT 2539.360 16.590 2542.260 16.730 ;
        RECT 2542.120 2.400 2542.260 16.590 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2254.990 245.380 2255.310 245.440 ;
        RECT 2259.590 245.380 2259.910 245.440 ;
        RECT 2254.990 245.240 2259.910 245.380 ;
        RECT 2254.990 245.180 2255.310 245.240 ;
        RECT 2259.590 245.180 2259.910 245.240 ;
        RECT 2259.590 72.320 2259.910 72.380 ;
        RECT 2559.970 72.320 2560.290 72.380 ;
        RECT 2259.590 72.180 2560.290 72.320 ;
        RECT 2259.590 72.120 2259.910 72.180 ;
        RECT 2559.970 72.120 2560.290 72.180 ;
      LAYER via ;
        RECT 2255.020 245.180 2255.280 245.440 ;
        RECT 2259.620 245.180 2259.880 245.440 ;
        RECT 2259.620 72.120 2259.880 72.380 ;
        RECT 2560.000 72.120 2560.260 72.380 ;
      LAYER met2 ;
        RECT 2254.970 260.000 2255.250 264.000 ;
        RECT 2255.080 245.470 2255.220 260.000 ;
        RECT 2255.020 245.150 2255.280 245.470 ;
        RECT 2259.620 245.150 2259.880 245.470 ;
        RECT 2259.680 72.410 2259.820 245.150 ;
        RECT 2259.620 72.090 2259.880 72.410 ;
        RECT 2560.000 72.090 2560.260 72.410 ;
        RECT 2560.060 2.400 2560.200 72.090 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2276.610 24.720 2276.930 24.780 ;
        RECT 2577.910 24.720 2578.230 24.780 ;
        RECT 2276.610 24.580 2578.230 24.720 ;
        RECT 2276.610 24.520 2276.930 24.580 ;
        RECT 2577.910 24.520 2578.230 24.580 ;
      LAYER via ;
        RECT 2276.640 24.520 2276.900 24.780 ;
        RECT 2577.940 24.520 2578.200 24.780 ;
      LAYER met2 ;
        RECT 2272.910 260.170 2273.190 264.000 ;
        RECT 2272.910 260.030 2276.840 260.170 ;
        RECT 2272.910 260.000 2273.190 260.030 ;
        RECT 2276.700 24.810 2276.840 260.030 ;
        RECT 2276.640 24.490 2276.900 24.810 ;
        RECT 2577.940 24.490 2578.200 24.810 ;
        RECT 2578.000 2.400 2578.140 24.490 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 502.850 30.840 503.170 30.900 ;
        RECT 811.510 30.840 811.830 30.900 ;
        RECT 502.850 30.700 811.830 30.840 ;
        RECT 502.850 30.640 503.170 30.700 ;
        RECT 811.510 30.640 811.830 30.700 ;
      LAYER via ;
        RECT 502.880 30.640 503.140 30.900 ;
        RECT 811.540 30.640 811.800 30.900 ;
      LAYER met2 ;
        RECT 503.290 260.170 503.570 264.000 ;
        RECT 502.940 260.030 503.570 260.170 ;
        RECT 502.940 30.930 503.080 260.030 ;
        RECT 503.290 260.000 503.570 260.030 ;
        RECT 502.880 30.610 503.140 30.930 ;
        RECT 811.540 30.610 811.800 30.930 ;
        RECT 811.600 2.400 811.740 30.610 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2290.870 243.680 2291.190 243.740 ;
        RECT 2297.310 243.680 2297.630 243.740 ;
        RECT 2290.870 243.540 2297.630 243.680 ;
        RECT 2290.870 243.480 2291.190 243.540 ;
        RECT 2297.310 243.480 2297.630 243.540 ;
        RECT 2297.310 24.380 2297.630 24.440 ;
        RECT 2595.390 24.380 2595.710 24.440 ;
        RECT 2297.310 24.240 2595.710 24.380 ;
        RECT 2297.310 24.180 2297.630 24.240 ;
        RECT 2595.390 24.180 2595.710 24.240 ;
      LAYER via ;
        RECT 2290.900 243.480 2291.160 243.740 ;
        RECT 2297.340 243.480 2297.600 243.740 ;
        RECT 2297.340 24.180 2297.600 24.440 ;
        RECT 2595.420 24.180 2595.680 24.440 ;
      LAYER met2 ;
        RECT 2290.850 260.000 2291.130 264.000 ;
        RECT 2290.960 243.770 2291.100 260.000 ;
        RECT 2290.900 243.450 2291.160 243.770 ;
        RECT 2297.340 243.450 2297.600 243.770 ;
        RECT 2297.400 24.470 2297.540 243.450 ;
        RECT 2297.340 24.150 2297.600 24.470 ;
        RECT 2595.420 24.150 2595.680 24.470 ;
        RECT 2595.480 2.400 2595.620 24.150 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2311.110 26.080 2311.430 26.140 ;
        RECT 2613.330 26.080 2613.650 26.140 ;
        RECT 2311.110 25.940 2613.650 26.080 ;
        RECT 2311.110 25.880 2311.430 25.940 ;
        RECT 2613.330 25.880 2613.650 25.940 ;
      LAYER via ;
        RECT 2311.140 25.880 2311.400 26.140 ;
        RECT 2613.360 25.880 2613.620 26.140 ;
      LAYER met2 ;
        RECT 2308.790 260.170 2309.070 264.000 ;
        RECT 2308.790 260.030 2311.340 260.170 ;
        RECT 2308.790 260.000 2309.070 260.030 ;
        RECT 2311.200 26.170 2311.340 260.030 ;
        RECT 2311.140 25.850 2311.400 26.170 ;
        RECT 2613.360 25.850 2613.620 26.170 ;
        RECT 2613.420 2.400 2613.560 25.850 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2326.750 244.020 2327.070 244.080 ;
        RECT 2331.810 244.020 2332.130 244.080 ;
        RECT 2326.750 243.880 2332.130 244.020 ;
        RECT 2326.750 243.820 2327.070 243.880 ;
        RECT 2331.810 243.820 2332.130 243.880 ;
        RECT 2331.810 25.060 2332.130 25.120 ;
        RECT 2631.270 25.060 2631.590 25.120 ;
        RECT 2331.810 24.920 2631.590 25.060 ;
        RECT 2331.810 24.860 2332.130 24.920 ;
        RECT 2631.270 24.860 2631.590 24.920 ;
      LAYER via ;
        RECT 2326.780 243.820 2327.040 244.080 ;
        RECT 2331.840 243.820 2332.100 244.080 ;
        RECT 2331.840 24.860 2332.100 25.120 ;
        RECT 2631.300 24.860 2631.560 25.120 ;
      LAYER met2 ;
        RECT 2326.730 260.000 2327.010 264.000 ;
        RECT 2326.840 244.110 2326.980 260.000 ;
        RECT 2326.780 243.790 2327.040 244.110 ;
        RECT 2331.840 243.790 2332.100 244.110 ;
        RECT 2331.900 25.150 2332.040 243.790 ;
        RECT 2331.840 24.830 2332.100 25.150 ;
        RECT 2631.300 24.830 2631.560 25.150 ;
        RECT 2631.360 2.400 2631.500 24.830 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 79.460 2345.930 79.520 ;
        RECT 2643.230 79.460 2643.550 79.520 ;
        RECT 2345.610 79.320 2643.550 79.460 ;
        RECT 2345.610 79.260 2345.930 79.320 ;
        RECT 2643.230 79.260 2643.550 79.320 ;
        RECT 2643.230 17.920 2643.550 17.980 ;
        RECT 2649.210 17.920 2649.530 17.980 ;
        RECT 2643.230 17.780 2649.530 17.920 ;
        RECT 2643.230 17.720 2643.550 17.780 ;
        RECT 2649.210 17.720 2649.530 17.780 ;
      LAYER via ;
        RECT 2345.640 79.260 2345.900 79.520 ;
        RECT 2643.260 79.260 2643.520 79.520 ;
        RECT 2643.260 17.720 2643.520 17.980 ;
        RECT 2649.240 17.720 2649.500 17.980 ;
      LAYER met2 ;
        RECT 2344.670 260.170 2344.950 264.000 ;
        RECT 2344.670 260.030 2345.840 260.170 ;
        RECT 2344.670 260.000 2344.950 260.030 ;
        RECT 2345.700 79.550 2345.840 260.030 ;
        RECT 2345.640 79.230 2345.900 79.550 ;
        RECT 2643.260 79.230 2643.520 79.550 ;
        RECT 2643.320 18.010 2643.460 79.230 ;
        RECT 2643.260 17.690 2643.520 18.010 ;
        RECT 2649.240 17.690 2649.500 18.010 ;
        RECT 2649.300 2.400 2649.440 17.690 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2362.170 243.680 2362.490 243.740 ;
        RECT 2369.990 243.680 2370.310 243.740 ;
        RECT 2362.170 243.540 2370.310 243.680 ;
        RECT 2362.170 243.480 2362.490 243.540 ;
        RECT 2369.990 243.480 2370.310 243.540 ;
        RECT 2369.990 93.060 2370.310 93.120 ;
        RECT 2663.470 93.060 2663.790 93.120 ;
        RECT 2369.990 92.920 2663.790 93.060 ;
        RECT 2369.990 92.860 2370.310 92.920 ;
        RECT 2663.470 92.860 2663.790 92.920 ;
      LAYER via ;
        RECT 2362.200 243.480 2362.460 243.740 ;
        RECT 2370.020 243.480 2370.280 243.740 ;
        RECT 2370.020 92.860 2370.280 93.120 ;
        RECT 2663.500 92.860 2663.760 93.120 ;
      LAYER met2 ;
        RECT 2362.150 260.000 2362.430 264.000 ;
        RECT 2362.260 243.770 2362.400 260.000 ;
        RECT 2362.200 243.450 2362.460 243.770 ;
        RECT 2370.020 243.450 2370.280 243.770 ;
        RECT 2370.080 93.150 2370.220 243.450 ;
        RECT 2370.020 92.830 2370.280 93.150 ;
        RECT 2663.500 92.830 2663.760 93.150 ;
        RECT 2663.560 17.410 2663.700 92.830 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2380.110 24.040 2380.430 24.100 ;
        RECT 2684.630 24.040 2684.950 24.100 ;
        RECT 2380.110 23.900 2684.950 24.040 ;
        RECT 2380.110 23.840 2380.430 23.900 ;
        RECT 2684.630 23.840 2684.950 23.900 ;
      LAYER via ;
        RECT 2380.140 23.840 2380.400 24.100 ;
        RECT 2684.660 23.840 2684.920 24.100 ;
      LAYER met2 ;
        RECT 2380.090 260.000 2380.370 264.000 ;
        RECT 2380.200 24.130 2380.340 260.000 ;
        RECT 2380.140 23.810 2380.400 24.130 ;
        RECT 2684.660 23.810 2684.920 24.130 ;
        RECT 2684.720 2.400 2684.860 23.810 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.810 224.300 2401.130 224.360 ;
        RECT 2697.970 224.300 2698.290 224.360 ;
        RECT 2400.810 224.160 2698.290 224.300 ;
        RECT 2400.810 224.100 2401.130 224.160 ;
        RECT 2697.970 224.100 2698.290 224.160 ;
      LAYER via ;
        RECT 2400.840 224.100 2401.100 224.360 ;
        RECT 2698.000 224.100 2698.260 224.360 ;
      LAYER met2 ;
        RECT 2398.030 260.170 2398.310 264.000 ;
        RECT 2398.030 260.030 2401.040 260.170 ;
        RECT 2398.030 260.000 2398.310 260.030 ;
        RECT 2400.900 224.390 2401.040 260.030 ;
        RECT 2400.840 224.070 2401.100 224.390 ;
        RECT 2698.000 224.070 2698.260 224.390 ;
        RECT 2698.060 17.410 2698.200 224.070 ;
        RECT 2698.060 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2415.990 244.020 2416.310 244.080 ;
        RECT 2421.510 244.020 2421.830 244.080 ;
        RECT 2415.990 243.880 2421.830 244.020 ;
        RECT 2415.990 243.820 2416.310 243.880 ;
        RECT 2421.510 243.820 2421.830 243.880 ;
        RECT 2421.510 25.400 2421.830 25.460 ;
        RECT 2720.510 25.400 2720.830 25.460 ;
        RECT 2421.510 25.260 2720.830 25.400 ;
        RECT 2421.510 25.200 2421.830 25.260 ;
        RECT 2720.510 25.200 2720.830 25.260 ;
      LAYER via ;
        RECT 2416.020 243.820 2416.280 244.080 ;
        RECT 2421.540 243.820 2421.800 244.080 ;
        RECT 2421.540 25.200 2421.800 25.460 ;
        RECT 2720.540 25.200 2720.800 25.460 ;
      LAYER met2 ;
        RECT 2415.970 260.000 2416.250 264.000 ;
        RECT 2416.080 244.110 2416.220 260.000 ;
        RECT 2416.020 243.790 2416.280 244.110 ;
        RECT 2421.540 243.790 2421.800 244.110 ;
        RECT 2421.600 25.490 2421.740 243.790 ;
        RECT 2421.540 25.170 2421.800 25.490 ;
        RECT 2720.540 25.170 2720.800 25.490 ;
        RECT 2720.600 2.400 2720.740 25.170 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2435.310 25.740 2435.630 25.800 ;
        RECT 2738.450 25.740 2738.770 25.800 ;
        RECT 2435.310 25.600 2738.770 25.740 ;
        RECT 2435.310 25.540 2435.630 25.600 ;
        RECT 2738.450 25.540 2738.770 25.600 ;
      LAYER via ;
        RECT 2435.340 25.540 2435.600 25.800 ;
        RECT 2738.480 25.540 2738.740 25.800 ;
      LAYER met2 ;
        RECT 2433.910 260.170 2434.190 264.000 ;
        RECT 2433.910 260.030 2435.540 260.170 ;
        RECT 2433.910 260.000 2434.190 260.030 ;
        RECT 2435.400 25.830 2435.540 260.030 ;
        RECT 2435.340 25.510 2435.600 25.830 ;
        RECT 2738.480 25.510 2738.740 25.830 ;
        RECT 2738.540 2.400 2738.680 25.510 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2451.870 237.900 2452.190 237.960 ;
        RECT 2753.170 237.900 2753.490 237.960 ;
        RECT 2451.870 237.760 2753.490 237.900 ;
        RECT 2451.870 237.700 2452.190 237.760 ;
        RECT 2753.170 237.700 2753.490 237.760 ;
      LAYER via ;
        RECT 2451.900 237.700 2452.160 237.960 ;
        RECT 2753.200 237.700 2753.460 237.960 ;
      LAYER met2 ;
        RECT 2451.850 260.000 2452.130 264.000 ;
        RECT 2451.960 237.990 2452.100 260.000 ;
        RECT 2451.900 237.670 2452.160 237.990 ;
        RECT 2753.200 237.670 2753.460 237.990 ;
        RECT 2753.260 17.410 2753.400 237.670 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 524.010 37.980 524.330 38.040 ;
        RECT 829.450 37.980 829.770 38.040 ;
        RECT 524.010 37.840 829.770 37.980 ;
        RECT 524.010 37.780 524.330 37.840 ;
        RECT 829.450 37.780 829.770 37.840 ;
      LAYER via ;
        RECT 524.040 37.780 524.300 38.040 ;
        RECT 829.480 37.780 829.740 38.040 ;
      LAYER met2 ;
        RECT 521.230 260.170 521.510 264.000 ;
        RECT 521.230 260.030 524.240 260.170 ;
        RECT 521.230 260.000 521.510 260.030 ;
        RECT 524.100 38.070 524.240 260.030 ;
        RECT 524.040 37.750 524.300 38.070 ;
        RECT 829.480 37.750 829.740 38.070 ;
        RECT 829.540 2.400 829.680 37.750 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2469.350 217.160 2469.670 217.220 ;
        RECT 2773.870 217.160 2774.190 217.220 ;
        RECT 2469.350 217.020 2774.190 217.160 ;
        RECT 2469.350 216.960 2469.670 217.020 ;
        RECT 2773.870 216.960 2774.190 217.020 ;
      LAYER via ;
        RECT 2469.380 216.960 2469.640 217.220 ;
        RECT 2773.900 216.960 2774.160 217.220 ;
      LAYER met2 ;
        RECT 2469.790 260.170 2470.070 264.000 ;
        RECT 2469.440 260.030 2470.070 260.170 ;
        RECT 2469.440 217.250 2469.580 260.030 ;
        RECT 2469.790 260.000 2470.070 260.030 ;
        RECT 2469.380 216.930 2469.640 217.250 ;
        RECT 2773.900 216.930 2774.160 217.250 ;
        RECT 2773.960 2.400 2774.100 216.930 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2490.510 210.360 2490.830 210.420 ;
        RECT 2787.670 210.360 2787.990 210.420 ;
        RECT 2490.510 210.220 2787.990 210.360 ;
        RECT 2490.510 210.160 2490.830 210.220 ;
        RECT 2787.670 210.160 2787.990 210.220 ;
      LAYER via ;
        RECT 2490.540 210.160 2490.800 210.420 ;
        RECT 2787.700 210.160 2787.960 210.420 ;
      LAYER met2 ;
        RECT 2487.270 260.170 2487.550 264.000 ;
        RECT 2487.270 260.030 2490.740 260.170 ;
        RECT 2487.270 260.000 2487.550 260.030 ;
        RECT 2490.600 210.450 2490.740 260.030 ;
        RECT 2490.540 210.130 2490.800 210.450 ;
        RECT 2787.700 210.130 2787.960 210.450 ;
        RECT 2787.760 17.410 2787.900 210.130 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2505.230 244.020 2505.550 244.080 ;
        RECT 2511.210 244.020 2511.530 244.080 ;
        RECT 2505.230 243.880 2511.530 244.020 ;
        RECT 2505.230 243.820 2505.550 243.880 ;
        RECT 2511.210 243.820 2511.530 243.880 ;
        RECT 2511.210 30.840 2511.530 30.900 ;
        RECT 2809.750 30.840 2810.070 30.900 ;
        RECT 2511.210 30.700 2810.070 30.840 ;
        RECT 2511.210 30.640 2511.530 30.700 ;
        RECT 2809.750 30.640 2810.070 30.700 ;
      LAYER via ;
        RECT 2505.260 243.820 2505.520 244.080 ;
        RECT 2511.240 243.820 2511.500 244.080 ;
        RECT 2511.240 30.640 2511.500 30.900 ;
        RECT 2809.780 30.640 2810.040 30.900 ;
      LAYER met2 ;
        RECT 2505.210 260.000 2505.490 264.000 ;
        RECT 2505.320 244.110 2505.460 260.000 ;
        RECT 2505.260 243.790 2505.520 244.110 ;
        RECT 2511.240 243.790 2511.500 244.110 ;
        RECT 2511.300 30.930 2511.440 243.790 ;
        RECT 2511.240 30.610 2511.500 30.930 ;
        RECT 2809.780 30.610 2810.040 30.930 ;
        RECT 2809.840 2.400 2809.980 30.610 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2523.170 231.100 2523.490 231.160 ;
        RECT 2822.170 231.100 2822.490 231.160 ;
        RECT 2523.170 230.960 2822.490 231.100 ;
        RECT 2523.170 230.900 2523.490 230.960 ;
        RECT 2822.170 230.900 2822.490 230.960 ;
      LAYER via ;
        RECT 2523.200 230.900 2523.460 231.160 ;
        RECT 2822.200 230.900 2822.460 231.160 ;
      LAYER met2 ;
        RECT 2523.150 260.000 2523.430 264.000 ;
        RECT 2523.260 231.190 2523.400 260.000 ;
        RECT 2523.200 230.870 2523.460 231.190 ;
        RECT 2822.200 230.870 2822.460 231.190 ;
        RECT 2822.260 17.410 2822.400 230.870 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2541.110 244.020 2541.430 244.080 ;
        RECT 2545.710 244.020 2546.030 244.080 ;
        RECT 2541.110 243.880 2546.030 244.020 ;
        RECT 2541.110 243.820 2541.430 243.880 ;
        RECT 2545.710 243.820 2546.030 243.880 ;
        RECT 2545.710 196.760 2546.030 196.820 ;
        RECT 2842.870 196.760 2843.190 196.820 ;
        RECT 2545.710 196.620 2843.190 196.760 ;
        RECT 2545.710 196.560 2546.030 196.620 ;
        RECT 2842.870 196.560 2843.190 196.620 ;
      LAYER via ;
        RECT 2541.140 243.820 2541.400 244.080 ;
        RECT 2545.740 243.820 2546.000 244.080 ;
        RECT 2545.740 196.560 2546.000 196.820 ;
        RECT 2842.900 196.560 2843.160 196.820 ;
      LAYER met2 ;
        RECT 2541.090 260.000 2541.370 264.000 ;
        RECT 2541.200 244.110 2541.340 260.000 ;
        RECT 2541.140 243.790 2541.400 244.110 ;
        RECT 2545.740 243.790 2546.000 244.110 ;
        RECT 2545.800 196.850 2545.940 243.790 ;
        RECT 2545.740 196.530 2546.000 196.850 ;
        RECT 2842.900 196.530 2843.160 196.850 ;
        RECT 2842.960 17.410 2843.100 196.530 ;
        RECT 2842.960 17.270 2845.400 17.410 ;
        RECT 2845.260 2.400 2845.400 17.270 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2559.050 189.620 2559.370 189.680 ;
        RECT 2857.130 189.620 2857.450 189.680 ;
        RECT 2559.050 189.480 2857.450 189.620 ;
        RECT 2559.050 189.420 2559.370 189.480 ;
        RECT 2857.130 189.420 2857.450 189.480 ;
        RECT 2857.130 17.580 2857.450 17.640 ;
        RECT 2863.110 17.580 2863.430 17.640 ;
        RECT 2857.130 17.440 2863.430 17.580 ;
        RECT 2857.130 17.380 2857.450 17.440 ;
        RECT 2863.110 17.380 2863.430 17.440 ;
      LAYER via ;
        RECT 2559.080 189.420 2559.340 189.680 ;
        RECT 2857.160 189.420 2857.420 189.680 ;
        RECT 2857.160 17.380 2857.420 17.640 ;
        RECT 2863.140 17.380 2863.400 17.640 ;
      LAYER met2 ;
        RECT 2559.030 260.000 2559.310 264.000 ;
        RECT 2559.140 189.710 2559.280 260.000 ;
        RECT 2559.080 189.390 2559.340 189.710 ;
        RECT 2857.160 189.390 2857.420 189.710 ;
        RECT 2857.220 17.670 2857.360 189.390 ;
        RECT 2857.160 17.350 2857.420 17.670 ;
        RECT 2863.140 17.350 2863.400 17.670 ;
        RECT 2863.200 2.400 2863.340 17.350 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2580.210 182.820 2580.530 182.880 ;
        RECT 2873.690 182.820 2874.010 182.880 ;
        RECT 2580.210 182.680 2874.010 182.820 ;
        RECT 2580.210 182.620 2580.530 182.680 ;
        RECT 2873.690 182.620 2874.010 182.680 ;
        RECT 2873.690 17.580 2874.010 17.640 ;
        RECT 2881.050 17.580 2881.370 17.640 ;
        RECT 2873.690 17.440 2881.370 17.580 ;
        RECT 2873.690 17.380 2874.010 17.440 ;
        RECT 2881.050 17.380 2881.370 17.440 ;
      LAYER via ;
        RECT 2580.240 182.620 2580.500 182.880 ;
        RECT 2873.720 182.620 2873.980 182.880 ;
        RECT 2873.720 17.380 2873.980 17.640 ;
        RECT 2881.080 17.380 2881.340 17.640 ;
      LAYER met2 ;
        RECT 2576.970 260.170 2577.250 264.000 ;
        RECT 2576.970 260.030 2580.440 260.170 ;
        RECT 2576.970 260.000 2577.250 260.030 ;
        RECT 2580.300 182.910 2580.440 260.030 ;
        RECT 2580.240 182.590 2580.500 182.910 ;
        RECT 2873.720 182.590 2873.980 182.910 ;
        RECT 2873.780 17.670 2873.920 182.590 ;
        RECT 2873.720 17.350 2873.980 17.670 ;
        RECT 2881.080 17.350 2881.340 17.670 ;
        RECT 2881.140 2.400 2881.280 17.350 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2594.930 244.020 2595.250 244.080 ;
        RECT 2600.450 244.020 2600.770 244.080 ;
        RECT 2594.930 243.880 2600.770 244.020 ;
        RECT 2594.930 243.820 2595.250 243.880 ;
        RECT 2600.450 243.820 2600.770 243.880 ;
        RECT 2600.450 37.980 2600.770 38.040 ;
        RECT 2898.990 37.980 2899.310 38.040 ;
        RECT 2600.450 37.840 2899.310 37.980 ;
        RECT 2600.450 37.780 2600.770 37.840 ;
        RECT 2898.990 37.780 2899.310 37.840 ;
      LAYER via ;
        RECT 2594.960 243.820 2595.220 244.080 ;
        RECT 2600.480 243.820 2600.740 244.080 ;
        RECT 2600.480 37.780 2600.740 38.040 ;
        RECT 2899.020 37.780 2899.280 38.040 ;
      LAYER met2 ;
        RECT 2594.910 260.000 2595.190 264.000 ;
        RECT 2595.020 244.110 2595.160 260.000 ;
        RECT 2594.960 243.790 2595.220 244.110 ;
        RECT 2600.480 243.790 2600.740 244.110 ;
        RECT 2600.540 38.070 2600.680 243.790 ;
        RECT 2600.480 37.750 2600.740 38.070 ;
        RECT 2899.020 37.750 2899.280 38.070 ;
        RECT 2899.080 2.400 2899.220 37.750 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 539.190 244.020 539.510 244.080 ;
        RECT 544.710 244.020 545.030 244.080 ;
        RECT 539.190 243.880 545.030 244.020 ;
        RECT 539.190 243.820 539.510 243.880 ;
        RECT 544.710 243.820 545.030 243.880 ;
        RECT 544.710 44.780 545.030 44.840 ;
        RECT 846.930 44.780 847.250 44.840 ;
        RECT 544.710 44.640 847.250 44.780 ;
        RECT 544.710 44.580 545.030 44.640 ;
        RECT 846.930 44.580 847.250 44.640 ;
      LAYER via ;
        RECT 539.220 243.820 539.480 244.080 ;
        RECT 544.740 243.820 545.000 244.080 ;
        RECT 544.740 44.580 545.000 44.840 ;
        RECT 846.960 44.580 847.220 44.840 ;
      LAYER met2 ;
        RECT 539.170 260.000 539.450 264.000 ;
        RECT 539.280 244.110 539.420 260.000 ;
        RECT 539.220 243.790 539.480 244.110 ;
        RECT 544.740 243.790 545.000 244.110 ;
        RECT 544.800 44.870 544.940 243.790 ;
        RECT 544.740 44.550 545.000 44.870 ;
        RECT 846.960 44.550 847.220 44.870 ;
        RECT 847.020 2.400 847.160 44.550 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.510 51.580 558.830 51.640 ;
        RECT 862.570 51.580 862.890 51.640 ;
        RECT 558.510 51.440 862.890 51.580 ;
        RECT 558.510 51.380 558.830 51.440 ;
        RECT 862.570 51.380 862.890 51.440 ;
      LAYER via ;
        RECT 558.540 51.380 558.800 51.640 ;
        RECT 862.600 51.380 862.860 51.640 ;
      LAYER met2 ;
        RECT 557.110 260.170 557.390 264.000 ;
        RECT 557.110 260.030 558.740 260.170 ;
        RECT 557.110 260.000 557.390 260.030 ;
        RECT 558.600 51.670 558.740 260.030 ;
        RECT 558.540 51.350 558.800 51.670 ;
        RECT 862.600 51.350 862.860 51.670 ;
        RECT 862.660 16.730 862.800 51.350 ;
        RECT 862.660 16.590 865.100 16.730 ;
        RECT 864.960 2.400 865.100 16.590 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 574.610 244.020 574.930 244.080 ;
        RECT 579.210 244.020 579.530 244.080 ;
        RECT 574.610 243.880 579.530 244.020 ;
        RECT 574.610 243.820 574.930 243.880 ;
        RECT 579.210 243.820 579.530 243.880 ;
        RECT 579.210 58.720 579.530 58.780 ;
        RECT 876.830 58.720 877.150 58.780 ;
        RECT 579.210 58.580 877.150 58.720 ;
        RECT 579.210 58.520 579.530 58.580 ;
        RECT 876.830 58.520 877.150 58.580 ;
        RECT 876.830 18.600 877.150 18.660 ;
        RECT 882.810 18.600 883.130 18.660 ;
        RECT 876.830 18.460 883.130 18.600 ;
        RECT 876.830 18.400 877.150 18.460 ;
        RECT 882.810 18.400 883.130 18.460 ;
      LAYER via ;
        RECT 574.640 243.820 574.900 244.080 ;
        RECT 579.240 243.820 579.500 244.080 ;
        RECT 579.240 58.520 579.500 58.780 ;
        RECT 876.860 58.520 877.120 58.780 ;
        RECT 876.860 18.400 877.120 18.660 ;
        RECT 882.840 18.400 883.100 18.660 ;
      LAYER met2 ;
        RECT 574.590 260.000 574.870 264.000 ;
        RECT 574.700 244.110 574.840 260.000 ;
        RECT 574.640 243.790 574.900 244.110 ;
        RECT 579.240 243.790 579.500 244.110 ;
        RECT 579.300 58.810 579.440 243.790 ;
        RECT 579.240 58.490 579.500 58.810 ;
        RECT 876.860 58.490 877.120 58.810 ;
        RECT 876.920 18.690 877.060 58.490 ;
        RECT 876.860 18.370 877.120 18.690 ;
        RECT 882.840 18.370 883.100 18.690 ;
        RECT 882.900 2.400 883.040 18.370 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 592.550 65.520 592.870 65.580 ;
        RECT 897.070 65.520 897.390 65.580 ;
        RECT 592.550 65.380 897.390 65.520 ;
        RECT 592.550 65.320 592.870 65.380 ;
        RECT 897.070 65.320 897.390 65.380 ;
      LAYER via ;
        RECT 592.580 65.320 592.840 65.580 ;
        RECT 897.100 65.320 897.360 65.580 ;
      LAYER met2 ;
        RECT 592.530 260.000 592.810 264.000 ;
        RECT 592.640 65.610 592.780 260.000 ;
        RECT 592.580 65.290 592.840 65.610 ;
        RECT 897.100 65.290 897.360 65.610 ;
        RECT 897.160 16.730 897.300 65.290 ;
        RECT 897.160 16.590 900.980 16.730 ;
        RECT 900.840 2.400 900.980 16.590 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 613.710 72.320 614.030 72.380 ;
        RECT 918.230 72.320 918.550 72.380 ;
        RECT 613.710 72.180 918.550 72.320 ;
        RECT 613.710 72.120 614.030 72.180 ;
        RECT 918.230 72.120 918.550 72.180 ;
      LAYER via ;
        RECT 613.740 72.120 614.000 72.380 ;
        RECT 918.260 72.120 918.520 72.380 ;
      LAYER met2 ;
        RECT 610.470 260.170 610.750 264.000 ;
        RECT 610.470 260.030 613.940 260.170 ;
        RECT 610.470 260.000 610.750 260.030 ;
        RECT 613.800 72.410 613.940 260.030 ;
        RECT 613.740 72.090 614.000 72.410 ;
        RECT 918.260 72.090 918.520 72.410 ;
        RECT 918.320 17.410 918.460 72.090 ;
        RECT 918.320 17.270 918.920 17.410 ;
        RECT 918.780 2.400 918.920 17.270 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 628.430 243.340 628.750 243.400 ;
        RECT 633.950 243.340 634.270 243.400 ;
        RECT 628.430 243.200 634.270 243.340 ;
        RECT 628.430 243.140 628.750 243.200 ;
        RECT 633.950 243.140 634.270 243.200 ;
        RECT 633.950 79.800 634.270 79.860 ;
        RECT 931.570 79.800 931.890 79.860 ;
        RECT 633.950 79.660 931.890 79.800 ;
        RECT 633.950 79.600 634.270 79.660 ;
        RECT 931.570 79.600 931.890 79.660 ;
      LAYER via ;
        RECT 628.460 243.140 628.720 243.400 ;
        RECT 633.980 243.140 634.240 243.400 ;
        RECT 633.980 79.600 634.240 79.860 ;
        RECT 931.600 79.600 931.860 79.860 ;
      LAYER met2 ;
        RECT 628.410 260.000 628.690 264.000 ;
        RECT 628.520 243.430 628.660 260.000 ;
        RECT 628.460 243.110 628.720 243.430 ;
        RECT 633.980 243.110 634.240 243.430 ;
        RECT 634.040 79.890 634.180 243.110 ;
        RECT 633.980 79.570 634.240 79.890 ;
        RECT 931.600 79.570 931.860 79.890 ;
        RECT 931.660 16.730 931.800 79.570 ;
        RECT 931.660 16.590 936.400 16.730 ;
        RECT 936.260 2.400 936.400 16.590 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 86.600 648.530 86.660 ;
        RECT 952.270 86.600 952.590 86.660 ;
        RECT 648.210 86.460 952.590 86.600 ;
        RECT 648.210 86.400 648.530 86.460 ;
        RECT 952.270 86.400 952.590 86.460 ;
      LAYER via ;
        RECT 648.240 86.400 648.500 86.660 ;
        RECT 952.300 86.400 952.560 86.660 ;
      LAYER met2 ;
        RECT 646.350 260.170 646.630 264.000 ;
        RECT 646.350 260.030 648.440 260.170 ;
        RECT 646.350 260.000 646.630 260.030 ;
        RECT 648.300 86.690 648.440 260.030 ;
        RECT 648.240 86.370 648.500 86.690 ;
        RECT 952.300 86.370 952.560 86.690 ;
        RECT 952.360 16.730 952.500 86.370 ;
        RECT 952.360 16.590 954.340 16.730 ;
        RECT 954.200 2.400 954.340 16.590 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 664.310 244.020 664.630 244.080 ;
        RECT 668.910 244.020 669.230 244.080 ;
        RECT 664.310 243.880 669.230 244.020 ;
        RECT 664.310 243.820 664.630 243.880 ;
        RECT 668.910 243.820 669.230 243.880 ;
        RECT 668.910 24.380 669.230 24.440 ;
        RECT 972.050 24.380 972.370 24.440 ;
        RECT 668.910 24.240 972.370 24.380 ;
        RECT 668.910 24.180 669.230 24.240 ;
        RECT 972.050 24.180 972.370 24.240 ;
      LAYER via ;
        RECT 664.340 243.820 664.600 244.080 ;
        RECT 668.940 243.820 669.200 244.080 ;
        RECT 668.940 24.180 669.200 24.440 ;
        RECT 972.080 24.180 972.340 24.440 ;
      LAYER met2 ;
        RECT 664.290 260.000 664.570 264.000 ;
        RECT 664.400 244.110 664.540 260.000 ;
        RECT 664.340 243.790 664.600 244.110 ;
        RECT 668.940 243.790 669.200 244.110 ;
        RECT 669.000 24.470 669.140 243.790 ;
        RECT 668.940 24.150 669.200 24.470 ;
        RECT 972.080 24.150 972.340 24.470 ;
        RECT 972.140 2.400 972.280 24.150 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 344.610 24.380 344.930 24.440 ;
        RECT 650.970 24.380 651.290 24.440 ;
        RECT 344.610 24.240 651.290 24.380 ;
        RECT 344.610 24.180 344.930 24.240 ;
        RECT 650.970 24.180 651.290 24.240 ;
      LAYER via ;
        RECT 344.640 24.180 344.900 24.440 ;
        RECT 651.000 24.180 651.260 24.440 ;
      LAYER met2 ;
        RECT 342.290 260.170 342.570 264.000 ;
        RECT 342.290 260.030 344.840 260.170 ;
        RECT 342.290 260.000 342.570 260.030 ;
        RECT 344.700 24.470 344.840 260.030 ;
        RECT 344.640 24.150 344.900 24.470 ;
        RECT 651.000 24.150 651.260 24.470 ;
        RECT 651.060 2.400 651.200 24.150 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 238.240 683.030 238.300 ;
        RECT 986.770 238.240 987.090 238.300 ;
        RECT 682.710 238.100 987.090 238.240 ;
        RECT 682.710 238.040 683.030 238.100 ;
        RECT 986.770 238.040 987.090 238.100 ;
      LAYER via ;
        RECT 682.740 238.040 683.000 238.300 ;
        RECT 986.800 238.040 987.060 238.300 ;
      LAYER met2 ;
        RECT 682.230 260.170 682.510 264.000 ;
        RECT 682.230 260.030 682.940 260.170 ;
        RECT 682.230 260.000 682.510 260.030 ;
        RECT 682.800 238.330 682.940 260.030 ;
        RECT 682.740 238.010 683.000 238.330 ;
        RECT 986.800 238.010 987.060 238.330 ;
        RECT 986.860 16.730 987.000 238.010 ;
        RECT 986.860 16.590 990.220 16.730 ;
        RECT 990.080 2.400 990.220 16.590 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 93.060 703.730 93.120 ;
        RECT 1007.930 93.060 1008.250 93.120 ;
        RECT 703.410 92.920 1008.250 93.060 ;
        RECT 703.410 92.860 703.730 92.920 ;
        RECT 1007.930 92.860 1008.250 92.920 ;
      LAYER via ;
        RECT 703.440 92.860 703.700 93.120 ;
        RECT 1007.960 92.860 1008.220 93.120 ;
      LAYER met2 ;
        RECT 699.710 260.170 699.990 264.000 ;
        RECT 699.710 260.030 703.640 260.170 ;
        RECT 699.710 260.000 699.990 260.030 ;
        RECT 703.500 93.150 703.640 260.030 ;
        RECT 703.440 92.830 703.700 93.150 ;
        RECT 1007.960 92.830 1008.220 93.150 ;
        RECT 1008.020 17.410 1008.160 92.830 ;
        RECT 1007.560 17.270 1008.160 17.410 ;
        RECT 1007.560 2.400 1007.700 17.270 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.670 244.020 717.990 244.080 ;
        RECT 724.110 244.020 724.430 244.080 ;
        RECT 717.670 243.880 724.430 244.020 ;
        RECT 717.670 243.820 717.990 243.880 ;
        RECT 724.110 243.820 724.430 243.880 ;
        RECT 724.110 99.860 724.430 99.920 ;
        RECT 1021.270 99.860 1021.590 99.920 ;
        RECT 724.110 99.720 1021.590 99.860 ;
        RECT 724.110 99.660 724.430 99.720 ;
        RECT 1021.270 99.660 1021.590 99.720 ;
      LAYER via ;
        RECT 717.700 243.820 717.960 244.080 ;
        RECT 724.140 243.820 724.400 244.080 ;
        RECT 724.140 99.660 724.400 99.920 ;
        RECT 1021.300 99.660 1021.560 99.920 ;
      LAYER met2 ;
        RECT 717.650 260.000 717.930 264.000 ;
        RECT 717.760 244.110 717.900 260.000 ;
        RECT 717.700 243.790 717.960 244.110 ;
        RECT 724.140 243.790 724.400 244.110 ;
        RECT 724.200 99.950 724.340 243.790 ;
        RECT 724.140 99.630 724.400 99.950 ;
        RECT 1021.300 99.630 1021.560 99.950 ;
        RECT 1021.360 16.730 1021.500 99.630 ;
        RECT 1021.360 16.590 1025.640 16.730 ;
        RECT 1025.500 2.400 1025.640 16.590 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 107.000 738.230 107.060 ;
        RECT 1041.970 107.000 1042.290 107.060 ;
        RECT 737.910 106.860 1042.290 107.000 ;
        RECT 737.910 106.800 738.230 106.860 ;
        RECT 1041.970 106.800 1042.290 106.860 ;
      LAYER via ;
        RECT 737.940 106.800 738.200 107.060 ;
        RECT 1042.000 106.800 1042.260 107.060 ;
      LAYER met2 ;
        RECT 735.590 260.170 735.870 264.000 ;
        RECT 735.590 260.030 738.140 260.170 ;
        RECT 735.590 260.000 735.870 260.030 ;
        RECT 738.000 107.090 738.140 260.030 ;
        RECT 737.940 106.770 738.200 107.090 ;
        RECT 1042.000 106.770 1042.260 107.090 ;
        RECT 1042.060 16.730 1042.200 106.770 ;
        RECT 1042.060 16.590 1043.580 16.730 ;
        RECT 1043.440 2.400 1043.580 16.590 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 753.550 244.020 753.870 244.080 ;
        RECT 758.610 244.020 758.930 244.080 ;
        RECT 753.550 243.880 758.930 244.020 ;
        RECT 753.550 243.820 753.870 243.880 ;
        RECT 758.610 243.820 758.930 243.880 ;
        RECT 758.610 113.800 758.930 113.860 ;
        RECT 1055.770 113.800 1056.090 113.860 ;
        RECT 758.610 113.660 1056.090 113.800 ;
        RECT 758.610 113.600 758.930 113.660 ;
        RECT 1055.770 113.600 1056.090 113.660 ;
      LAYER via ;
        RECT 753.580 243.820 753.840 244.080 ;
        RECT 758.640 243.820 758.900 244.080 ;
        RECT 758.640 113.600 758.900 113.860 ;
        RECT 1055.800 113.600 1056.060 113.860 ;
      LAYER met2 ;
        RECT 753.530 260.000 753.810 264.000 ;
        RECT 753.640 244.110 753.780 260.000 ;
        RECT 753.580 243.790 753.840 244.110 ;
        RECT 758.640 243.790 758.900 244.110 ;
        RECT 758.700 113.890 758.840 243.790 ;
        RECT 758.640 113.570 758.900 113.890 ;
        RECT 1055.800 113.570 1056.060 113.890 ;
        RECT 1055.860 16.730 1056.000 113.570 ;
        RECT 1055.860 16.590 1061.520 16.730 ;
        RECT 1061.380 2.400 1061.520 16.590 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 772.410 120.600 772.730 120.660 ;
        RECT 1076.470 120.600 1076.790 120.660 ;
        RECT 772.410 120.460 1076.790 120.600 ;
        RECT 772.410 120.400 772.730 120.460 ;
        RECT 1076.470 120.400 1076.790 120.460 ;
      LAYER via ;
        RECT 772.440 120.400 772.700 120.660 ;
        RECT 1076.500 120.400 1076.760 120.660 ;
      LAYER met2 ;
        RECT 771.470 260.170 771.750 264.000 ;
        RECT 771.470 260.030 772.640 260.170 ;
        RECT 771.470 260.000 771.750 260.030 ;
        RECT 772.500 120.690 772.640 260.030 ;
        RECT 772.440 120.370 772.700 120.690 ;
        RECT 1076.500 120.370 1076.760 120.690 ;
        RECT 1076.560 16.730 1076.700 120.370 ;
        RECT 1076.560 16.590 1079.460 16.730 ;
        RECT 1079.320 2.400 1079.460 16.590 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 789.430 244.020 789.750 244.080 ;
        RECT 793.110 244.020 793.430 244.080 ;
        RECT 789.430 243.880 793.430 244.020 ;
        RECT 789.430 243.820 789.750 243.880 ;
        RECT 793.110 243.820 793.430 243.880 ;
        RECT 793.110 127.740 793.430 127.800 ;
        RECT 1090.270 127.740 1090.590 127.800 ;
        RECT 793.110 127.600 1090.590 127.740 ;
        RECT 793.110 127.540 793.430 127.600 ;
        RECT 1090.270 127.540 1090.590 127.600 ;
        RECT 1090.270 16.560 1090.590 16.620 ;
        RECT 1096.710 16.560 1097.030 16.620 ;
        RECT 1090.270 16.420 1097.030 16.560 ;
        RECT 1090.270 16.360 1090.590 16.420 ;
        RECT 1096.710 16.360 1097.030 16.420 ;
      LAYER via ;
        RECT 789.460 243.820 789.720 244.080 ;
        RECT 793.140 243.820 793.400 244.080 ;
        RECT 793.140 127.540 793.400 127.800 ;
        RECT 1090.300 127.540 1090.560 127.800 ;
        RECT 1090.300 16.360 1090.560 16.620 ;
        RECT 1096.740 16.360 1097.000 16.620 ;
      LAYER met2 ;
        RECT 789.410 260.000 789.690 264.000 ;
        RECT 789.520 244.110 789.660 260.000 ;
        RECT 789.460 243.790 789.720 244.110 ;
        RECT 793.140 243.790 793.400 244.110 ;
        RECT 793.200 127.830 793.340 243.790 ;
        RECT 793.140 127.510 793.400 127.830 ;
        RECT 1090.300 127.510 1090.560 127.830 ;
        RECT 1090.360 16.650 1090.500 127.510 ;
        RECT 1090.300 16.330 1090.560 16.650 ;
        RECT 1096.740 16.330 1097.000 16.650 ;
        RECT 1096.800 2.400 1096.940 16.330 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 807.370 243.680 807.690 243.740 ;
        RECT 838.190 243.680 838.510 243.740 ;
        RECT 807.370 243.540 838.510 243.680 ;
        RECT 807.370 243.480 807.690 243.540 ;
        RECT 838.190 243.480 838.510 243.540 ;
        RECT 838.190 31.520 838.510 31.580 ;
        RECT 1114.650 31.520 1114.970 31.580 ;
        RECT 838.190 31.380 1114.970 31.520 ;
        RECT 838.190 31.320 838.510 31.380 ;
        RECT 1114.650 31.320 1114.970 31.380 ;
      LAYER via ;
        RECT 807.400 243.480 807.660 243.740 ;
        RECT 838.220 243.480 838.480 243.740 ;
        RECT 838.220 31.320 838.480 31.580 ;
        RECT 1114.680 31.320 1114.940 31.580 ;
      LAYER met2 ;
        RECT 807.350 260.000 807.630 264.000 ;
        RECT 807.460 243.770 807.600 260.000 ;
        RECT 807.400 243.450 807.660 243.770 ;
        RECT 838.220 243.450 838.480 243.770 ;
        RECT 838.280 31.610 838.420 243.450 ;
        RECT 838.220 31.290 838.480 31.610 ;
        RECT 1114.680 31.290 1114.940 31.610 ;
        RECT 1114.740 2.400 1114.880 31.290 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 134.540 827.930 134.600 ;
        RECT 1131.670 134.540 1131.990 134.600 ;
        RECT 827.610 134.400 1131.990 134.540 ;
        RECT 827.610 134.340 827.930 134.400 ;
        RECT 1131.670 134.340 1131.990 134.400 ;
      LAYER via ;
        RECT 827.640 134.340 827.900 134.600 ;
        RECT 1131.700 134.340 1131.960 134.600 ;
      LAYER met2 ;
        RECT 824.830 260.170 825.110 264.000 ;
        RECT 824.830 260.030 827.840 260.170 ;
        RECT 824.830 260.000 825.110 260.030 ;
        RECT 827.700 134.630 827.840 260.030 ;
        RECT 827.640 134.310 827.900 134.630 ;
        RECT 1131.700 134.310 1131.960 134.630 ;
        RECT 1131.760 16.730 1131.900 134.310 ;
        RECT 1131.760 16.590 1132.820 16.730 ;
        RECT 1132.680 2.400 1132.820 16.590 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 842.790 244.020 843.110 244.080 ;
        RECT 848.310 244.020 848.630 244.080 ;
        RECT 842.790 243.880 848.630 244.020 ;
        RECT 842.790 243.820 843.110 243.880 ;
        RECT 848.310 243.820 848.630 243.880 ;
        RECT 848.310 37.980 848.630 38.040 ;
        RECT 1150.530 37.980 1150.850 38.040 ;
        RECT 848.310 37.840 1150.850 37.980 ;
        RECT 848.310 37.780 848.630 37.840 ;
        RECT 1150.530 37.780 1150.850 37.840 ;
      LAYER via ;
        RECT 842.820 243.820 843.080 244.080 ;
        RECT 848.340 243.820 848.600 244.080 ;
        RECT 848.340 37.780 848.600 38.040 ;
        RECT 1150.560 37.780 1150.820 38.040 ;
      LAYER met2 ;
        RECT 842.770 260.000 843.050 264.000 ;
        RECT 842.880 244.110 843.020 260.000 ;
        RECT 842.820 243.790 843.080 244.110 ;
        RECT 848.340 243.790 848.600 244.110 ;
        RECT 848.400 38.070 848.540 243.790 ;
        RECT 848.340 37.750 848.600 38.070 ;
        RECT 1150.560 37.750 1150.820 38.070 ;
        RECT 1150.620 2.400 1150.760 37.750 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 360.250 244.020 360.570 244.080 ;
        RECT 365.310 244.020 365.630 244.080 ;
        RECT 360.250 243.880 365.630 244.020 ;
        RECT 360.250 243.820 360.570 243.880 ;
        RECT 365.310 243.820 365.630 243.880 ;
        RECT 365.310 93.060 365.630 93.120 ;
        RECT 662.930 93.060 663.250 93.120 ;
        RECT 365.310 92.920 663.250 93.060 ;
        RECT 365.310 92.860 365.630 92.920 ;
        RECT 662.930 92.860 663.250 92.920 ;
        RECT 662.930 17.580 663.250 17.640 ;
        RECT 668.910 17.580 669.230 17.640 ;
        RECT 662.930 17.440 669.230 17.580 ;
        RECT 662.930 17.380 663.250 17.440 ;
        RECT 668.910 17.380 669.230 17.440 ;
      LAYER via ;
        RECT 360.280 243.820 360.540 244.080 ;
        RECT 365.340 243.820 365.600 244.080 ;
        RECT 365.340 92.860 365.600 93.120 ;
        RECT 662.960 92.860 663.220 93.120 ;
        RECT 662.960 17.380 663.220 17.640 ;
        RECT 668.940 17.380 669.200 17.640 ;
      LAYER met2 ;
        RECT 360.230 260.000 360.510 264.000 ;
        RECT 360.340 244.110 360.480 260.000 ;
        RECT 360.280 243.790 360.540 244.110 ;
        RECT 365.340 243.790 365.600 244.110 ;
        RECT 365.400 93.150 365.540 243.790 ;
        RECT 365.340 92.830 365.600 93.150 ;
        RECT 662.960 92.830 663.220 93.150 ;
        RECT 663.020 17.670 663.160 92.830 ;
        RECT 662.960 17.350 663.220 17.670 ;
        RECT 668.940 17.350 669.200 17.670 ;
        RECT 669.000 2.400 669.140 17.350 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 44.780 862.430 44.840 ;
        RECT 1168.470 44.780 1168.790 44.840 ;
        RECT 862.110 44.640 1168.790 44.780 ;
        RECT 862.110 44.580 862.430 44.640 ;
        RECT 1168.470 44.580 1168.790 44.640 ;
      LAYER via ;
        RECT 862.140 44.580 862.400 44.840 ;
        RECT 1168.500 44.580 1168.760 44.840 ;
      LAYER met2 ;
        RECT 860.710 260.170 860.990 264.000 ;
        RECT 860.710 260.030 862.340 260.170 ;
        RECT 860.710 260.000 860.990 260.030 ;
        RECT 862.200 44.870 862.340 260.030 ;
        RECT 862.140 44.550 862.400 44.870 ;
        RECT 1168.500 44.550 1168.760 44.870 ;
        RECT 1168.560 2.400 1168.700 44.550 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 878.670 243.000 878.990 243.060 ;
        RECT 882.810 243.000 883.130 243.060 ;
        RECT 878.670 242.860 883.130 243.000 ;
        RECT 878.670 242.800 878.990 242.860 ;
        RECT 882.810 242.800 883.130 242.860 ;
        RECT 882.810 51.920 883.130 51.980 ;
        RECT 1180.430 51.920 1180.750 51.980 ;
        RECT 882.810 51.780 1180.750 51.920 ;
        RECT 882.810 51.720 883.130 51.780 ;
        RECT 1180.430 51.720 1180.750 51.780 ;
      LAYER via ;
        RECT 878.700 242.800 878.960 243.060 ;
        RECT 882.840 242.800 883.100 243.060 ;
        RECT 882.840 51.720 883.100 51.980 ;
        RECT 1180.460 51.720 1180.720 51.980 ;
      LAYER met2 ;
        RECT 878.650 260.000 878.930 264.000 ;
        RECT 878.760 243.090 878.900 260.000 ;
        RECT 878.700 242.770 878.960 243.090 ;
        RECT 882.840 242.770 883.100 243.090 ;
        RECT 882.900 52.010 883.040 242.770 ;
        RECT 882.840 51.690 883.100 52.010 ;
        RECT 1180.460 51.690 1180.720 52.010 ;
        RECT 1180.520 17.410 1180.660 51.690 ;
        RECT 1180.520 17.270 1186.180 17.410 ;
        RECT 1186.040 2.400 1186.180 17.270 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.150 58.720 896.470 58.780 ;
        RECT 1200.670 58.720 1200.990 58.780 ;
        RECT 896.150 58.580 1200.990 58.720 ;
        RECT 896.150 58.520 896.470 58.580 ;
        RECT 1200.670 58.520 1200.990 58.580 ;
      LAYER via ;
        RECT 896.180 58.520 896.440 58.780 ;
        RECT 1200.700 58.520 1200.960 58.780 ;
      LAYER met2 ;
        RECT 896.590 260.170 896.870 264.000 ;
        RECT 896.240 260.030 896.870 260.170 ;
        RECT 896.240 58.810 896.380 260.030 ;
        RECT 896.590 260.000 896.870 260.030 ;
        RECT 896.180 58.490 896.440 58.810 ;
        RECT 1200.700 58.490 1200.960 58.810 ;
        RECT 1200.760 16.730 1200.900 58.490 ;
        RECT 1200.760 16.590 1204.120 16.730 ;
        RECT 1203.980 2.400 1204.120 16.590 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 65.520 917.630 65.580 ;
        RECT 1221.830 65.520 1222.150 65.580 ;
        RECT 917.310 65.380 1222.150 65.520 ;
        RECT 917.310 65.320 917.630 65.380 ;
        RECT 1221.830 65.320 1222.150 65.380 ;
      LAYER via ;
        RECT 917.340 65.320 917.600 65.580 ;
        RECT 1221.860 65.320 1222.120 65.580 ;
      LAYER met2 ;
        RECT 914.530 260.170 914.810 264.000 ;
        RECT 914.530 260.030 917.540 260.170 ;
        RECT 914.530 260.000 914.810 260.030 ;
        RECT 917.400 65.610 917.540 260.030 ;
        RECT 917.340 65.290 917.600 65.610 ;
        RECT 1221.860 65.290 1222.120 65.610 ;
        RECT 1221.920 2.400 1222.060 65.290 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 932.490 244.020 932.810 244.080 ;
        RECT 938.010 244.020 938.330 244.080 ;
        RECT 932.490 243.880 938.330 244.020 ;
        RECT 932.490 243.820 932.810 243.880 ;
        RECT 938.010 243.820 938.330 243.880 ;
        RECT 938.010 72.660 938.330 72.720 ;
        RECT 1235.170 72.660 1235.490 72.720 ;
        RECT 938.010 72.520 1235.490 72.660 ;
        RECT 938.010 72.460 938.330 72.520 ;
        RECT 1235.170 72.460 1235.490 72.520 ;
        RECT 1235.170 62.120 1235.490 62.180 ;
        RECT 1239.770 62.120 1240.090 62.180 ;
        RECT 1235.170 61.980 1240.090 62.120 ;
        RECT 1235.170 61.920 1235.490 61.980 ;
        RECT 1239.770 61.920 1240.090 61.980 ;
      LAYER via ;
        RECT 932.520 243.820 932.780 244.080 ;
        RECT 938.040 243.820 938.300 244.080 ;
        RECT 938.040 72.460 938.300 72.720 ;
        RECT 1235.200 72.460 1235.460 72.720 ;
        RECT 1235.200 61.920 1235.460 62.180 ;
        RECT 1239.800 61.920 1240.060 62.180 ;
      LAYER met2 ;
        RECT 932.470 260.000 932.750 264.000 ;
        RECT 932.580 244.110 932.720 260.000 ;
        RECT 932.520 243.790 932.780 244.110 ;
        RECT 938.040 243.790 938.300 244.110 ;
        RECT 938.100 72.750 938.240 243.790 ;
        RECT 938.040 72.430 938.300 72.750 ;
        RECT 1235.200 72.430 1235.460 72.750 ;
        RECT 1235.260 62.210 1235.400 72.430 ;
        RECT 1235.200 61.890 1235.460 62.210 ;
        RECT 1239.800 61.890 1240.060 62.210 ;
        RECT 1239.860 2.400 1240.000 61.890 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 24.040 952.130 24.100 ;
        RECT 1257.250 24.040 1257.570 24.100 ;
        RECT 951.810 23.900 1257.570 24.040 ;
        RECT 951.810 23.840 952.130 23.900 ;
        RECT 1257.250 23.840 1257.570 23.900 ;
      LAYER via ;
        RECT 951.840 23.840 952.100 24.100 ;
        RECT 1257.280 23.840 1257.540 24.100 ;
      LAYER met2 ;
        RECT 950.410 260.170 950.690 264.000 ;
        RECT 950.410 260.030 952.040 260.170 ;
        RECT 950.410 260.000 950.690 260.030 ;
        RECT 951.900 24.130 952.040 260.030 ;
        RECT 951.840 23.810 952.100 24.130 ;
        RECT 1257.280 23.810 1257.540 24.130 ;
        RECT 1257.340 2.400 1257.480 23.810 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 967.910 244.020 968.230 244.080 ;
        RECT 972.510 244.020 972.830 244.080 ;
        RECT 967.910 243.880 972.830 244.020 ;
        RECT 967.910 243.820 968.230 243.880 ;
        RECT 972.510 243.820 972.830 243.880 ;
        RECT 972.510 79.460 972.830 79.520 ;
        RECT 1269.670 79.460 1269.990 79.520 ;
        RECT 972.510 79.320 1269.990 79.460 ;
        RECT 972.510 79.260 972.830 79.320 ;
        RECT 1269.670 79.260 1269.990 79.320 ;
        RECT 1269.670 62.120 1269.990 62.180 ;
        RECT 1275.190 62.120 1275.510 62.180 ;
        RECT 1269.670 61.980 1275.510 62.120 ;
        RECT 1269.670 61.920 1269.990 61.980 ;
        RECT 1275.190 61.920 1275.510 61.980 ;
      LAYER via ;
        RECT 967.940 243.820 968.200 244.080 ;
        RECT 972.540 243.820 972.800 244.080 ;
        RECT 972.540 79.260 972.800 79.520 ;
        RECT 1269.700 79.260 1269.960 79.520 ;
        RECT 1269.700 61.920 1269.960 62.180 ;
        RECT 1275.220 61.920 1275.480 62.180 ;
      LAYER met2 ;
        RECT 967.890 260.000 968.170 264.000 ;
        RECT 968.000 244.110 968.140 260.000 ;
        RECT 967.940 243.790 968.200 244.110 ;
        RECT 972.540 243.790 972.800 244.110 ;
        RECT 972.600 79.550 972.740 243.790 ;
        RECT 972.540 79.230 972.800 79.550 ;
        RECT 1269.700 79.230 1269.960 79.550 ;
        RECT 1269.760 62.210 1269.900 79.230 ;
        RECT 1269.700 61.890 1269.960 62.210 ;
        RECT 1275.220 61.890 1275.480 62.210 ;
        RECT 1275.280 2.400 1275.420 61.890 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 985.850 86.260 986.170 86.320 ;
        RECT 1290.370 86.260 1290.690 86.320 ;
        RECT 985.850 86.120 1290.690 86.260 ;
        RECT 985.850 86.060 986.170 86.120 ;
        RECT 1290.370 86.060 1290.690 86.120 ;
        RECT 1290.370 62.120 1290.690 62.180 ;
        RECT 1293.130 62.120 1293.450 62.180 ;
        RECT 1290.370 61.980 1293.450 62.120 ;
        RECT 1290.370 61.920 1290.690 61.980 ;
        RECT 1293.130 61.920 1293.450 61.980 ;
      LAYER via ;
        RECT 985.880 86.060 986.140 86.320 ;
        RECT 1290.400 86.060 1290.660 86.320 ;
        RECT 1290.400 61.920 1290.660 62.180 ;
        RECT 1293.160 61.920 1293.420 62.180 ;
      LAYER met2 ;
        RECT 985.830 260.000 986.110 264.000 ;
        RECT 985.940 86.350 986.080 260.000 ;
        RECT 985.880 86.030 986.140 86.350 ;
        RECT 1290.400 86.030 1290.660 86.350 ;
        RECT 1290.460 62.210 1290.600 86.030 ;
        RECT 1290.400 61.890 1290.660 62.210 ;
        RECT 1293.160 61.890 1293.420 62.210 ;
        RECT 1293.220 2.400 1293.360 61.890 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 93.400 1007.330 93.460 ;
        RECT 1311.530 93.400 1311.850 93.460 ;
        RECT 1007.010 93.260 1311.850 93.400 ;
        RECT 1007.010 93.200 1007.330 93.260 ;
        RECT 1311.530 93.200 1311.850 93.260 ;
      LAYER via ;
        RECT 1007.040 93.200 1007.300 93.460 ;
        RECT 1311.560 93.200 1311.820 93.460 ;
      LAYER met2 ;
        RECT 1003.770 260.170 1004.050 264.000 ;
        RECT 1003.770 260.030 1007.240 260.170 ;
        RECT 1003.770 260.000 1004.050 260.030 ;
        RECT 1007.100 93.490 1007.240 260.030 ;
        RECT 1007.040 93.170 1007.300 93.490 ;
        RECT 1311.560 93.170 1311.820 93.490 ;
        RECT 1311.620 37.130 1311.760 93.170 ;
        RECT 1311.160 36.990 1311.760 37.130 ;
        RECT 1311.160 2.400 1311.300 36.990 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.730 244.020 1022.050 244.080 ;
        RECT 1027.710 244.020 1028.030 244.080 ;
        RECT 1021.730 243.880 1028.030 244.020 ;
        RECT 1021.730 243.820 1022.050 243.880 ;
        RECT 1027.710 243.820 1028.030 243.880 ;
        RECT 1027.710 99.860 1028.030 99.920 ;
        RECT 1324.870 99.860 1325.190 99.920 ;
        RECT 1027.710 99.720 1325.190 99.860 ;
        RECT 1027.710 99.660 1028.030 99.720 ;
        RECT 1324.870 99.660 1325.190 99.720 ;
        RECT 1324.870 62.120 1325.190 62.180 ;
        RECT 1329.010 62.120 1329.330 62.180 ;
        RECT 1324.870 61.980 1329.330 62.120 ;
        RECT 1324.870 61.920 1325.190 61.980 ;
        RECT 1329.010 61.920 1329.330 61.980 ;
      LAYER via ;
        RECT 1021.760 243.820 1022.020 244.080 ;
        RECT 1027.740 243.820 1028.000 244.080 ;
        RECT 1027.740 99.660 1028.000 99.920 ;
        RECT 1324.900 99.660 1325.160 99.920 ;
        RECT 1324.900 61.920 1325.160 62.180 ;
        RECT 1329.040 61.920 1329.300 62.180 ;
      LAYER met2 ;
        RECT 1021.710 260.000 1021.990 264.000 ;
        RECT 1021.820 244.110 1021.960 260.000 ;
        RECT 1021.760 243.790 1022.020 244.110 ;
        RECT 1027.740 243.790 1028.000 244.110 ;
        RECT 1027.800 99.950 1027.940 243.790 ;
        RECT 1027.740 99.630 1028.000 99.950 ;
        RECT 1324.900 99.630 1325.160 99.950 ;
        RECT 1324.960 62.210 1325.100 99.630 ;
        RECT 1324.900 61.890 1325.160 62.210 ;
        RECT 1329.040 61.890 1329.300 62.210 ;
        RECT 1329.100 2.400 1329.240 61.890 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 379.110 99.860 379.430 99.920 ;
        RECT 683.170 99.860 683.490 99.920 ;
        RECT 379.110 99.720 683.490 99.860 ;
        RECT 379.110 99.660 379.430 99.720 ;
        RECT 683.170 99.660 683.490 99.720 ;
      LAYER via ;
        RECT 379.140 99.660 379.400 99.920 ;
        RECT 683.200 99.660 683.460 99.920 ;
      LAYER met2 ;
        RECT 378.170 260.170 378.450 264.000 ;
        RECT 378.170 260.030 379.340 260.170 ;
        RECT 378.170 260.000 378.450 260.030 ;
        RECT 379.200 99.950 379.340 260.030 ;
        RECT 379.140 99.630 379.400 99.950 ;
        RECT 683.200 99.630 683.460 99.950 ;
        RECT 683.260 16.730 683.400 99.630 ;
        RECT 683.260 16.590 686.620 16.730 ;
        RECT 686.480 2.400 686.620 16.590 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1345.645 48.365 1345.815 96.475 ;
      LAYER mcon ;
        RECT 1345.645 96.305 1345.815 96.475 ;
      LAYER met1 ;
        RECT 1041.510 141.340 1041.830 141.400 ;
        RECT 1345.570 141.340 1345.890 141.400 ;
        RECT 1041.510 141.200 1345.890 141.340 ;
        RECT 1041.510 141.140 1041.830 141.200 ;
        RECT 1345.570 141.140 1345.890 141.200 ;
        RECT 1345.570 96.460 1345.890 96.520 ;
        RECT 1345.375 96.320 1345.890 96.460 ;
        RECT 1345.570 96.260 1345.890 96.320 ;
        RECT 1345.585 48.520 1345.875 48.565 ;
        RECT 1346.490 48.520 1346.810 48.580 ;
        RECT 1345.585 48.380 1346.810 48.520 ;
        RECT 1345.585 48.335 1345.875 48.380 ;
        RECT 1346.490 48.320 1346.810 48.380 ;
      LAYER via ;
        RECT 1041.540 141.140 1041.800 141.400 ;
        RECT 1345.600 141.140 1345.860 141.400 ;
        RECT 1345.600 96.260 1345.860 96.520 ;
        RECT 1346.520 48.320 1346.780 48.580 ;
      LAYER met2 ;
        RECT 1039.650 260.170 1039.930 264.000 ;
        RECT 1039.650 260.030 1041.740 260.170 ;
        RECT 1039.650 260.000 1039.930 260.030 ;
        RECT 1041.600 141.430 1041.740 260.030 ;
        RECT 1041.540 141.110 1041.800 141.430 ;
        RECT 1345.600 141.110 1345.860 141.430 ;
        RECT 1345.660 96.550 1345.800 141.110 ;
        RECT 1345.600 96.230 1345.860 96.550 ;
        RECT 1346.520 48.290 1346.780 48.610 ;
        RECT 1346.580 2.400 1346.720 48.290 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1057.610 241.640 1057.930 241.700 ;
        RECT 1062.210 241.640 1062.530 241.700 ;
        RECT 1057.610 241.500 1062.530 241.640 ;
        RECT 1057.610 241.440 1057.930 241.500 ;
        RECT 1062.210 241.440 1062.530 241.500 ;
        RECT 1062.210 107.000 1062.530 107.060 ;
        RECT 1359.370 107.000 1359.690 107.060 ;
        RECT 1062.210 106.860 1359.690 107.000 ;
        RECT 1062.210 106.800 1062.530 106.860 ;
        RECT 1359.370 106.800 1359.690 106.860 ;
        RECT 1359.370 62.120 1359.690 62.180 ;
        RECT 1364.430 62.120 1364.750 62.180 ;
        RECT 1359.370 61.980 1364.750 62.120 ;
        RECT 1359.370 61.920 1359.690 61.980 ;
        RECT 1364.430 61.920 1364.750 61.980 ;
      LAYER via ;
        RECT 1057.640 241.440 1057.900 241.700 ;
        RECT 1062.240 241.440 1062.500 241.700 ;
        RECT 1062.240 106.800 1062.500 107.060 ;
        RECT 1359.400 106.800 1359.660 107.060 ;
        RECT 1359.400 61.920 1359.660 62.180 ;
        RECT 1364.460 61.920 1364.720 62.180 ;
      LAYER met2 ;
        RECT 1057.590 260.000 1057.870 264.000 ;
        RECT 1057.700 241.730 1057.840 260.000 ;
        RECT 1057.640 241.410 1057.900 241.730 ;
        RECT 1062.240 241.410 1062.500 241.730 ;
        RECT 1062.300 107.090 1062.440 241.410 ;
        RECT 1062.240 106.770 1062.500 107.090 ;
        RECT 1359.400 106.770 1359.660 107.090 ;
        RECT 1359.460 62.210 1359.600 106.770 ;
        RECT 1359.400 61.890 1359.660 62.210 ;
        RECT 1364.460 61.890 1364.720 62.210 ;
        RECT 1364.520 2.400 1364.660 61.890 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1075.550 113.800 1075.870 113.860 ;
        RECT 1380.070 113.800 1380.390 113.860 ;
        RECT 1075.550 113.660 1380.390 113.800 ;
        RECT 1075.550 113.600 1075.870 113.660 ;
        RECT 1380.070 113.600 1380.390 113.660 ;
        RECT 1380.070 62.260 1380.390 62.520 ;
        RECT 1380.160 61.780 1380.300 62.260 ;
        RECT 1382.370 61.780 1382.690 61.840 ;
        RECT 1380.160 61.640 1382.690 61.780 ;
        RECT 1382.370 61.580 1382.690 61.640 ;
        RECT 1382.370 47.980 1382.690 48.240 ;
        RECT 1382.460 47.560 1382.600 47.980 ;
        RECT 1382.370 47.300 1382.690 47.560 ;
      LAYER via ;
        RECT 1075.580 113.600 1075.840 113.860 ;
        RECT 1380.100 113.600 1380.360 113.860 ;
        RECT 1380.100 62.260 1380.360 62.520 ;
        RECT 1382.400 61.580 1382.660 61.840 ;
        RECT 1382.400 47.980 1382.660 48.240 ;
        RECT 1382.400 47.300 1382.660 47.560 ;
      LAYER met2 ;
        RECT 1075.530 260.000 1075.810 264.000 ;
        RECT 1075.640 113.890 1075.780 260.000 ;
        RECT 1075.580 113.570 1075.840 113.890 ;
        RECT 1380.100 113.570 1380.360 113.890 ;
        RECT 1380.160 62.550 1380.300 113.570 ;
        RECT 1380.100 62.230 1380.360 62.550 ;
        RECT 1382.400 61.550 1382.660 61.870 ;
        RECT 1382.460 48.270 1382.600 61.550 ;
        RECT 1382.400 47.950 1382.660 48.270 ;
        RECT 1382.400 47.270 1382.660 47.590 ;
        RECT 1382.460 2.400 1382.600 47.270 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1093.030 244.020 1093.350 244.080 ;
        RECT 1096.710 244.020 1097.030 244.080 ;
        RECT 1093.030 243.880 1097.030 244.020 ;
        RECT 1093.030 243.820 1093.350 243.880 ;
        RECT 1096.710 243.820 1097.030 243.880 ;
        RECT 1096.710 31.180 1097.030 31.240 ;
        RECT 1399.850 31.180 1400.170 31.240 ;
        RECT 1096.710 31.040 1400.170 31.180 ;
        RECT 1096.710 30.980 1097.030 31.040 ;
        RECT 1399.850 30.980 1400.170 31.040 ;
      LAYER via ;
        RECT 1093.060 243.820 1093.320 244.080 ;
        RECT 1096.740 243.820 1097.000 244.080 ;
        RECT 1096.740 30.980 1097.000 31.240 ;
        RECT 1399.880 30.980 1400.140 31.240 ;
      LAYER met2 ;
        RECT 1093.010 260.000 1093.290 264.000 ;
        RECT 1093.120 244.110 1093.260 260.000 ;
        RECT 1093.060 243.790 1093.320 244.110 ;
        RECT 1096.740 243.790 1097.000 244.110 ;
        RECT 1096.800 31.270 1096.940 243.790 ;
        RECT 1096.740 30.950 1097.000 31.270 ;
        RECT 1399.880 30.950 1400.140 31.270 ;
        RECT 1399.940 30.330 1400.080 30.950 ;
        RECT 1399.940 30.190 1400.540 30.330 ;
        RECT 1400.400 2.400 1400.540 30.190 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.970 244.020 1111.290 244.080 ;
        RECT 1117.410 244.020 1117.730 244.080 ;
        RECT 1110.970 243.880 1117.730 244.020 ;
        RECT 1110.970 243.820 1111.290 243.880 ;
        RECT 1117.410 243.820 1117.730 243.880 ;
        RECT 1117.410 38.320 1117.730 38.380 ;
        RECT 1418.250 38.320 1418.570 38.380 ;
        RECT 1117.410 38.180 1418.570 38.320 ;
        RECT 1117.410 38.120 1117.730 38.180 ;
        RECT 1418.250 38.120 1418.570 38.180 ;
      LAYER via ;
        RECT 1111.000 243.820 1111.260 244.080 ;
        RECT 1117.440 243.820 1117.700 244.080 ;
        RECT 1117.440 38.120 1117.700 38.380 ;
        RECT 1418.280 38.120 1418.540 38.380 ;
      LAYER met2 ;
        RECT 1110.950 260.000 1111.230 264.000 ;
        RECT 1111.060 244.110 1111.200 260.000 ;
        RECT 1111.000 243.790 1111.260 244.110 ;
        RECT 1117.440 243.790 1117.700 244.110 ;
        RECT 1117.500 38.410 1117.640 243.790 ;
        RECT 1117.440 38.090 1117.700 38.410 ;
        RECT 1418.280 38.090 1418.540 38.410 ;
        RECT 1418.340 2.400 1418.480 38.090 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 120.600 1131.530 120.660 ;
        RECT 1435.730 120.600 1436.050 120.660 ;
        RECT 1131.210 120.460 1436.050 120.600 ;
        RECT 1131.210 120.400 1131.530 120.460 ;
        RECT 1435.730 120.400 1436.050 120.460 ;
      LAYER via ;
        RECT 1131.240 120.400 1131.500 120.660 ;
        RECT 1435.760 120.400 1436.020 120.660 ;
      LAYER met2 ;
        RECT 1128.890 260.170 1129.170 264.000 ;
        RECT 1128.890 260.030 1131.440 260.170 ;
        RECT 1128.890 260.000 1129.170 260.030 ;
        RECT 1131.300 120.690 1131.440 260.030 ;
        RECT 1131.240 120.370 1131.500 120.690 ;
        RECT 1435.760 120.370 1436.020 120.690 ;
        RECT 1435.820 2.400 1435.960 120.370 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1146.850 244.020 1147.170 244.080 ;
        RECT 1151.910 244.020 1152.230 244.080 ;
        RECT 1146.850 243.880 1152.230 244.020 ;
        RECT 1146.850 243.820 1147.170 243.880 ;
        RECT 1151.910 243.820 1152.230 243.880 ;
        RECT 1151.910 45.460 1152.230 45.520 ;
        RECT 1453.670 45.460 1453.990 45.520 ;
        RECT 1151.910 45.320 1453.990 45.460 ;
        RECT 1151.910 45.260 1152.230 45.320 ;
        RECT 1453.670 45.260 1453.990 45.320 ;
      LAYER via ;
        RECT 1146.880 243.820 1147.140 244.080 ;
        RECT 1151.940 243.820 1152.200 244.080 ;
        RECT 1151.940 45.260 1152.200 45.520 ;
        RECT 1453.700 45.260 1453.960 45.520 ;
      LAYER met2 ;
        RECT 1146.830 260.000 1147.110 264.000 ;
        RECT 1146.940 244.110 1147.080 260.000 ;
        RECT 1146.880 243.790 1147.140 244.110 ;
        RECT 1151.940 243.790 1152.200 244.110 ;
        RECT 1152.000 45.550 1152.140 243.790 ;
        RECT 1151.940 45.230 1152.200 45.550 ;
        RECT 1453.700 45.230 1453.960 45.550 ;
        RECT 1453.760 2.400 1453.900 45.230 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 51.580 1166.030 51.640 ;
        RECT 1471.610 51.580 1471.930 51.640 ;
        RECT 1165.710 51.440 1471.930 51.580 ;
        RECT 1165.710 51.380 1166.030 51.440 ;
        RECT 1471.610 51.380 1471.930 51.440 ;
      LAYER via ;
        RECT 1165.740 51.380 1166.000 51.640 ;
        RECT 1471.640 51.380 1471.900 51.640 ;
      LAYER met2 ;
        RECT 1164.770 260.170 1165.050 264.000 ;
        RECT 1164.770 260.030 1165.940 260.170 ;
        RECT 1164.770 260.000 1165.050 260.030 ;
        RECT 1165.800 51.670 1165.940 260.030 ;
        RECT 1165.740 51.350 1166.000 51.670 ;
        RECT 1471.640 51.350 1471.900 51.670 ;
        RECT 1471.700 2.400 1471.840 51.350 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 59.060 1186.730 59.120 ;
        RECT 1489.550 59.060 1489.870 59.120 ;
        RECT 1186.410 58.920 1489.870 59.060 ;
        RECT 1186.410 58.860 1186.730 58.920 ;
        RECT 1489.550 58.860 1489.870 58.920 ;
      LAYER via ;
        RECT 1186.440 58.860 1186.700 59.120 ;
        RECT 1489.580 58.860 1489.840 59.120 ;
      LAYER met2 ;
        RECT 1182.710 260.170 1182.990 264.000 ;
        RECT 1182.710 260.030 1186.640 260.170 ;
        RECT 1182.710 260.000 1182.990 260.030 ;
        RECT 1186.500 59.150 1186.640 260.030 ;
        RECT 1186.440 58.830 1186.700 59.150 ;
        RECT 1489.580 58.830 1489.840 59.150 ;
        RECT 1489.640 2.400 1489.780 58.830 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1507.105 48.365 1507.275 65.875 ;
      LAYER mcon ;
        RECT 1507.105 65.705 1507.275 65.875 ;
      LAYER met1 ;
        RECT 1200.670 244.020 1200.990 244.080 ;
        RECT 1207.110 244.020 1207.430 244.080 ;
        RECT 1200.670 243.880 1207.430 244.020 ;
        RECT 1200.670 243.820 1200.990 243.880 ;
        RECT 1207.110 243.820 1207.430 243.880 ;
        RECT 1207.110 65.860 1207.430 65.920 ;
        RECT 1507.045 65.860 1507.335 65.905 ;
        RECT 1207.110 65.720 1507.335 65.860 ;
        RECT 1207.110 65.660 1207.430 65.720 ;
        RECT 1507.045 65.675 1507.335 65.720 ;
        RECT 1507.030 48.520 1507.350 48.580 ;
        RECT 1506.835 48.380 1507.350 48.520 ;
        RECT 1507.030 48.320 1507.350 48.380 ;
        RECT 1506.570 2.960 1506.890 3.020 ;
        RECT 1507.030 2.960 1507.350 3.020 ;
        RECT 1506.570 2.820 1507.350 2.960 ;
        RECT 1506.570 2.760 1506.890 2.820 ;
        RECT 1507.030 2.760 1507.350 2.820 ;
      LAYER via ;
        RECT 1200.700 243.820 1200.960 244.080 ;
        RECT 1207.140 243.820 1207.400 244.080 ;
        RECT 1207.140 65.660 1207.400 65.920 ;
        RECT 1507.060 48.320 1507.320 48.580 ;
        RECT 1506.600 2.760 1506.860 3.020 ;
        RECT 1507.060 2.760 1507.320 3.020 ;
      LAYER met2 ;
        RECT 1200.650 260.000 1200.930 264.000 ;
        RECT 1200.760 244.110 1200.900 260.000 ;
        RECT 1200.700 243.790 1200.960 244.110 ;
        RECT 1207.140 243.790 1207.400 244.110 ;
        RECT 1207.200 65.950 1207.340 243.790 ;
        RECT 1207.140 65.630 1207.400 65.950 ;
        RECT 1507.060 48.290 1507.320 48.610 ;
        RECT 1507.120 48.010 1507.260 48.290 ;
        RECT 1506.660 47.870 1507.260 48.010 ;
        RECT 1506.660 3.050 1506.800 47.870 ;
        RECT 1506.600 2.730 1506.860 3.050 ;
        RECT 1507.060 2.730 1507.320 3.050 ;
        RECT 1507.120 2.400 1507.260 2.730 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 399.810 107.000 400.130 107.060 ;
        RECT 704.330 107.000 704.650 107.060 ;
        RECT 399.810 106.860 704.650 107.000 ;
        RECT 399.810 106.800 400.130 106.860 ;
        RECT 704.330 106.800 704.650 106.860 ;
      LAYER via ;
        RECT 399.840 106.800 400.100 107.060 ;
        RECT 704.360 106.800 704.620 107.060 ;
      LAYER met2 ;
        RECT 396.110 260.170 396.390 264.000 ;
        RECT 396.110 260.030 400.040 260.170 ;
        RECT 396.110 260.000 396.390 260.030 ;
        RECT 399.900 107.090 400.040 260.030 ;
        RECT 399.840 106.770 400.100 107.090 ;
        RECT 704.360 106.770 704.620 107.090 ;
        RECT 704.420 2.400 704.560 106.770 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 72.320 1221.230 72.380 ;
        RECT 1525.430 72.320 1525.750 72.380 ;
        RECT 1220.910 72.180 1525.750 72.320 ;
        RECT 1220.910 72.120 1221.230 72.180 ;
        RECT 1525.430 72.120 1525.750 72.180 ;
      LAYER via ;
        RECT 1220.940 72.120 1221.200 72.380 ;
        RECT 1525.460 72.120 1525.720 72.380 ;
      LAYER met2 ;
        RECT 1218.130 260.170 1218.410 264.000 ;
        RECT 1218.130 260.030 1221.140 260.170 ;
        RECT 1218.130 260.000 1218.410 260.030 ;
        RECT 1221.000 72.410 1221.140 260.030 ;
        RECT 1220.940 72.090 1221.200 72.410 ;
        RECT 1525.460 72.090 1525.720 72.410 ;
        RECT 1525.520 7.210 1525.660 72.090 ;
        RECT 1525.060 7.070 1525.660 7.210 ;
        RECT 1525.060 2.400 1525.200 7.070 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1249.045 25.245 1249.215 26.095 ;
        RECT 1296.885 24.905 1297.055 26.095 ;
        RECT 1304.245 24.905 1304.415 25.755 ;
        RECT 1352.545 24.905 1352.715 25.755 ;
        RECT 1393.945 24.225 1394.115 25.755 ;
        RECT 1435.345 23.545 1435.515 24.395 ;
        RECT 1483.185 23.545 1483.355 25.075 ;
      LAYER mcon ;
        RECT 1249.045 25.925 1249.215 26.095 ;
        RECT 1296.885 25.925 1297.055 26.095 ;
        RECT 1304.245 25.585 1304.415 25.755 ;
        RECT 1352.545 25.585 1352.715 25.755 ;
        RECT 1393.945 25.585 1394.115 25.755 ;
        RECT 1483.185 24.905 1483.355 25.075 ;
        RECT 1435.345 24.225 1435.515 24.395 ;
      LAYER met1 ;
        RECT 1236.090 244.020 1236.410 244.080 ;
        RECT 1241.610 244.020 1241.930 244.080 ;
        RECT 1236.090 243.880 1241.930 244.020 ;
        RECT 1236.090 243.820 1236.410 243.880 ;
        RECT 1241.610 243.820 1241.930 243.880 ;
        RECT 1248.985 26.080 1249.275 26.125 ;
        RECT 1296.825 26.080 1297.115 26.125 ;
        RECT 1248.985 25.940 1297.115 26.080 ;
        RECT 1248.985 25.895 1249.275 25.940 ;
        RECT 1296.825 25.895 1297.115 25.940 ;
        RECT 1304.185 25.740 1304.475 25.785 ;
        RECT 1352.485 25.740 1352.775 25.785 ;
        RECT 1393.885 25.740 1394.175 25.785 ;
        RECT 1304.185 25.600 1312.220 25.740 ;
        RECT 1304.185 25.555 1304.475 25.600 ;
        RECT 1241.610 25.400 1241.930 25.460 ;
        RECT 1248.985 25.400 1249.275 25.445 ;
        RECT 1241.610 25.260 1249.275 25.400 ;
        RECT 1241.610 25.200 1241.930 25.260 ;
        RECT 1248.985 25.215 1249.275 25.260 ;
        RECT 1296.825 25.060 1297.115 25.105 ;
        RECT 1304.185 25.060 1304.475 25.105 ;
        RECT 1296.825 24.920 1304.475 25.060 ;
        RECT 1312.080 25.060 1312.220 25.600 ;
        RECT 1352.485 25.600 1394.175 25.740 ;
        RECT 1352.485 25.555 1352.775 25.600 ;
        RECT 1393.885 25.555 1394.175 25.600 ;
        RECT 1352.485 25.060 1352.775 25.105 ;
        RECT 1312.080 24.920 1352.775 25.060 ;
        RECT 1296.825 24.875 1297.115 24.920 ;
        RECT 1304.185 24.875 1304.475 24.920 ;
        RECT 1352.485 24.875 1352.775 24.920 ;
        RECT 1483.125 25.060 1483.415 25.105 ;
        RECT 1483.125 24.920 1490.240 25.060 ;
        RECT 1483.125 24.875 1483.415 24.920 ;
        RECT 1490.100 24.720 1490.240 24.920 ;
        RECT 1542.910 24.720 1543.230 24.780 ;
        RECT 1490.100 24.580 1543.230 24.720 ;
        RECT 1542.910 24.520 1543.230 24.580 ;
        RECT 1393.885 24.380 1394.175 24.425 ;
        RECT 1435.285 24.380 1435.575 24.425 ;
        RECT 1393.885 24.240 1435.575 24.380 ;
        RECT 1393.885 24.195 1394.175 24.240 ;
        RECT 1435.285 24.195 1435.575 24.240 ;
        RECT 1435.285 23.700 1435.575 23.745 ;
        RECT 1483.125 23.700 1483.415 23.745 ;
        RECT 1435.285 23.560 1483.415 23.700 ;
        RECT 1435.285 23.515 1435.575 23.560 ;
        RECT 1483.125 23.515 1483.415 23.560 ;
      LAYER via ;
        RECT 1236.120 243.820 1236.380 244.080 ;
        RECT 1241.640 243.820 1241.900 244.080 ;
        RECT 1241.640 25.200 1241.900 25.460 ;
        RECT 1542.940 24.520 1543.200 24.780 ;
      LAYER met2 ;
        RECT 1236.070 260.000 1236.350 264.000 ;
        RECT 1236.180 244.110 1236.320 260.000 ;
        RECT 1236.120 243.790 1236.380 244.110 ;
        RECT 1241.640 243.790 1241.900 244.110 ;
        RECT 1241.700 25.490 1241.840 243.790 ;
        RECT 1241.640 25.170 1241.900 25.490 ;
        RECT 1542.940 24.490 1543.200 24.810 ;
        RECT 1543.000 2.400 1543.140 24.490 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 127.740 1255.730 127.800 ;
        RECT 1559.470 127.740 1559.790 127.800 ;
        RECT 1255.410 127.600 1559.790 127.740 ;
        RECT 1255.410 127.540 1255.730 127.600 ;
        RECT 1559.470 127.540 1559.790 127.600 ;
      LAYER via ;
        RECT 1255.440 127.540 1255.700 127.800 ;
        RECT 1559.500 127.540 1559.760 127.800 ;
      LAYER met2 ;
        RECT 1254.010 260.170 1254.290 264.000 ;
        RECT 1254.010 260.030 1255.640 260.170 ;
        RECT 1254.010 260.000 1254.290 260.030 ;
        RECT 1255.500 127.830 1255.640 260.030 ;
        RECT 1255.440 127.510 1255.700 127.830 ;
        RECT 1559.500 127.510 1559.760 127.830 ;
        RECT 1559.560 16.730 1559.700 127.510 ;
        RECT 1559.560 16.590 1561.080 16.730 ;
        RECT 1560.940 2.400 1561.080 16.590 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1271.970 244.020 1272.290 244.080 ;
        RECT 1276.110 244.020 1276.430 244.080 ;
        RECT 1271.970 243.880 1276.430 244.020 ;
        RECT 1271.970 243.820 1272.290 243.880 ;
        RECT 1276.110 243.820 1276.430 243.880 ;
        RECT 1276.110 79.800 1276.430 79.860 ;
        RECT 1573.270 79.800 1573.590 79.860 ;
        RECT 1276.110 79.660 1573.590 79.800 ;
        RECT 1276.110 79.600 1276.430 79.660 ;
        RECT 1573.270 79.600 1573.590 79.660 ;
      LAYER via ;
        RECT 1272.000 243.820 1272.260 244.080 ;
        RECT 1276.140 243.820 1276.400 244.080 ;
        RECT 1276.140 79.600 1276.400 79.860 ;
        RECT 1573.300 79.600 1573.560 79.860 ;
      LAYER met2 ;
        RECT 1271.950 260.000 1272.230 264.000 ;
        RECT 1272.060 244.110 1272.200 260.000 ;
        RECT 1272.000 243.790 1272.260 244.110 ;
        RECT 1276.140 243.790 1276.400 244.110 ;
        RECT 1276.200 79.890 1276.340 243.790 ;
        RECT 1276.140 79.570 1276.400 79.890 ;
        RECT 1573.300 79.570 1573.560 79.890 ;
        RECT 1573.360 16.730 1573.500 79.570 ;
        RECT 1573.360 16.590 1579.020 16.730 ;
        RECT 1578.880 2.400 1579.020 16.590 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.450 134.540 1289.770 134.600 ;
        RECT 1593.970 134.540 1594.290 134.600 ;
        RECT 1289.450 134.400 1594.290 134.540 ;
        RECT 1289.450 134.340 1289.770 134.400 ;
        RECT 1593.970 134.340 1594.290 134.400 ;
      LAYER via ;
        RECT 1289.480 134.340 1289.740 134.600 ;
        RECT 1594.000 134.340 1594.260 134.600 ;
      LAYER met2 ;
        RECT 1289.890 260.170 1290.170 264.000 ;
        RECT 1289.540 260.030 1290.170 260.170 ;
        RECT 1289.540 134.630 1289.680 260.030 ;
        RECT 1289.890 260.000 1290.170 260.030 ;
        RECT 1289.480 134.310 1289.740 134.630 ;
        RECT 1594.000 134.310 1594.260 134.630 ;
        RECT 1594.060 16.730 1594.200 134.310 ;
        RECT 1594.060 16.590 1596.500 16.730 ;
        RECT 1596.360 2.400 1596.500 16.590 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 86.260 1310.930 86.320 ;
        RECT 1608.230 86.260 1608.550 86.320 ;
        RECT 1310.610 86.120 1608.550 86.260 ;
        RECT 1310.610 86.060 1310.930 86.120 ;
        RECT 1608.230 86.060 1608.550 86.120 ;
        RECT 1608.230 17.920 1608.550 17.980 ;
        RECT 1614.210 17.920 1614.530 17.980 ;
        RECT 1608.230 17.780 1614.530 17.920 ;
        RECT 1608.230 17.720 1608.550 17.780 ;
        RECT 1614.210 17.720 1614.530 17.780 ;
      LAYER via ;
        RECT 1310.640 86.060 1310.900 86.320 ;
        RECT 1608.260 86.060 1608.520 86.320 ;
        RECT 1608.260 17.720 1608.520 17.980 ;
        RECT 1614.240 17.720 1614.500 17.980 ;
      LAYER met2 ;
        RECT 1307.830 260.170 1308.110 264.000 ;
        RECT 1307.830 260.030 1310.840 260.170 ;
        RECT 1307.830 260.000 1308.110 260.030 ;
        RECT 1310.700 86.350 1310.840 260.030 ;
        RECT 1310.640 86.030 1310.900 86.350 ;
        RECT 1608.260 86.030 1608.520 86.350 ;
        RECT 1608.320 18.010 1608.460 86.030 ;
        RECT 1608.260 17.690 1608.520 18.010 ;
        RECT 1614.240 17.690 1614.500 18.010 ;
        RECT 1614.300 2.400 1614.440 17.690 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1325.790 244.020 1326.110 244.080 ;
        RECT 1331.310 244.020 1331.630 244.080 ;
        RECT 1325.790 243.880 1331.630 244.020 ;
        RECT 1325.790 243.820 1326.110 243.880 ;
        RECT 1331.310 243.820 1331.630 243.880 ;
        RECT 1331.310 93.400 1331.630 93.460 ;
        RECT 1628.470 93.400 1628.790 93.460 ;
        RECT 1331.310 93.260 1628.790 93.400 ;
        RECT 1331.310 93.200 1331.630 93.260 ;
        RECT 1628.470 93.200 1628.790 93.260 ;
      LAYER via ;
        RECT 1325.820 243.820 1326.080 244.080 ;
        RECT 1331.340 243.820 1331.600 244.080 ;
        RECT 1331.340 93.200 1331.600 93.460 ;
        RECT 1628.500 93.200 1628.760 93.460 ;
      LAYER met2 ;
        RECT 1325.770 260.000 1326.050 264.000 ;
        RECT 1325.880 244.110 1326.020 260.000 ;
        RECT 1325.820 243.790 1326.080 244.110 ;
        RECT 1331.340 243.790 1331.600 244.110 ;
        RECT 1331.400 93.490 1331.540 243.790 ;
        RECT 1331.340 93.170 1331.600 93.490 ;
        RECT 1628.500 93.170 1628.760 93.490 ;
        RECT 1628.560 16.730 1628.700 93.170 ;
        RECT 1628.560 16.590 1632.380 16.730 ;
        RECT 1632.240 2.400 1632.380 16.590 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 99.860 1345.430 99.920 ;
        RECT 1649.170 99.860 1649.490 99.920 ;
        RECT 1345.110 99.720 1649.490 99.860 ;
        RECT 1345.110 99.660 1345.430 99.720 ;
        RECT 1649.170 99.660 1649.490 99.720 ;
      LAYER via ;
        RECT 1345.140 99.660 1345.400 99.920 ;
        RECT 1649.200 99.660 1649.460 99.920 ;
      LAYER met2 ;
        RECT 1343.250 260.170 1343.530 264.000 ;
        RECT 1343.250 260.030 1345.340 260.170 ;
        RECT 1343.250 260.000 1343.530 260.030 ;
        RECT 1345.200 99.950 1345.340 260.030 ;
        RECT 1345.140 99.630 1345.400 99.950 ;
        RECT 1649.200 99.630 1649.460 99.950 ;
        RECT 1649.260 16.730 1649.400 99.630 ;
        RECT 1649.260 16.590 1650.320 16.730 ;
        RECT 1650.180 2.400 1650.320 16.590 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.210 244.020 1361.530 244.080 ;
        RECT 1365.810 244.020 1366.130 244.080 ;
        RECT 1361.210 243.880 1366.130 244.020 ;
        RECT 1361.210 243.820 1361.530 243.880 ;
        RECT 1365.810 243.820 1366.130 243.880 ;
        RECT 1365.810 107.000 1366.130 107.060 ;
        RECT 1662.970 107.000 1663.290 107.060 ;
        RECT 1365.810 106.860 1663.290 107.000 ;
        RECT 1365.810 106.800 1366.130 106.860 ;
        RECT 1662.970 106.800 1663.290 106.860 ;
      LAYER via ;
        RECT 1361.240 243.820 1361.500 244.080 ;
        RECT 1365.840 243.820 1366.100 244.080 ;
        RECT 1365.840 106.800 1366.100 107.060 ;
        RECT 1663.000 106.800 1663.260 107.060 ;
      LAYER met2 ;
        RECT 1361.190 260.000 1361.470 264.000 ;
        RECT 1361.300 244.110 1361.440 260.000 ;
        RECT 1361.240 243.790 1361.500 244.110 ;
        RECT 1365.840 243.790 1366.100 244.110 ;
        RECT 1365.900 107.090 1366.040 243.790 ;
        RECT 1365.840 106.770 1366.100 107.090 ;
        RECT 1663.000 106.770 1663.260 107.090 ;
        RECT 1663.060 16.730 1663.200 106.770 ;
        RECT 1663.060 16.590 1668.260 16.730 ;
        RECT 1668.120 2.400 1668.260 16.590 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.150 238.240 1379.470 238.300 ;
        RECT 1683.670 238.240 1683.990 238.300 ;
        RECT 1379.150 238.100 1683.990 238.240 ;
        RECT 1379.150 238.040 1379.470 238.100 ;
        RECT 1683.670 238.040 1683.990 238.100 ;
      LAYER via ;
        RECT 1379.180 238.040 1379.440 238.300 ;
        RECT 1683.700 238.040 1683.960 238.300 ;
      LAYER met2 ;
        RECT 1379.130 260.000 1379.410 264.000 ;
        RECT 1379.240 238.330 1379.380 260.000 ;
        RECT 1379.180 238.010 1379.440 238.330 ;
        RECT 1683.700 238.010 1683.960 238.330 ;
        RECT 1683.760 16.730 1683.900 238.010 ;
        RECT 1683.760 16.590 1685.740 16.730 ;
        RECT 1685.600 2.400 1685.740 16.590 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 414.070 248.440 414.390 248.500 ;
        RECT 424.190 248.440 424.510 248.500 ;
        RECT 414.070 248.300 424.510 248.440 ;
        RECT 414.070 248.240 414.390 248.300 ;
        RECT 424.190 248.240 424.510 248.300 ;
        RECT 424.190 113.800 424.510 113.860 ;
        RECT 717.670 113.800 717.990 113.860 ;
        RECT 424.190 113.660 717.990 113.800 ;
        RECT 424.190 113.600 424.510 113.660 ;
        RECT 717.670 113.600 717.990 113.660 ;
      LAYER via ;
        RECT 414.100 248.240 414.360 248.500 ;
        RECT 424.220 248.240 424.480 248.500 ;
        RECT 424.220 113.600 424.480 113.860 ;
        RECT 717.700 113.600 717.960 113.860 ;
      LAYER met2 ;
        RECT 414.050 260.000 414.330 264.000 ;
        RECT 414.160 248.530 414.300 260.000 ;
        RECT 414.100 248.210 414.360 248.530 ;
        RECT 424.220 248.210 424.480 248.530 ;
        RECT 424.280 113.890 424.420 248.210 ;
        RECT 424.220 113.570 424.480 113.890 ;
        RECT 717.700 113.570 717.960 113.890 ;
        RECT 717.760 16.730 717.900 113.570 ;
        RECT 717.760 16.590 722.500 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 31.180 1400.630 31.240 ;
        RECT 1703.450 31.180 1703.770 31.240 ;
        RECT 1400.310 31.040 1703.770 31.180 ;
        RECT 1400.310 30.980 1400.630 31.040 ;
        RECT 1703.450 30.980 1703.770 31.040 ;
      LAYER via ;
        RECT 1400.340 30.980 1400.600 31.240 ;
        RECT 1703.480 30.980 1703.740 31.240 ;
      LAYER met2 ;
        RECT 1397.070 260.170 1397.350 264.000 ;
        RECT 1397.070 260.030 1400.540 260.170 ;
        RECT 1397.070 260.000 1397.350 260.030 ;
        RECT 1400.400 31.270 1400.540 260.030 ;
        RECT 1400.340 30.950 1400.600 31.270 ;
        RECT 1703.480 30.950 1703.740 31.270 ;
        RECT 1703.540 2.400 1703.680 30.950 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1415.030 244.020 1415.350 244.080 ;
        RECT 1421.010 244.020 1421.330 244.080 ;
        RECT 1415.030 243.880 1421.330 244.020 ;
        RECT 1415.030 243.820 1415.350 243.880 ;
        RECT 1421.010 243.820 1421.330 243.880 ;
        RECT 1421.010 39.000 1421.330 39.060 ;
        RECT 1421.010 38.860 1442.400 39.000 ;
        RECT 1421.010 38.800 1421.330 38.860 ;
        RECT 1442.260 38.320 1442.400 38.860 ;
        RECT 1721.390 38.320 1721.710 38.380 ;
        RECT 1442.260 38.180 1721.710 38.320 ;
        RECT 1721.390 38.120 1721.710 38.180 ;
      LAYER via ;
        RECT 1415.060 243.820 1415.320 244.080 ;
        RECT 1421.040 243.820 1421.300 244.080 ;
        RECT 1421.040 38.800 1421.300 39.060 ;
        RECT 1721.420 38.120 1721.680 38.380 ;
      LAYER met2 ;
        RECT 1415.010 260.000 1415.290 264.000 ;
        RECT 1415.120 244.110 1415.260 260.000 ;
        RECT 1415.060 243.790 1415.320 244.110 ;
        RECT 1421.040 243.790 1421.300 244.110 ;
        RECT 1421.100 39.090 1421.240 243.790 ;
        RECT 1421.040 38.770 1421.300 39.090 ;
        RECT 1721.420 38.090 1721.680 38.410 ;
        RECT 1721.480 2.400 1721.620 38.090 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 113.800 1435.130 113.860 ;
        RECT 1739.330 113.800 1739.650 113.860 ;
        RECT 1434.810 113.660 1739.650 113.800 ;
        RECT 1434.810 113.600 1435.130 113.660 ;
        RECT 1739.330 113.600 1739.650 113.660 ;
      LAYER via ;
        RECT 1434.840 113.600 1435.100 113.860 ;
        RECT 1739.360 113.600 1739.620 113.860 ;
      LAYER met2 ;
        RECT 1432.950 260.170 1433.230 264.000 ;
        RECT 1432.950 260.030 1435.040 260.170 ;
        RECT 1432.950 260.000 1433.230 260.030 ;
        RECT 1434.900 113.890 1435.040 260.030 ;
        RECT 1434.840 113.570 1435.100 113.890 ;
        RECT 1739.360 113.570 1739.620 113.890 ;
        RECT 1739.420 2.400 1739.560 113.570 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1450.910 244.020 1451.230 244.080 ;
        RECT 1455.510 244.020 1455.830 244.080 ;
        RECT 1450.910 243.880 1455.830 244.020 ;
        RECT 1450.910 243.820 1451.230 243.880 ;
        RECT 1455.510 243.820 1455.830 243.880 ;
        RECT 1455.510 45.460 1455.830 45.520 ;
        RECT 1756.810 45.460 1757.130 45.520 ;
        RECT 1455.510 45.320 1757.130 45.460 ;
        RECT 1455.510 45.260 1455.830 45.320 ;
        RECT 1756.810 45.260 1757.130 45.320 ;
      LAYER via ;
        RECT 1450.940 243.820 1451.200 244.080 ;
        RECT 1455.540 243.820 1455.800 244.080 ;
        RECT 1455.540 45.260 1455.800 45.520 ;
        RECT 1756.840 45.260 1757.100 45.520 ;
      LAYER met2 ;
        RECT 1450.890 260.000 1451.170 264.000 ;
        RECT 1451.000 244.110 1451.140 260.000 ;
        RECT 1450.940 243.790 1451.200 244.110 ;
        RECT 1455.540 243.790 1455.800 244.110 ;
        RECT 1455.600 45.550 1455.740 243.790 ;
        RECT 1455.540 45.230 1455.800 45.550 ;
        RECT 1756.840 45.230 1757.100 45.550 ;
        RECT 1756.900 2.400 1757.040 45.230 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1468.390 241.980 1468.710 242.040 ;
        RECT 1472.990 241.980 1473.310 242.040 ;
        RECT 1468.390 241.840 1473.310 241.980 ;
        RECT 1468.390 241.780 1468.710 241.840 ;
        RECT 1472.990 241.780 1473.310 241.840 ;
        RECT 1472.990 51.580 1473.310 51.640 ;
        RECT 1773.370 51.580 1773.690 51.640 ;
        RECT 1472.990 51.440 1773.690 51.580 ;
        RECT 1472.990 51.380 1473.310 51.440 ;
        RECT 1773.370 51.380 1773.690 51.440 ;
        RECT 1773.370 2.960 1773.690 3.020 ;
        RECT 1774.750 2.960 1775.070 3.020 ;
        RECT 1773.370 2.820 1775.070 2.960 ;
        RECT 1773.370 2.760 1773.690 2.820 ;
        RECT 1774.750 2.760 1775.070 2.820 ;
      LAYER via ;
        RECT 1468.420 241.780 1468.680 242.040 ;
        RECT 1473.020 241.780 1473.280 242.040 ;
        RECT 1473.020 51.380 1473.280 51.640 ;
        RECT 1773.400 51.380 1773.660 51.640 ;
        RECT 1773.400 2.760 1773.660 3.020 ;
        RECT 1774.780 2.760 1775.040 3.020 ;
      LAYER met2 ;
        RECT 1468.370 260.000 1468.650 264.000 ;
        RECT 1468.480 242.070 1468.620 260.000 ;
        RECT 1468.420 241.750 1468.680 242.070 ;
        RECT 1473.020 241.750 1473.280 242.070 ;
        RECT 1473.080 51.670 1473.220 241.750 ;
        RECT 1473.020 51.350 1473.280 51.670 ;
        RECT 1773.400 51.350 1773.660 51.670 ;
        RECT 1773.460 3.050 1773.600 51.350 ;
        RECT 1773.400 2.730 1773.660 3.050 ;
        RECT 1774.780 2.730 1775.040 3.050 ;
        RECT 1774.840 2.400 1774.980 2.730 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 59.060 1490.330 59.120 ;
        RECT 1787.170 59.060 1787.490 59.120 ;
        RECT 1490.010 58.920 1787.490 59.060 ;
        RECT 1490.010 58.860 1490.330 58.920 ;
        RECT 1787.170 58.860 1787.490 58.920 ;
        RECT 1787.170 2.960 1787.490 3.020 ;
        RECT 1792.690 2.960 1793.010 3.020 ;
        RECT 1787.170 2.820 1793.010 2.960 ;
        RECT 1787.170 2.760 1787.490 2.820 ;
        RECT 1792.690 2.760 1793.010 2.820 ;
      LAYER via ;
        RECT 1490.040 58.860 1490.300 59.120 ;
        RECT 1787.200 58.860 1787.460 59.120 ;
        RECT 1787.200 2.760 1787.460 3.020 ;
        RECT 1792.720 2.760 1792.980 3.020 ;
      LAYER met2 ;
        RECT 1486.310 260.170 1486.590 264.000 ;
        RECT 1486.310 260.030 1490.240 260.170 ;
        RECT 1486.310 260.000 1486.590 260.030 ;
        RECT 1490.100 59.150 1490.240 260.030 ;
        RECT 1490.040 58.830 1490.300 59.150 ;
        RECT 1787.200 58.830 1787.460 59.150 ;
        RECT 1787.260 3.050 1787.400 58.830 ;
        RECT 1787.200 2.730 1787.460 3.050 ;
        RECT 1792.720 2.730 1792.980 3.050 ;
        RECT 1792.780 2.400 1792.920 2.730 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1504.270 242.660 1504.590 242.720 ;
        RECT 1510.710 242.660 1511.030 242.720 ;
        RECT 1504.270 242.520 1511.030 242.660 ;
        RECT 1504.270 242.460 1504.590 242.520 ;
        RECT 1510.710 242.460 1511.030 242.520 ;
        RECT 1510.710 65.520 1511.030 65.580 ;
        RECT 1807.870 65.520 1808.190 65.580 ;
        RECT 1510.710 65.380 1808.190 65.520 ;
        RECT 1510.710 65.320 1511.030 65.380 ;
        RECT 1807.870 65.320 1808.190 65.380 ;
        RECT 1807.870 2.960 1808.190 3.020 ;
        RECT 1810.630 2.960 1810.950 3.020 ;
        RECT 1807.870 2.820 1810.950 2.960 ;
        RECT 1807.870 2.760 1808.190 2.820 ;
        RECT 1810.630 2.760 1810.950 2.820 ;
      LAYER via ;
        RECT 1504.300 242.460 1504.560 242.720 ;
        RECT 1510.740 242.460 1511.000 242.720 ;
        RECT 1510.740 65.320 1511.000 65.580 ;
        RECT 1807.900 65.320 1808.160 65.580 ;
        RECT 1807.900 2.760 1808.160 3.020 ;
        RECT 1810.660 2.760 1810.920 3.020 ;
      LAYER met2 ;
        RECT 1504.250 260.000 1504.530 264.000 ;
        RECT 1504.360 242.750 1504.500 260.000 ;
        RECT 1504.300 242.430 1504.560 242.750 ;
        RECT 1510.740 242.430 1511.000 242.750 ;
        RECT 1510.800 65.610 1510.940 242.430 ;
        RECT 1510.740 65.290 1511.000 65.610 ;
        RECT 1807.900 65.290 1808.160 65.610 ;
        RECT 1807.960 3.050 1808.100 65.290 ;
        RECT 1807.900 2.730 1808.160 3.050 ;
        RECT 1810.660 2.730 1810.920 3.050 ;
        RECT 1810.720 2.400 1810.860 2.730 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 72.660 1524.830 72.720 ;
        RECT 1829.030 72.660 1829.350 72.720 ;
        RECT 1524.510 72.520 1829.350 72.660 ;
        RECT 1524.510 72.460 1524.830 72.520 ;
        RECT 1829.030 72.460 1829.350 72.520 ;
      LAYER via ;
        RECT 1524.540 72.460 1524.800 72.720 ;
        RECT 1829.060 72.460 1829.320 72.720 ;
      LAYER met2 ;
        RECT 1522.190 260.170 1522.470 264.000 ;
        RECT 1522.190 260.030 1524.740 260.170 ;
        RECT 1522.190 260.000 1522.470 260.030 ;
        RECT 1524.600 72.750 1524.740 260.030 ;
        RECT 1524.540 72.430 1524.800 72.750 ;
        RECT 1829.060 72.430 1829.320 72.750 ;
        RECT 1829.120 7.210 1829.260 72.430 ;
        RECT 1828.660 7.070 1829.260 7.210 ;
        RECT 1828.660 2.400 1828.800 7.070 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1540.150 244.020 1540.470 244.080 ;
        RECT 1545.210 244.020 1545.530 244.080 ;
        RECT 1540.150 243.880 1545.530 244.020 ;
        RECT 1540.150 243.820 1540.470 243.880 ;
        RECT 1545.210 243.820 1545.530 243.880 ;
        RECT 1545.210 121.280 1545.530 121.340 ;
        RECT 1842.370 121.280 1842.690 121.340 ;
        RECT 1545.210 121.140 1842.690 121.280 ;
        RECT 1545.210 121.080 1545.530 121.140 ;
        RECT 1842.370 121.080 1842.690 121.140 ;
      LAYER via ;
        RECT 1540.180 243.820 1540.440 244.080 ;
        RECT 1545.240 243.820 1545.500 244.080 ;
        RECT 1545.240 121.080 1545.500 121.340 ;
        RECT 1842.400 121.080 1842.660 121.340 ;
      LAYER met2 ;
        RECT 1540.130 260.000 1540.410 264.000 ;
        RECT 1540.240 244.110 1540.380 260.000 ;
        RECT 1540.180 243.790 1540.440 244.110 ;
        RECT 1545.240 243.790 1545.500 244.110 ;
        RECT 1545.300 121.370 1545.440 243.790 ;
        RECT 1545.240 121.050 1545.500 121.370 ;
        RECT 1842.400 121.050 1842.660 121.370 ;
        RECT 1842.460 16.730 1842.600 121.050 ;
        RECT 1842.460 16.590 1846.280 16.730 ;
        RECT 1846.140 2.400 1846.280 16.590 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 141.340 1559.330 141.400 ;
        RECT 1863.070 141.340 1863.390 141.400 ;
        RECT 1559.010 141.200 1863.390 141.340 ;
        RECT 1559.010 141.140 1559.330 141.200 ;
        RECT 1863.070 141.140 1863.390 141.200 ;
      LAYER via ;
        RECT 1559.040 141.140 1559.300 141.400 ;
        RECT 1863.100 141.140 1863.360 141.400 ;
      LAYER met2 ;
        RECT 1558.070 260.170 1558.350 264.000 ;
        RECT 1558.070 260.030 1559.240 260.170 ;
        RECT 1558.070 260.000 1558.350 260.030 ;
        RECT 1559.100 141.430 1559.240 260.030 ;
        RECT 1559.040 141.110 1559.300 141.430 ;
        RECT 1863.100 141.110 1863.360 141.430 ;
        RECT 1863.160 16.730 1863.300 141.110 ;
        RECT 1863.160 16.590 1864.220 16.730 ;
        RECT 1864.080 2.400 1864.220 16.590 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 434.310 120.600 434.630 120.660 ;
        RECT 738.370 120.600 738.690 120.660 ;
        RECT 434.310 120.460 738.690 120.600 ;
        RECT 434.310 120.400 434.630 120.460 ;
        RECT 738.370 120.400 738.690 120.460 ;
      LAYER via ;
        RECT 434.340 120.400 434.600 120.660 ;
        RECT 738.400 120.400 738.660 120.660 ;
      LAYER met2 ;
        RECT 431.990 260.170 432.270 264.000 ;
        RECT 431.990 260.030 434.540 260.170 ;
        RECT 431.990 260.000 432.270 260.030 ;
        RECT 434.400 120.690 434.540 260.030 ;
        RECT 434.340 120.370 434.600 120.690 ;
        RECT 738.400 120.370 738.660 120.690 ;
        RECT 738.460 16.730 738.600 120.370 ;
        RECT 738.460 16.590 740.440 16.730 ;
        RECT 740.300 2.400 740.440 16.590 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1576.030 243.000 1576.350 243.060 ;
        RECT 1579.710 243.000 1580.030 243.060 ;
        RECT 1576.030 242.860 1580.030 243.000 ;
        RECT 1576.030 242.800 1576.350 242.860 ;
        RECT 1579.710 242.800 1580.030 242.860 ;
        RECT 1579.710 79.800 1580.030 79.860 ;
        RECT 1876.870 79.800 1877.190 79.860 ;
        RECT 1579.710 79.660 1877.190 79.800 ;
        RECT 1579.710 79.600 1580.030 79.660 ;
        RECT 1876.870 79.600 1877.190 79.660 ;
      LAYER via ;
        RECT 1576.060 242.800 1576.320 243.060 ;
        RECT 1579.740 242.800 1580.000 243.060 ;
        RECT 1579.740 79.600 1580.000 79.860 ;
        RECT 1876.900 79.600 1877.160 79.860 ;
      LAYER met2 ;
        RECT 1576.010 260.000 1576.290 264.000 ;
        RECT 1576.120 243.090 1576.260 260.000 ;
        RECT 1576.060 242.770 1576.320 243.090 ;
        RECT 1579.740 242.770 1580.000 243.090 ;
        RECT 1579.800 79.890 1579.940 242.770 ;
        RECT 1579.740 79.570 1580.000 79.890 ;
        RECT 1876.900 79.570 1877.160 79.890 ;
        RECT 1876.960 16.730 1877.100 79.570 ;
        RECT 1876.960 16.590 1882.160 16.730 ;
        RECT 1882.020 2.400 1882.160 16.590 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 245.040 1593.830 245.100 ;
        RECT 1873.190 245.040 1873.510 245.100 ;
        RECT 1593.510 244.900 1873.510 245.040 ;
        RECT 1593.510 244.840 1593.830 244.900 ;
        RECT 1873.190 244.840 1873.510 244.900 ;
        RECT 1873.190 27.780 1873.510 27.840 ;
        RECT 1899.870 27.780 1900.190 27.840 ;
        RECT 1873.190 27.640 1900.190 27.780 ;
        RECT 1873.190 27.580 1873.510 27.640 ;
        RECT 1899.870 27.580 1900.190 27.640 ;
      LAYER via ;
        RECT 1593.540 244.840 1593.800 245.100 ;
        RECT 1873.220 244.840 1873.480 245.100 ;
        RECT 1873.220 27.580 1873.480 27.840 ;
        RECT 1899.900 27.580 1900.160 27.840 ;
      LAYER met2 ;
        RECT 1593.490 260.000 1593.770 264.000 ;
        RECT 1593.600 245.130 1593.740 260.000 ;
        RECT 1593.540 244.810 1593.800 245.130 ;
        RECT 1873.220 244.810 1873.480 245.130 ;
        RECT 1873.280 27.870 1873.420 244.810 ;
        RECT 1873.220 27.550 1873.480 27.870 ;
        RECT 1899.900 27.550 1900.160 27.870 ;
        RECT 1899.960 2.400 1900.100 27.550 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 86.260 1614.530 86.320 ;
        RECT 1911.830 86.260 1912.150 86.320 ;
        RECT 1614.210 86.120 1912.150 86.260 ;
        RECT 1614.210 86.060 1614.530 86.120 ;
        RECT 1911.830 86.060 1912.150 86.120 ;
        RECT 1911.830 18.260 1912.150 18.320 ;
        RECT 1917.810 18.260 1918.130 18.320 ;
        RECT 1911.830 18.120 1918.130 18.260 ;
        RECT 1911.830 18.060 1912.150 18.120 ;
        RECT 1917.810 18.060 1918.130 18.120 ;
      LAYER via ;
        RECT 1614.240 86.060 1614.500 86.320 ;
        RECT 1911.860 86.060 1912.120 86.320 ;
        RECT 1911.860 18.060 1912.120 18.320 ;
        RECT 1917.840 18.060 1918.100 18.320 ;
      LAYER met2 ;
        RECT 1611.430 260.170 1611.710 264.000 ;
        RECT 1611.430 260.030 1614.440 260.170 ;
        RECT 1611.430 260.000 1611.710 260.030 ;
        RECT 1614.300 86.350 1614.440 260.030 ;
        RECT 1614.240 86.030 1614.500 86.350 ;
        RECT 1911.860 86.030 1912.120 86.350 ;
        RECT 1911.920 18.350 1912.060 86.030 ;
        RECT 1911.860 18.030 1912.120 18.350 ;
        RECT 1917.840 18.030 1918.100 18.350 ;
        RECT 1917.900 2.400 1918.040 18.030 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1629.390 244.020 1629.710 244.080 ;
        RECT 1634.910 244.020 1635.230 244.080 ;
        RECT 1629.390 243.880 1635.230 244.020 ;
        RECT 1629.390 243.820 1629.710 243.880 ;
        RECT 1634.910 243.820 1635.230 243.880 ;
        RECT 1634.910 93.400 1635.230 93.460 ;
        RECT 1932.070 93.400 1932.390 93.460 ;
        RECT 1634.910 93.260 1932.390 93.400 ;
        RECT 1634.910 93.200 1635.230 93.260 ;
        RECT 1932.070 93.200 1932.390 93.260 ;
      LAYER via ;
        RECT 1629.420 243.820 1629.680 244.080 ;
        RECT 1634.940 243.820 1635.200 244.080 ;
        RECT 1634.940 93.200 1635.200 93.460 ;
        RECT 1932.100 93.200 1932.360 93.460 ;
      LAYER met2 ;
        RECT 1629.370 260.000 1629.650 264.000 ;
        RECT 1629.480 244.110 1629.620 260.000 ;
        RECT 1629.420 243.790 1629.680 244.110 ;
        RECT 1634.940 243.790 1635.200 244.110 ;
        RECT 1635.000 93.490 1635.140 243.790 ;
        RECT 1634.940 93.170 1635.200 93.490 ;
        RECT 1932.100 93.170 1932.360 93.490 ;
        RECT 1932.160 16.730 1932.300 93.170 ;
        RECT 1932.160 16.590 1935.520 16.730 ;
        RECT 1935.380 2.400 1935.520 16.590 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1647.330 244.020 1647.650 244.080 ;
        RECT 1652.390 244.020 1652.710 244.080 ;
        RECT 1647.330 243.880 1652.710 244.020 ;
        RECT 1647.330 243.820 1647.650 243.880 ;
        RECT 1652.390 243.820 1652.710 243.880 ;
        RECT 1652.390 99.860 1652.710 99.920 ;
        RECT 1953.230 99.860 1953.550 99.920 ;
        RECT 1652.390 99.720 1953.550 99.860 ;
        RECT 1652.390 99.660 1652.710 99.720 ;
        RECT 1953.230 99.660 1953.550 99.720 ;
      LAYER via ;
        RECT 1647.360 243.820 1647.620 244.080 ;
        RECT 1652.420 243.820 1652.680 244.080 ;
        RECT 1652.420 99.660 1652.680 99.920 ;
        RECT 1953.260 99.660 1953.520 99.920 ;
      LAYER met2 ;
        RECT 1647.310 260.000 1647.590 264.000 ;
        RECT 1647.420 244.110 1647.560 260.000 ;
        RECT 1647.360 243.790 1647.620 244.110 ;
        RECT 1652.420 243.790 1652.680 244.110 ;
        RECT 1652.480 99.950 1652.620 243.790 ;
        RECT 1652.420 99.630 1652.680 99.950 ;
        RECT 1953.260 99.630 1953.520 99.950 ;
        RECT 1953.320 2.400 1953.460 99.630 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1665.270 244.020 1665.590 244.080 ;
        RECT 1669.410 244.020 1669.730 244.080 ;
        RECT 1665.270 243.880 1669.730 244.020 ;
        RECT 1665.270 243.820 1665.590 243.880 ;
        RECT 1669.410 243.820 1669.730 243.880 ;
        RECT 1669.410 107.000 1669.730 107.060 ;
        RECT 1966.570 107.000 1966.890 107.060 ;
        RECT 1669.410 106.860 1966.890 107.000 ;
        RECT 1669.410 106.800 1669.730 106.860 ;
        RECT 1966.570 106.800 1966.890 106.860 ;
      LAYER via ;
        RECT 1665.300 243.820 1665.560 244.080 ;
        RECT 1669.440 243.820 1669.700 244.080 ;
        RECT 1669.440 106.800 1669.700 107.060 ;
        RECT 1966.600 106.800 1966.860 107.060 ;
      LAYER met2 ;
        RECT 1665.250 260.000 1665.530 264.000 ;
        RECT 1665.360 244.110 1665.500 260.000 ;
        RECT 1665.300 243.790 1665.560 244.110 ;
        RECT 1669.440 243.790 1669.700 244.110 ;
        RECT 1669.500 107.090 1669.640 243.790 ;
        RECT 1669.440 106.770 1669.700 107.090 ;
        RECT 1966.600 106.770 1966.860 107.090 ;
        RECT 1966.660 16.730 1966.800 106.770 ;
        RECT 1966.660 16.590 1971.400 16.730 ;
        RECT 1971.260 2.400 1971.400 16.590 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1684.130 237.900 1684.450 237.960 ;
        RECT 1987.270 237.900 1987.590 237.960 ;
        RECT 1684.130 237.760 1987.590 237.900 ;
        RECT 1684.130 237.700 1684.450 237.760 ;
        RECT 1987.270 237.700 1987.590 237.760 ;
      LAYER via ;
        RECT 1684.160 237.700 1684.420 237.960 ;
        RECT 1987.300 237.700 1987.560 237.960 ;
      LAYER met2 ;
        RECT 1683.190 260.000 1683.470 264.000 ;
        RECT 1683.300 244.530 1683.440 260.000 ;
        RECT 1683.300 244.390 1684.360 244.530 ;
        RECT 1684.220 237.990 1684.360 244.390 ;
        RECT 1684.160 237.670 1684.420 237.990 ;
        RECT 1987.300 237.670 1987.560 237.990 ;
        RECT 1987.360 16.730 1987.500 237.670 ;
        RECT 1987.360 16.590 1989.340 16.730 ;
        RECT 1989.200 2.400 1989.340 16.590 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 30.840 1704.230 30.900 ;
        RECT 2006.590 30.840 2006.910 30.900 ;
        RECT 1703.910 30.700 2006.910 30.840 ;
        RECT 1703.910 30.640 1704.230 30.700 ;
        RECT 2006.590 30.640 2006.910 30.700 ;
      LAYER via ;
        RECT 1703.940 30.640 1704.200 30.900 ;
        RECT 2006.620 30.640 2006.880 30.900 ;
      LAYER met2 ;
        RECT 1701.130 260.170 1701.410 264.000 ;
        RECT 1701.130 260.030 1704.140 260.170 ;
        RECT 1701.130 260.000 1701.410 260.030 ;
        RECT 1704.000 30.930 1704.140 260.030 ;
        RECT 1703.940 30.610 1704.200 30.930 ;
        RECT 2006.620 30.610 2006.880 30.930 ;
        RECT 2006.680 2.400 2006.820 30.610 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1718.630 244.020 1718.950 244.080 ;
        RECT 1724.610 244.020 1724.930 244.080 ;
        RECT 1718.630 243.880 1724.930 244.020 ;
        RECT 1718.630 243.820 1718.950 243.880 ;
        RECT 1724.610 243.820 1724.930 243.880 ;
        RECT 1724.610 37.980 1724.930 38.040 ;
        RECT 2024.530 37.980 2024.850 38.040 ;
        RECT 1724.610 37.840 2024.850 37.980 ;
        RECT 1724.610 37.780 1724.930 37.840 ;
        RECT 2024.530 37.780 2024.850 37.840 ;
      LAYER via ;
        RECT 1718.660 243.820 1718.920 244.080 ;
        RECT 1724.640 243.820 1724.900 244.080 ;
        RECT 1724.640 37.780 1724.900 38.040 ;
        RECT 2024.560 37.780 2024.820 38.040 ;
      LAYER met2 ;
        RECT 1718.610 260.000 1718.890 264.000 ;
        RECT 1718.720 244.110 1718.860 260.000 ;
        RECT 1718.660 243.790 1718.920 244.110 ;
        RECT 1724.640 243.790 1724.900 244.110 ;
        RECT 1724.700 38.070 1724.840 243.790 ;
        RECT 1724.640 37.750 1724.900 38.070 ;
        RECT 2024.560 37.750 2024.820 38.070 ;
        RECT 2024.620 2.400 2024.760 37.750 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1736.570 244.020 1736.890 244.080 ;
        RECT 1742.090 244.020 1742.410 244.080 ;
        RECT 1736.570 243.880 1742.410 244.020 ;
        RECT 1736.570 243.820 1736.890 243.880 ;
        RECT 1742.090 243.820 1742.410 243.880 ;
        RECT 1742.090 113.800 1742.410 113.860 ;
        RECT 2042.930 113.800 2043.250 113.860 ;
        RECT 1742.090 113.660 2043.250 113.800 ;
        RECT 1742.090 113.600 1742.410 113.660 ;
        RECT 2042.930 113.600 2043.250 113.660 ;
      LAYER via ;
        RECT 1736.600 243.820 1736.860 244.080 ;
        RECT 1742.120 243.820 1742.380 244.080 ;
        RECT 1742.120 113.600 1742.380 113.860 ;
        RECT 2042.960 113.600 2043.220 113.860 ;
      LAYER met2 ;
        RECT 1736.550 260.000 1736.830 264.000 ;
        RECT 1736.660 244.110 1736.800 260.000 ;
        RECT 1736.600 243.790 1736.860 244.110 ;
        RECT 1742.120 243.790 1742.380 244.110 ;
        RECT 1742.180 113.890 1742.320 243.790 ;
        RECT 1742.120 113.570 1742.380 113.890 ;
        RECT 2042.960 113.570 2043.220 113.890 ;
        RECT 2043.020 17.410 2043.160 113.570 ;
        RECT 2042.560 17.270 2043.160 17.410 ;
        RECT 2042.560 2.400 2042.700 17.270 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 449.490 244.020 449.810 244.080 ;
        RECT 455.010 244.020 455.330 244.080 ;
        RECT 449.490 243.880 455.330 244.020 ;
        RECT 449.490 243.820 449.810 243.880 ;
        RECT 455.010 243.820 455.330 243.880 ;
        RECT 455.010 127.740 455.330 127.800 ;
        RECT 752.630 127.740 752.950 127.800 ;
        RECT 455.010 127.600 752.950 127.740 ;
        RECT 455.010 127.540 455.330 127.600 ;
        RECT 752.630 127.540 752.950 127.600 ;
        RECT 752.630 19.620 752.950 19.680 ;
        RECT 757.690 19.620 758.010 19.680 ;
        RECT 752.630 19.480 758.010 19.620 ;
        RECT 752.630 19.420 752.950 19.480 ;
        RECT 757.690 19.420 758.010 19.480 ;
      LAYER via ;
        RECT 449.520 243.820 449.780 244.080 ;
        RECT 455.040 243.820 455.300 244.080 ;
        RECT 455.040 127.540 455.300 127.800 ;
        RECT 752.660 127.540 752.920 127.800 ;
        RECT 752.660 19.420 752.920 19.680 ;
        RECT 757.720 19.420 757.980 19.680 ;
      LAYER met2 ;
        RECT 449.470 260.000 449.750 264.000 ;
        RECT 449.580 244.110 449.720 260.000 ;
        RECT 449.520 243.790 449.780 244.110 ;
        RECT 455.040 243.790 455.300 244.110 ;
        RECT 455.100 127.830 455.240 243.790 ;
        RECT 455.040 127.510 455.300 127.830 ;
        RECT 752.660 127.510 752.920 127.830 ;
        RECT 752.720 19.710 752.860 127.510 ;
        RECT 752.660 19.390 752.920 19.710 ;
        RECT 757.720 19.390 757.980 19.710 ;
        RECT 757.780 2.400 757.920 19.390 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.510 244.020 1754.830 244.080 ;
        RECT 1759.110 244.020 1759.430 244.080 ;
        RECT 1754.510 243.880 1759.430 244.020 ;
        RECT 1754.510 243.820 1754.830 243.880 ;
        RECT 1759.110 243.820 1759.430 243.880 ;
        RECT 1759.110 45.120 1759.430 45.180 ;
        RECT 2060.410 45.120 2060.730 45.180 ;
        RECT 1759.110 44.980 2060.730 45.120 ;
        RECT 1759.110 44.920 1759.430 44.980 ;
        RECT 2060.410 44.920 2060.730 44.980 ;
      LAYER via ;
        RECT 1754.540 243.820 1754.800 244.080 ;
        RECT 1759.140 243.820 1759.400 244.080 ;
        RECT 1759.140 44.920 1759.400 45.180 ;
        RECT 2060.440 44.920 2060.700 45.180 ;
      LAYER met2 ;
        RECT 1754.490 260.000 1754.770 264.000 ;
        RECT 1754.600 244.110 1754.740 260.000 ;
        RECT 1754.540 243.790 1754.800 244.110 ;
        RECT 1759.140 243.790 1759.400 244.110 ;
        RECT 1759.200 45.210 1759.340 243.790 ;
        RECT 1759.140 44.890 1759.400 45.210 ;
        RECT 2060.440 44.890 2060.700 45.210 ;
        RECT 2060.500 2.400 2060.640 44.890 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.450 248.440 1772.770 248.500 ;
        RECT 1776.590 248.440 1776.910 248.500 ;
        RECT 1772.450 248.300 1776.910 248.440 ;
        RECT 1772.450 248.240 1772.770 248.300 ;
        RECT 1776.590 248.240 1776.910 248.300 ;
        RECT 1776.590 51.580 1776.910 51.640 ;
        RECT 2076.970 51.580 2077.290 51.640 ;
        RECT 1776.590 51.440 2077.290 51.580 ;
        RECT 1776.590 51.380 1776.910 51.440 ;
        RECT 2076.970 51.380 2077.290 51.440 ;
      LAYER via ;
        RECT 1772.480 248.240 1772.740 248.500 ;
        RECT 1776.620 248.240 1776.880 248.500 ;
        RECT 1776.620 51.380 1776.880 51.640 ;
        RECT 2077.000 51.380 2077.260 51.640 ;
      LAYER met2 ;
        RECT 1772.430 260.000 1772.710 264.000 ;
        RECT 1772.540 248.530 1772.680 260.000 ;
        RECT 1772.480 248.210 1772.740 248.530 ;
        RECT 1776.620 248.210 1776.880 248.530 ;
        RECT 1776.680 51.670 1776.820 248.210 ;
        RECT 1776.620 51.350 1776.880 51.670 ;
        RECT 2077.000 51.350 2077.260 51.670 ;
        RECT 2077.060 3.130 2077.200 51.350 ;
        RECT 2077.060 2.990 2078.580 3.130 ;
        RECT 2078.440 2.400 2078.580 2.990 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 25.060 1793.930 25.120 ;
        RECT 1793.610 24.920 1845.820 25.060 ;
        RECT 1793.610 24.860 1793.930 24.920 ;
        RECT 1845.680 24.720 1845.820 24.920 ;
        RECT 2095.830 24.720 2096.150 24.780 ;
        RECT 1845.680 24.580 2096.150 24.720 ;
        RECT 2095.830 24.520 2096.150 24.580 ;
      LAYER via ;
        RECT 1793.640 24.860 1793.900 25.120 ;
        RECT 2095.860 24.520 2096.120 24.780 ;
      LAYER met2 ;
        RECT 1790.370 260.170 1790.650 264.000 ;
        RECT 1790.370 260.030 1793.840 260.170 ;
        RECT 1790.370 260.000 1790.650 260.030 ;
        RECT 1793.700 25.150 1793.840 260.030 ;
        RECT 1793.640 24.830 1793.900 25.150 ;
        RECT 2095.860 24.490 2096.120 24.810 ;
        RECT 2095.920 2.400 2096.060 24.490 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1808.330 244.020 1808.650 244.080 ;
        RECT 1814.310 244.020 1814.630 244.080 ;
        RECT 1808.330 243.880 1814.630 244.020 ;
        RECT 1808.330 243.820 1808.650 243.880 ;
        RECT 1814.310 243.820 1814.630 243.880 ;
        RECT 1814.310 26.420 1814.630 26.480 ;
        RECT 2113.770 26.420 2114.090 26.480 ;
        RECT 1814.310 26.280 2114.090 26.420 ;
        RECT 1814.310 26.220 1814.630 26.280 ;
        RECT 2113.770 26.220 2114.090 26.280 ;
      LAYER via ;
        RECT 1808.360 243.820 1808.620 244.080 ;
        RECT 1814.340 243.820 1814.600 244.080 ;
        RECT 1814.340 26.220 1814.600 26.480 ;
        RECT 2113.800 26.220 2114.060 26.480 ;
      LAYER met2 ;
        RECT 1808.310 260.000 1808.590 264.000 ;
        RECT 1808.420 244.110 1808.560 260.000 ;
        RECT 1808.360 243.790 1808.620 244.110 ;
        RECT 1814.340 243.790 1814.600 244.110 ;
        RECT 1814.400 26.510 1814.540 243.790 ;
        RECT 1814.340 26.190 1814.600 26.510 ;
        RECT 2113.800 26.190 2114.060 26.510 ;
        RECT 2113.860 2.400 2114.000 26.190 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1826.270 243.340 1826.590 243.400 ;
        RECT 1838.690 243.340 1839.010 243.400 ;
        RECT 1826.270 243.200 1839.010 243.340 ;
        RECT 1826.270 243.140 1826.590 243.200 ;
        RECT 1838.690 243.140 1839.010 243.200 ;
        RECT 1838.690 59.060 1839.010 59.120 ;
        RECT 2125.270 59.060 2125.590 59.120 ;
        RECT 1838.690 58.920 2125.590 59.060 ;
        RECT 1838.690 58.860 1839.010 58.920 ;
        RECT 2125.270 58.860 2125.590 58.920 ;
        RECT 2125.270 16.900 2125.590 16.960 ;
        RECT 2131.710 16.900 2132.030 16.960 ;
        RECT 2125.270 16.760 2132.030 16.900 ;
        RECT 2125.270 16.700 2125.590 16.760 ;
        RECT 2131.710 16.700 2132.030 16.760 ;
      LAYER via ;
        RECT 1826.300 243.140 1826.560 243.400 ;
        RECT 1838.720 243.140 1838.980 243.400 ;
        RECT 1838.720 58.860 1838.980 59.120 ;
        RECT 2125.300 58.860 2125.560 59.120 ;
        RECT 2125.300 16.700 2125.560 16.960 ;
        RECT 2131.740 16.700 2132.000 16.960 ;
      LAYER met2 ;
        RECT 1826.250 260.000 1826.530 264.000 ;
        RECT 1826.360 243.430 1826.500 260.000 ;
        RECT 1826.300 243.110 1826.560 243.430 ;
        RECT 1838.720 243.110 1838.980 243.430 ;
        RECT 1838.780 59.150 1838.920 243.110 ;
        RECT 1838.720 58.830 1838.980 59.150 ;
        RECT 2125.300 58.830 2125.560 59.150 ;
        RECT 2125.360 16.990 2125.500 58.830 ;
        RECT 2125.300 16.670 2125.560 16.990 ;
        RECT 2131.740 16.670 2132.000 16.990 ;
        RECT 2131.800 2.400 2131.940 16.670 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1844.210 241.640 1844.530 241.700 ;
        RECT 1848.810 241.640 1849.130 241.700 ;
        RECT 1844.210 241.500 1849.130 241.640 ;
        RECT 1844.210 241.440 1844.530 241.500 ;
        RECT 1848.810 241.440 1849.130 241.500 ;
        RECT 1848.810 25.060 1849.130 25.120 ;
        RECT 2149.650 25.060 2149.970 25.120 ;
        RECT 1848.810 24.920 2149.970 25.060 ;
        RECT 1848.810 24.860 1849.130 24.920 ;
        RECT 2149.650 24.860 2149.970 24.920 ;
      LAYER via ;
        RECT 1844.240 241.440 1844.500 241.700 ;
        RECT 1848.840 241.440 1849.100 241.700 ;
        RECT 1848.840 24.860 1849.100 25.120 ;
        RECT 2149.680 24.860 2149.940 25.120 ;
      LAYER met2 ;
        RECT 1844.190 260.000 1844.470 264.000 ;
        RECT 1844.300 241.730 1844.440 260.000 ;
        RECT 1844.240 241.410 1844.500 241.730 ;
        RECT 1848.840 241.410 1849.100 241.730 ;
        RECT 1848.900 25.150 1849.040 241.410 ;
        RECT 1848.840 24.830 1849.100 25.150 ;
        RECT 2149.680 24.830 2149.940 25.150 ;
        RECT 2149.740 2.400 2149.880 24.830 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 24.040 1862.930 24.100 ;
        RECT 2167.590 24.040 2167.910 24.100 ;
        RECT 1862.610 23.900 2167.910 24.040 ;
        RECT 1862.610 23.840 1862.930 23.900 ;
        RECT 2167.590 23.840 2167.910 23.900 ;
      LAYER via ;
        RECT 1862.640 23.840 1862.900 24.100 ;
        RECT 2167.620 23.840 2167.880 24.100 ;
      LAYER met2 ;
        RECT 1861.670 260.170 1861.950 264.000 ;
        RECT 1861.670 260.030 1862.840 260.170 ;
        RECT 1861.670 260.000 1861.950 260.030 ;
        RECT 1862.700 24.130 1862.840 260.030 ;
        RECT 1862.640 23.810 1862.900 24.130 ;
        RECT 2167.620 23.810 2167.880 24.130 ;
        RECT 2167.680 2.400 2167.820 23.810 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2185.145 2.805 2185.315 48.195 ;
      LAYER mcon ;
        RECT 2185.145 48.025 2185.315 48.195 ;
      LAYER met1 ;
        RECT 1879.630 244.020 1879.950 244.080 ;
        RECT 1883.310 244.020 1883.630 244.080 ;
        RECT 1879.630 243.880 1883.630 244.020 ;
        RECT 1879.630 243.820 1879.950 243.880 ;
        RECT 1883.310 243.820 1883.630 243.880 ;
        RECT 1883.310 65.520 1883.630 65.580 ;
        RECT 2180.470 65.520 2180.790 65.580 ;
        RECT 1883.310 65.380 2180.790 65.520 ;
        RECT 1883.310 65.320 1883.630 65.380 ;
        RECT 2180.470 65.320 2180.790 65.380 ;
        RECT 2180.470 48.180 2180.790 48.240 ;
        RECT 2185.085 48.180 2185.375 48.225 ;
        RECT 2180.470 48.040 2185.375 48.180 ;
        RECT 2180.470 47.980 2180.790 48.040 ;
        RECT 2185.085 47.995 2185.375 48.040 ;
        RECT 2185.070 2.960 2185.390 3.020 ;
        RECT 2184.875 2.820 2185.390 2.960 ;
        RECT 2185.070 2.760 2185.390 2.820 ;
      LAYER via ;
        RECT 1879.660 243.820 1879.920 244.080 ;
        RECT 1883.340 243.820 1883.600 244.080 ;
        RECT 1883.340 65.320 1883.600 65.580 ;
        RECT 2180.500 65.320 2180.760 65.580 ;
        RECT 2180.500 47.980 2180.760 48.240 ;
        RECT 2185.100 2.760 2185.360 3.020 ;
      LAYER met2 ;
        RECT 1879.610 260.000 1879.890 264.000 ;
        RECT 1879.720 244.110 1879.860 260.000 ;
        RECT 1879.660 243.790 1879.920 244.110 ;
        RECT 1883.340 243.790 1883.600 244.110 ;
        RECT 1883.400 65.610 1883.540 243.790 ;
        RECT 1883.340 65.290 1883.600 65.610 ;
        RECT 2180.500 65.290 2180.760 65.610 ;
        RECT 2180.560 48.270 2180.700 65.290 ;
        RECT 2180.500 47.950 2180.760 48.270 ;
        RECT 2185.100 2.730 2185.360 3.050 ;
        RECT 2185.160 2.400 2185.300 2.730 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1897.570 244.020 1897.890 244.080 ;
        RECT 1904.010 244.020 1904.330 244.080 ;
        RECT 1897.570 243.880 1904.330 244.020 ;
        RECT 1897.570 243.820 1897.890 243.880 ;
        RECT 1904.010 243.820 1904.330 243.880 ;
        RECT 1904.010 26.080 1904.330 26.140 ;
        RECT 2203.010 26.080 2203.330 26.140 ;
        RECT 1904.010 25.940 2203.330 26.080 ;
        RECT 1904.010 25.880 1904.330 25.940 ;
        RECT 2203.010 25.880 2203.330 25.940 ;
      LAYER via ;
        RECT 1897.600 243.820 1897.860 244.080 ;
        RECT 1904.040 243.820 1904.300 244.080 ;
        RECT 1904.040 25.880 1904.300 26.140 ;
        RECT 2203.040 25.880 2203.300 26.140 ;
      LAYER met2 ;
        RECT 1897.550 260.000 1897.830 264.000 ;
        RECT 1897.660 244.110 1897.800 260.000 ;
        RECT 1897.600 243.790 1897.860 244.110 ;
        RECT 1904.040 243.790 1904.300 244.110 ;
        RECT 1904.100 26.170 1904.240 243.790 ;
        RECT 1904.040 25.850 1904.300 26.170 ;
        RECT 2203.040 25.850 2203.300 26.170 ;
        RECT 2203.100 2.400 2203.240 25.850 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1915.510 248.440 1915.830 248.500 ;
        RECT 1921.490 248.440 1921.810 248.500 ;
        RECT 1915.510 248.300 1921.810 248.440 ;
        RECT 1915.510 248.240 1915.830 248.300 ;
        RECT 1921.490 248.240 1921.810 248.300 ;
        RECT 1921.490 72.320 1921.810 72.380 ;
        RECT 2215.430 72.320 2215.750 72.380 ;
        RECT 1921.490 72.180 2215.750 72.320 ;
        RECT 1921.490 72.120 1921.810 72.180 ;
        RECT 2215.430 72.120 2215.750 72.180 ;
      LAYER via ;
        RECT 1915.540 248.240 1915.800 248.500 ;
        RECT 1921.520 248.240 1921.780 248.500 ;
        RECT 1921.520 72.120 1921.780 72.380 ;
        RECT 2215.460 72.120 2215.720 72.380 ;
      LAYER met2 ;
        RECT 1915.490 260.000 1915.770 264.000 ;
        RECT 1915.600 248.530 1915.740 260.000 ;
        RECT 1915.540 248.210 1915.800 248.530 ;
        RECT 1921.520 248.210 1921.780 248.530 ;
        RECT 1921.580 72.410 1921.720 248.210 ;
        RECT 1921.520 72.090 1921.780 72.410 ;
        RECT 2215.460 72.090 2215.720 72.410 ;
        RECT 2215.520 16.730 2215.660 72.090 ;
        RECT 2215.520 16.590 2221.180 16.730 ;
        RECT 2221.040 2.400 2221.180 16.590 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 468.810 134.540 469.130 134.600 ;
        RECT 772.870 134.540 773.190 134.600 ;
        RECT 468.810 134.400 773.190 134.540 ;
        RECT 468.810 134.340 469.130 134.400 ;
        RECT 772.870 134.340 773.190 134.400 ;
      LAYER via ;
        RECT 468.840 134.340 469.100 134.600 ;
        RECT 772.900 134.340 773.160 134.600 ;
      LAYER met2 ;
        RECT 467.410 260.170 467.690 264.000 ;
        RECT 467.410 260.030 469.040 260.170 ;
        RECT 467.410 260.000 467.690 260.030 ;
        RECT 468.900 134.630 469.040 260.030 ;
        RECT 468.840 134.310 469.100 134.630 ;
        RECT 772.900 134.310 773.160 134.630 ;
        RECT 772.960 16.730 773.100 134.310 ;
        RECT 772.960 16.590 775.860 16.730 ;
        RECT 775.720 2.400 775.860 16.590 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1933.450 244.020 1933.770 244.080 ;
        RECT 1938.510 244.020 1938.830 244.080 ;
        RECT 1933.450 243.880 1938.830 244.020 ;
        RECT 1933.450 243.820 1933.770 243.880 ;
        RECT 1938.510 243.820 1938.830 243.880 ;
        RECT 1938.510 25.400 1938.830 25.460 ;
        RECT 2238.890 25.400 2239.210 25.460 ;
        RECT 1938.510 25.260 2239.210 25.400 ;
        RECT 1938.510 25.200 1938.830 25.260 ;
        RECT 2238.890 25.200 2239.210 25.260 ;
      LAYER via ;
        RECT 1933.480 243.820 1933.740 244.080 ;
        RECT 1938.540 243.820 1938.800 244.080 ;
        RECT 1938.540 25.200 1938.800 25.460 ;
        RECT 2238.920 25.200 2239.180 25.460 ;
      LAYER met2 ;
        RECT 1933.430 260.000 1933.710 264.000 ;
        RECT 1933.540 244.110 1933.680 260.000 ;
        RECT 1933.480 243.790 1933.740 244.110 ;
        RECT 1938.540 243.790 1938.800 244.110 ;
        RECT 1938.600 25.490 1938.740 243.790 ;
        RECT 1938.540 25.170 1938.800 25.490 ;
        RECT 2238.920 25.170 2239.180 25.490 ;
        RECT 2238.980 2.400 2239.120 25.170 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1966.645 23.545 1966.815 24.395 ;
        RECT 2014.945 23.545 2015.115 24.395 ;
        RECT 2096.365 23.545 2096.535 24.735 ;
        RECT 2125.345 23.205 2125.515 24.735 ;
        RECT 2173.185 23.205 2173.355 24.395 ;
        RECT 2173.645 23.545 2173.815 24.735 ;
        RECT 2221.485 23.545 2221.655 24.395 ;
        RECT 2225.625 14.705 2225.795 24.395 ;
      LAYER mcon ;
        RECT 2096.365 24.565 2096.535 24.735 ;
        RECT 1966.645 24.225 1966.815 24.395 ;
        RECT 2014.945 24.225 2015.115 24.395 ;
        RECT 2125.345 24.565 2125.515 24.735 ;
        RECT 2173.645 24.565 2173.815 24.735 ;
        RECT 2173.185 24.225 2173.355 24.395 ;
        RECT 2221.485 24.225 2221.655 24.395 ;
        RECT 2225.625 24.225 2225.795 24.395 ;
      LAYER met1 ;
        RECT 2096.305 24.720 2096.595 24.765 ;
        RECT 2125.285 24.720 2125.575 24.765 ;
        RECT 2173.585 24.720 2173.875 24.765 ;
        RECT 2096.305 24.580 2125.575 24.720 ;
        RECT 2096.305 24.535 2096.595 24.580 ;
        RECT 2125.285 24.535 2125.575 24.580 ;
        RECT 2173.200 24.580 2173.875 24.720 ;
        RECT 2173.200 24.425 2173.340 24.580 ;
        RECT 2173.585 24.535 2173.875 24.580 ;
        RECT 1966.585 24.380 1966.875 24.425 ;
        RECT 2014.885 24.380 2015.175 24.425 ;
        RECT 1966.585 24.240 2015.175 24.380 ;
        RECT 1966.585 24.195 1966.875 24.240 ;
        RECT 2014.885 24.195 2015.175 24.240 ;
        RECT 2173.125 24.195 2173.415 24.425 ;
        RECT 2221.425 24.380 2221.715 24.425 ;
        RECT 2225.565 24.380 2225.855 24.425 ;
        RECT 2221.425 24.240 2225.855 24.380 ;
        RECT 2221.425 24.195 2221.715 24.240 ;
        RECT 2225.565 24.195 2225.855 24.240 ;
        RECT 1952.310 23.700 1952.630 23.760 ;
        RECT 1966.585 23.700 1966.875 23.745 ;
        RECT 1952.310 23.560 1966.875 23.700 ;
        RECT 1952.310 23.500 1952.630 23.560 ;
        RECT 1966.585 23.515 1966.875 23.560 ;
        RECT 2014.885 23.700 2015.175 23.745 ;
        RECT 2096.305 23.700 2096.595 23.745 ;
        RECT 2014.885 23.560 2096.595 23.700 ;
        RECT 2014.885 23.515 2015.175 23.560 ;
        RECT 2096.305 23.515 2096.595 23.560 ;
        RECT 2173.585 23.700 2173.875 23.745 ;
        RECT 2221.425 23.700 2221.715 23.745 ;
        RECT 2173.585 23.560 2221.715 23.700 ;
        RECT 2173.585 23.515 2173.875 23.560 ;
        RECT 2221.425 23.515 2221.715 23.560 ;
        RECT 2125.285 23.360 2125.575 23.405 ;
        RECT 2173.125 23.360 2173.415 23.405 ;
        RECT 2125.285 23.220 2173.415 23.360 ;
        RECT 2125.285 23.175 2125.575 23.220 ;
        RECT 2173.125 23.175 2173.415 23.220 ;
        RECT 2225.565 14.860 2225.855 14.905 ;
        RECT 2256.370 14.860 2256.690 14.920 ;
        RECT 2225.565 14.720 2256.690 14.860 ;
        RECT 2225.565 14.675 2225.855 14.720 ;
        RECT 2256.370 14.660 2256.690 14.720 ;
      LAYER via ;
        RECT 1952.340 23.500 1952.600 23.760 ;
        RECT 2256.400 14.660 2256.660 14.920 ;
      LAYER met2 ;
        RECT 1951.370 260.170 1951.650 264.000 ;
        RECT 1951.370 260.030 1952.540 260.170 ;
        RECT 1951.370 260.000 1951.650 260.030 ;
        RECT 1952.400 23.790 1952.540 260.030 ;
        RECT 1952.340 23.470 1952.600 23.790 ;
        RECT 2256.400 14.630 2256.660 14.950 ;
        RECT 2256.460 2.400 2256.600 14.630 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.010 25.740 1973.330 25.800 ;
        RECT 2274.310 25.740 2274.630 25.800 ;
        RECT 1973.010 25.600 2274.630 25.740 ;
        RECT 1973.010 25.540 1973.330 25.600 ;
        RECT 2274.310 25.540 2274.630 25.600 ;
      LAYER via ;
        RECT 1973.040 25.540 1973.300 25.800 ;
        RECT 2274.340 25.540 2274.600 25.800 ;
      LAYER met2 ;
        RECT 1969.310 260.170 1969.590 264.000 ;
        RECT 1969.310 260.030 1973.240 260.170 ;
        RECT 1969.310 260.000 1969.590 260.030 ;
        RECT 1973.100 25.830 1973.240 260.030 ;
        RECT 1973.040 25.510 1973.300 25.830 ;
        RECT 2274.340 25.510 2274.600 25.830 ;
        RECT 2274.400 2.400 2274.540 25.510 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.810 79.460 1987.130 79.520 ;
        RECT 2290.870 79.460 2291.190 79.520 ;
        RECT 1986.810 79.320 2291.190 79.460 ;
        RECT 1986.810 79.260 1987.130 79.320 ;
        RECT 2290.870 79.260 2291.190 79.320 ;
      LAYER via ;
        RECT 1986.840 79.260 1987.100 79.520 ;
        RECT 2290.900 79.260 2291.160 79.520 ;
      LAYER met2 ;
        RECT 1986.790 260.000 1987.070 264.000 ;
        RECT 1986.900 79.550 1987.040 260.000 ;
        RECT 1986.840 79.230 1987.100 79.550 ;
        RECT 2290.900 79.230 2291.160 79.550 ;
        RECT 2290.960 3.130 2291.100 79.230 ;
        RECT 2290.960 2.990 2292.020 3.130 ;
        RECT 2291.880 2.960 2292.020 2.990 ;
        RECT 2291.880 2.820 2292.480 2.960 ;
        RECT 2292.340 2.400 2292.480 2.820 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2004.750 248.440 2005.070 248.500 ;
        RECT 2018.090 248.440 2018.410 248.500 ;
        RECT 2004.750 248.300 2018.410 248.440 ;
        RECT 2004.750 248.240 2005.070 248.300 ;
        RECT 2018.090 248.240 2018.410 248.300 ;
        RECT 2018.090 86.600 2018.410 86.660 ;
        RECT 2304.670 86.600 2304.990 86.660 ;
        RECT 2018.090 86.460 2304.990 86.600 ;
        RECT 2018.090 86.400 2018.410 86.460 ;
        RECT 2304.670 86.400 2304.990 86.460 ;
        RECT 2305.130 2.960 2305.450 3.020 ;
        RECT 2310.190 2.960 2310.510 3.020 ;
        RECT 2305.130 2.820 2310.510 2.960 ;
        RECT 2305.130 2.760 2305.450 2.820 ;
        RECT 2310.190 2.760 2310.510 2.820 ;
      LAYER via ;
        RECT 2004.780 248.240 2005.040 248.500 ;
        RECT 2018.120 248.240 2018.380 248.500 ;
        RECT 2018.120 86.400 2018.380 86.660 ;
        RECT 2304.700 86.400 2304.960 86.660 ;
        RECT 2305.160 2.760 2305.420 3.020 ;
        RECT 2310.220 2.760 2310.480 3.020 ;
      LAYER met2 ;
        RECT 2004.730 260.000 2005.010 264.000 ;
        RECT 2004.840 248.530 2004.980 260.000 ;
        RECT 2004.780 248.210 2005.040 248.530 ;
        RECT 2018.120 248.210 2018.380 248.530 ;
        RECT 2018.180 86.690 2018.320 248.210 ;
        RECT 2018.120 86.370 2018.380 86.690 ;
        RECT 2304.700 86.370 2304.960 86.690 ;
        RECT 2304.760 20.130 2304.900 86.370 ;
        RECT 2304.760 19.990 2305.360 20.130 ;
        RECT 2305.220 3.050 2305.360 19.990 ;
        RECT 2305.160 2.730 2305.420 3.050 ;
        RECT 2310.220 2.730 2310.480 3.050 ;
        RECT 2310.280 2.400 2310.420 2.730 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2022.690 244.020 2023.010 244.080 ;
        RECT 2028.210 244.020 2028.530 244.080 ;
        RECT 2022.690 243.880 2028.530 244.020 ;
        RECT 2022.690 243.820 2023.010 243.880 ;
        RECT 2028.210 243.820 2028.530 243.880 ;
        RECT 2028.210 93.060 2028.530 93.120 ;
        RECT 2325.370 93.060 2325.690 93.120 ;
        RECT 2028.210 92.920 2325.690 93.060 ;
        RECT 2028.210 92.860 2028.530 92.920 ;
        RECT 2325.370 92.860 2325.690 92.920 ;
        RECT 2325.370 2.960 2325.690 3.020 ;
        RECT 2328.130 2.960 2328.450 3.020 ;
        RECT 2325.370 2.820 2328.450 2.960 ;
        RECT 2325.370 2.760 2325.690 2.820 ;
        RECT 2328.130 2.760 2328.450 2.820 ;
      LAYER via ;
        RECT 2022.720 243.820 2022.980 244.080 ;
        RECT 2028.240 243.820 2028.500 244.080 ;
        RECT 2028.240 92.860 2028.500 93.120 ;
        RECT 2325.400 92.860 2325.660 93.120 ;
        RECT 2325.400 2.760 2325.660 3.020 ;
        RECT 2328.160 2.760 2328.420 3.020 ;
      LAYER met2 ;
        RECT 2022.670 260.000 2022.950 264.000 ;
        RECT 2022.780 244.110 2022.920 260.000 ;
        RECT 2022.720 243.790 2022.980 244.110 ;
        RECT 2028.240 243.790 2028.500 244.110 ;
        RECT 2028.300 93.150 2028.440 243.790 ;
        RECT 2028.240 92.830 2028.500 93.150 ;
        RECT 2325.400 92.830 2325.660 93.150 ;
        RECT 2325.460 3.050 2325.600 92.830 ;
        RECT 2325.400 2.730 2325.660 3.050 ;
        RECT 2328.160 2.730 2328.420 3.050 ;
        RECT 2328.220 2.400 2328.360 2.730 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 99.860 2042.330 99.920 ;
        RECT 2339.170 99.860 2339.490 99.920 ;
        RECT 2042.010 99.720 2339.490 99.860 ;
        RECT 2042.010 99.660 2042.330 99.720 ;
        RECT 2339.170 99.660 2339.490 99.720 ;
        RECT 2339.170 17.920 2339.490 17.980 ;
        RECT 2345.610 17.920 2345.930 17.980 ;
        RECT 2339.170 17.780 2345.930 17.920 ;
        RECT 2339.170 17.720 2339.490 17.780 ;
        RECT 2345.610 17.720 2345.930 17.780 ;
      LAYER via ;
        RECT 2042.040 99.660 2042.300 99.920 ;
        RECT 2339.200 99.660 2339.460 99.920 ;
        RECT 2339.200 17.720 2339.460 17.980 ;
        RECT 2345.640 17.720 2345.900 17.980 ;
      LAYER met2 ;
        RECT 2040.610 260.170 2040.890 264.000 ;
        RECT 2040.610 260.030 2042.240 260.170 ;
        RECT 2040.610 260.000 2040.890 260.030 ;
        RECT 2042.100 99.950 2042.240 260.030 ;
        RECT 2042.040 99.630 2042.300 99.950 ;
        RECT 2339.200 99.630 2339.460 99.950 ;
        RECT 2339.260 18.010 2339.400 99.630 ;
        RECT 2339.200 17.690 2339.460 18.010 ;
        RECT 2345.640 17.690 2345.900 18.010 ;
        RECT 2345.700 2.400 2345.840 17.690 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2058.570 242.320 2058.890 242.380 ;
        RECT 2062.710 242.320 2063.030 242.380 ;
        RECT 2058.570 242.180 2063.030 242.320 ;
        RECT 2058.570 242.120 2058.890 242.180 ;
        RECT 2062.710 242.120 2063.030 242.180 ;
        RECT 2062.710 107.000 2063.030 107.060 ;
        RECT 2359.870 107.000 2360.190 107.060 ;
        RECT 2062.710 106.860 2360.190 107.000 ;
        RECT 2062.710 106.800 2063.030 106.860 ;
        RECT 2359.870 106.800 2360.190 106.860 ;
      LAYER via ;
        RECT 2058.600 242.120 2058.860 242.380 ;
        RECT 2062.740 242.120 2063.000 242.380 ;
        RECT 2062.740 106.800 2063.000 107.060 ;
        RECT 2359.900 106.800 2360.160 107.060 ;
      LAYER met2 ;
        RECT 2058.550 260.000 2058.830 264.000 ;
        RECT 2058.660 242.410 2058.800 260.000 ;
        RECT 2058.600 242.090 2058.860 242.410 ;
        RECT 2062.740 242.090 2063.000 242.410 ;
        RECT 2062.800 107.090 2062.940 242.090 ;
        RECT 2062.740 106.770 2063.000 107.090 ;
        RECT 2359.900 106.770 2360.160 107.090 ;
        RECT 2359.960 16.730 2360.100 106.770 ;
        RECT 2359.960 16.590 2363.780 16.730 ;
        RECT 2363.640 2.400 2363.780 16.590 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.050 224.300 2076.370 224.360 ;
        RECT 2380.570 224.300 2380.890 224.360 ;
        RECT 2076.050 224.160 2380.890 224.300 ;
        RECT 2076.050 224.100 2076.370 224.160 ;
        RECT 2380.570 224.100 2380.890 224.160 ;
      LAYER via ;
        RECT 2076.080 224.100 2076.340 224.360 ;
        RECT 2380.600 224.100 2380.860 224.360 ;
      LAYER met2 ;
        RECT 2076.490 260.170 2076.770 264.000 ;
        RECT 2076.140 260.030 2076.770 260.170 ;
        RECT 2076.140 224.390 2076.280 260.030 ;
        RECT 2076.490 260.000 2076.770 260.030 ;
        RECT 2076.080 224.070 2076.340 224.390 ;
        RECT 2380.600 224.070 2380.860 224.390 ;
        RECT 2380.660 16.730 2380.800 224.070 ;
        RECT 2380.660 16.590 2381.720 16.730 ;
        RECT 2381.580 2.400 2381.720 16.590 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2097.210 210.360 2097.530 210.420 ;
        RECT 2394.370 210.360 2394.690 210.420 ;
        RECT 2097.210 210.220 2394.690 210.360 ;
        RECT 2097.210 210.160 2097.530 210.220 ;
        RECT 2394.370 210.160 2394.690 210.220 ;
      LAYER via ;
        RECT 2097.240 210.160 2097.500 210.420 ;
        RECT 2394.400 210.160 2394.660 210.420 ;
      LAYER met2 ;
        RECT 2094.430 260.170 2094.710 264.000 ;
        RECT 2094.430 260.030 2097.440 260.170 ;
        RECT 2094.430 260.000 2094.710 260.030 ;
        RECT 2097.300 210.450 2097.440 260.030 ;
        RECT 2097.240 210.130 2097.500 210.450 ;
        RECT 2394.400 210.130 2394.660 210.450 ;
        RECT 2394.460 16.730 2394.600 210.130 ;
        RECT 2394.460 16.590 2399.660 16.730 ;
        RECT 2399.520 2.400 2399.660 16.590 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 485.370 244.020 485.690 244.080 ;
        RECT 489.510 244.020 489.830 244.080 ;
        RECT 485.370 243.880 489.830 244.020 ;
        RECT 485.370 243.820 485.690 243.880 ;
        RECT 489.510 243.820 489.830 243.880 ;
        RECT 489.510 141.680 489.830 141.740 ;
        RECT 794.030 141.680 794.350 141.740 ;
        RECT 489.510 141.540 794.350 141.680 ;
        RECT 489.510 141.480 489.830 141.540 ;
        RECT 794.030 141.480 794.350 141.540 ;
      LAYER via ;
        RECT 485.400 243.820 485.660 244.080 ;
        RECT 489.540 243.820 489.800 244.080 ;
        RECT 489.540 141.480 489.800 141.740 ;
        RECT 794.060 141.480 794.320 141.740 ;
      LAYER met2 ;
        RECT 485.350 260.000 485.630 264.000 ;
        RECT 485.460 244.110 485.600 260.000 ;
        RECT 485.400 243.790 485.660 244.110 ;
        RECT 489.540 243.790 489.800 244.110 ;
        RECT 489.600 141.770 489.740 243.790 ;
        RECT 489.540 141.450 489.800 141.770 ;
        RECT 794.060 141.450 794.320 141.770 ;
        RECT 794.120 17.410 794.260 141.450 ;
        RECT 793.660 17.270 794.260 17.410 ;
        RECT 793.660 2.400 793.800 17.270 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 330.350 244.020 330.670 244.080 ;
        RECT 334.490 244.020 334.810 244.080 ;
        RECT 330.350 243.880 334.810 244.020 ;
        RECT 330.350 243.820 330.670 243.880 ;
        RECT 334.490 243.820 334.810 243.880 ;
        RECT 334.490 79.460 334.810 79.520 ;
        RECT 634.870 79.460 635.190 79.520 ;
        RECT 334.490 79.320 635.190 79.460 ;
        RECT 334.490 79.260 334.810 79.320 ;
        RECT 634.870 79.260 635.190 79.320 ;
      LAYER via ;
        RECT 330.380 243.820 330.640 244.080 ;
        RECT 334.520 243.820 334.780 244.080 ;
        RECT 334.520 79.260 334.780 79.520 ;
        RECT 634.900 79.260 635.160 79.520 ;
      LAYER met2 ;
        RECT 330.330 260.000 330.610 264.000 ;
        RECT 330.440 244.110 330.580 260.000 ;
        RECT 330.380 243.790 330.640 244.110 ;
        RECT 334.520 243.790 334.780 244.110 ;
        RECT 334.580 79.550 334.720 243.790 ;
        RECT 334.520 79.230 334.780 79.550 ;
        RECT 634.900 79.230 635.160 79.550 ;
        RECT 634.960 17.410 635.100 79.230 ;
        RECT 634.960 17.270 639.240 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2117.450 113.800 2117.770 113.860 ;
        RECT 2421.970 113.800 2422.290 113.860 ;
        RECT 2117.450 113.660 2422.290 113.800 ;
        RECT 2117.450 113.600 2117.770 113.660 ;
        RECT 2421.970 113.600 2422.290 113.660 ;
      LAYER via ;
        RECT 2117.480 113.600 2117.740 113.860 ;
        RECT 2422.000 113.600 2422.260 113.860 ;
      LAYER met2 ;
        RECT 2117.890 260.170 2118.170 264.000 ;
        RECT 2117.540 260.030 2118.170 260.170 ;
        RECT 2117.540 113.890 2117.680 260.030 ;
        RECT 2117.890 260.000 2118.170 260.030 ;
        RECT 2117.480 113.570 2117.740 113.890 ;
        RECT 2422.000 113.570 2422.260 113.890 ;
        RECT 2422.060 16.730 2422.200 113.570 ;
        RECT 2422.060 16.590 2423.120 16.730 ;
        RECT 2422.980 2.400 2423.120 16.590 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.610 120.600 2138.930 120.660 ;
        RECT 2435.770 120.600 2436.090 120.660 ;
        RECT 2138.610 120.460 2436.090 120.600 ;
        RECT 2138.610 120.400 2138.930 120.460 ;
        RECT 2435.770 120.400 2436.090 120.460 ;
      LAYER via ;
        RECT 2138.640 120.400 2138.900 120.660 ;
        RECT 2435.800 120.400 2436.060 120.660 ;
      LAYER met2 ;
        RECT 2135.830 260.170 2136.110 264.000 ;
        RECT 2135.830 260.030 2138.840 260.170 ;
        RECT 2135.830 260.000 2136.110 260.030 ;
        RECT 2138.700 120.690 2138.840 260.030 ;
        RECT 2138.640 120.370 2138.900 120.690 ;
        RECT 2435.800 120.370 2436.060 120.690 ;
        RECT 2435.860 16.730 2436.000 120.370 ;
        RECT 2435.860 16.590 2441.060 16.730 ;
        RECT 2440.920 2.400 2441.060 16.590 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2153.790 244.020 2154.110 244.080 ;
        RECT 2159.310 244.020 2159.630 244.080 ;
        RECT 2153.790 243.880 2159.630 244.020 ;
        RECT 2153.790 243.820 2154.110 243.880 ;
        RECT 2159.310 243.820 2159.630 243.880 ;
        RECT 2159.310 128.080 2159.630 128.140 ;
        RECT 2456.470 128.080 2456.790 128.140 ;
        RECT 2159.310 127.940 2456.790 128.080 ;
        RECT 2159.310 127.880 2159.630 127.940 ;
        RECT 2456.470 127.880 2456.790 127.940 ;
      LAYER via ;
        RECT 2153.820 243.820 2154.080 244.080 ;
        RECT 2159.340 243.820 2159.600 244.080 ;
        RECT 2159.340 127.880 2159.600 128.140 ;
        RECT 2456.500 127.880 2456.760 128.140 ;
      LAYER met2 ;
        RECT 2153.770 260.000 2154.050 264.000 ;
        RECT 2153.880 244.110 2154.020 260.000 ;
        RECT 2153.820 243.790 2154.080 244.110 ;
        RECT 2159.340 243.790 2159.600 244.110 ;
        RECT 2159.400 128.170 2159.540 243.790 ;
        RECT 2159.340 127.850 2159.600 128.170 ;
        RECT 2456.500 127.850 2456.760 128.170 ;
        RECT 2456.560 17.410 2456.700 127.850 ;
        RECT 2456.560 17.270 2459.000 17.410 ;
        RECT 2458.860 2.400 2459.000 17.270 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2173.110 134.540 2173.430 134.600 ;
        RECT 2470.270 134.540 2470.590 134.600 ;
        RECT 2173.110 134.400 2470.590 134.540 ;
        RECT 2173.110 134.340 2173.430 134.400 ;
        RECT 2470.270 134.340 2470.590 134.400 ;
        RECT 2470.270 17.580 2470.590 17.640 ;
        RECT 2476.710 17.580 2477.030 17.640 ;
        RECT 2470.270 17.440 2477.030 17.580 ;
        RECT 2470.270 17.380 2470.590 17.440 ;
        RECT 2476.710 17.380 2477.030 17.440 ;
      LAYER via ;
        RECT 2173.140 134.340 2173.400 134.600 ;
        RECT 2470.300 134.340 2470.560 134.600 ;
        RECT 2470.300 17.380 2470.560 17.640 ;
        RECT 2476.740 17.380 2477.000 17.640 ;
      LAYER met2 ;
        RECT 2171.710 260.170 2171.990 264.000 ;
        RECT 2171.710 260.030 2173.340 260.170 ;
        RECT 2171.710 260.000 2171.990 260.030 ;
        RECT 2173.200 134.630 2173.340 260.030 ;
        RECT 2173.140 134.310 2173.400 134.630 ;
        RECT 2470.300 134.310 2470.560 134.630 ;
        RECT 2470.360 17.670 2470.500 134.310 ;
        RECT 2470.300 17.350 2470.560 17.670 ;
        RECT 2476.740 17.350 2477.000 17.670 ;
        RECT 2476.800 2.400 2476.940 17.350 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2189.670 244.020 2189.990 244.080 ;
        RECT 2193.810 244.020 2194.130 244.080 ;
        RECT 2189.670 243.880 2194.130 244.020 ;
        RECT 2189.670 243.820 2189.990 243.880 ;
        RECT 2193.810 243.820 2194.130 243.880 ;
        RECT 2193.810 148.140 2194.130 148.200 ;
        RECT 2490.970 148.140 2491.290 148.200 ;
        RECT 2193.810 148.000 2491.290 148.140 ;
        RECT 2193.810 147.940 2194.130 148.000 ;
        RECT 2490.970 147.940 2491.290 148.000 ;
      LAYER via ;
        RECT 2189.700 243.820 2189.960 244.080 ;
        RECT 2193.840 243.820 2194.100 244.080 ;
        RECT 2193.840 147.940 2194.100 148.200 ;
        RECT 2491.000 147.940 2491.260 148.200 ;
      LAYER met2 ;
        RECT 2189.650 260.000 2189.930 264.000 ;
        RECT 2189.760 244.110 2189.900 260.000 ;
        RECT 2189.700 243.790 2189.960 244.110 ;
        RECT 2193.840 243.790 2194.100 244.110 ;
        RECT 2193.900 148.230 2194.040 243.790 ;
        RECT 2193.840 147.910 2194.100 148.230 ;
        RECT 2491.000 147.910 2491.260 148.230 ;
        RECT 2491.060 17.410 2491.200 147.910 ;
        RECT 2491.060 17.270 2494.880 17.410 ;
        RECT 2494.740 2.400 2494.880 17.270 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2207.610 169.220 2207.930 169.280 ;
        RECT 2512.130 169.220 2512.450 169.280 ;
        RECT 2207.610 169.080 2512.450 169.220 ;
        RECT 2207.610 169.020 2207.930 169.080 ;
        RECT 2512.130 169.020 2512.450 169.080 ;
      LAYER via ;
        RECT 2207.640 169.020 2207.900 169.280 ;
        RECT 2512.160 169.020 2512.420 169.280 ;
      LAYER met2 ;
        RECT 2207.590 260.000 2207.870 264.000 ;
        RECT 2207.700 169.310 2207.840 260.000 ;
        RECT 2207.640 168.990 2207.900 169.310 ;
        RECT 2512.160 168.990 2512.420 169.310 ;
        RECT 2512.220 2.400 2512.360 168.990 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2228.310 141.340 2228.630 141.400 ;
        RECT 2525.470 141.340 2525.790 141.400 ;
        RECT 2228.310 141.200 2525.790 141.340 ;
        RECT 2228.310 141.140 2228.630 141.200 ;
        RECT 2525.470 141.140 2525.790 141.200 ;
      LAYER via ;
        RECT 2228.340 141.140 2228.600 141.400 ;
        RECT 2525.500 141.140 2525.760 141.400 ;
      LAYER met2 ;
        RECT 2225.530 260.170 2225.810 264.000 ;
        RECT 2225.530 260.030 2228.540 260.170 ;
        RECT 2225.530 260.000 2225.810 260.030 ;
        RECT 2228.400 141.430 2228.540 260.030 ;
        RECT 2228.340 141.110 2228.600 141.430 ;
        RECT 2525.500 141.110 2525.760 141.430 ;
        RECT 2525.560 16.730 2525.700 141.110 ;
        RECT 2525.560 16.590 2530.300 16.730 ;
        RECT 2530.160 2.400 2530.300 16.590 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2243.030 244.020 2243.350 244.080 ;
        RECT 2248.550 244.020 2248.870 244.080 ;
        RECT 2243.030 243.880 2248.870 244.020 ;
        RECT 2243.030 243.820 2243.350 243.880 ;
        RECT 2248.550 243.820 2248.870 243.880 ;
        RECT 2248.550 155.280 2248.870 155.340 ;
        RECT 2546.170 155.280 2546.490 155.340 ;
        RECT 2248.550 155.140 2546.490 155.280 ;
        RECT 2248.550 155.080 2248.870 155.140 ;
        RECT 2546.170 155.080 2546.490 155.140 ;
      LAYER via ;
        RECT 2243.060 243.820 2243.320 244.080 ;
        RECT 2248.580 243.820 2248.840 244.080 ;
        RECT 2248.580 155.080 2248.840 155.340 ;
        RECT 2546.200 155.080 2546.460 155.340 ;
      LAYER met2 ;
        RECT 2243.010 260.000 2243.290 264.000 ;
        RECT 2243.120 244.110 2243.260 260.000 ;
        RECT 2243.060 243.790 2243.320 244.110 ;
        RECT 2248.580 243.790 2248.840 244.110 ;
        RECT 2248.640 155.370 2248.780 243.790 ;
        RECT 2248.580 155.050 2248.840 155.370 ;
        RECT 2546.200 155.050 2546.460 155.370 ;
        RECT 2546.260 16.730 2546.400 155.050 ;
        RECT 2546.260 16.590 2548.240 16.730 ;
        RECT 2548.100 2.400 2548.240 16.590 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2262.810 37.980 2263.130 38.040 ;
        RECT 2565.950 37.980 2566.270 38.040 ;
        RECT 2262.810 37.840 2566.270 37.980 ;
        RECT 2262.810 37.780 2263.130 37.840 ;
        RECT 2565.950 37.780 2566.270 37.840 ;
      LAYER via ;
        RECT 2262.840 37.780 2263.100 38.040 ;
        RECT 2565.980 37.780 2566.240 38.040 ;
      LAYER met2 ;
        RECT 2260.950 260.170 2261.230 264.000 ;
        RECT 2260.950 260.030 2263.040 260.170 ;
        RECT 2260.950 260.000 2261.230 260.030 ;
        RECT 2262.900 38.070 2263.040 260.030 ;
        RECT 2262.840 37.750 2263.100 38.070 ;
        RECT 2565.980 37.750 2566.240 38.070 ;
        RECT 2566.040 2.400 2566.180 37.750 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2278.910 244.020 2279.230 244.080 ;
        RECT 2283.510 244.020 2283.830 244.080 ;
        RECT 2278.910 243.880 2283.830 244.020 ;
        RECT 2278.910 243.820 2279.230 243.880 ;
        RECT 2283.510 243.820 2283.830 243.880 ;
        RECT 2283.510 86.260 2283.830 86.320 ;
        RECT 2580.670 86.260 2580.990 86.320 ;
        RECT 2283.510 86.120 2580.990 86.260 ;
        RECT 2283.510 86.060 2283.830 86.120 ;
        RECT 2580.670 86.060 2580.990 86.120 ;
      LAYER via ;
        RECT 2278.940 243.820 2279.200 244.080 ;
        RECT 2283.540 243.820 2283.800 244.080 ;
        RECT 2283.540 86.060 2283.800 86.320 ;
        RECT 2580.700 86.060 2580.960 86.320 ;
      LAYER met2 ;
        RECT 2278.890 260.000 2279.170 264.000 ;
        RECT 2279.000 244.110 2279.140 260.000 ;
        RECT 2278.940 243.790 2279.200 244.110 ;
        RECT 2283.540 243.790 2283.800 244.110 ;
        RECT 2283.600 86.350 2283.740 243.790 ;
        RECT 2283.540 86.030 2283.800 86.350 ;
        RECT 2580.700 86.030 2580.960 86.350 ;
        RECT 2580.760 16.730 2580.900 86.030 ;
        RECT 2580.760 16.590 2584.120 16.730 ;
        RECT 2583.980 2.400 2584.120 16.590 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 510.210 148.140 510.530 148.200 ;
        RECT 814.270 148.140 814.590 148.200 ;
        RECT 510.210 148.000 814.590 148.140 ;
        RECT 510.210 147.940 510.530 148.000 ;
        RECT 814.270 147.940 814.590 148.000 ;
      LAYER via ;
        RECT 510.240 147.940 510.500 148.200 ;
        RECT 814.300 147.940 814.560 148.200 ;
      LAYER met2 ;
        RECT 509.270 260.170 509.550 264.000 ;
        RECT 509.270 260.030 510.440 260.170 ;
        RECT 509.270 260.000 509.550 260.030 ;
        RECT 510.300 148.230 510.440 260.030 ;
        RECT 510.240 147.910 510.500 148.230 ;
        RECT 814.300 147.910 814.560 148.230 ;
        RECT 814.360 17.410 814.500 147.910 ;
        RECT 814.360 17.270 817.720 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2296.850 244.020 2297.170 244.080 ;
        RECT 2300.990 244.020 2301.310 244.080 ;
        RECT 2296.850 243.880 2301.310 244.020 ;
        RECT 2296.850 243.820 2297.170 243.880 ;
        RECT 2300.990 243.820 2301.310 243.880 ;
        RECT 2300.990 176.020 2301.310 176.080 ;
        RECT 2601.830 176.020 2602.150 176.080 ;
        RECT 2300.990 175.880 2602.150 176.020 ;
        RECT 2300.990 175.820 2301.310 175.880 ;
        RECT 2601.830 175.820 2602.150 175.880 ;
      LAYER via ;
        RECT 2296.880 243.820 2297.140 244.080 ;
        RECT 2301.020 243.820 2301.280 244.080 ;
        RECT 2301.020 175.820 2301.280 176.080 ;
        RECT 2601.860 175.820 2602.120 176.080 ;
      LAYER met2 ;
        RECT 2296.830 260.000 2297.110 264.000 ;
        RECT 2296.940 244.110 2297.080 260.000 ;
        RECT 2296.880 243.790 2297.140 244.110 ;
        RECT 2301.020 243.790 2301.280 244.110 ;
        RECT 2301.080 176.110 2301.220 243.790 ;
        RECT 2301.020 175.790 2301.280 176.110 ;
        RECT 2601.860 175.790 2602.120 176.110 ;
        RECT 2601.920 17.410 2602.060 175.790 ;
        RECT 2601.460 17.270 2602.060 17.410 ;
        RECT 2601.460 2.400 2601.600 17.270 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 26.420 2318.330 26.480 ;
        RECT 2619.310 26.420 2619.630 26.480 ;
        RECT 2318.010 26.280 2619.630 26.420 ;
        RECT 2318.010 26.220 2318.330 26.280 ;
        RECT 2619.310 26.220 2619.630 26.280 ;
      LAYER via ;
        RECT 2318.040 26.220 2318.300 26.480 ;
        RECT 2619.340 26.220 2619.600 26.480 ;
      LAYER met2 ;
        RECT 2314.770 260.170 2315.050 264.000 ;
        RECT 2314.770 260.030 2318.240 260.170 ;
        RECT 2314.770 260.000 2315.050 260.030 ;
        RECT 2318.100 26.510 2318.240 260.030 ;
        RECT 2318.040 26.190 2318.300 26.510 ;
        RECT 2619.340 26.190 2619.600 26.510 ;
        RECT 2619.400 2.400 2619.540 26.190 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2332.730 244.020 2333.050 244.080 ;
        RECT 2338.710 244.020 2339.030 244.080 ;
        RECT 2332.730 243.880 2339.030 244.020 ;
        RECT 2332.730 243.820 2333.050 243.880 ;
        RECT 2338.710 243.820 2339.030 243.880 ;
        RECT 2338.710 162.080 2339.030 162.140 ;
        RECT 2635.870 162.080 2636.190 162.140 ;
        RECT 2338.710 161.940 2636.190 162.080 ;
        RECT 2338.710 161.880 2339.030 161.940 ;
        RECT 2635.870 161.880 2636.190 161.940 ;
      LAYER via ;
        RECT 2332.760 243.820 2333.020 244.080 ;
        RECT 2338.740 243.820 2339.000 244.080 ;
        RECT 2338.740 161.880 2339.000 162.140 ;
        RECT 2635.900 161.880 2636.160 162.140 ;
      LAYER met2 ;
        RECT 2332.710 260.000 2332.990 264.000 ;
        RECT 2332.820 244.110 2332.960 260.000 ;
        RECT 2332.760 243.790 2333.020 244.110 ;
        RECT 2338.740 243.790 2339.000 244.110 ;
        RECT 2338.800 162.170 2338.940 243.790 ;
        RECT 2338.740 161.850 2339.000 162.170 ;
        RECT 2635.900 161.850 2636.160 162.170 ;
        RECT 2635.960 16.730 2636.100 161.850 ;
        RECT 2635.960 16.590 2637.480 16.730 ;
        RECT 2637.340 2.400 2637.480 16.590 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2352.510 99.860 2352.830 99.920 ;
        RECT 2649.670 99.860 2649.990 99.920 ;
        RECT 2352.510 99.720 2649.990 99.860 ;
        RECT 2352.510 99.660 2352.830 99.720 ;
        RECT 2649.670 99.660 2649.990 99.720 ;
      LAYER via ;
        RECT 2352.540 99.660 2352.800 99.920 ;
        RECT 2649.700 99.660 2649.960 99.920 ;
      LAYER met2 ;
        RECT 2350.650 260.170 2350.930 264.000 ;
        RECT 2350.650 260.030 2352.740 260.170 ;
        RECT 2350.650 260.000 2350.930 260.030 ;
        RECT 2352.600 99.950 2352.740 260.030 ;
        RECT 2352.540 99.630 2352.800 99.950 ;
        RECT 2649.700 99.630 2649.960 99.950 ;
        RECT 2649.760 17.410 2649.900 99.630 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2368.150 244.020 2368.470 244.080 ;
        RECT 2373.210 244.020 2373.530 244.080 ;
        RECT 2368.150 243.880 2373.530 244.020 ;
        RECT 2368.150 243.820 2368.470 243.880 ;
        RECT 2373.210 243.820 2373.530 243.880 ;
        RECT 2373.210 107.000 2373.530 107.060 ;
        RECT 2670.370 107.000 2670.690 107.060 ;
        RECT 2373.210 106.860 2670.690 107.000 ;
        RECT 2373.210 106.800 2373.530 106.860 ;
        RECT 2670.370 106.800 2670.690 106.860 ;
      LAYER via ;
        RECT 2368.180 243.820 2368.440 244.080 ;
        RECT 2373.240 243.820 2373.500 244.080 ;
        RECT 2373.240 106.800 2373.500 107.060 ;
        RECT 2670.400 106.800 2670.660 107.060 ;
      LAYER met2 ;
        RECT 2368.130 260.000 2368.410 264.000 ;
        RECT 2368.240 244.110 2368.380 260.000 ;
        RECT 2368.180 243.790 2368.440 244.110 ;
        RECT 2373.240 243.790 2373.500 244.110 ;
        RECT 2373.300 107.090 2373.440 243.790 ;
        RECT 2373.240 106.770 2373.500 107.090 ;
        RECT 2670.400 106.770 2670.660 107.090 ;
        RECT 2670.460 17.410 2670.600 106.770 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2386.090 248.440 2386.410 248.500 ;
        RECT 2411.390 248.440 2411.710 248.500 ;
        RECT 2386.090 248.300 2411.710 248.440 ;
        RECT 2386.090 248.240 2386.410 248.300 ;
        RECT 2411.390 248.240 2411.710 248.300 ;
        RECT 2411.390 114.140 2411.710 114.200 ;
        RECT 2684.170 114.140 2684.490 114.200 ;
        RECT 2411.390 114.000 2684.490 114.140 ;
        RECT 2411.390 113.940 2411.710 114.000 ;
        RECT 2684.170 113.940 2684.490 114.000 ;
        RECT 2684.170 17.920 2684.490 17.980 ;
        RECT 2690.610 17.920 2690.930 17.980 ;
        RECT 2684.170 17.780 2690.930 17.920 ;
        RECT 2684.170 17.720 2684.490 17.780 ;
        RECT 2690.610 17.720 2690.930 17.780 ;
      LAYER via ;
        RECT 2386.120 248.240 2386.380 248.500 ;
        RECT 2411.420 248.240 2411.680 248.500 ;
        RECT 2411.420 113.940 2411.680 114.200 ;
        RECT 2684.200 113.940 2684.460 114.200 ;
        RECT 2684.200 17.720 2684.460 17.980 ;
        RECT 2690.640 17.720 2690.900 17.980 ;
      LAYER met2 ;
        RECT 2386.070 260.000 2386.350 264.000 ;
        RECT 2386.180 248.530 2386.320 260.000 ;
        RECT 2386.120 248.210 2386.380 248.530 ;
        RECT 2411.420 248.210 2411.680 248.530 ;
        RECT 2411.480 114.230 2411.620 248.210 ;
        RECT 2411.420 113.910 2411.680 114.230 ;
        RECT 2684.200 113.910 2684.460 114.230 ;
        RECT 2684.260 18.010 2684.400 113.910 ;
        RECT 2684.200 17.690 2684.460 18.010 ;
        RECT 2690.640 17.690 2690.900 18.010 ;
        RECT 2690.700 2.400 2690.840 17.690 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2404.030 244.020 2404.350 244.080 ;
        RECT 2407.710 244.020 2408.030 244.080 ;
        RECT 2404.030 243.880 2408.030 244.020 ;
        RECT 2404.030 243.820 2404.350 243.880 ;
        RECT 2407.710 243.820 2408.030 243.880 ;
        RECT 2407.710 120.940 2408.030 121.000 ;
        RECT 2704.870 120.940 2705.190 121.000 ;
        RECT 2407.710 120.800 2705.190 120.940 ;
        RECT 2407.710 120.740 2408.030 120.800 ;
        RECT 2704.870 120.740 2705.190 120.800 ;
      LAYER via ;
        RECT 2404.060 243.820 2404.320 244.080 ;
        RECT 2407.740 243.820 2408.000 244.080 ;
        RECT 2407.740 120.740 2408.000 121.000 ;
        RECT 2704.900 120.740 2705.160 121.000 ;
      LAYER met2 ;
        RECT 2404.010 260.000 2404.290 264.000 ;
        RECT 2404.120 244.110 2404.260 260.000 ;
        RECT 2404.060 243.790 2404.320 244.110 ;
        RECT 2407.740 243.790 2408.000 244.110 ;
        RECT 2407.800 121.030 2407.940 243.790 ;
        RECT 2407.740 120.710 2408.000 121.030 ;
        RECT 2704.900 120.710 2705.160 121.030 ;
        RECT 2704.960 17.410 2705.100 120.710 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2421.970 244.020 2422.290 244.080 ;
        RECT 2427.950 244.020 2428.270 244.080 ;
        RECT 2421.970 243.880 2428.270 244.020 ;
        RECT 2421.970 243.820 2422.290 243.880 ;
        RECT 2427.950 243.820 2428.270 243.880 ;
        RECT 2427.950 127.740 2428.270 127.800 ;
        RECT 2725.570 127.740 2725.890 127.800 ;
        RECT 2427.950 127.600 2725.890 127.740 ;
        RECT 2427.950 127.540 2428.270 127.600 ;
        RECT 2725.570 127.540 2725.890 127.600 ;
      LAYER via ;
        RECT 2422.000 243.820 2422.260 244.080 ;
        RECT 2427.980 243.820 2428.240 244.080 ;
        RECT 2427.980 127.540 2428.240 127.800 ;
        RECT 2725.600 127.540 2725.860 127.800 ;
      LAYER met2 ;
        RECT 2421.950 260.000 2422.230 264.000 ;
        RECT 2422.060 244.110 2422.200 260.000 ;
        RECT 2422.000 243.790 2422.260 244.110 ;
        RECT 2427.980 243.790 2428.240 244.110 ;
        RECT 2428.040 127.830 2428.180 243.790 ;
        RECT 2427.980 127.510 2428.240 127.830 ;
        RECT 2725.600 127.510 2725.860 127.830 ;
        RECT 2725.660 17.410 2725.800 127.510 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2439.910 243.680 2440.230 243.740 ;
        RECT 2445.890 243.680 2446.210 243.740 ;
        RECT 2439.910 243.540 2446.210 243.680 ;
        RECT 2439.910 243.480 2440.230 243.540 ;
        RECT 2445.890 243.480 2446.210 243.540 ;
        RECT 2445.890 45.120 2446.210 45.180 ;
        RECT 2744.430 45.120 2744.750 45.180 ;
        RECT 2445.890 44.980 2744.750 45.120 ;
        RECT 2445.890 44.920 2446.210 44.980 ;
        RECT 2744.430 44.920 2744.750 44.980 ;
      LAYER via ;
        RECT 2439.940 243.480 2440.200 243.740 ;
        RECT 2445.920 243.480 2446.180 243.740 ;
        RECT 2445.920 44.920 2446.180 45.180 ;
        RECT 2744.460 44.920 2744.720 45.180 ;
      LAYER met2 ;
        RECT 2439.890 260.000 2440.170 264.000 ;
        RECT 2440.000 243.770 2440.140 260.000 ;
        RECT 2439.940 243.450 2440.200 243.770 ;
        RECT 2445.920 243.450 2446.180 243.770 ;
        RECT 2445.980 45.210 2446.120 243.450 ;
        RECT 2445.920 44.890 2446.180 45.210 ;
        RECT 2744.460 44.890 2744.720 45.210 ;
        RECT 2744.520 2.400 2744.660 44.890 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2457.850 244.020 2458.170 244.080 ;
        RECT 2462.910 244.020 2463.230 244.080 ;
        RECT 2457.850 243.880 2463.230 244.020 ;
        RECT 2457.850 243.820 2458.170 243.880 ;
        RECT 2462.910 243.820 2463.230 243.880 ;
        RECT 2462.910 134.880 2463.230 134.940 ;
        RECT 2760.070 134.880 2760.390 134.940 ;
        RECT 2462.910 134.740 2760.390 134.880 ;
        RECT 2462.910 134.680 2463.230 134.740 ;
        RECT 2760.070 134.680 2760.390 134.740 ;
      LAYER via ;
        RECT 2457.880 243.820 2458.140 244.080 ;
        RECT 2462.940 243.820 2463.200 244.080 ;
        RECT 2462.940 134.680 2463.200 134.940 ;
        RECT 2760.100 134.680 2760.360 134.940 ;
      LAYER met2 ;
        RECT 2457.830 260.000 2458.110 264.000 ;
        RECT 2457.940 244.110 2458.080 260.000 ;
        RECT 2457.880 243.790 2458.140 244.110 ;
        RECT 2462.940 243.790 2463.200 244.110 ;
        RECT 2463.000 134.970 2463.140 243.790 ;
        RECT 2462.940 134.650 2463.200 134.970 ;
        RECT 2760.100 134.650 2760.360 134.970 ;
        RECT 2760.160 17.410 2760.300 134.650 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 527.230 244.020 527.550 244.080 ;
        RECT 530.910 244.020 531.230 244.080 ;
        RECT 527.230 243.880 531.230 244.020 ;
        RECT 527.230 243.820 527.550 243.880 ;
        RECT 530.910 243.820 531.230 243.880 ;
        RECT 530.910 155.280 531.230 155.340 ;
        RECT 835.430 155.280 835.750 155.340 ;
        RECT 530.910 155.140 835.750 155.280 ;
        RECT 530.910 155.080 531.230 155.140 ;
        RECT 835.430 155.080 835.750 155.140 ;
      LAYER via ;
        RECT 527.260 243.820 527.520 244.080 ;
        RECT 530.940 243.820 531.200 244.080 ;
        RECT 530.940 155.080 531.200 155.340 ;
        RECT 835.460 155.080 835.720 155.340 ;
      LAYER met2 ;
        RECT 527.210 260.000 527.490 264.000 ;
        RECT 527.320 244.110 527.460 260.000 ;
        RECT 527.260 243.790 527.520 244.110 ;
        RECT 530.940 243.790 531.200 244.110 ;
        RECT 531.000 155.370 531.140 243.790 ;
        RECT 530.940 155.050 531.200 155.370 ;
        RECT 835.460 155.050 835.720 155.370 ;
        RECT 835.520 2.400 835.660 155.050 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2475.790 244.020 2476.110 244.080 ;
        RECT 2480.390 244.020 2480.710 244.080 ;
        RECT 2475.790 243.880 2480.710 244.020 ;
        RECT 2475.790 243.820 2476.110 243.880 ;
        RECT 2480.390 243.820 2480.710 243.880 ;
        RECT 2480.390 51.580 2480.710 51.640 ;
        RECT 2774.330 51.580 2774.650 51.640 ;
        RECT 2480.390 51.440 2774.650 51.580 ;
        RECT 2480.390 51.380 2480.710 51.440 ;
        RECT 2774.330 51.380 2774.650 51.440 ;
      LAYER via ;
        RECT 2475.820 243.820 2476.080 244.080 ;
        RECT 2480.420 243.820 2480.680 244.080 ;
        RECT 2480.420 51.380 2480.680 51.640 ;
        RECT 2774.360 51.380 2774.620 51.640 ;
      LAYER met2 ;
        RECT 2475.770 260.000 2476.050 264.000 ;
        RECT 2475.880 244.110 2476.020 260.000 ;
        RECT 2475.820 243.790 2476.080 244.110 ;
        RECT 2480.420 243.790 2480.680 244.110 ;
        RECT 2480.480 51.670 2480.620 243.790 ;
        RECT 2480.420 51.350 2480.680 51.670 ;
        RECT 2774.360 51.350 2774.620 51.670 ;
        RECT 2774.420 17.410 2774.560 51.350 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2493.270 244.020 2493.590 244.080 ;
        RECT 2497.410 244.020 2497.730 244.080 ;
        RECT 2493.270 243.880 2497.730 244.020 ;
        RECT 2493.270 243.820 2493.590 243.880 ;
        RECT 2497.410 243.820 2497.730 243.880 ;
        RECT 2497.410 58.720 2497.730 58.780 ;
        RECT 2794.570 58.720 2794.890 58.780 ;
        RECT 2497.410 58.580 2794.890 58.720 ;
        RECT 2497.410 58.520 2497.730 58.580 ;
        RECT 2794.570 58.520 2794.890 58.580 ;
      LAYER via ;
        RECT 2493.300 243.820 2493.560 244.080 ;
        RECT 2497.440 243.820 2497.700 244.080 ;
        RECT 2497.440 58.520 2497.700 58.780 ;
        RECT 2794.600 58.520 2794.860 58.780 ;
      LAYER met2 ;
        RECT 2493.250 260.000 2493.530 264.000 ;
        RECT 2493.360 244.110 2493.500 260.000 ;
        RECT 2493.300 243.790 2493.560 244.110 ;
        RECT 2497.440 243.790 2497.700 244.110 ;
        RECT 2497.500 58.810 2497.640 243.790 ;
        RECT 2497.440 58.490 2497.700 58.810 ;
        RECT 2794.600 58.490 2794.860 58.810 ;
        RECT 2794.660 17.410 2794.800 58.490 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2510.750 168.880 2511.070 168.940 ;
        RECT 2815.730 168.880 2816.050 168.940 ;
        RECT 2510.750 168.740 2816.050 168.880 ;
        RECT 2510.750 168.680 2511.070 168.740 ;
        RECT 2815.730 168.680 2816.050 168.740 ;
      LAYER via ;
        RECT 2510.780 168.680 2511.040 168.940 ;
        RECT 2815.760 168.680 2816.020 168.940 ;
      LAYER met2 ;
        RECT 2511.190 260.170 2511.470 264.000 ;
        RECT 2510.840 260.030 2511.470 260.170 ;
        RECT 2510.840 168.970 2510.980 260.030 ;
        RECT 2511.190 260.000 2511.470 260.030 ;
        RECT 2510.780 168.650 2511.040 168.970 ;
        RECT 2815.760 168.650 2816.020 168.970 ;
        RECT 2815.820 2.400 2815.960 168.650 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2531.910 65.860 2532.230 65.920 ;
        RECT 2829.070 65.860 2829.390 65.920 ;
        RECT 2531.910 65.720 2829.390 65.860 ;
        RECT 2531.910 65.660 2532.230 65.720 ;
        RECT 2829.070 65.660 2829.390 65.720 ;
      LAYER via ;
        RECT 2531.940 65.660 2532.200 65.920 ;
        RECT 2829.100 65.660 2829.360 65.920 ;
      LAYER met2 ;
        RECT 2529.130 260.170 2529.410 264.000 ;
        RECT 2529.130 260.030 2532.140 260.170 ;
        RECT 2529.130 260.000 2529.410 260.030 ;
        RECT 2532.000 65.950 2532.140 260.030 ;
        RECT 2531.940 65.630 2532.200 65.950 ;
        RECT 2829.100 65.630 2829.360 65.950 ;
        RECT 2829.160 17.410 2829.300 65.630 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2547.090 244.020 2547.410 244.080 ;
        RECT 2552.610 244.020 2552.930 244.080 ;
        RECT 2547.090 243.880 2552.930 244.020 ;
        RECT 2547.090 243.820 2547.410 243.880 ;
        RECT 2552.610 243.820 2552.930 243.880 ;
        RECT 2552.610 155.280 2552.930 155.340 ;
        RECT 2849.770 155.280 2850.090 155.340 ;
        RECT 2552.610 155.140 2850.090 155.280 ;
        RECT 2552.610 155.080 2552.930 155.140 ;
        RECT 2849.770 155.080 2850.090 155.140 ;
      LAYER via ;
        RECT 2547.120 243.820 2547.380 244.080 ;
        RECT 2552.640 243.820 2552.900 244.080 ;
        RECT 2552.640 155.080 2552.900 155.340 ;
        RECT 2849.800 155.080 2850.060 155.340 ;
      LAYER met2 ;
        RECT 2547.070 260.000 2547.350 264.000 ;
        RECT 2547.180 244.110 2547.320 260.000 ;
        RECT 2547.120 243.790 2547.380 244.110 ;
        RECT 2552.640 243.790 2552.900 244.110 ;
        RECT 2552.700 155.370 2552.840 243.790 ;
        RECT 2552.640 155.050 2552.900 155.370 ;
        RECT 2849.800 155.050 2850.060 155.370 ;
        RECT 2849.860 17.410 2850.000 155.050 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2566.410 15.880 2566.730 15.940 ;
        RECT 2869.090 15.880 2869.410 15.940 ;
        RECT 2566.410 15.740 2869.410 15.880 ;
        RECT 2566.410 15.680 2566.730 15.740 ;
        RECT 2869.090 15.680 2869.410 15.740 ;
      LAYER via ;
        RECT 2566.440 15.680 2566.700 15.940 ;
        RECT 2869.120 15.680 2869.380 15.940 ;
      LAYER met2 ;
        RECT 2565.010 260.170 2565.290 264.000 ;
        RECT 2565.010 260.030 2566.640 260.170 ;
        RECT 2565.010 260.000 2565.290 260.030 ;
        RECT 2566.500 15.970 2566.640 260.030 ;
        RECT 2566.440 15.650 2566.700 15.970 ;
        RECT 2869.120 15.650 2869.380 15.970 ;
        RECT 2869.180 2.400 2869.320 15.650 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2582.970 244.020 2583.290 244.080 ;
        RECT 2587.110 244.020 2587.430 244.080 ;
        RECT 2582.970 243.880 2587.430 244.020 ;
        RECT 2582.970 243.820 2583.290 243.880 ;
        RECT 2587.110 243.820 2587.430 243.880 ;
        RECT 2587.110 16.900 2587.430 16.960 ;
        RECT 2887.030 16.900 2887.350 16.960 ;
        RECT 2587.110 16.760 2887.350 16.900 ;
        RECT 2587.110 16.700 2587.430 16.760 ;
        RECT 2887.030 16.700 2887.350 16.760 ;
      LAYER via ;
        RECT 2583.000 243.820 2583.260 244.080 ;
        RECT 2587.140 243.820 2587.400 244.080 ;
        RECT 2587.140 16.700 2587.400 16.960 ;
        RECT 2887.060 16.700 2887.320 16.960 ;
      LAYER met2 ;
        RECT 2582.950 260.000 2583.230 264.000 ;
        RECT 2583.060 244.110 2583.200 260.000 ;
        RECT 2583.000 243.790 2583.260 244.110 ;
        RECT 2587.140 243.790 2587.400 244.110 ;
        RECT 2587.200 16.990 2587.340 243.790 ;
        RECT 2587.140 16.670 2587.400 16.990 ;
        RECT 2887.060 16.670 2887.320 16.990 ;
        RECT 2887.120 2.400 2887.260 16.670 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2600.890 260.000 2601.170 264.000 ;
        RECT 2601.000 16.845 2601.140 260.000 ;
        RECT 2600.930 16.475 2601.210 16.845 ;
        RECT 2904.990 16.475 2905.270 16.845 ;
        RECT 2905.060 2.400 2905.200 16.475 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2600.930 16.520 2601.210 16.800 ;
        RECT 2904.990 16.520 2905.270 16.800 ;
      LAYER met3 ;
        RECT 2600.905 16.810 2601.235 16.825 ;
        RECT 2904.965 16.810 2905.295 16.825 ;
        RECT 2600.905 16.510 2905.295 16.810 ;
        RECT 2600.905 16.495 2601.235 16.510 ;
        RECT 2904.965 16.495 2905.295 16.510 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 545.170 244.020 545.490 244.080 ;
        RECT 551.150 244.020 551.470 244.080 ;
        RECT 545.170 243.880 551.470 244.020 ;
        RECT 545.170 243.820 545.490 243.880 ;
        RECT 551.150 243.820 551.470 243.880 ;
        RECT 551.150 31.180 551.470 31.240 ;
        RECT 852.910 31.180 853.230 31.240 ;
        RECT 551.150 31.040 853.230 31.180 ;
        RECT 551.150 30.980 551.470 31.040 ;
        RECT 852.910 30.980 853.230 31.040 ;
      LAYER via ;
        RECT 545.200 243.820 545.460 244.080 ;
        RECT 551.180 243.820 551.440 244.080 ;
        RECT 551.180 30.980 551.440 31.240 ;
        RECT 852.940 30.980 853.200 31.240 ;
      LAYER met2 ;
        RECT 545.150 260.000 545.430 264.000 ;
        RECT 545.260 244.110 545.400 260.000 ;
        RECT 545.200 243.790 545.460 244.110 ;
        RECT 551.180 243.790 551.440 244.110 ;
        RECT 551.240 31.270 551.380 243.790 ;
        RECT 551.180 30.950 551.440 31.270 ;
        RECT 852.940 30.950 853.200 31.270 ;
        RECT 853.000 2.400 853.140 30.950 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 563.110 231.100 563.430 231.160 ;
        RECT 869.470 231.100 869.790 231.160 ;
        RECT 563.110 230.960 869.790 231.100 ;
        RECT 563.110 230.900 563.430 230.960 ;
        RECT 869.470 230.900 869.790 230.960 ;
      LAYER via ;
        RECT 563.140 230.900 563.400 231.160 ;
        RECT 869.500 230.900 869.760 231.160 ;
      LAYER met2 ;
        RECT 563.090 260.000 563.370 264.000 ;
        RECT 563.200 231.190 563.340 260.000 ;
        RECT 563.140 230.870 563.400 231.190 ;
        RECT 869.500 230.870 869.760 231.190 ;
        RECT 869.560 16.730 869.700 230.870 ;
        RECT 869.560 16.590 871.080 16.730 ;
        RECT 870.940 2.400 871.080 16.590 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 580.590 244.020 580.910 244.080 ;
        RECT 586.110 244.020 586.430 244.080 ;
        RECT 580.590 243.880 586.430 244.020 ;
        RECT 580.590 243.820 580.910 243.880 ;
        RECT 586.110 243.820 586.430 243.880 ;
        RECT 586.110 224.300 586.430 224.360 ;
        RECT 883.270 224.300 883.590 224.360 ;
        RECT 586.110 224.160 883.590 224.300 ;
        RECT 586.110 224.100 586.430 224.160 ;
        RECT 883.270 224.100 883.590 224.160 ;
      LAYER via ;
        RECT 580.620 243.820 580.880 244.080 ;
        RECT 586.140 243.820 586.400 244.080 ;
        RECT 586.140 224.100 586.400 224.360 ;
        RECT 883.300 224.100 883.560 224.360 ;
      LAYER met2 ;
        RECT 580.570 260.000 580.850 264.000 ;
        RECT 580.680 244.110 580.820 260.000 ;
        RECT 580.620 243.790 580.880 244.110 ;
        RECT 586.140 243.790 586.400 244.110 ;
        RECT 586.200 224.390 586.340 243.790 ;
        RECT 586.140 224.070 586.400 224.390 ;
        RECT 883.300 224.070 883.560 224.390 ;
        RECT 883.360 16.730 883.500 224.070 ;
        RECT 883.360 16.590 889.020 16.730 ;
        RECT 888.880 2.400 889.020 16.590 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 599.910 162.080 600.230 162.140 ;
        RECT 903.970 162.080 904.290 162.140 ;
        RECT 599.910 161.940 904.290 162.080 ;
        RECT 599.910 161.880 600.230 161.940 ;
        RECT 903.970 161.880 904.290 161.940 ;
      LAYER via ;
        RECT 599.940 161.880 600.200 162.140 ;
        RECT 904.000 161.880 904.260 162.140 ;
      LAYER met2 ;
        RECT 598.510 260.170 598.790 264.000 ;
        RECT 598.510 260.030 600.140 260.170 ;
        RECT 598.510 260.000 598.790 260.030 ;
        RECT 600.000 162.170 600.140 260.030 ;
        RECT 599.940 161.850 600.200 162.170 ;
        RECT 904.000 161.850 904.260 162.170 ;
        RECT 904.060 16.730 904.200 161.850 ;
        RECT 904.060 16.590 906.960 16.730 ;
        RECT 906.820 2.400 906.960 16.590 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 616.470 243.680 616.790 243.740 ;
        RECT 620.610 243.680 620.930 243.740 ;
        RECT 616.470 243.540 620.930 243.680 ;
        RECT 616.470 243.480 616.790 243.540 ;
        RECT 620.610 243.480 620.930 243.540 ;
        RECT 620.610 169.220 620.930 169.280 ;
        RECT 917.770 169.220 918.090 169.280 ;
        RECT 620.610 169.080 918.090 169.220 ;
        RECT 620.610 169.020 620.930 169.080 ;
        RECT 917.770 169.020 918.090 169.080 ;
        RECT 917.770 18.260 918.090 18.320 ;
        RECT 924.210 18.260 924.530 18.320 ;
        RECT 917.770 18.120 924.530 18.260 ;
        RECT 917.770 18.060 918.090 18.120 ;
        RECT 924.210 18.060 924.530 18.120 ;
      LAYER via ;
        RECT 616.500 243.480 616.760 243.740 ;
        RECT 620.640 243.480 620.900 243.740 ;
        RECT 620.640 169.020 620.900 169.280 ;
        RECT 917.800 169.020 918.060 169.280 ;
        RECT 917.800 18.060 918.060 18.320 ;
        RECT 924.240 18.060 924.500 18.320 ;
      LAYER met2 ;
        RECT 616.450 260.000 616.730 264.000 ;
        RECT 616.560 243.770 616.700 260.000 ;
        RECT 616.500 243.450 616.760 243.770 ;
        RECT 620.640 243.450 620.900 243.770 ;
        RECT 620.700 169.310 620.840 243.450 ;
        RECT 620.640 168.990 620.900 169.310 ;
        RECT 917.800 168.990 918.060 169.310 ;
        RECT 917.860 18.350 918.000 168.990 ;
        RECT 917.800 18.030 918.060 18.350 ;
        RECT 924.240 18.030 924.500 18.350 ;
        RECT 924.300 2.400 924.440 18.030 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 634.410 24.040 634.730 24.100 ;
        RECT 942.150 24.040 942.470 24.100 ;
        RECT 634.410 23.900 942.470 24.040 ;
        RECT 634.410 23.840 634.730 23.900 ;
        RECT 942.150 23.840 942.470 23.900 ;
      LAYER via ;
        RECT 634.440 23.840 634.700 24.100 ;
        RECT 942.180 23.840 942.440 24.100 ;
      LAYER met2 ;
        RECT 634.390 260.000 634.670 264.000 ;
        RECT 634.500 24.130 634.640 260.000 ;
        RECT 634.440 23.810 634.700 24.130 ;
        RECT 942.180 23.810 942.440 24.130 ;
        RECT 942.240 2.400 942.380 23.810 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 655.110 176.020 655.430 176.080 ;
        RECT 959.170 176.020 959.490 176.080 ;
        RECT 655.110 175.880 959.490 176.020 ;
        RECT 655.110 175.820 655.430 175.880 ;
        RECT 959.170 175.820 959.490 175.880 ;
      LAYER via ;
        RECT 655.140 175.820 655.400 176.080 ;
        RECT 959.200 175.820 959.460 176.080 ;
      LAYER met2 ;
        RECT 652.330 260.170 652.610 264.000 ;
        RECT 652.330 260.030 655.340 260.170 ;
        RECT 652.330 260.000 652.610 260.030 ;
        RECT 655.200 176.110 655.340 260.030 ;
        RECT 655.140 175.790 655.400 176.110 ;
        RECT 959.200 175.790 959.460 176.110 ;
        RECT 959.260 16.730 959.400 175.790 ;
        RECT 959.260 16.590 960.320 16.730 ;
        RECT 960.180 2.400 960.320 16.590 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 670.290 244.020 670.610 244.080 ;
        RECT 675.810 244.020 676.130 244.080 ;
        RECT 670.290 243.880 676.130 244.020 ;
        RECT 670.290 243.820 670.610 243.880 ;
        RECT 675.810 243.820 676.130 243.880 ;
        RECT 675.810 217.500 676.130 217.560 ;
        RECT 972.970 217.500 973.290 217.560 ;
        RECT 675.810 217.360 973.290 217.500 ;
        RECT 675.810 217.300 676.130 217.360 ;
        RECT 972.970 217.300 973.290 217.360 ;
      LAYER via ;
        RECT 670.320 243.820 670.580 244.080 ;
        RECT 675.840 243.820 676.100 244.080 ;
        RECT 675.840 217.300 676.100 217.560 ;
        RECT 973.000 217.300 973.260 217.560 ;
      LAYER met2 ;
        RECT 670.270 260.000 670.550 264.000 ;
        RECT 670.380 244.110 670.520 260.000 ;
        RECT 670.320 243.790 670.580 244.110 ;
        RECT 675.840 243.790 676.100 244.110 ;
        RECT 675.900 217.590 676.040 243.790 ;
        RECT 675.840 217.270 676.100 217.590 ;
        RECT 973.000 217.270 973.260 217.590 ;
        RECT 973.060 16.730 973.200 217.270 ;
        RECT 973.060 16.590 978.260 16.730 ;
        RECT 978.120 2.400 978.260 16.590 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 351.510 86.260 351.830 86.320 ;
        RECT 655.570 86.260 655.890 86.320 ;
        RECT 351.510 86.120 655.890 86.260 ;
        RECT 351.510 86.060 351.830 86.120 ;
        RECT 655.570 86.060 655.890 86.120 ;
      LAYER via ;
        RECT 351.540 86.060 351.800 86.320 ;
        RECT 655.600 86.060 655.860 86.320 ;
      LAYER met2 ;
        RECT 348.270 260.170 348.550 264.000 ;
        RECT 348.270 260.030 351.740 260.170 ;
        RECT 348.270 260.000 348.550 260.030 ;
        RECT 351.600 86.350 351.740 260.030 ;
        RECT 351.540 86.030 351.800 86.350 ;
        RECT 655.600 86.030 655.860 86.350 ;
        RECT 655.660 17.410 655.800 86.030 ;
        RECT 655.660 17.270 657.180 17.410 ;
        RECT 657.040 2.400 657.180 17.270 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.610 182.820 689.930 182.880 ;
        RECT 993.670 182.820 993.990 182.880 ;
        RECT 689.610 182.680 993.990 182.820 ;
        RECT 689.610 182.620 689.930 182.680 ;
        RECT 993.670 182.620 993.990 182.680 ;
      LAYER via ;
        RECT 689.640 182.620 689.900 182.880 ;
        RECT 993.700 182.620 993.960 182.880 ;
      LAYER met2 ;
        RECT 688.210 260.170 688.490 264.000 ;
        RECT 688.210 260.030 689.840 260.170 ;
        RECT 688.210 260.000 688.490 260.030 ;
        RECT 689.700 182.910 689.840 260.030 ;
        RECT 689.640 182.590 689.900 182.910 ;
        RECT 993.700 182.590 993.960 182.910 ;
        RECT 993.760 16.730 993.900 182.590 ;
        RECT 993.760 16.590 996.200 16.730 ;
        RECT 996.060 2.400 996.200 16.590 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 705.710 244.020 706.030 244.080 ;
        RECT 710.310 244.020 710.630 244.080 ;
        RECT 705.710 243.880 710.630 244.020 ;
        RECT 705.710 243.820 706.030 243.880 ;
        RECT 710.310 243.820 710.630 243.880 ;
        RECT 710.310 189.960 710.630 190.020 ;
        RECT 1007.470 189.960 1007.790 190.020 ;
        RECT 710.310 189.820 1007.790 189.960 ;
        RECT 710.310 189.760 710.630 189.820 ;
        RECT 1007.470 189.760 1007.790 189.820 ;
        RECT 1007.470 19.280 1007.790 19.340 ;
        RECT 1013.450 19.280 1013.770 19.340 ;
        RECT 1007.470 19.140 1013.770 19.280 ;
        RECT 1007.470 19.080 1007.790 19.140 ;
        RECT 1013.450 19.080 1013.770 19.140 ;
      LAYER via ;
        RECT 705.740 243.820 706.000 244.080 ;
        RECT 710.340 243.820 710.600 244.080 ;
        RECT 710.340 189.760 710.600 190.020 ;
        RECT 1007.500 189.760 1007.760 190.020 ;
        RECT 1007.500 19.080 1007.760 19.340 ;
        RECT 1013.480 19.080 1013.740 19.340 ;
      LAYER met2 ;
        RECT 705.690 260.000 705.970 264.000 ;
        RECT 705.800 244.110 705.940 260.000 ;
        RECT 705.740 243.790 706.000 244.110 ;
        RECT 710.340 243.790 710.600 244.110 ;
        RECT 710.400 190.050 710.540 243.790 ;
        RECT 710.340 189.730 710.600 190.050 ;
        RECT 1007.500 189.730 1007.760 190.050 ;
        RECT 1007.560 19.370 1007.700 189.730 ;
        RECT 1007.500 19.050 1007.760 19.370 ;
        RECT 1013.480 19.050 1013.740 19.370 ;
        RECT 1013.540 2.400 1013.680 19.050 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 723.650 141.340 723.970 141.400 ;
        RECT 1028.170 141.340 1028.490 141.400 ;
        RECT 723.650 141.200 1028.490 141.340 ;
        RECT 723.650 141.140 723.970 141.200 ;
        RECT 1028.170 141.140 1028.490 141.200 ;
      LAYER via ;
        RECT 723.680 141.140 723.940 141.400 ;
        RECT 1028.200 141.140 1028.460 141.400 ;
      LAYER met2 ;
        RECT 723.630 260.000 723.910 264.000 ;
        RECT 723.740 141.430 723.880 260.000 ;
        RECT 723.680 141.110 723.940 141.430 ;
        RECT 1028.200 141.110 1028.460 141.430 ;
        RECT 1028.260 16.730 1028.400 141.110 ;
        RECT 1028.260 16.590 1031.620 16.730 ;
        RECT 1031.480 2.400 1031.620 16.590 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 744.810 210.360 745.130 210.420 ;
        RECT 1049.330 210.360 1049.650 210.420 ;
        RECT 744.810 210.220 1049.650 210.360 ;
        RECT 744.810 210.160 745.130 210.220 ;
        RECT 1049.330 210.160 1049.650 210.220 ;
      LAYER via ;
        RECT 744.840 210.160 745.100 210.420 ;
        RECT 1049.360 210.160 1049.620 210.420 ;
      LAYER met2 ;
        RECT 741.570 260.170 741.850 264.000 ;
        RECT 741.570 260.030 745.040 260.170 ;
        RECT 741.570 260.000 741.850 260.030 ;
        RECT 744.900 210.450 745.040 260.030 ;
        RECT 744.840 210.130 745.100 210.450 ;
        RECT 1049.360 210.130 1049.620 210.450 ;
        RECT 1049.420 2.400 1049.560 210.130 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 759.530 244.020 759.850 244.080 ;
        RECT 769.190 244.020 769.510 244.080 ;
        RECT 759.530 243.880 769.510 244.020 ;
        RECT 759.530 243.820 759.850 243.880 ;
        RECT 769.190 243.820 769.510 243.880 ;
        RECT 769.190 196.760 769.510 196.820 ;
        RECT 1062.670 196.760 1062.990 196.820 ;
        RECT 769.190 196.620 1062.990 196.760 ;
        RECT 769.190 196.560 769.510 196.620 ;
        RECT 1062.670 196.560 1062.990 196.620 ;
      LAYER via ;
        RECT 759.560 243.820 759.820 244.080 ;
        RECT 769.220 243.820 769.480 244.080 ;
        RECT 769.220 196.560 769.480 196.820 ;
        RECT 1062.700 196.560 1062.960 196.820 ;
      LAYER met2 ;
        RECT 759.510 260.000 759.790 264.000 ;
        RECT 759.620 244.110 759.760 260.000 ;
        RECT 759.560 243.790 759.820 244.110 ;
        RECT 769.220 243.790 769.480 244.110 ;
        RECT 769.280 196.850 769.420 243.790 ;
        RECT 769.220 196.530 769.480 196.850 ;
        RECT 1062.700 196.530 1062.960 196.850 ;
        RECT 1062.760 16.730 1062.900 196.530 ;
        RECT 1062.760 16.590 1067.500 16.730 ;
        RECT 1067.360 2.400 1067.500 16.590 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 779.310 148.480 779.630 148.540 ;
        RECT 1083.370 148.480 1083.690 148.540 ;
        RECT 779.310 148.340 1083.690 148.480 ;
        RECT 779.310 148.280 779.630 148.340 ;
        RECT 1083.370 148.280 1083.690 148.340 ;
      LAYER via ;
        RECT 779.340 148.280 779.600 148.540 ;
        RECT 1083.400 148.280 1083.660 148.540 ;
      LAYER met2 ;
        RECT 777.450 260.170 777.730 264.000 ;
        RECT 777.450 260.030 779.540 260.170 ;
        RECT 777.450 260.000 777.730 260.030 ;
        RECT 779.400 148.570 779.540 260.030 ;
        RECT 779.340 148.250 779.600 148.570 ;
        RECT 1083.400 148.250 1083.660 148.570 ;
        RECT 1083.460 16.730 1083.600 148.250 ;
        RECT 1083.460 16.590 1085.440 16.730 ;
        RECT 1085.300 2.400 1085.440 16.590 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 795.410 244.020 795.730 244.080 ;
        RECT 800.010 244.020 800.330 244.080 ;
        RECT 795.410 243.880 800.330 244.020 ;
        RECT 795.410 243.820 795.730 243.880 ;
        RECT 800.010 243.820 800.330 243.880 ;
        RECT 800.010 155.620 800.330 155.680 ;
        RECT 1097.170 155.620 1097.490 155.680 ;
        RECT 800.010 155.480 1097.490 155.620 ;
        RECT 800.010 155.420 800.330 155.480 ;
        RECT 1097.170 155.420 1097.490 155.480 ;
      LAYER via ;
        RECT 795.440 243.820 795.700 244.080 ;
        RECT 800.040 243.820 800.300 244.080 ;
        RECT 800.040 155.420 800.300 155.680 ;
        RECT 1097.200 155.420 1097.460 155.680 ;
      LAYER met2 ;
        RECT 795.390 260.000 795.670 264.000 ;
        RECT 795.500 244.110 795.640 260.000 ;
        RECT 795.440 243.790 795.700 244.110 ;
        RECT 800.040 243.790 800.300 244.110 ;
        RECT 800.100 155.710 800.240 243.790 ;
        RECT 800.040 155.390 800.300 155.710 ;
        RECT 1097.200 155.390 1097.460 155.710 ;
        RECT 1097.260 16.730 1097.400 155.390 ;
        RECT 1097.260 16.590 1102.920 16.730 ;
        RECT 1102.780 2.400 1102.920 16.590 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 813.810 203.560 814.130 203.620 ;
        RECT 1117.870 203.560 1118.190 203.620 ;
        RECT 813.810 203.420 1118.190 203.560 ;
        RECT 813.810 203.360 814.130 203.420 ;
        RECT 1117.870 203.360 1118.190 203.420 ;
      LAYER via ;
        RECT 813.840 203.360 814.100 203.620 ;
        RECT 1117.900 203.360 1118.160 203.620 ;
      LAYER met2 ;
        RECT 813.330 260.170 813.610 264.000 ;
        RECT 813.330 260.030 814.040 260.170 ;
        RECT 813.330 260.000 813.610 260.030 ;
        RECT 813.900 203.650 814.040 260.030 ;
        RECT 813.840 203.330 814.100 203.650 ;
        RECT 1117.900 203.330 1118.160 203.650 ;
        RECT 1117.960 16.730 1118.100 203.330 ;
        RECT 1117.960 16.590 1120.860 16.730 ;
        RECT 1120.720 2.400 1120.860 16.590 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 830.830 244.020 831.150 244.080 ;
        RECT 838.650 244.020 838.970 244.080 ;
        RECT 830.830 243.880 838.970 244.020 ;
        RECT 830.830 243.820 831.150 243.880 ;
        RECT 838.650 243.820 838.970 243.880 ;
        RECT 838.650 162.420 838.970 162.480 ;
        RECT 1139.030 162.420 1139.350 162.480 ;
        RECT 838.650 162.280 1139.350 162.420 ;
        RECT 838.650 162.220 838.970 162.280 ;
        RECT 1139.030 162.220 1139.350 162.280 ;
      LAYER via ;
        RECT 830.860 243.820 831.120 244.080 ;
        RECT 838.680 243.820 838.940 244.080 ;
        RECT 838.680 162.220 838.940 162.480 ;
        RECT 1139.060 162.220 1139.320 162.480 ;
      LAYER met2 ;
        RECT 830.810 260.000 831.090 264.000 ;
        RECT 830.920 244.110 831.060 260.000 ;
        RECT 830.860 243.790 831.120 244.110 ;
        RECT 838.680 243.790 838.940 244.110 ;
        RECT 838.740 162.510 838.880 243.790 ;
        RECT 838.680 162.190 838.940 162.510 ;
        RECT 1139.060 162.190 1139.320 162.510 ;
        RECT 1139.120 17.410 1139.260 162.190 ;
        RECT 1138.660 17.270 1139.260 17.410 ;
        RECT 1138.660 2.400 1138.800 17.270 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 848.770 248.440 849.090 248.500 ;
        RECT 861.650 248.440 861.970 248.500 ;
        RECT 848.770 248.300 861.970 248.440 ;
        RECT 848.770 248.240 849.090 248.300 ;
        RECT 861.650 248.240 861.970 248.300 ;
        RECT 861.650 231.440 861.970 231.500 ;
        RECT 1152.370 231.440 1152.690 231.500 ;
        RECT 861.650 231.300 1152.690 231.440 ;
        RECT 861.650 231.240 861.970 231.300 ;
        RECT 1152.370 231.240 1152.690 231.300 ;
      LAYER via ;
        RECT 848.800 248.240 849.060 248.500 ;
        RECT 861.680 248.240 861.940 248.500 ;
        RECT 861.680 231.240 861.940 231.500 ;
        RECT 1152.400 231.240 1152.660 231.500 ;
      LAYER met2 ;
        RECT 848.750 260.000 849.030 264.000 ;
        RECT 848.860 248.530 849.000 260.000 ;
        RECT 848.800 248.210 849.060 248.530 ;
        RECT 861.680 248.210 861.940 248.530 ;
        RECT 861.740 231.530 861.880 248.210 ;
        RECT 861.680 231.210 861.940 231.530 ;
        RECT 1152.400 231.210 1152.660 231.530 ;
        RECT 1152.460 17.410 1152.600 231.210 ;
        RECT 1152.460 17.270 1156.740 17.410 ;
        RECT 1156.600 2.400 1156.740 17.270 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 366.230 244.020 366.550 244.080 ;
        RECT 372.210 244.020 372.530 244.080 ;
        RECT 366.230 243.880 372.530 244.020 ;
        RECT 366.230 243.820 366.550 243.880 ;
        RECT 372.210 243.820 372.530 243.880 ;
        RECT 372.210 72.660 372.530 72.720 ;
        RECT 669.370 72.660 669.690 72.720 ;
        RECT 372.210 72.520 669.690 72.660 ;
        RECT 372.210 72.460 372.530 72.520 ;
        RECT 669.370 72.460 669.690 72.520 ;
      LAYER via ;
        RECT 366.260 243.820 366.520 244.080 ;
        RECT 372.240 243.820 372.500 244.080 ;
        RECT 372.240 72.460 372.500 72.720 ;
        RECT 669.400 72.460 669.660 72.720 ;
      LAYER met2 ;
        RECT 366.210 260.000 366.490 264.000 ;
        RECT 366.320 244.110 366.460 260.000 ;
        RECT 366.260 243.790 366.520 244.110 ;
        RECT 372.240 243.790 372.500 244.110 ;
        RECT 372.300 72.750 372.440 243.790 ;
        RECT 372.240 72.430 372.500 72.750 ;
        RECT 669.400 72.430 669.660 72.750 ;
        RECT 669.460 16.730 669.600 72.430 ;
        RECT 669.460 16.590 674.660 16.730 ;
        RECT 674.520 2.400 674.660 16.590 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 869.010 168.880 869.330 168.940 ;
        RECT 1173.070 168.880 1173.390 168.940 ;
        RECT 869.010 168.740 1173.390 168.880 ;
        RECT 869.010 168.680 869.330 168.740 ;
        RECT 1173.070 168.680 1173.390 168.740 ;
      LAYER via ;
        RECT 869.040 168.680 869.300 168.940 ;
        RECT 1173.100 168.680 1173.360 168.940 ;
      LAYER met2 ;
        RECT 866.690 260.170 866.970 264.000 ;
        RECT 866.690 260.030 869.240 260.170 ;
        RECT 866.690 260.000 866.970 260.030 ;
        RECT 869.100 168.970 869.240 260.030 ;
        RECT 869.040 168.650 869.300 168.970 ;
        RECT 1173.100 168.650 1173.360 168.970 ;
        RECT 1173.160 17.410 1173.300 168.650 ;
        RECT 1173.160 17.270 1174.220 17.410 ;
        RECT 1174.080 2.400 1174.220 17.270 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 884.650 244.020 884.970 244.080 ;
        RECT 889.710 244.020 890.030 244.080 ;
        RECT 884.650 243.880 890.030 244.020 ;
        RECT 884.650 243.820 884.970 243.880 ;
        RECT 889.710 243.820 890.030 243.880 ;
        RECT 889.710 224.300 890.030 224.360 ;
        RECT 1186.870 224.300 1187.190 224.360 ;
        RECT 889.710 224.160 1187.190 224.300 ;
        RECT 889.710 224.100 890.030 224.160 ;
        RECT 1186.870 224.100 1187.190 224.160 ;
      LAYER via ;
        RECT 884.680 243.820 884.940 244.080 ;
        RECT 889.740 243.820 890.000 244.080 ;
        RECT 889.740 224.100 890.000 224.360 ;
        RECT 1186.900 224.100 1187.160 224.360 ;
      LAYER met2 ;
        RECT 884.630 260.000 884.910 264.000 ;
        RECT 884.740 244.110 884.880 260.000 ;
        RECT 884.680 243.790 884.940 244.110 ;
        RECT 889.740 243.790 890.000 244.110 ;
        RECT 889.800 224.390 889.940 243.790 ;
        RECT 889.740 224.070 890.000 224.390 ;
        RECT 1186.900 224.070 1187.160 224.390 ;
        RECT 1186.960 17.410 1187.100 224.070 ;
        RECT 1186.960 17.270 1192.160 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 903.510 30.840 903.830 30.900 ;
        RECT 1209.870 30.840 1210.190 30.900 ;
        RECT 903.510 30.700 1210.190 30.840 ;
        RECT 903.510 30.640 903.830 30.700 ;
        RECT 1209.870 30.640 1210.190 30.700 ;
      LAYER via ;
        RECT 903.540 30.640 903.800 30.900 ;
        RECT 1209.900 30.640 1210.160 30.900 ;
      LAYER met2 ;
        RECT 902.570 260.170 902.850 264.000 ;
        RECT 902.570 260.030 903.740 260.170 ;
        RECT 902.570 260.000 902.850 260.030 ;
        RECT 903.600 30.930 903.740 260.030 ;
        RECT 903.540 30.610 903.800 30.930 ;
        RECT 1209.900 30.610 1210.160 30.930 ;
        RECT 1209.960 2.400 1210.100 30.610 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 176.360 924.530 176.420 ;
        RECT 1221.370 176.360 1221.690 176.420 ;
        RECT 924.210 176.220 1221.690 176.360 ;
        RECT 924.210 176.160 924.530 176.220 ;
        RECT 1221.370 176.160 1221.690 176.220 ;
        RECT 1221.370 37.640 1221.690 37.700 ;
        RECT 1227.810 37.640 1228.130 37.700 ;
        RECT 1221.370 37.500 1228.130 37.640 ;
        RECT 1221.370 37.440 1221.690 37.500 ;
        RECT 1227.810 37.440 1228.130 37.500 ;
      LAYER via ;
        RECT 924.240 176.160 924.500 176.420 ;
        RECT 1221.400 176.160 1221.660 176.420 ;
        RECT 1221.400 37.440 1221.660 37.700 ;
        RECT 1227.840 37.440 1228.100 37.700 ;
      LAYER met2 ;
        RECT 920.510 260.170 920.790 264.000 ;
        RECT 920.510 260.030 924.440 260.170 ;
        RECT 920.510 260.000 920.790 260.030 ;
        RECT 924.300 176.450 924.440 260.030 ;
        RECT 924.240 176.130 924.500 176.450 ;
        RECT 1221.400 176.130 1221.660 176.450 ;
        RECT 1221.460 37.730 1221.600 176.130 ;
        RECT 1221.400 37.410 1221.660 37.730 ;
        RECT 1227.840 37.410 1228.100 37.730 ;
        RECT 1227.900 2.400 1228.040 37.410 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1242.145 48.365 1242.315 96.475 ;
      LAYER mcon ;
        RECT 1242.145 96.305 1242.315 96.475 ;
      LAYER met1 ;
        RECT 938.470 244.020 938.790 244.080 ;
        RECT 948.590 244.020 948.910 244.080 ;
        RECT 938.470 243.880 948.910 244.020 ;
        RECT 938.470 243.820 938.790 243.880 ;
        RECT 948.590 243.820 948.910 243.880 ;
        RECT 948.590 183.160 948.910 183.220 ;
        RECT 1242.070 183.160 1242.390 183.220 ;
        RECT 948.590 183.020 1242.390 183.160 ;
        RECT 948.590 182.960 948.910 183.020 ;
        RECT 1242.070 182.960 1242.390 183.020 ;
        RECT 1242.070 144.740 1242.390 144.800 ;
        RECT 1242.530 144.740 1242.850 144.800 ;
        RECT 1242.070 144.600 1242.850 144.740 ;
        RECT 1242.070 144.540 1242.390 144.600 ;
        RECT 1242.530 144.540 1242.850 144.600 ;
        RECT 1242.070 96.460 1242.390 96.520 ;
        RECT 1241.875 96.320 1242.390 96.460 ;
        RECT 1242.070 96.260 1242.390 96.320 ;
        RECT 1242.085 48.520 1242.375 48.565 ;
        RECT 1245.750 48.520 1246.070 48.580 ;
        RECT 1242.085 48.380 1246.070 48.520 ;
        RECT 1242.085 48.335 1242.375 48.380 ;
        RECT 1245.750 48.320 1246.070 48.380 ;
      LAYER via ;
        RECT 938.500 243.820 938.760 244.080 ;
        RECT 948.620 243.820 948.880 244.080 ;
        RECT 948.620 182.960 948.880 183.220 ;
        RECT 1242.100 182.960 1242.360 183.220 ;
        RECT 1242.100 144.540 1242.360 144.800 ;
        RECT 1242.560 144.540 1242.820 144.800 ;
        RECT 1242.100 96.260 1242.360 96.520 ;
        RECT 1245.780 48.320 1246.040 48.580 ;
      LAYER met2 ;
        RECT 938.450 260.000 938.730 264.000 ;
        RECT 938.560 244.110 938.700 260.000 ;
        RECT 938.500 243.790 938.760 244.110 ;
        RECT 948.620 243.790 948.880 244.110 ;
        RECT 948.680 183.250 948.820 243.790 ;
        RECT 948.620 182.930 948.880 183.250 ;
        RECT 1242.100 182.930 1242.360 183.250 ;
        RECT 1242.160 144.830 1242.300 182.930 ;
        RECT 1242.100 144.510 1242.360 144.830 ;
        RECT 1242.560 144.510 1242.820 144.830 ;
        RECT 1242.620 96.970 1242.760 144.510 ;
        RECT 1242.160 96.830 1242.760 96.970 ;
        RECT 1242.160 96.550 1242.300 96.830 ;
        RECT 1242.100 96.230 1242.360 96.550 ;
        RECT 1245.780 48.290 1246.040 48.610 ;
        RECT 1245.840 2.400 1245.980 48.290 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 958.710 217.160 959.030 217.220 ;
        RECT 1263.230 217.160 1263.550 217.220 ;
        RECT 958.710 217.020 1263.550 217.160 ;
        RECT 958.710 216.960 959.030 217.020 ;
        RECT 1263.230 216.960 1263.550 217.020 ;
      LAYER via ;
        RECT 958.740 216.960 959.000 217.220 ;
        RECT 1263.260 216.960 1263.520 217.220 ;
      LAYER met2 ;
        RECT 955.930 260.170 956.210 264.000 ;
        RECT 955.930 260.030 958.940 260.170 ;
        RECT 955.930 260.000 956.210 260.030 ;
        RECT 958.800 217.250 958.940 260.030 ;
        RECT 958.740 216.930 959.000 217.250 ;
        RECT 1263.260 216.930 1263.520 217.250 ;
        RECT 1263.320 2.400 1263.460 216.930 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 973.890 238.580 974.210 238.640 ;
        RECT 1276.570 238.580 1276.890 238.640 ;
        RECT 973.890 238.440 1276.890 238.580 ;
        RECT 973.890 238.380 974.210 238.440 ;
        RECT 1276.570 238.380 1276.890 238.440 ;
        RECT 1276.570 62.120 1276.890 62.180 ;
        RECT 1281.170 62.120 1281.490 62.180 ;
        RECT 1276.570 61.980 1281.490 62.120 ;
        RECT 1276.570 61.920 1276.890 61.980 ;
        RECT 1281.170 61.920 1281.490 61.980 ;
      LAYER via ;
        RECT 973.920 238.380 974.180 238.640 ;
        RECT 1276.600 238.380 1276.860 238.640 ;
        RECT 1276.600 61.920 1276.860 62.180 ;
        RECT 1281.200 61.920 1281.460 62.180 ;
      LAYER met2 ;
        RECT 973.870 260.000 974.150 264.000 ;
        RECT 973.980 238.670 974.120 260.000 ;
        RECT 973.920 238.350 974.180 238.670 ;
        RECT 1276.600 238.350 1276.860 238.670 ;
        RECT 1276.660 62.210 1276.800 238.350 ;
        RECT 1276.600 61.890 1276.860 62.210 ;
        RECT 1281.200 61.890 1281.460 62.210 ;
        RECT 1281.260 2.400 1281.400 61.890 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1297.345 48.365 1297.515 96.475 ;
      LAYER mcon ;
        RECT 1297.345 96.305 1297.515 96.475 ;
      LAYER met1 ;
        RECT 993.210 189.620 993.530 189.680 ;
        RECT 1297.270 189.620 1297.590 189.680 ;
        RECT 993.210 189.480 1297.590 189.620 ;
        RECT 993.210 189.420 993.530 189.480 ;
        RECT 1297.270 189.420 1297.590 189.480 ;
        RECT 1297.270 96.460 1297.590 96.520 ;
        RECT 1297.075 96.320 1297.590 96.460 ;
        RECT 1297.270 96.260 1297.590 96.320 ;
        RECT 1297.285 48.520 1297.575 48.565 ;
        RECT 1299.110 48.520 1299.430 48.580 ;
        RECT 1297.285 48.380 1299.430 48.520 ;
        RECT 1297.285 48.335 1297.575 48.380 ;
        RECT 1299.110 48.320 1299.430 48.380 ;
      LAYER via ;
        RECT 993.240 189.420 993.500 189.680 ;
        RECT 1297.300 189.420 1297.560 189.680 ;
        RECT 1297.300 96.260 1297.560 96.520 ;
        RECT 1299.140 48.320 1299.400 48.580 ;
      LAYER met2 ;
        RECT 991.810 260.170 992.090 264.000 ;
        RECT 991.810 260.030 993.440 260.170 ;
        RECT 991.810 260.000 992.090 260.030 ;
        RECT 993.300 189.710 993.440 260.030 ;
        RECT 993.240 189.390 993.500 189.710 ;
        RECT 1297.300 189.390 1297.560 189.710 ;
        RECT 1297.360 96.550 1297.500 189.390 ;
        RECT 1297.300 96.230 1297.560 96.550 ;
        RECT 1299.140 48.290 1299.400 48.610 ;
        RECT 1299.200 2.400 1299.340 48.290 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1009.770 244.020 1010.090 244.080 ;
        RECT 1013.910 244.020 1014.230 244.080 ;
        RECT 1009.770 243.880 1014.230 244.020 ;
        RECT 1009.770 243.820 1010.090 243.880 ;
        RECT 1013.910 243.820 1014.230 243.880 ;
        RECT 1013.910 210.700 1014.230 210.760 ;
        RECT 1311.070 210.700 1311.390 210.760 ;
        RECT 1013.910 210.560 1311.390 210.700 ;
        RECT 1013.910 210.500 1014.230 210.560 ;
        RECT 1311.070 210.500 1311.390 210.560 ;
        RECT 1311.070 37.640 1311.390 37.700 ;
        RECT 1317.050 37.640 1317.370 37.700 ;
        RECT 1311.070 37.500 1317.370 37.640 ;
        RECT 1311.070 37.440 1311.390 37.500 ;
        RECT 1317.050 37.440 1317.370 37.500 ;
      LAYER via ;
        RECT 1009.800 243.820 1010.060 244.080 ;
        RECT 1013.940 243.820 1014.200 244.080 ;
        RECT 1013.940 210.500 1014.200 210.760 ;
        RECT 1311.100 210.500 1311.360 210.760 ;
        RECT 1311.100 37.440 1311.360 37.700 ;
        RECT 1317.080 37.440 1317.340 37.700 ;
      LAYER met2 ;
        RECT 1009.750 260.000 1010.030 264.000 ;
        RECT 1009.860 244.110 1010.000 260.000 ;
        RECT 1009.800 243.790 1010.060 244.110 ;
        RECT 1013.940 243.790 1014.200 244.110 ;
        RECT 1014.000 210.790 1014.140 243.790 ;
        RECT 1013.940 210.470 1014.200 210.790 ;
        RECT 1311.100 210.470 1311.360 210.790 ;
        RECT 1311.160 37.730 1311.300 210.470 ;
        RECT 1311.100 37.410 1311.360 37.730 ;
        RECT 1317.080 37.410 1317.340 37.730 ;
        RECT 1317.140 2.400 1317.280 37.410 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1027.250 148.140 1027.570 148.200 ;
        RECT 1331.770 148.140 1332.090 148.200 ;
        RECT 1027.250 148.000 1332.090 148.140 ;
        RECT 1027.250 147.940 1027.570 148.000 ;
        RECT 1331.770 147.940 1332.090 148.000 ;
        RECT 1331.770 62.120 1332.090 62.180 ;
        RECT 1334.990 62.120 1335.310 62.180 ;
        RECT 1331.770 61.980 1335.310 62.120 ;
        RECT 1331.770 61.920 1332.090 61.980 ;
        RECT 1334.990 61.920 1335.310 61.980 ;
      LAYER via ;
        RECT 1027.280 147.940 1027.540 148.200 ;
        RECT 1331.800 147.940 1332.060 148.200 ;
        RECT 1331.800 61.920 1332.060 62.180 ;
        RECT 1335.020 61.920 1335.280 62.180 ;
      LAYER met2 ;
        RECT 1027.690 260.170 1027.970 264.000 ;
        RECT 1027.340 260.030 1027.970 260.170 ;
        RECT 1027.340 148.230 1027.480 260.030 ;
        RECT 1027.690 260.000 1027.970 260.030 ;
        RECT 1027.280 147.910 1027.540 148.230 ;
        RECT 1331.800 147.910 1332.060 148.230 ;
        RECT 1331.860 62.210 1332.000 147.910 ;
        RECT 1331.800 61.890 1332.060 62.210 ;
        RECT 1335.020 61.890 1335.280 62.210 ;
        RECT 1335.080 2.400 1335.220 61.890 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 384.170 244.020 384.490 244.080 ;
        RECT 389.690 244.020 390.010 244.080 ;
        RECT 384.170 243.880 390.010 244.020 ;
        RECT 384.170 243.820 384.490 243.880 ;
        RECT 389.690 243.820 390.010 243.880 ;
        RECT 389.690 189.620 390.010 189.680 ;
        RECT 690.070 189.620 690.390 189.680 ;
        RECT 389.690 189.480 690.390 189.620 ;
        RECT 389.690 189.420 390.010 189.480 ;
        RECT 690.070 189.420 690.390 189.480 ;
      LAYER via ;
        RECT 384.200 243.820 384.460 244.080 ;
        RECT 389.720 243.820 389.980 244.080 ;
        RECT 389.720 189.420 389.980 189.680 ;
        RECT 690.100 189.420 690.360 189.680 ;
      LAYER met2 ;
        RECT 384.150 260.000 384.430 264.000 ;
        RECT 384.260 244.110 384.400 260.000 ;
        RECT 384.200 243.790 384.460 244.110 ;
        RECT 389.720 243.790 389.980 244.110 ;
        RECT 389.780 189.710 389.920 243.790 ;
        RECT 389.720 189.390 389.980 189.710 ;
        RECT 690.100 189.390 690.360 189.710 ;
        RECT 690.160 16.730 690.300 189.390 ;
        RECT 690.160 16.590 692.600 16.730 ;
        RECT 692.460 2.400 692.600 16.590 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1048.410 24.380 1048.730 24.440 ;
        RECT 1352.930 24.380 1353.250 24.440 ;
        RECT 1048.410 24.240 1353.250 24.380 ;
        RECT 1048.410 24.180 1048.730 24.240 ;
        RECT 1352.930 24.180 1353.250 24.240 ;
      LAYER via ;
        RECT 1048.440 24.180 1048.700 24.440 ;
        RECT 1352.960 24.180 1353.220 24.440 ;
      LAYER met2 ;
        RECT 1045.630 260.170 1045.910 264.000 ;
        RECT 1045.630 260.030 1048.640 260.170 ;
        RECT 1045.630 260.000 1045.910 260.030 ;
        RECT 1048.500 24.470 1048.640 260.030 ;
        RECT 1048.440 24.150 1048.700 24.470 ;
        RECT 1352.960 24.150 1353.220 24.470 ;
        RECT 1353.020 13.330 1353.160 24.150 ;
        RECT 1352.560 13.190 1353.160 13.330 ;
        RECT 1352.560 2.400 1352.700 13.190 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1063.590 244.020 1063.910 244.080 ;
        RECT 1069.110 244.020 1069.430 244.080 ;
        RECT 1063.590 243.880 1069.430 244.020 ;
        RECT 1063.590 243.820 1063.910 243.880 ;
        RECT 1069.110 243.820 1069.430 243.880 ;
        RECT 1069.110 196.760 1069.430 196.820 ;
        RECT 1366.270 196.760 1366.590 196.820 ;
        RECT 1069.110 196.620 1366.590 196.760 ;
        RECT 1069.110 196.560 1069.430 196.620 ;
        RECT 1366.270 196.560 1366.590 196.620 ;
        RECT 1366.270 62.120 1366.590 62.180 ;
        RECT 1370.410 62.120 1370.730 62.180 ;
        RECT 1366.270 61.980 1370.730 62.120 ;
        RECT 1366.270 61.920 1366.590 61.980 ;
        RECT 1370.410 61.920 1370.730 61.980 ;
      LAYER via ;
        RECT 1063.620 243.820 1063.880 244.080 ;
        RECT 1069.140 243.820 1069.400 244.080 ;
        RECT 1069.140 196.560 1069.400 196.820 ;
        RECT 1366.300 196.560 1366.560 196.820 ;
        RECT 1366.300 61.920 1366.560 62.180 ;
        RECT 1370.440 61.920 1370.700 62.180 ;
      LAYER met2 ;
        RECT 1063.570 260.000 1063.850 264.000 ;
        RECT 1063.680 244.110 1063.820 260.000 ;
        RECT 1063.620 243.790 1063.880 244.110 ;
        RECT 1069.140 243.790 1069.400 244.110 ;
        RECT 1069.200 196.850 1069.340 243.790 ;
        RECT 1069.140 196.530 1069.400 196.850 ;
        RECT 1366.300 196.530 1366.560 196.850 ;
        RECT 1366.360 62.210 1366.500 196.530 ;
        RECT 1366.300 61.890 1366.560 62.210 ;
        RECT 1370.440 61.890 1370.700 62.210 ;
        RECT 1370.500 2.400 1370.640 61.890 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1082.910 155.280 1083.230 155.340 ;
        RECT 1386.970 155.280 1387.290 155.340 ;
        RECT 1082.910 155.140 1387.290 155.280 ;
        RECT 1082.910 155.080 1083.230 155.140 ;
        RECT 1386.970 155.080 1387.290 155.140 ;
        RECT 1386.970 96.460 1387.290 96.520 ;
        RECT 1388.810 96.460 1389.130 96.520 ;
        RECT 1386.970 96.320 1389.130 96.460 ;
        RECT 1386.970 96.260 1387.290 96.320 ;
        RECT 1388.810 96.260 1389.130 96.320 ;
      LAYER via ;
        RECT 1082.940 155.080 1083.200 155.340 ;
        RECT 1387.000 155.080 1387.260 155.340 ;
        RECT 1387.000 96.260 1387.260 96.520 ;
        RECT 1388.840 96.260 1389.100 96.520 ;
      LAYER met2 ;
        RECT 1081.050 260.170 1081.330 264.000 ;
        RECT 1081.050 260.030 1083.140 260.170 ;
        RECT 1081.050 260.000 1081.330 260.030 ;
        RECT 1083.000 155.370 1083.140 260.030 ;
        RECT 1082.940 155.050 1083.200 155.370 ;
        RECT 1387.000 155.050 1387.260 155.370 ;
        RECT 1387.060 96.550 1387.200 155.050 ;
        RECT 1387.000 96.230 1387.260 96.550 ;
        RECT 1388.840 96.230 1389.100 96.550 ;
        RECT 1388.900 24.380 1389.040 96.230 ;
        RECT 1388.440 24.240 1389.040 24.380 ;
        RECT 1388.440 2.400 1388.580 24.240 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1099.010 244.020 1099.330 244.080 ;
        RECT 1103.610 244.020 1103.930 244.080 ;
        RECT 1099.010 243.880 1103.930 244.020 ;
        RECT 1099.010 243.820 1099.330 243.880 ;
        RECT 1103.610 243.820 1103.930 243.880 ;
        RECT 1103.610 203.900 1103.930 203.960 ;
        RECT 1400.770 203.900 1401.090 203.960 ;
        RECT 1103.610 203.760 1401.090 203.900 ;
        RECT 1103.610 203.700 1103.930 203.760 ;
        RECT 1400.770 203.700 1401.090 203.760 ;
        RECT 1400.770 62.120 1401.090 62.180 ;
        RECT 1406.290 62.120 1406.610 62.180 ;
        RECT 1400.770 61.980 1406.610 62.120 ;
        RECT 1400.770 61.920 1401.090 61.980 ;
        RECT 1406.290 61.920 1406.610 61.980 ;
      LAYER via ;
        RECT 1099.040 243.820 1099.300 244.080 ;
        RECT 1103.640 243.820 1103.900 244.080 ;
        RECT 1103.640 203.700 1103.900 203.960 ;
        RECT 1400.800 203.700 1401.060 203.960 ;
        RECT 1400.800 61.920 1401.060 62.180 ;
        RECT 1406.320 61.920 1406.580 62.180 ;
      LAYER met2 ;
        RECT 1098.990 260.000 1099.270 264.000 ;
        RECT 1099.100 244.110 1099.240 260.000 ;
        RECT 1099.040 243.790 1099.300 244.110 ;
        RECT 1103.640 243.790 1103.900 244.110 ;
        RECT 1103.700 203.990 1103.840 243.790 ;
        RECT 1103.640 203.670 1103.900 203.990 ;
        RECT 1400.800 203.670 1401.060 203.990 ;
        RECT 1400.860 62.210 1401.000 203.670 ;
        RECT 1400.800 61.890 1401.060 62.210 ;
        RECT 1406.320 61.890 1406.580 62.210 ;
        RECT 1406.380 2.400 1406.520 61.890 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1421.545 48.365 1421.715 96.475 ;
      LAYER mcon ;
        RECT 1421.545 96.305 1421.715 96.475 ;
      LAYER met1 ;
        RECT 1116.950 162.080 1117.270 162.140 ;
        RECT 1421.470 162.080 1421.790 162.140 ;
        RECT 1116.950 161.940 1421.790 162.080 ;
        RECT 1116.950 161.880 1117.270 161.940 ;
        RECT 1421.470 161.880 1421.790 161.940 ;
        RECT 1421.470 96.460 1421.790 96.520 ;
        RECT 1421.275 96.320 1421.790 96.460 ;
        RECT 1421.470 96.260 1421.790 96.320 ;
        RECT 1421.485 48.520 1421.775 48.565 ;
        RECT 1423.770 48.520 1424.090 48.580 ;
        RECT 1421.485 48.380 1424.090 48.520 ;
        RECT 1421.485 48.335 1421.775 48.380 ;
        RECT 1423.770 48.320 1424.090 48.380 ;
      LAYER via ;
        RECT 1116.980 161.880 1117.240 162.140 ;
        RECT 1421.500 161.880 1421.760 162.140 ;
        RECT 1421.500 96.260 1421.760 96.520 ;
        RECT 1423.800 48.320 1424.060 48.580 ;
      LAYER met2 ;
        RECT 1116.930 260.000 1117.210 264.000 ;
        RECT 1117.040 162.170 1117.180 260.000 ;
        RECT 1116.980 161.850 1117.240 162.170 ;
        RECT 1421.500 161.850 1421.760 162.170 ;
        RECT 1421.560 96.550 1421.700 161.850 ;
        RECT 1421.500 96.230 1421.760 96.550 ;
        RECT 1423.800 48.290 1424.060 48.610 ;
        RECT 1423.860 2.400 1424.000 48.290 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1138.110 169.220 1138.430 169.280 ;
        RECT 1435.270 169.220 1435.590 169.280 ;
        RECT 1138.110 169.080 1435.590 169.220 ;
        RECT 1138.110 169.020 1138.430 169.080 ;
        RECT 1435.270 169.020 1435.590 169.080 ;
        RECT 1435.270 38.320 1435.590 38.380 ;
        RECT 1441.710 38.320 1442.030 38.380 ;
        RECT 1435.270 38.180 1442.030 38.320 ;
        RECT 1435.270 38.120 1435.590 38.180 ;
        RECT 1441.710 38.120 1442.030 38.180 ;
      LAYER via ;
        RECT 1138.140 169.020 1138.400 169.280 ;
        RECT 1435.300 169.020 1435.560 169.280 ;
        RECT 1435.300 38.120 1435.560 38.380 ;
        RECT 1441.740 38.120 1442.000 38.380 ;
      LAYER met2 ;
        RECT 1134.870 260.170 1135.150 264.000 ;
        RECT 1134.870 260.030 1138.340 260.170 ;
        RECT 1134.870 260.000 1135.150 260.030 ;
        RECT 1138.200 169.310 1138.340 260.030 ;
        RECT 1138.140 168.990 1138.400 169.310 ;
        RECT 1435.300 168.990 1435.560 169.310 ;
        RECT 1435.360 38.410 1435.500 168.990 ;
        RECT 1435.300 38.090 1435.560 38.410 ;
        RECT 1441.740 38.090 1442.000 38.410 ;
        RECT 1441.800 2.400 1441.940 38.090 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1152.830 231.100 1153.150 231.160 ;
        RECT 1455.970 231.100 1456.290 231.160 ;
        RECT 1152.830 230.960 1456.290 231.100 ;
        RECT 1152.830 230.900 1153.150 230.960 ;
        RECT 1455.970 230.900 1456.290 230.960 ;
        RECT 1455.970 62.120 1456.290 62.180 ;
        RECT 1459.650 62.120 1459.970 62.180 ;
        RECT 1455.970 61.980 1459.970 62.120 ;
        RECT 1455.970 61.920 1456.290 61.980 ;
        RECT 1459.650 61.920 1459.970 61.980 ;
      LAYER via ;
        RECT 1152.860 230.900 1153.120 231.160 ;
        RECT 1456.000 230.900 1456.260 231.160 ;
        RECT 1456.000 61.920 1456.260 62.180 ;
        RECT 1459.680 61.920 1459.940 62.180 ;
      LAYER met2 ;
        RECT 1152.810 260.000 1153.090 264.000 ;
        RECT 1152.920 231.190 1153.060 260.000 ;
        RECT 1152.860 230.870 1153.120 231.190 ;
        RECT 1456.000 230.870 1456.260 231.190 ;
        RECT 1456.060 62.210 1456.200 230.870 ;
        RECT 1456.000 61.890 1456.260 62.210 ;
        RECT 1459.680 61.890 1459.940 62.210 ;
        RECT 1459.740 2.400 1459.880 61.890 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1172.610 37.980 1172.930 38.040 ;
        RECT 1477.590 37.980 1477.910 38.040 ;
        RECT 1172.610 37.840 1477.910 37.980 ;
        RECT 1172.610 37.780 1172.930 37.840 ;
        RECT 1477.590 37.780 1477.910 37.840 ;
      LAYER via ;
        RECT 1172.640 37.780 1172.900 38.040 ;
        RECT 1477.620 37.780 1477.880 38.040 ;
      LAYER met2 ;
        RECT 1170.750 260.170 1171.030 264.000 ;
        RECT 1170.750 260.030 1172.840 260.170 ;
        RECT 1170.750 260.000 1171.030 260.030 ;
        RECT 1172.700 38.070 1172.840 260.030 ;
        RECT 1172.640 37.750 1172.900 38.070 ;
        RECT 1477.620 37.750 1477.880 38.070 ;
        RECT 1477.680 2.400 1477.820 37.750 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1188.710 244.020 1189.030 244.080 ;
        RECT 1193.310 244.020 1193.630 244.080 ;
        RECT 1188.710 243.880 1193.630 244.020 ;
        RECT 1188.710 243.820 1189.030 243.880 ;
        RECT 1193.310 243.820 1193.630 243.880 ;
        RECT 1193.310 224.640 1193.630 224.700 ;
        RECT 1490.470 224.640 1490.790 224.700 ;
        RECT 1193.310 224.500 1490.790 224.640 ;
        RECT 1193.310 224.440 1193.630 224.500 ;
        RECT 1490.470 224.440 1490.790 224.500 ;
        RECT 1490.470 62.120 1490.790 62.180 ;
        RECT 1495.530 62.120 1495.850 62.180 ;
        RECT 1490.470 61.980 1495.850 62.120 ;
        RECT 1490.470 61.920 1490.790 61.980 ;
        RECT 1495.530 61.920 1495.850 61.980 ;
      LAYER via ;
        RECT 1188.740 243.820 1189.000 244.080 ;
        RECT 1193.340 243.820 1193.600 244.080 ;
        RECT 1193.340 224.440 1193.600 224.700 ;
        RECT 1490.500 224.440 1490.760 224.700 ;
        RECT 1490.500 61.920 1490.760 62.180 ;
        RECT 1495.560 61.920 1495.820 62.180 ;
      LAYER met2 ;
        RECT 1188.690 260.000 1188.970 264.000 ;
        RECT 1188.800 244.110 1188.940 260.000 ;
        RECT 1188.740 243.790 1189.000 244.110 ;
        RECT 1193.340 243.790 1193.600 244.110 ;
        RECT 1193.400 224.730 1193.540 243.790 ;
        RECT 1193.340 224.410 1193.600 224.730 ;
        RECT 1490.500 224.410 1490.760 224.730 ;
        RECT 1490.560 62.210 1490.700 224.410 ;
        RECT 1490.500 61.890 1490.760 62.210 ;
        RECT 1495.560 61.890 1495.820 62.210 ;
        RECT 1495.620 2.400 1495.760 61.890 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1206.650 176.020 1206.970 176.080 ;
        RECT 1511.170 176.020 1511.490 176.080 ;
        RECT 1206.650 175.880 1511.490 176.020 ;
        RECT 1206.650 175.820 1206.970 175.880 ;
        RECT 1511.170 175.820 1511.490 175.880 ;
      LAYER via ;
        RECT 1206.680 175.820 1206.940 176.080 ;
        RECT 1511.200 175.820 1511.460 176.080 ;
      LAYER met2 ;
        RECT 1206.630 260.000 1206.910 264.000 ;
        RECT 1206.740 176.110 1206.880 260.000 ;
        RECT 1206.680 175.790 1206.940 176.110 ;
        RECT 1511.200 175.790 1511.460 176.110 ;
        RECT 1511.260 17.410 1511.400 175.790 ;
        RECT 1511.260 17.270 1513.240 17.410 ;
        RECT 1513.100 2.400 1513.240 17.270 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 402.110 244.020 402.430 244.080 ;
        RECT 410.390 244.020 410.710 244.080 ;
        RECT 402.110 243.880 410.710 244.020 ;
        RECT 402.110 243.820 402.430 243.880 ;
        RECT 410.390 243.820 410.710 243.880 ;
        RECT 410.390 196.760 410.710 196.820 ;
        RECT 703.870 196.760 704.190 196.820 ;
        RECT 410.390 196.620 704.190 196.760 ;
        RECT 410.390 196.560 410.710 196.620 ;
        RECT 703.870 196.560 704.190 196.620 ;
        RECT 703.870 17.240 704.190 17.300 ;
        RECT 710.310 17.240 710.630 17.300 ;
        RECT 703.870 17.100 710.630 17.240 ;
        RECT 703.870 17.040 704.190 17.100 ;
        RECT 710.310 17.040 710.630 17.100 ;
      LAYER via ;
        RECT 402.140 243.820 402.400 244.080 ;
        RECT 410.420 243.820 410.680 244.080 ;
        RECT 410.420 196.560 410.680 196.820 ;
        RECT 703.900 196.560 704.160 196.820 ;
        RECT 703.900 17.040 704.160 17.300 ;
        RECT 710.340 17.040 710.600 17.300 ;
      LAYER met2 ;
        RECT 402.090 260.000 402.370 264.000 ;
        RECT 402.200 244.110 402.340 260.000 ;
        RECT 402.140 243.790 402.400 244.110 ;
        RECT 410.420 243.790 410.680 244.110 ;
        RECT 410.480 196.850 410.620 243.790 ;
        RECT 410.420 196.530 410.680 196.850 ;
        RECT 703.900 196.530 704.160 196.850 ;
        RECT 703.960 17.330 704.100 196.530 ;
        RECT 703.900 17.010 704.160 17.330 ;
        RECT 710.340 17.010 710.600 17.330 ;
        RECT 710.400 2.400 710.540 17.010 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 182.820 1228.130 182.880 ;
        RECT 1524.970 182.820 1525.290 182.880 ;
        RECT 1227.810 182.680 1525.290 182.820 ;
        RECT 1227.810 182.620 1228.130 182.680 ;
        RECT 1524.970 182.620 1525.290 182.680 ;
        RECT 1524.970 17.580 1525.290 17.640 ;
        RECT 1530.950 17.580 1531.270 17.640 ;
        RECT 1524.970 17.440 1531.270 17.580 ;
        RECT 1524.970 17.380 1525.290 17.440 ;
        RECT 1530.950 17.380 1531.270 17.440 ;
      LAYER via ;
        RECT 1227.840 182.620 1228.100 182.880 ;
        RECT 1525.000 182.620 1525.260 182.880 ;
        RECT 1525.000 17.380 1525.260 17.640 ;
        RECT 1530.980 17.380 1531.240 17.640 ;
      LAYER met2 ;
        RECT 1224.110 260.170 1224.390 264.000 ;
        RECT 1224.110 260.030 1228.040 260.170 ;
        RECT 1224.110 260.000 1224.390 260.030 ;
        RECT 1227.900 182.910 1228.040 260.030 ;
        RECT 1227.840 182.590 1228.100 182.910 ;
        RECT 1525.000 182.590 1525.260 182.910 ;
        RECT 1525.060 17.670 1525.200 182.590 ;
        RECT 1525.000 17.350 1525.260 17.670 ;
        RECT 1530.980 17.350 1531.240 17.670 ;
        RECT 1531.040 2.400 1531.180 17.350 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1242.070 242.660 1242.390 242.720 ;
        RECT 1248.050 242.660 1248.370 242.720 ;
        RECT 1242.070 242.520 1248.370 242.660 ;
        RECT 1242.070 242.460 1242.390 242.520 ;
        RECT 1248.050 242.460 1248.370 242.520 ;
        RECT 1248.050 217.500 1248.370 217.560 ;
        RECT 1545.670 217.500 1545.990 217.560 ;
        RECT 1248.050 217.360 1545.990 217.500 ;
        RECT 1248.050 217.300 1248.370 217.360 ;
        RECT 1545.670 217.300 1545.990 217.360 ;
      LAYER via ;
        RECT 1242.100 242.460 1242.360 242.720 ;
        RECT 1248.080 242.460 1248.340 242.720 ;
        RECT 1248.080 217.300 1248.340 217.560 ;
        RECT 1545.700 217.300 1545.960 217.560 ;
      LAYER met2 ;
        RECT 1242.050 260.000 1242.330 264.000 ;
        RECT 1242.160 242.750 1242.300 260.000 ;
        RECT 1242.100 242.430 1242.360 242.750 ;
        RECT 1248.080 242.430 1248.340 242.750 ;
        RECT 1248.140 217.590 1248.280 242.430 ;
        RECT 1248.080 217.270 1248.340 217.590 ;
        RECT 1545.700 217.270 1545.960 217.590 ;
        RECT 1545.760 16.730 1545.900 217.270 ;
        RECT 1545.760 16.590 1549.120 16.730 ;
        RECT 1548.980 2.400 1549.120 16.590 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1262.310 30.840 1262.630 30.900 ;
        RECT 1566.830 30.840 1567.150 30.900 ;
        RECT 1262.310 30.700 1567.150 30.840 ;
        RECT 1262.310 30.640 1262.630 30.700 ;
        RECT 1566.830 30.640 1567.150 30.700 ;
      LAYER via ;
        RECT 1262.340 30.640 1262.600 30.900 ;
        RECT 1566.860 30.640 1567.120 30.900 ;
      LAYER met2 ;
        RECT 1259.990 260.170 1260.270 264.000 ;
        RECT 1259.990 260.030 1262.540 260.170 ;
        RECT 1259.990 260.000 1260.270 260.030 ;
        RECT 1262.400 30.930 1262.540 260.030 ;
        RECT 1262.340 30.610 1262.600 30.930 ;
        RECT 1566.860 30.610 1567.120 30.930 ;
        RECT 1566.920 2.400 1567.060 30.610 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1277.950 244.020 1278.270 244.080 ;
        RECT 1283.010 244.020 1283.330 244.080 ;
        RECT 1277.950 243.880 1283.330 244.020 ;
        RECT 1277.950 243.820 1278.270 243.880 ;
        RECT 1283.010 243.820 1283.330 243.880 ;
        RECT 1283.010 189.960 1283.330 190.020 ;
        RECT 1580.170 189.960 1580.490 190.020 ;
        RECT 1283.010 189.820 1580.490 189.960 ;
        RECT 1283.010 189.760 1283.330 189.820 ;
        RECT 1580.170 189.760 1580.490 189.820 ;
      LAYER via ;
        RECT 1277.980 243.820 1278.240 244.080 ;
        RECT 1283.040 243.820 1283.300 244.080 ;
        RECT 1283.040 189.760 1283.300 190.020 ;
        RECT 1580.200 189.760 1580.460 190.020 ;
      LAYER met2 ;
        RECT 1277.930 260.000 1278.210 264.000 ;
        RECT 1278.040 244.110 1278.180 260.000 ;
        RECT 1277.980 243.790 1278.240 244.110 ;
        RECT 1283.040 243.790 1283.300 244.110 ;
        RECT 1283.100 190.050 1283.240 243.790 ;
        RECT 1283.040 189.730 1283.300 190.050 ;
        RECT 1580.200 189.730 1580.460 190.050 ;
        RECT 1580.260 16.730 1580.400 189.730 ;
        RECT 1580.260 16.590 1585.000 16.730 ;
        RECT 1584.860 2.400 1585.000 16.590 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1296.810 148.480 1297.130 148.540 ;
        RECT 1600.870 148.480 1601.190 148.540 ;
        RECT 1296.810 148.340 1601.190 148.480 ;
        RECT 1296.810 148.280 1297.130 148.340 ;
        RECT 1600.870 148.280 1601.190 148.340 ;
      LAYER via ;
        RECT 1296.840 148.280 1297.100 148.540 ;
        RECT 1600.900 148.280 1601.160 148.540 ;
      LAYER met2 ;
        RECT 1295.870 260.170 1296.150 264.000 ;
        RECT 1295.870 260.030 1297.040 260.170 ;
        RECT 1295.870 260.000 1296.150 260.030 ;
        RECT 1296.900 148.570 1297.040 260.030 ;
        RECT 1296.840 148.250 1297.100 148.570 ;
        RECT 1600.900 148.250 1601.160 148.570 ;
        RECT 1600.960 16.730 1601.100 148.250 ;
        RECT 1600.960 16.590 1602.480 16.730 ;
        RECT 1602.340 2.400 1602.480 16.590 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1313.830 243.680 1314.150 243.740 ;
        RECT 1317.510 243.680 1317.830 243.740 ;
        RECT 1313.830 243.540 1317.830 243.680 ;
        RECT 1313.830 243.480 1314.150 243.540 ;
        RECT 1317.510 243.480 1317.830 243.540 ;
        RECT 1317.510 210.700 1317.830 210.760 ;
        RECT 1614.670 210.700 1614.990 210.760 ;
        RECT 1317.510 210.560 1614.990 210.700 ;
        RECT 1317.510 210.500 1317.830 210.560 ;
        RECT 1614.670 210.500 1614.990 210.560 ;
      LAYER via ;
        RECT 1313.860 243.480 1314.120 243.740 ;
        RECT 1317.540 243.480 1317.800 243.740 ;
        RECT 1317.540 210.500 1317.800 210.760 ;
        RECT 1614.700 210.500 1614.960 210.760 ;
      LAYER met2 ;
        RECT 1313.810 260.000 1314.090 264.000 ;
        RECT 1313.920 243.770 1314.060 260.000 ;
        RECT 1313.860 243.450 1314.120 243.770 ;
        RECT 1317.540 243.450 1317.800 243.770 ;
        RECT 1317.600 210.790 1317.740 243.450 ;
        RECT 1317.540 210.470 1317.800 210.790 ;
        RECT 1614.700 210.470 1614.960 210.790 ;
        RECT 1614.760 16.730 1614.900 210.470 ;
        RECT 1614.760 16.590 1620.420 16.730 ;
        RECT 1620.280 2.400 1620.420 16.590 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1331.770 244.020 1332.090 244.080 ;
        RECT 1337.750 244.020 1338.070 244.080 ;
        RECT 1331.770 243.880 1338.070 244.020 ;
        RECT 1331.770 243.820 1332.090 243.880 ;
        RECT 1337.750 243.820 1338.070 243.880 ;
        RECT 1337.750 155.620 1338.070 155.680 ;
        RECT 1635.370 155.620 1635.690 155.680 ;
        RECT 1337.750 155.480 1635.690 155.620 ;
        RECT 1337.750 155.420 1338.070 155.480 ;
        RECT 1635.370 155.420 1635.690 155.480 ;
      LAYER via ;
        RECT 1331.800 243.820 1332.060 244.080 ;
        RECT 1337.780 243.820 1338.040 244.080 ;
        RECT 1337.780 155.420 1338.040 155.680 ;
        RECT 1635.400 155.420 1635.660 155.680 ;
      LAYER met2 ;
        RECT 1331.750 260.000 1332.030 264.000 ;
        RECT 1331.860 244.110 1332.000 260.000 ;
        RECT 1331.800 243.790 1332.060 244.110 ;
        RECT 1337.780 243.790 1338.040 244.110 ;
        RECT 1337.840 155.710 1337.980 243.790 ;
        RECT 1337.780 155.390 1338.040 155.710 ;
        RECT 1635.400 155.390 1635.660 155.710 ;
        RECT 1635.460 16.730 1635.600 155.390 ;
        RECT 1635.460 16.590 1638.360 16.730 ;
        RECT 1638.220 2.400 1638.360 16.590 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.010 24.040 1352.330 24.100 ;
        RECT 1656.530 24.040 1656.850 24.100 ;
        RECT 1352.010 23.900 1656.850 24.040 ;
        RECT 1352.010 23.840 1352.330 23.900 ;
        RECT 1656.530 23.840 1656.850 23.900 ;
      LAYER via ;
        RECT 1352.040 23.840 1352.300 24.100 ;
        RECT 1656.560 23.840 1656.820 24.100 ;
      LAYER met2 ;
        RECT 1349.230 260.170 1349.510 264.000 ;
        RECT 1349.230 260.030 1352.240 260.170 ;
        RECT 1349.230 260.000 1349.510 260.030 ;
        RECT 1352.100 24.130 1352.240 260.030 ;
        RECT 1352.040 23.810 1352.300 24.130 ;
        RECT 1656.560 23.810 1656.820 24.130 ;
        RECT 1656.620 16.730 1656.760 23.810 ;
        RECT 1656.160 16.590 1656.760 16.730 ;
        RECT 1656.160 2.400 1656.300 16.590 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1367.190 244.020 1367.510 244.080 ;
        RECT 1372.710 244.020 1373.030 244.080 ;
        RECT 1367.190 243.880 1373.030 244.020 ;
        RECT 1367.190 243.820 1367.510 243.880 ;
        RECT 1372.710 243.820 1373.030 243.880 ;
        RECT 1372.710 197.100 1373.030 197.160 ;
        RECT 1669.870 197.100 1670.190 197.160 ;
        RECT 1372.710 196.960 1670.190 197.100 ;
        RECT 1372.710 196.900 1373.030 196.960 ;
        RECT 1669.870 196.900 1670.190 196.960 ;
      LAYER via ;
        RECT 1367.220 243.820 1367.480 244.080 ;
        RECT 1372.740 243.820 1373.000 244.080 ;
        RECT 1372.740 196.900 1373.000 197.160 ;
        RECT 1669.900 196.900 1670.160 197.160 ;
      LAYER met2 ;
        RECT 1367.170 260.000 1367.450 264.000 ;
        RECT 1367.280 244.110 1367.420 260.000 ;
        RECT 1367.220 243.790 1367.480 244.110 ;
        RECT 1372.740 243.790 1373.000 244.110 ;
        RECT 1372.800 197.190 1372.940 243.790 ;
        RECT 1372.740 196.870 1373.000 197.190 ;
        RECT 1669.900 196.870 1670.160 197.190 ;
        RECT 1669.960 16.730 1670.100 196.870 ;
        RECT 1669.960 16.590 1673.780 16.730 ;
        RECT 1673.640 2.400 1673.780 16.590 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1386.510 203.560 1386.830 203.620 ;
        RECT 1690.570 203.560 1690.890 203.620 ;
        RECT 1386.510 203.420 1690.890 203.560 ;
        RECT 1386.510 203.360 1386.830 203.420 ;
        RECT 1690.570 203.360 1690.890 203.420 ;
      LAYER via ;
        RECT 1386.540 203.360 1386.800 203.620 ;
        RECT 1690.600 203.360 1690.860 203.620 ;
      LAYER met2 ;
        RECT 1385.110 260.170 1385.390 264.000 ;
        RECT 1385.110 260.030 1386.740 260.170 ;
        RECT 1385.110 260.000 1385.390 260.030 ;
        RECT 1386.600 203.650 1386.740 260.030 ;
        RECT 1386.540 203.330 1386.800 203.650 ;
        RECT 1690.600 203.330 1690.860 203.650 ;
        RECT 1690.660 16.730 1690.800 203.330 ;
        RECT 1690.660 16.590 1691.720 16.730 ;
        RECT 1691.580 2.400 1691.720 16.590 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 420.510 210.360 420.830 210.420 ;
        RECT 724.570 210.360 724.890 210.420 ;
        RECT 420.510 210.220 724.890 210.360 ;
        RECT 420.510 210.160 420.830 210.220 ;
        RECT 724.570 210.160 724.890 210.220 ;
      LAYER via ;
        RECT 420.540 210.160 420.800 210.420 ;
        RECT 724.600 210.160 724.860 210.420 ;
      LAYER met2 ;
        RECT 420.030 260.170 420.310 264.000 ;
        RECT 420.030 260.030 420.740 260.170 ;
        RECT 420.030 260.000 420.310 260.030 ;
        RECT 420.600 210.450 420.740 260.030 ;
        RECT 420.540 210.130 420.800 210.450 ;
        RECT 724.600 210.130 724.860 210.450 ;
        RECT 724.660 16.730 724.800 210.130 ;
        RECT 724.660 16.590 728.480 16.730 ;
        RECT 728.340 2.400 728.480 16.590 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1403.070 244.020 1403.390 244.080 ;
        RECT 1407.210 244.020 1407.530 244.080 ;
        RECT 1403.070 243.880 1407.530 244.020 ;
        RECT 1403.070 243.820 1403.390 243.880 ;
        RECT 1407.210 243.820 1407.530 243.880 ;
        RECT 1407.210 162.420 1407.530 162.480 ;
        RECT 1704.370 162.420 1704.690 162.480 ;
        RECT 1407.210 162.280 1704.690 162.420 ;
        RECT 1407.210 162.220 1407.530 162.280 ;
        RECT 1704.370 162.220 1704.690 162.280 ;
      LAYER via ;
        RECT 1403.100 243.820 1403.360 244.080 ;
        RECT 1407.240 243.820 1407.500 244.080 ;
        RECT 1407.240 162.220 1407.500 162.480 ;
        RECT 1704.400 162.220 1704.660 162.480 ;
      LAYER met2 ;
        RECT 1403.050 260.000 1403.330 264.000 ;
        RECT 1403.160 244.110 1403.300 260.000 ;
        RECT 1403.100 243.790 1403.360 244.110 ;
        RECT 1407.240 243.790 1407.500 244.110 ;
        RECT 1407.300 162.510 1407.440 243.790 ;
        RECT 1407.240 162.190 1407.500 162.510 ;
        RECT 1704.400 162.190 1704.660 162.510 ;
        RECT 1704.460 16.730 1704.600 162.190 ;
        RECT 1704.460 16.590 1709.660 16.730 ;
        RECT 1709.520 2.400 1709.660 16.590 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1420.550 168.880 1420.870 168.940 ;
        RECT 1725.070 168.880 1725.390 168.940 ;
        RECT 1420.550 168.740 1725.390 168.880 ;
        RECT 1420.550 168.680 1420.870 168.740 ;
        RECT 1725.070 168.680 1725.390 168.740 ;
      LAYER via ;
        RECT 1420.580 168.680 1420.840 168.940 ;
        RECT 1725.100 168.680 1725.360 168.940 ;
      LAYER met2 ;
        RECT 1420.990 260.170 1421.270 264.000 ;
        RECT 1420.640 260.030 1421.270 260.170 ;
        RECT 1420.640 168.970 1420.780 260.030 ;
        RECT 1420.990 260.000 1421.270 260.030 ;
        RECT 1420.580 168.650 1420.840 168.970 ;
        RECT 1725.100 168.650 1725.360 168.970 ;
        RECT 1725.160 17.410 1725.300 168.650 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 176.360 1442.030 176.420 ;
        RECT 1738.870 176.360 1739.190 176.420 ;
        RECT 1441.710 176.220 1739.190 176.360 ;
        RECT 1441.710 176.160 1442.030 176.220 ;
        RECT 1738.870 176.160 1739.190 176.220 ;
        RECT 1738.870 17.580 1739.190 17.640 ;
        RECT 1745.310 17.580 1745.630 17.640 ;
        RECT 1738.870 17.440 1745.630 17.580 ;
        RECT 1738.870 17.380 1739.190 17.440 ;
        RECT 1745.310 17.380 1745.630 17.440 ;
      LAYER via ;
        RECT 1441.740 176.160 1442.000 176.420 ;
        RECT 1738.900 176.160 1739.160 176.420 ;
        RECT 1738.900 17.380 1739.160 17.640 ;
        RECT 1745.340 17.380 1745.600 17.640 ;
      LAYER met2 ;
        RECT 1438.930 260.170 1439.210 264.000 ;
        RECT 1438.930 260.030 1441.940 260.170 ;
        RECT 1438.930 260.000 1439.210 260.030 ;
        RECT 1441.800 176.450 1441.940 260.030 ;
        RECT 1441.740 176.130 1442.000 176.450 ;
        RECT 1738.900 176.130 1739.160 176.450 ;
        RECT 1738.960 17.670 1739.100 176.130 ;
        RECT 1738.900 17.350 1739.160 17.670 ;
        RECT 1745.340 17.350 1745.600 17.670 ;
        RECT 1745.400 2.400 1745.540 17.350 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1456.890 231.440 1457.210 231.500 ;
        RECT 1759.570 231.440 1759.890 231.500 ;
        RECT 1456.890 231.300 1759.890 231.440 ;
        RECT 1456.890 231.240 1457.210 231.300 ;
        RECT 1759.570 231.240 1759.890 231.300 ;
      LAYER via ;
        RECT 1456.920 231.240 1457.180 231.500 ;
        RECT 1759.600 231.240 1759.860 231.500 ;
      LAYER met2 ;
        RECT 1456.870 260.000 1457.150 264.000 ;
        RECT 1456.980 231.530 1457.120 260.000 ;
        RECT 1456.920 231.210 1457.180 231.530 ;
        RECT 1759.600 231.210 1759.860 231.530 ;
        RECT 1759.660 17.410 1759.800 231.210 ;
        RECT 1759.660 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1476.210 224.300 1476.530 224.360 ;
        RECT 1780.270 224.300 1780.590 224.360 ;
        RECT 1476.210 224.160 1780.590 224.300 ;
        RECT 1476.210 224.100 1476.530 224.160 ;
        RECT 1780.270 224.100 1780.590 224.160 ;
      LAYER via ;
        RECT 1476.240 224.100 1476.500 224.360 ;
        RECT 1780.300 224.100 1780.560 224.360 ;
      LAYER met2 ;
        RECT 1474.350 260.170 1474.630 264.000 ;
        RECT 1474.350 260.030 1476.440 260.170 ;
        RECT 1474.350 260.000 1474.630 260.030 ;
        RECT 1476.300 224.390 1476.440 260.030 ;
        RECT 1476.240 224.070 1476.500 224.390 ;
        RECT 1780.300 224.070 1780.560 224.390 ;
        RECT 1780.360 3.130 1780.500 224.070 ;
        RECT 1780.360 2.990 1780.960 3.130 ;
        RECT 1780.820 2.400 1780.960 2.990 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1492.310 244.020 1492.630 244.080 ;
        RECT 1496.910 244.020 1497.230 244.080 ;
        RECT 1492.310 243.880 1497.230 244.020 ;
        RECT 1492.310 243.820 1492.630 243.880 ;
        RECT 1496.910 243.820 1497.230 243.880 ;
        RECT 1496.910 183.160 1497.230 183.220 ;
        RECT 1794.070 183.160 1794.390 183.220 ;
        RECT 1496.910 183.020 1794.390 183.160 ;
        RECT 1496.910 182.960 1497.230 183.020 ;
        RECT 1794.070 182.960 1794.390 183.020 ;
        RECT 1794.070 2.960 1794.390 3.020 ;
        RECT 1798.670 2.960 1798.990 3.020 ;
        RECT 1794.070 2.820 1798.990 2.960 ;
        RECT 1794.070 2.760 1794.390 2.820 ;
        RECT 1798.670 2.760 1798.990 2.820 ;
      LAYER via ;
        RECT 1492.340 243.820 1492.600 244.080 ;
        RECT 1496.940 243.820 1497.200 244.080 ;
        RECT 1496.940 182.960 1497.200 183.220 ;
        RECT 1794.100 182.960 1794.360 183.220 ;
        RECT 1794.100 2.760 1794.360 3.020 ;
        RECT 1798.700 2.760 1798.960 3.020 ;
      LAYER met2 ;
        RECT 1492.290 260.000 1492.570 264.000 ;
        RECT 1492.400 244.110 1492.540 260.000 ;
        RECT 1492.340 243.790 1492.600 244.110 ;
        RECT 1496.940 243.790 1497.200 244.110 ;
        RECT 1497.000 183.250 1497.140 243.790 ;
        RECT 1496.940 182.930 1497.200 183.250 ;
        RECT 1794.100 182.930 1794.360 183.250 ;
        RECT 1794.160 3.050 1794.300 182.930 ;
        RECT 1794.100 2.730 1794.360 3.050 ;
        RECT 1798.700 2.730 1798.960 3.050 ;
        RECT 1798.760 2.400 1798.900 2.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1510.250 217.160 1510.570 217.220 ;
        RECT 1814.770 217.160 1815.090 217.220 ;
        RECT 1510.250 217.020 1815.090 217.160 ;
        RECT 1510.250 216.960 1510.570 217.020 ;
        RECT 1814.770 216.960 1815.090 217.020 ;
      LAYER via ;
        RECT 1510.280 216.960 1510.540 217.220 ;
        RECT 1814.800 216.960 1815.060 217.220 ;
      LAYER met2 ;
        RECT 1510.230 260.000 1510.510 264.000 ;
        RECT 1510.340 217.250 1510.480 260.000 ;
        RECT 1510.280 216.930 1510.540 217.250 ;
        RECT 1814.800 216.930 1815.060 217.250 ;
        RECT 1814.860 3.130 1815.000 216.930 ;
        RECT 1814.860 2.990 1816.840 3.130 ;
        RECT 1816.700 2.400 1816.840 2.990 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1531.410 128.080 1531.730 128.140 ;
        RECT 1828.570 128.080 1828.890 128.140 ;
        RECT 1531.410 127.940 1828.890 128.080 ;
        RECT 1531.410 127.880 1531.730 127.940 ;
        RECT 1828.570 127.880 1828.890 127.940 ;
        RECT 1828.570 16.220 1828.890 16.280 ;
        RECT 1834.550 16.220 1834.870 16.280 ;
        RECT 1828.570 16.080 1834.870 16.220 ;
        RECT 1828.570 16.020 1828.890 16.080 ;
        RECT 1834.550 16.020 1834.870 16.080 ;
      LAYER via ;
        RECT 1531.440 127.880 1531.700 128.140 ;
        RECT 1828.600 127.880 1828.860 128.140 ;
        RECT 1828.600 16.020 1828.860 16.280 ;
        RECT 1834.580 16.020 1834.840 16.280 ;
      LAYER met2 ;
        RECT 1528.170 260.170 1528.450 264.000 ;
        RECT 1528.170 260.030 1531.640 260.170 ;
        RECT 1528.170 260.000 1528.450 260.030 ;
        RECT 1531.500 128.170 1531.640 260.030 ;
        RECT 1531.440 127.850 1531.700 128.170 ;
        RECT 1828.600 127.850 1828.860 128.170 ;
        RECT 1828.660 16.310 1828.800 127.850 ;
        RECT 1828.600 15.990 1828.860 16.310 ;
        RECT 1834.580 15.990 1834.840 16.310 ;
        RECT 1834.640 2.400 1834.780 15.990 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1546.130 246.060 1546.450 246.120 ;
        RECT 1597.190 246.060 1597.510 246.120 ;
        RECT 1546.130 245.920 1597.510 246.060 ;
        RECT 1546.130 245.860 1546.450 245.920 ;
        RECT 1597.190 245.860 1597.510 245.920 ;
        RECT 1597.190 134.880 1597.510 134.940 ;
        RECT 1849.270 134.880 1849.590 134.940 ;
        RECT 1597.190 134.740 1849.590 134.880 ;
        RECT 1597.190 134.680 1597.510 134.740 ;
        RECT 1849.270 134.680 1849.590 134.740 ;
      LAYER via ;
        RECT 1546.160 245.860 1546.420 246.120 ;
        RECT 1597.220 245.860 1597.480 246.120 ;
        RECT 1597.220 134.680 1597.480 134.940 ;
        RECT 1849.300 134.680 1849.560 134.940 ;
      LAYER met2 ;
        RECT 1546.110 260.000 1546.390 264.000 ;
        RECT 1546.220 246.150 1546.360 260.000 ;
        RECT 1546.160 245.830 1546.420 246.150 ;
        RECT 1597.220 245.830 1597.480 246.150 ;
        RECT 1597.280 134.970 1597.420 245.830 ;
        RECT 1597.220 134.650 1597.480 134.970 ;
        RECT 1849.300 134.650 1849.560 134.970 ;
        RECT 1849.360 11.290 1849.500 134.650 ;
        RECT 1849.360 11.150 1852.260 11.290 ;
        RECT 1852.120 2.400 1852.260 11.150 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1565.910 189.620 1566.230 189.680 ;
        RECT 1870.430 189.620 1870.750 189.680 ;
        RECT 1565.910 189.480 1870.750 189.620 ;
        RECT 1565.910 189.420 1566.230 189.480 ;
        RECT 1870.430 189.420 1870.750 189.480 ;
      LAYER via ;
        RECT 1565.940 189.420 1566.200 189.680 ;
        RECT 1870.460 189.420 1870.720 189.680 ;
      LAYER met2 ;
        RECT 1564.050 260.170 1564.330 264.000 ;
        RECT 1564.050 260.030 1566.140 260.170 ;
        RECT 1564.050 260.000 1564.330 260.030 ;
        RECT 1566.000 189.710 1566.140 260.030 ;
        RECT 1565.940 189.390 1566.200 189.710 ;
        RECT 1870.460 189.390 1870.720 189.710 ;
        RECT 1870.520 7.210 1870.660 189.390 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 441.210 203.560 441.530 203.620 ;
        RECT 745.270 203.560 745.590 203.620 ;
        RECT 441.210 203.420 745.590 203.560 ;
        RECT 441.210 203.360 441.530 203.420 ;
        RECT 745.270 203.360 745.590 203.420 ;
      LAYER via ;
        RECT 441.240 203.360 441.500 203.620 ;
        RECT 745.300 203.360 745.560 203.620 ;
      LAYER met2 ;
        RECT 437.970 260.170 438.250 264.000 ;
        RECT 437.970 260.030 441.440 260.170 ;
        RECT 437.970 260.000 438.250 260.030 ;
        RECT 441.300 203.650 441.440 260.030 ;
        RECT 441.240 203.330 441.500 203.650 ;
        RECT 745.300 203.330 745.560 203.650 ;
        RECT 745.360 17.240 745.500 203.330 ;
        RECT 745.360 17.100 746.420 17.240 ;
        RECT 746.280 2.400 746.420 17.100 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1582.010 244.020 1582.330 244.080 ;
        RECT 1586.610 244.020 1586.930 244.080 ;
        RECT 1582.010 243.880 1586.930 244.020 ;
        RECT 1582.010 243.820 1582.330 243.880 ;
        RECT 1586.610 243.820 1586.930 243.880 ;
        RECT 1586.610 148.140 1586.930 148.200 ;
        RECT 1883.770 148.140 1884.090 148.200 ;
        RECT 1586.610 148.000 1884.090 148.140 ;
        RECT 1586.610 147.940 1586.930 148.000 ;
        RECT 1883.770 147.940 1884.090 148.000 ;
      LAYER via ;
        RECT 1582.040 243.820 1582.300 244.080 ;
        RECT 1586.640 243.820 1586.900 244.080 ;
        RECT 1586.640 147.940 1586.900 148.200 ;
        RECT 1883.800 147.940 1884.060 148.200 ;
      LAYER met2 ;
        RECT 1581.990 260.000 1582.270 264.000 ;
        RECT 1582.100 244.110 1582.240 260.000 ;
        RECT 1582.040 243.790 1582.300 244.110 ;
        RECT 1586.640 243.790 1586.900 244.110 ;
        RECT 1586.700 148.230 1586.840 243.790 ;
        RECT 1586.640 147.910 1586.900 148.230 ;
        RECT 1883.800 147.910 1884.060 148.230 ;
        RECT 1883.860 16.730 1884.000 147.910 ;
        RECT 1883.860 16.590 1888.140 16.730 ;
        RECT 1888.000 2.400 1888.140 16.590 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1600.410 210.360 1600.730 210.420 ;
        RECT 1904.470 210.360 1904.790 210.420 ;
        RECT 1600.410 210.220 1904.790 210.360 ;
        RECT 1600.410 210.160 1600.730 210.220 ;
        RECT 1904.470 210.160 1904.790 210.220 ;
      LAYER via ;
        RECT 1600.440 210.160 1600.700 210.420 ;
        RECT 1904.500 210.160 1904.760 210.420 ;
      LAYER met2 ;
        RECT 1599.470 260.170 1599.750 264.000 ;
        RECT 1599.470 260.030 1600.640 260.170 ;
        RECT 1599.470 260.000 1599.750 260.030 ;
        RECT 1600.500 210.450 1600.640 260.030 ;
        RECT 1600.440 210.130 1600.700 210.450 ;
        RECT 1904.500 210.130 1904.760 210.450 ;
        RECT 1904.560 16.730 1904.700 210.130 ;
        RECT 1904.560 16.590 1906.080 16.730 ;
        RECT 1905.940 2.400 1906.080 16.590 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1617.430 244.020 1617.750 244.080 ;
        RECT 1621.110 244.020 1621.430 244.080 ;
        RECT 1617.430 243.880 1621.430 244.020 ;
        RECT 1617.430 243.820 1617.750 243.880 ;
        RECT 1621.110 243.820 1621.430 243.880 ;
        RECT 1621.110 155.280 1621.430 155.340 ;
        RECT 1918.270 155.280 1918.590 155.340 ;
        RECT 1621.110 155.140 1918.590 155.280 ;
        RECT 1621.110 155.080 1621.430 155.140 ;
        RECT 1918.270 155.080 1918.590 155.140 ;
      LAYER via ;
        RECT 1617.460 243.820 1617.720 244.080 ;
        RECT 1621.140 243.820 1621.400 244.080 ;
        RECT 1621.140 155.080 1621.400 155.340 ;
        RECT 1918.300 155.080 1918.560 155.340 ;
      LAYER met2 ;
        RECT 1617.410 260.000 1617.690 264.000 ;
        RECT 1617.520 244.110 1617.660 260.000 ;
        RECT 1617.460 243.790 1617.720 244.110 ;
        RECT 1621.140 243.790 1621.400 244.110 ;
        RECT 1621.200 155.370 1621.340 243.790 ;
        RECT 1621.140 155.050 1621.400 155.370 ;
        RECT 1918.300 155.050 1918.560 155.370 ;
        RECT 1918.360 16.730 1918.500 155.050 ;
        RECT 1918.360 16.590 1923.560 16.730 ;
        RECT 1923.420 2.400 1923.560 16.590 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1635.370 244.020 1635.690 244.080 ;
        RECT 1641.350 244.020 1641.670 244.080 ;
        RECT 1635.370 243.880 1641.670 244.020 ;
        RECT 1635.370 243.820 1635.690 243.880 ;
        RECT 1641.350 243.820 1641.670 243.880 ;
        RECT 1641.350 196.760 1641.670 196.820 ;
        RECT 1938.970 196.760 1939.290 196.820 ;
        RECT 1641.350 196.620 1939.290 196.760 ;
        RECT 1641.350 196.560 1641.670 196.620 ;
        RECT 1938.970 196.560 1939.290 196.620 ;
      LAYER via ;
        RECT 1635.400 243.820 1635.660 244.080 ;
        RECT 1641.380 243.820 1641.640 244.080 ;
        RECT 1641.380 196.560 1641.640 196.820 ;
        RECT 1939.000 196.560 1939.260 196.820 ;
      LAYER met2 ;
        RECT 1635.350 260.000 1635.630 264.000 ;
        RECT 1635.460 244.110 1635.600 260.000 ;
        RECT 1635.400 243.790 1635.660 244.110 ;
        RECT 1641.380 243.790 1641.640 244.110 ;
        RECT 1641.440 196.850 1641.580 243.790 ;
        RECT 1641.380 196.530 1641.640 196.850 ;
        RECT 1939.000 196.530 1939.260 196.850 ;
        RECT 1939.060 16.730 1939.200 196.530 ;
        RECT 1939.060 16.590 1941.500 16.730 ;
        RECT 1941.360 2.400 1941.500 16.590 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.610 203.900 1655.930 203.960 ;
        RECT 1952.770 203.900 1953.090 203.960 ;
        RECT 1655.610 203.760 1953.090 203.900 ;
        RECT 1655.610 203.700 1655.930 203.760 ;
        RECT 1952.770 203.700 1953.090 203.760 ;
        RECT 1952.770 18.260 1953.090 18.320 ;
        RECT 1959.210 18.260 1959.530 18.320 ;
        RECT 1952.770 18.120 1959.530 18.260 ;
        RECT 1952.770 18.060 1953.090 18.120 ;
        RECT 1959.210 18.060 1959.530 18.120 ;
      LAYER via ;
        RECT 1655.640 203.700 1655.900 203.960 ;
        RECT 1952.800 203.700 1953.060 203.960 ;
        RECT 1952.800 18.060 1953.060 18.320 ;
        RECT 1959.240 18.060 1959.500 18.320 ;
      LAYER met2 ;
        RECT 1653.290 260.170 1653.570 264.000 ;
        RECT 1653.290 260.030 1655.840 260.170 ;
        RECT 1653.290 260.000 1653.570 260.030 ;
        RECT 1655.700 203.990 1655.840 260.030 ;
        RECT 1655.640 203.670 1655.900 203.990 ;
        RECT 1952.800 203.670 1953.060 203.990 ;
        RECT 1952.860 18.350 1953.000 203.670 ;
        RECT 1952.800 18.030 1953.060 18.350 ;
        RECT 1959.240 18.030 1959.500 18.350 ;
        RECT 1959.300 2.400 1959.440 18.030 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1671.250 243.680 1671.570 243.740 ;
        RECT 1676.310 243.680 1676.630 243.740 ;
        RECT 1671.250 243.540 1676.630 243.680 ;
        RECT 1671.250 243.480 1671.570 243.540 ;
        RECT 1676.310 243.480 1676.630 243.540 ;
        RECT 1676.310 162.080 1676.630 162.140 ;
        RECT 1973.470 162.080 1973.790 162.140 ;
        RECT 1676.310 161.940 1973.790 162.080 ;
        RECT 1676.310 161.880 1676.630 161.940 ;
        RECT 1973.470 161.880 1973.790 161.940 ;
      LAYER via ;
        RECT 1671.280 243.480 1671.540 243.740 ;
        RECT 1676.340 243.480 1676.600 243.740 ;
        RECT 1676.340 161.880 1676.600 162.140 ;
        RECT 1973.500 161.880 1973.760 162.140 ;
      LAYER met2 ;
        RECT 1671.230 260.000 1671.510 264.000 ;
        RECT 1671.340 243.770 1671.480 260.000 ;
        RECT 1671.280 243.450 1671.540 243.770 ;
        RECT 1676.340 243.450 1676.600 243.770 ;
        RECT 1676.400 162.170 1676.540 243.450 ;
        RECT 1676.340 161.850 1676.600 162.170 ;
        RECT 1973.500 161.850 1973.760 162.170 ;
        RECT 1973.560 16.730 1973.700 161.850 ;
        RECT 1973.560 16.590 1977.380 16.730 ;
        RECT 1977.240 2.400 1977.380 16.590 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1690.110 169.220 1690.430 169.280 ;
        RECT 1994.170 169.220 1994.490 169.280 ;
        RECT 1690.110 169.080 1994.490 169.220 ;
        RECT 1690.110 169.020 1690.430 169.080 ;
        RECT 1994.170 169.020 1994.490 169.080 ;
      LAYER via ;
        RECT 1690.140 169.020 1690.400 169.280 ;
        RECT 1994.200 169.020 1994.460 169.280 ;
      LAYER met2 ;
        RECT 1689.170 260.170 1689.450 264.000 ;
        RECT 1689.170 260.030 1690.340 260.170 ;
        RECT 1689.170 260.000 1689.450 260.030 ;
        RECT 1690.200 169.310 1690.340 260.030 ;
        RECT 1690.140 168.990 1690.400 169.310 ;
        RECT 1994.200 168.990 1994.460 169.310 ;
        RECT 1994.260 16.730 1994.400 168.990 ;
        RECT 1994.260 16.590 1995.320 16.730 ;
        RECT 1995.180 2.400 1995.320 16.590 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1710.810 176.020 1711.130 176.080 ;
        RECT 2007.970 176.020 2008.290 176.080 ;
        RECT 1710.810 175.880 2008.290 176.020 ;
        RECT 1710.810 175.820 1711.130 175.880 ;
        RECT 2007.970 175.820 2008.290 175.880 ;
      LAYER via ;
        RECT 1710.840 175.820 1711.100 176.080 ;
        RECT 2008.000 175.820 2008.260 176.080 ;
      LAYER met2 ;
        RECT 1707.110 260.170 1707.390 264.000 ;
        RECT 1707.110 260.030 1711.040 260.170 ;
        RECT 1707.110 260.000 1707.390 260.030 ;
        RECT 1710.900 176.110 1711.040 260.030 ;
        RECT 1710.840 175.790 1711.100 176.110 ;
        RECT 2008.000 175.790 2008.260 176.110 ;
        RECT 2008.060 16.730 2008.200 175.790 ;
        RECT 2008.060 16.590 2012.800 16.730 ;
        RECT 2012.660 2.400 2012.800 16.590 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.150 231.100 1724.470 231.160 ;
        RECT 2028.670 231.100 2028.990 231.160 ;
        RECT 1724.150 230.960 2028.990 231.100 ;
        RECT 1724.150 230.900 1724.470 230.960 ;
        RECT 2028.670 230.900 2028.990 230.960 ;
      LAYER via ;
        RECT 1724.180 230.900 1724.440 231.160 ;
        RECT 2028.700 230.900 2028.960 231.160 ;
      LAYER met2 ;
        RECT 1724.590 260.170 1724.870 264.000 ;
        RECT 1724.240 260.030 1724.870 260.170 ;
        RECT 1724.240 231.190 1724.380 260.030 ;
        RECT 1724.590 260.000 1724.870 260.030 ;
        RECT 1724.180 230.870 1724.440 231.190 ;
        RECT 2028.700 230.870 2028.960 231.190 ;
        RECT 2028.760 16.730 2028.900 230.870 ;
        RECT 2028.760 16.590 2030.740 16.730 ;
        RECT 2030.600 2.400 2030.740 16.590 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1745.310 224.640 1745.630 224.700 ;
        RECT 2042.470 224.640 2042.790 224.700 ;
        RECT 1745.310 224.500 2042.790 224.640 ;
        RECT 1745.310 224.440 1745.630 224.500 ;
        RECT 2042.470 224.440 2042.790 224.500 ;
        RECT 2042.470 18.260 2042.790 18.320 ;
        RECT 2048.450 18.260 2048.770 18.320 ;
        RECT 2042.470 18.120 2048.770 18.260 ;
        RECT 2042.470 18.060 2042.790 18.120 ;
        RECT 2048.450 18.060 2048.770 18.120 ;
      LAYER via ;
        RECT 1745.340 224.440 1745.600 224.700 ;
        RECT 2042.500 224.440 2042.760 224.700 ;
        RECT 2042.500 18.060 2042.760 18.320 ;
        RECT 2048.480 18.060 2048.740 18.320 ;
      LAYER met2 ;
        RECT 1742.530 260.170 1742.810 264.000 ;
        RECT 1742.530 260.030 1745.540 260.170 ;
        RECT 1742.530 260.000 1742.810 260.030 ;
        RECT 1745.400 224.730 1745.540 260.030 ;
        RECT 1745.340 224.410 1745.600 224.730 ;
        RECT 2042.500 224.410 2042.760 224.730 ;
        RECT 2042.560 18.350 2042.700 224.410 ;
        RECT 2042.500 18.030 2042.760 18.350 ;
        RECT 2048.480 18.030 2048.740 18.350 ;
        RECT 2048.540 2.400 2048.680 18.030 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 455.470 244.020 455.790 244.080 ;
        RECT 461.450 244.020 461.770 244.080 ;
        RECT 455.470 243.880 461.770 244.020 ;
        RECT 455.470 243.820 455.790 243.880 ;
        RECT 461.450 243.820 461.770 243.880 ;
        RECT 461.450 65.860 461.770 65.920 ;
        RECT 759.070 65.860 759.390 65.920 ;
        RECT 461.450 65.720 759.390 65.860 ;
        RECT 461.450 65.660 461.770 65.720 ;
        RECT 759.070 65.660 759.390 65.720 ;
      LAYER via ;
        RECT 455.500 243.820 455.760 244.080 ;
        RECT 461.480 243.820 461.740 244.080 ;
        RECT 461.480 65.660 461.740 65.920 ;
        RECT 759.100 65.660 759.360 65.920 ;
      LAYER met2 ;
        RECT 455.450 260.000 455.730 264.000 ;
        RECT 455.560 244.110 455.700 260.000 ;
        RECT 455.500 243.790 455.760 244.110 ;
        RECT 461.480 243.790 461.740 244.110 ;
        RECT 461.540 65.950 461.680 243.790 ;
        RECT 461.480 65.630 461.740 65.950 ;
        RECT 759.100 65.630 759.360 65.950 ;
        RECT 759.160 16.730 759.300 65.630 ;
        RECT 759.160 16.590 763.900 16.730 ;
        RECT 763.760 2.400 763.900 16.590 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1760.490 242.320 1760.810 242.380 ;
        RECT 1766.010 242.320 1766.330 242.380 ;
        RECT 1760.490 242.180 1766.330 242.320 ;
        RECT 1760.490 242.120 1760.810 242.180 ;
        RECT 1766.010 242.120 1766.330 242.180 ;
        RECT 1766.010 183.500 1766.330 183.560 ;
        RECT 2063.170 183.500 2063.490 183.560 ;
        RECT 1766.010 183.360 2063.490 183.500 ;
        RECT 1766.010 183.300 1766.330 183.360 ;
        RECT 2063.170 183.300 2063.490 183.360 ;
      LAYER via ;
        RECT 1760.520 242.120 1760.780 242.380 ;
        RECT 1766.040 242.120 1766.300 242.380 ;
        RECT 1766.040 183.300 1766.300 183.560 ;
        RECT 2063.200 183.300 2063.460 183.560 ;
      LAYER met2 ;
        RECT 1760.470 260.000 1760.750 264.000 ;
        RECT 1760.580 242.410 1760.720 260.000 ;
        RECT 1760.520 242.090 1760.780 242.410 ;
        RECT 1766.040 242.090 1766.300 242.410 ;
        RECT 1766.100 183.590 1766.240 242.090 ;
        RECT 1766.040 183.270 1766.300 183.590 ;
        RECT 2063.200 183.270 2063.460 183.590 ;
        RECT 2063.260 16.730 2063.400 183.270 ;
        RECT 2063.260 16.590 2066.620 16.730 ;
        RECT 2066.480 2.400 2066.620 16.590 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.810 217.500 1780.130 217.560 ;
        RECT 2084.330 217.500 2084.650 217.560 ;
        RECT 1779.810 217.360 2084.650 217.500 ;
        RECT 1779.810 217.300 1780.130 217.360 ;
        RECT 2084.330 217.300 2084.650 217.360 ;
      LAYER via ;
        RECT 1779.840 217.300 1780.100 217.560 ;
        RECT 2084.360 217.300 2084.620 217.560 ;
      LAYER met2 ;
        RECT 1778.410 260.170 1778.690 264.000 ;
        RECT 1778.410 260.030 1780.040 260.170 ;
        RECT 1778.410 260.000 1778.690 260.030 ;
        RECT 1779.900 217.590 1780.040 260.030 ;
        RECT 1779.840 217.270 1780.100 217.590 ;
        RECT 2084.360 217.270 2084.620 217.590 ;
        RECT 2084.420 2.400 2084.560 217.270 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1796.370 244.020 1796.690 244.080 ;
        RECT 1800.510 244.020 1800.830 244.080 ;
        RECT 1796.370 243.880 1800.830 244.020 ;
        RECT 1796.370 243.820 1796.690 243.880 ;
        RECT 1800.510 243.820 1800.830 243.880 ;
        RECT 1800.510 127.740 1800.830 127.800 ;
        RECT 2097.670 127.740 2097.990 127.800 ;
        RECT 1800.510 127.600 2097.990 127.740 ;
        RECT 1800.510 127.540 1800.830 127.600 ;
        RECT 2097.670 127.540 2097.990 127.600 ;
      LAYER via ;
        RECT 1796.400 243.820 1796.660 244.080 ;
        RECT 1800.540 243.820 1800.800 244.080 ;
        RECT 1800.540 127.540 1800.800 127.800 ;
        RECT 2097.700 127.540 2097.960 127.800 ;
      LAYER met2 ;
        RECT 1796.350 260.000 1796.630 264.000 ;
        RECT 1796.460 244.110 1796.600 260.000 ;
        RECT 1796.400 243.790 1796.660 244.110 ;
        RECT 1800.540 243.790 1800.800 244.110 ;
        RECT 1800.600 127.830 1800.740 243.790 ;
        RECT 1800.540 127.510 1800.800 127.830 ;
        RECT 2097.700 127.510 2097.960 127.830 ;
        RECT 2097.760 16.730 2097.900 127.510 ;
        RECT 2097.760 16.590 2102.040 16.730 ;
        RECT 2101.900 2.400 2102.040 16.590 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1813.850 120.600 1814.170 120.660 ;
        RECT 2118.370 120.600 2118.690 120.660 ;
        RECT 1813.850 120.460 2118.690 120.600 ;
        RECT 1813.850 120.400 1814.170 120.460 ;
        RECT 2118.370 120.400 2118.690 120.460 ;
      LAYER via ;
        RECT 1813.880 120.400 1814.140 120.660 ;
        RECT 2118.400 120.400 2118.660 120.660 ;
      LAYER met2 ;
        RECT 1814.290 260.170 1814.570 264.000 ;
        RECT 1813.940 260.030 1814.570 260.170 ;
        RECT 1813.940 120.690 1814.080 260.030 ;
        RECT 1814.290 260.000 1814.570 260.030 ;
        RECT 1813.880 120.370 1814.140 120.690 ;
        RECT 2118.400 120.370 2118.660 120.690 ;
        RECT 2118.460 16.730 2118.600 120.370 ;
        RECT 2118.460 16.590 2119.980 16.730 ;
        RECT 2119.840 2.400 2119.980 16.590 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.010 134.540 1835.330 134.600 ;
        RECT 2132.170 134.540 2132.490 134.600 ;
        RECT 1835.010 134.400 2132.490 134.540 ;
        RECT 1835.010 134.340 1835.330 134.400 ;
        RECT 2132.170 134.340 2132.490 134.400 ;
      LAYER via ;
        RECT 1835.040 134.340 1835.300 134.600 ;
        RECT 2132.200 134.340 2132.460 134.600 ;
      LAYER met2 ;
        RECT 1832.230 260.170 1832.510 264.000 ;
        RECT 1832.230 260.030 1835.240 260.170 ;
        RECT 1832.230 260.000 1832.510 260.030 ;
        RECT 1835.100 134.630 1835.240 260.030 ;
        RECT 1835.040 134.310 1835.300 134.630 ;
        RECT 2132.200 134.310 2132.460 134.630 ;
        RECT 2132.260 16.730 2132.400 134.310 ;
        RECT 2132.260 16.590 2137.920 16.730 ;
        RECT 2137.780 2.400 2137.920 16.590 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2155.705 2.805 2155.875 48.195 ;
      LAYER mcon ;
        RECT 2155.705 48.025 2155.875 48.195 ;
      LAYER met1 ;
        RECT 1849.730 244.020 1850.050 244.080 ;
        RECT 1855.250 244.020 1855.570 244.080 ;
        RECT 1849.730 243.880 1855.570 244.020 ;
        RECT 1849.730 243.820 1850.050 243.880 ;
        RECT 1855.250 243.820 1855.570 243.880 ;
        RECT 1855.250 141.680 1855.570 141.740 ;
        RECT 2152.870 141.680 2153.190 141.740 ;
        RECT 1855.250 141.540 2153.190 141.680 ;
        RECT 1855.250 141.480 1855.570 141.540 ;
        RECT 2152.870 141.480 2153.190 141.540 ;
        RECT 2152.870 48.180 2153.190 48.240 ;
        RECT 2155.645 48.180 2155.935 48.225 ;
        RECT 2152.870 48.040 2155.935 48.180 ;
        RECT 2152.870 47.980 2153.190 48.040 ;
        RECT 2155.645 47.995 2155.935 48.040 ;
        RECT 2155.630 2.960 2155.950 3.020 ;
        RECT 2155.435 2.820 2155.950 2.960 ;
        RECT 2155.630 2.760 2155.950 2.820 ;
      LAYER via ;
        RECT 1849.760 243.820 1850.020 244.080 ;
        RECT 1855.280 243.820 1855.540 244.080 ;
        RECT 1855.280 141.480 1855.540 141.740 ;
        RECT 2152.900 141.480 2153.160 141.740 ;
        RECT 2152.900 47.980 2153.160 48.240 ;
        RECT 2155.660 2.760 2155.920 3.020 ;
      LAYER met2 ;
        RECT 1849.710 260.000 1849.990 264.000 ;
        RECT 1849.820 244.110 1849.960 260.000 ;
        RECT 1849.760 243.790 1850.020 244.110 ;
        RECT 1855.280 243.790 1855.540 244.110 ;
        RECT 1855.340 141.770 1855.480 243.790 ;
        RECT 1855.280 141.450 1855.540 141.770 ;
        RECT 2152.900 141.450 2153.160 141.770 ;
        RECT 2152.960 48.270 2153.100 141.450 ;
        RECT 2152.900 47.950 2153.160 48.270 ;
        RECT 2155.660 2.730 2155.920 3.050 ;
        RECT 2155.720 2.400 2155.860 2.730 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1869.510 148.480 1869.830 148.540 ;
        RECT 2166.670 148.480 2166.990 148.540 ;
        RECT 1869.510 148.340 2166.990 148.480 ;
        RECT 1869.510 148.280 1869.830 148.340 ;
        RECT 2166.670 148.280 2166.990 148.340 ;
        RECT 2166.670 37.980 2166.990 38.040 ;
        RECT 2173.110 37.980 2173.430 38.040 ;
        RECT 2166.670 37.840 2173.430 37.980 ;
        RECT 2166.670 37.780 2166.990 37.840 ;
        RECT 2173.110 37.780 2173.430 37.840 ;
      LAYER via ;
        RECT 1869.540 148.280 1869.800 148.540 ;
        RECT 2166.700 148.280 2166.960 148.540 ;
        RECT 2166.700 37.780 2166.960 38.040 ;
        RECT 2173.140 37.780 2173.400 38.040 ;
      LAYER met2 ;
        RECT 1867.650 260.170 1867.930 264.000 ;
        RECT 1867.650 260.030 1869.740 260.170 ;
        RECT 1867.650 260.000 1867.930 260.030 ;
        RECT 1869.600 148.570 1869.740 260.030 ;
        RECT 1869.540 148.250 1869.800 148.570 ;
        RECT 2166.700 148.250 2166.960 148.570 ;
        RECT 2166.760 38.070 2166.900 148.250 ;
        RECT 2166.700 37.750 2166.960 38.070 ;
        RECT 2173.140 37.750 2173.400 38.070 ;
        RECT 2173.200 2.400 2173.340 37.750 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1885.610 241.640 1885.930 241.700 ;
        RECT 1890.210 241.640 1890.530 241.700 ;
        RECT 1885.610 241.500 1890.530 241.640 ;
        RECT 1885.610 241.440 1885.930 241.500 ;
        RECT 1890.210 241.440 1890.530 241.500 ;
        RECT 1890.210 155.620 1890.530 155.680 ;
        RECT 2187.370 155.620 2187.690 155.680 ;
        RECT 1890.210 155.480 2187.690 155.620 ;
        RECT 1890.210 155.420 1890.530 155.480 ;
        RECT 2187.370 155.420 2187.690 155.480 ;
      LAYER via ;
        RECT 1885.640 241.440 1885.900 241.700 ;
        RECT 1890.240 241.440 1890.500 241.700 ;
        RECT 1890.240 155.420 1890.500 155.680 ;
        RECT 2187.400 155.420 2187.660 155.680 ;
      LAYER met2 ;
        RECT 1885.590 260.000 1885.870 264.000 ;
        RECT 1885.700 241.730 1885.840 260.000 ;
        RECT 1885.640 241.410 1885.900 241.730 ;
        RECT 1890.240 241.410 1890.500 241.730 ;
        RECT 1890.300 155.710 1890.440 241.410 ;
        RECT 1890.240 155.390 1890.500 155.710 ;
        RECT 2187.400 155.390 2187.660 155.710 ;
        RECT 2187.460 16.730 2187.600 155.390 ;
        RECT 2187.460 16.590 2191.280 16.730 ;
        RECT 2191.140 2.400 2191.280 16.590 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1903.550 189.620 1903.870 189.680 ;
        RECT 2208.070 189.620 2208.390 189.680 ;
        RECT 1903.550 189.480 2208.390 189.620 ;
        RECT 1903.550 189.420 1903.870 189.480 ;
        RECT 2208.070 189.420 2208.390 189.480 ;
      LAYER via ;
        RECT 1903.580 189.420 1903.840 189.680 ;
        RECT 2208.100 189.420 2208.360 189.680 ;
      LAYER met2 ;
        RECT 1903.530 260.000 1903.810 264.000 ;
        RECT 1903.640 189.710 1903.780 260.000 ;
        RECT 1903.580 189.390 1903.840 189.710 ;
        RECT 2208.100 189.390 2208.360 189.710 ;
        RECT 2208.160 16.730 2208.300 189.390 ;
        RECT 2208.160 16.590 2209.220 16.730 ;
        RECT 2209.080 2.400 2209.220 16.590 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 197.100 1925.030 197.160 ;
        RECT 2221.870 197.100 2222.190 197.160 ;
        RECT 1924.710 196.960 2222.190 197.100 ;
        RECT 1924.710 196.900 1925.030 196.960 ;
        RECT 2221.870 196.900 2222.190 196.960 ;
      LAYER via ;
        RECT 1924.740 196.900 1925.000 197.160 ;
        RECT 2221.900 196.900 2222.160 197.160 ;
      LAYER met2 ;
        RECT 1921.470 260.170 1921.750 264.000 ;
        RECT 1921.470 260.030 1924.940 260.170 ;
        RECT 1921.470 260.000 1921.750 260.030 ;
        RECT 1924.800 197.190 1924.940 260.030 ;
        RECT 1924.740 196.870 1925.000 197.190 ;
        RECT 2221.900 196.870 2222.160 197.190 ;
        RECT 2221.960 16.730 2222.100 196.870 ;
        RECT 2221.960 16.590 2227.160 16.730 ;
        RECT 2227.020 2.400 2227.160 16.590 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 473.410 237.900 473.730 237.960 ;
        RECT 779.770 237.900 780.090 237.960 ;
        RECT 473.410 237.760 780.090 237.900 ;
        RECT 473.410 237.700 473.730 237.760 ;
        RECT 779.770 237.700 780.090 237.760 ;
      LAYER via ;
        RECT 473.440 237.700 473.700 237.960 ;
        RECT 779.800 237.700 780.060 237.960 ;
      LAYER met2 ;
        RECT 473.390 260.000 473.670 264.000 ;
        RECT 473.500 237.990 473.640 260.000 ;
        RECT 473.440 237.670 473.700 237.990 ;
        RECT 779.800 237.670 780.060 237.990 ;
        RECT 779.860 16.730 780.000 237.670 ;
        RECT 779.860 16.590 781.840 16.730 ;
        RECT 781.700 2.400 781.840 16.590 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1939.430 244.020 1939.750 244.080 ;
        RECT 1945.410 244.020 1945.730 244.080 ;
        RECT 1939.430 243.880 1945.730 244.020 ;
        RECT 1939.430 243.820 1939.750 243.880 ;
        RECT 1945.410 243.820 1945.730 243.880 ;
        RECT 1945.410 162.420 1945.730 162.480 ;
        RECT 2242.570 162.420 2242.890 162.480 ;
        RECT 1945.410 162.280 2242.890 162.420 ;
        RECT 1945.410 162.220 1945.730 162.280 ;
        RECT 2242.570 162.220 2242.890 162.280 ;
      LAYER via ;
        RECT 1939.460 243.820 1939.720 244.080 ;
        RECT 1945.440 243.820 1945.700 244.080 ;
        RECT 1945.440 162.220 1945.700 162.480 ;
        RECT 2242.600 162.220 2242.860 162.480 ;
      LAYER met2 ;
        RECT 1939.410 260.000 1939.690 264.000 ;
        RECT 1939.520 244.110 1939.660 260.000 ;
        RECT 1939.460 243.790 1939.720 244.110 ;
        RECT 1945.440 243.790 1945.700 244.110 ;
        RECT 1945.500 162.510 1945.640 243.790 ;
        RECT 1945.440 162.190 1945.700 162.510 ;
        RECT 2242.600 162.190 2242.860 162.510 ;
        RECT 2242.660 16.730 2242.800 162.190 ;
        RECT 2242.660 16.590 2245.100 16.730 ;
        RECT 2244.960 2.400 2245.100 16.590 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1959.210 203.560 1959.530 203.620 ;
        RECT 2256.370 203.560 2256.690 203.620 ;
        RECT 1959.210 203.420 2256.690 203.560 ;
        RECT 1959.210 203.360 1959.530 203.420 ;
        RECT 2256.370 203.360 2256.690 203.420 ;
        RECT 2256.370 17.920 2256.690 17.980 ;
        RECT 2262.350 17.920 2262.670 17.980 ;
        RECT 2256.370 17.780 2262.670 17.920 ;
        RECT 2256.370 17.720 2256.690 17.780 ;
        RECT 2262.350 17.720 2262.670 17.780 ;
      LAYER via ;
        RECT 1959.240 203.360 1959.500 203.620 ;
        RECT 2256.400 203.360 2256.660 203.620 ;
        RECT 2256.400 17.720 2256.660 17.980 ;
        RECT 2262.380 17.720 2262.640 17.980 ;
      LAYER met2 ;
        RECT 1957.350 260.170 1957.630 264.000 ;
        RECT 1957.350 260.030 1959.440 260.170 ;
        RECT 1957.350 260.000 1957.630 260.030 ;
        RECT 1959.300 203.650 1959.440 260.030 ;
        RECT 1959.240 203.330 1959.500 203.650 ;
        RECT 2256.400 203.330 2256.660 203.650 ;
        RECT 2256.460 18.010 2256.600 203.330 ;
        RECT 2256.400 17.690 2256.660 18.010 ;
        RECT 2262.380 17.690 2262.640 18.010 ;
        RECT 2262.440 2.400 2262.580 17.690 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1974.850 244.020 1975.170 244.080 ;
        RECT 1979.910 244.020 1980.230 244.080 ;
        RECT 1974.850 243.880 1980.230 244.020 ;
        RECT 1974.850 243.820 1975.170 243.880 ;
        RECT 1979.910 243.820 1980.230 243.880 ;
        RECT 1979.910 176.360 1980.230 176.420 ;
        RECT 2277.070 176.360 2277.390 176.420 ;
        RECT 1979.910 176.220 2277.390 176.360 ;
        RECT 1979.910 176.160 1980.230 176.220 ;
        RECT 2277.070 176.160 2277.390 176.220 ;
      LAYER via ;
        RECT 1974.880 243.820 1975.140 244.080 ;
        RECT 1979.940 243.820 1980.200 244.080 ;
        RECT 1979.940 176.160 1980.200 176.420 ;
        RECT 2277.100 176.160 2277.360 176.420 ;
      LAYER met2 ;
        RECT 1974.830 260.000 1975.110 264.000 ;
        RECT 1974.940 244.110 1975.080 260.000 ;
        RECT 1974.880 243.790 1975.140 244.110 ;
        RECT 1979.940 243.790 1980.200 244.110 ;
        RECT 1980.000 176.450 1980.140 243.790 ;
        RECT 1979.940 176.130 1980.200 176.450 ;
        RECT 2277.100 176.130 2277.360 176.450 ;
        RECT 2277.160 3.130 2277.300 176.130 ;
        RECT 2277.160 2.990 2280.060 3.130 ;
        RECT 2279.920 2.960 2280.060 2.990 ;
        RECT 2279.920 2.820 2280.520 2.960 ;
        RECT 2280.380 2.400 2280.520 2.820 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1993.710 182.820 1994.030 182.880 ;
        RECT 2298.230 182.820 2298.550 182.880 ;
        RECT 1993.710 182.680 2298.550 182.820 ;
        RECT 1993.710 182.620 1994.030 182.680 ;
        RECT 2298.230 182.620 2298.550 182.680 ;
      LAYER via ;
        RECT 1993.740 182.620 1994.000 182.880 ;
        RECT 2298.260 182.620 2298.520 182.880 ;
      LAYER met2 ;
        RECT 1992.770 260.170 1993.050 264.000 ;
        RECT 1992.770 260.030 1993.940 260.170 ;
        RECT 1992.770 260.000 1993.050 260.030 ;
        RECT 1993.800 182.910 1993.940 260.030 ;
        RECT 1993.740 182.590 1994.000 182.910 ;
        RECT 2298.260 182.590 2298.520 182.910 ;
        RECT 2298.320 2.400 2298.460 182.590 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2014.410 217.160 2014.730 217.220 ;
        RECT 2311.570 217.160 2311.890 217.220 ;
        RECT 2014.410 217.020 2311.890 217.160 ;
        RECT 2014.410 216.960 2014.730 217.020 ;
        RECT 2311.570 216.960 2311.890 217.020 ;
        RECT 2311.570 2.960 2311.890 3.020 ;
        RECT 2316.170 2.960 2316.490 3.020 ;
        RECT 2311.570 2.820 2316.490 2.960 ;
        RECT 2311.570 2.760 2311.890 2.820 ;
        RECT 2316.170 2.760 2316.490 2.820 ;
      LAYER via ;
        RECT 2014.440 216.960 2014.700 217.220 ;
        RECT 2311.600 216.960 2311.860 217.220 ;
        RECT 2311.600 2.760 2311.860 3.020 ;
        RECT 2316.200 2.760 2316.460 3.020 ;
      LAYER met2 ;
        RECT 2010.710 260.170 2010.990 264.000 ;
        RECT 2010.710 260.030 2014.640 260.170 ;
        RECT 2010.710 260.000 2010.990 260.030 ;
        RECT 2014.500 217.250 2014.640 260.030 ;
        RECT 2014.440 216.930 2014.700 217.250 ;
        RECT 2311.600 216.930 2311.860 217.250 ;
        RECT 2311.660 3.050 2311.800 216.930 ;
        RECT 2311.600 2.730 2311.860 3.050 ;
        RECT 2316.200 2.730 2316.460 3.050 ;
        RECT 2316.260 2.400 2316.400 2.730 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2030.050 231.100 2030.370 231.160 ;
        RECT 2332.270 231.100 2332.590 231.160 ;
        RECT 2030.050 230.960 2332.590 231.100 ;
        RECT 2030.050 230.900 2030.370 230.960 ;
        RECT 2332.270 230.900 2332.590 230.960 ;
        RECT 2332.270 2.960 2332.590 3.020 ;
        RECT 2334.110 2.960 2334.430 3.020 ;
        RECT 2332.270 2.820 2334.430 2.960 ;
        RECT 2332.270 2.760 2332.590 2.820 ;
        RECT 2334.110 2.760 2334.430 2.820 ;
      LAYER via ;
        RECT 2030.080 230.900 2030.340 231.160 ;
        RECT 2332.300 230.900 2332.560 231.160 ;
        RECT 2332.300 2.760 2332.560 3.020 ;
        RECT 2334.140 2.760 2334.400 3.020 ;
      LAYER met2 ;
        RECT 2028.650 260.170 2028.930 264.000 ;
        RECT 2028.650 260.030 2030.280 260.170 ;
        RECT 2028.650 260.000 2028.930 260.030 ;
        RECT 2030.140 231.190 2030.280 260.030 ;
        RECT 2030.080 230.870 2030.340 231.190 ;
        RECT 2332.300 230.870 2332.560 231.190 ;
        RECT 2332.360 3.050 2332.500 230.870 ;
        RECT 2332.300 2.730 2332.560 3.050 ;
        RECT 2334.140 2.730 2334.400 3.050 ;
        RECT 2334.200 2.400 2334.340 2.730 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2048.910 168.880 2049.230 168.940 ;
        RECT 2346.070 168.880 2346.390 168.940 ;
        RECT 2048.910 168.740 2346.390 168.880 ;
        RECT 2048.910 168.680 2049.230 168.740 ;
        RECT 2346.070 168.680 2346.390 168.740 ;
        RECT 2346.070 2.960 2346.390 3.020 ;
        RECT 2351.590 2.960 2351.910 3.020 ;
        RECT 2346.070 2.820 2351.910 2.960 ;
        RECT 2346.070 2.760 2346.390 2.820 ;
        RECT 2351.590 2.760 2351.910 2.820 ;
      LAYER via ;
        RECT 2048.940 168.680 2049.200 168.940 ;
        RECT 2346.100 168.680 2346.360 168.940 ;
        RECT 2346.100 2.760 2346.360 3.020 ;
        RECT 2351.620 2.760 2351.880 3.020 ;
      LAYER met2 ;
        RECT 2046.590 260.170 2046.870 264.000 ;
        RECT 2046.590 260.030 2049.140 260.170 ;
        RECT 2046.590 260.000 2046.870 260.030 ;
        RECT 2049.000 168.970 2049.140 260.030 ;
        RECT 2048.940 168.650 2049.200 168.970 ;
        RECT 2346.100 168.650 2346.360 168.970 ;
        RECT 2346.160 3.050 2346.300 168.650 ;
        RECT 2346.100 2.730 2346.360 3.050 ;
        RECT 2351.620 2.730 2351.880 3.050 ;
        RECT 2351.680 2.400 2351.820 2.730 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2064.550 244.020 2064.870 244.080 ;
        RECT 2069.610 244.020 2069.930 244.080 ;
        RECT 2064.550 243.880 2069.930 244.020 ;
        RECT 2064.550 243.820 2064.870 243.880 ;
        RECT 2069.610 243.820 2069.930 243.880 ;
        RECT 2069.610 189.960 2069.930 190.020 ;
        RECT 2366.770 189.960 2367.090 190.020 ;
        RECT 2069.610 189.820 2367.090 189.960 ;
        RECT 2069.610 189.760 2069.930 189.820 ;
        RECT 2366.770 189.760 2367.090 189.820 ;
      LAYER via ;
        RECT 2064.580 243.820 2064.840 244.080 ;
        RECT 2069.640 243.820 2069.900 244.080 ;
        RECT 2069.640 189.760 2069.900 190.020 ;
        RECT 2366.800 189.760 2367.060 190.020 ;
      LAYER met2 ;
        RECT 2064.530 260.000 2064.810 264.000 ;
        RECT 2064.640 244.110 2064.780 260.000 ;
        RECT 2064.580 243.790 2064.840 244.110 ;
        RECT 2069.640 243.790 2069.900 244.110 ;
        RECT 2069.700 190.050 2069.840 243.790 ;
        RECT 2069.640 189.730 2069.900 190.050 ;
        RECT 2366.800 189.730 2367.060 190.050 ;
        RECT 2366.860 16.730 2367.000 189.730 ;
        RECT 2366.860 16.590 2369.760 16.730 ;
        RECT 2369.620 2.400 2369.760 16.590 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2083.410 51.580 2083.730 51.640 ;
        RECT 2387.930 51.580 2388.250 51.640 ;
        RECT 2083.410 51.440 2388.250 51.580 ;
        RECT 2083.410 51.380 2083.730 51.440 ;
        RECT 2387.930 51.380 2388.250 51.440 ;
      LAYER via ;
        RECT 2083.440 51.380 2083.700 51.640 ;
        RECT 2387.960 51.380 2388.220 51.640 ;
      LAYER met2 ;
        RECT 2082.470 260.170 2082.750 264.000 ;
        RECT 2082.470 260.030 2083.640 260.170 ;
        RECT 2082.470 260.000 2082.750 260.030 ;
        RECT 2083.500 51.670 2083.640 260.030 ;
        RECT 2083.440 51.350 2083.700 51.670 ;
        RECT 2387.960 51.350 2388.220 51.670 ;
        RECT 2388.020 17.410 2388.160 51.350 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2100.430 244.020 2100.750 244.080 ;
        RECT 2104.110 244.020 2104.430 244.080 ;
        RECT 2100.430 243.880 2104.430 244.020 ;
        RECT 2100.430 243.820 2100.750 243.880 ;
        RECT 2104.110 243.820 2104.430 243.880 ;
        RECT 2104.110 196.760 2104.430 196.820 ;
        RECT 2401.270 196.760 2401.590 196.820 ;
        RECT 2104.110 196.620 2401.590 196.760 ;
        RECT 2104.110 196.560 2104.430 196.620 ;
        RECT 2401.270 196.560 2401.590 196.620 ;
      LAYER via ;
        RECT 2100.460 243.820 2100.720 244.080 ;
        RECT 2104.140 243.820 2104.400 244.080 ;
        RECT 2104.140 196.560 2104.400 196.820 ;
        RECT 2401.300 196.560 2401.560 196.820 ;
      LAYER met2 ;
        RECT 2100.410 260.000 2100.690 264.000 ;
        RECT 2100.520 244.110 2100.660 260.000 ;
        RECT 2100.460 243.790 2100.720 244.110 ;
        RECT 2104.140 243.790 2104.400 244.110 ;
        RECT 2104.200 196.850 2104.340 243.790 ;
        RECT 2104.140 196.530 2104.400 196.850 ;
        RECT 2401.300 196.530 2401.560 196.850 ;
        RECT 2401.360 16.730 2401.500 196.530 ;
        RECT 2401.360 16.590 2405.640 16.730 ;
        RECT 2405.500 2.400 2405.640 16.590 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 491.350 244.020 491.670 244.080 ;
        RECT 496.410 244.020 496.730 244.080 ;
        RECT 491.350 243.880 496.730 244.020 ;
        RECT 491.350 243.820 491.670 243.880 ;
        RECT 496.410 243.820 496.730 243.880 ;
        RECT 496.410 15.200 496.730 15.260 ;
        RECT 799.550 15.200 799.870 15.260 ;
        RECT 496.410 15.060 799.870 15.200 ;
        RECT 496.410 15.000 496.730 15.060 ;
        RECT 799.550 15.000 799.870 15.060 ;
      LAYER via ;
        RECT 491.380 243.820 491.640 244.080 ;
        RECT 496.440 243.820 496.700 244.080 ;
        RECT 496.440 15.000 496.700 15.260 ;
        RECT 799.580 15.000 799.840 15.260 ;
      LAYER met2 ;
        RECT 491.330 260.000 491.610 264.000 ;
        RECT 491.440 244.110 491.580 260.000 ;
        RECT 491.380 243.790 491.640 244.110 ;
        RECT 496.440 243.790 496.700 244.110 ;
        RECT 496.500 15.290 496.640 243.790 ;
        RECT 496.440 14.970 496.700 15.290 ;
        RECT 799.580 14.970 799.840 15.290 ;
        RECT 799.640 2.400 799.780 14.970 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 336.330 245.040 336.650 245.100 ;
        RECT 642.230 245.040 642.550 245.100 ;
        RECT 336.330 244.900 642.550 245.040 ;
        RECT 336.330 244.840 336.650 244.900 ;
        RECT 642.230 244.840 642.550 244.900 ;
      LAYER via ;
        RECT 336.360 244.840 336.620 245.100 ;
        RECT 642.260 244.840 642.520 245.100 ;
      LAYER met2 ;
        RECT 336.310 260.000 336.590 264.000 ;
        RECT 336.420 245.130 336.560 260.000 ;
        RECT 336.360 244.810 336.620 245.130 ;
        RECT 642.260 244.810 642.520 245.130 ;
        RECT 642.320 17.410 642.460 244.810 ;
        RECT 642.320 17.270 645.220 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2124.810 58.720 2125.130 58.780 ;
        RECT 2429.330 58.720 2429.650 58.780 ;
        RECT 2124.810 58.580 2429.650 58.720 ;
        RECT 2124.810 58.520 2125.130 58.580 ;
        RECT 2429.330 58.520 2429.650 58.580 ;
      LAYER via ;
        RECT 2124.840 58.520 2125.100 58.780 ;
        RECT 2429.360 58.520 2429.620 58.780 ;
      LAYER met2 ;
        RECT 2123.870 260.170 2124.150 264.000 ;
        RECT 2123.870 260.030 2125.040 260.170 ;
        RECT 2123.870 260.000 2124.150 260.030 ;
        RECT 2124.900 58.810 2125.040 260.030 ;
        RECT 2124.840 58.490 2125.100 58.810 ;
        RECT 2429.360 58.490 2429.620 58.810 ;
        RECT 2429.420 17.410 2429.560 58.490 ;
        RECT 2428.960 17.270 2429.560 17.410 ;
        RECT 2428.960 2.400 2429.100 17.270 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2141.830 244.020 2142.150 244.080 ;
        RECT 2145.510 244.020 2145.830 244.080 ;
        RECT 2141.830 243.880 2145.830 244.020 ;
        RECT 2141.830 243.820 2142.150 243.880 ;
        RECT 2145.510 243.820 2145.830 243.880 ;
        RECT 2145.510 19.620 2145.830 19.680 ;
        RECT 2446.810 19.620 2447.130 19.680 ;
        RECT 2145.510 19.480 2447.130 19.620 ;
        RECT 2145.510 19.420 2145.830 19.480 ;
        RECT 2446.810 19.420 2447.130 19.480 ;
      LAYER via ;
        RECT 2141.860 243.820 2142.120 244.080 ;
        RECT 2145.540 243.820 2145.800 244.080 ;
        RECT 2145.540 19.420 2145.800 19.680 ;
        RECT 2446.840 19.420 2447.100 19.680 ;
      LAYER met2 ;
        RECT 2141.810 260.000 2142.090 264.000 ;
        RECT 2141.920 244.110 2142.060 260.000 ;
        RECT 2141.860 243.790 2142.120 244.110 ;
        RECT 2145.540 243.790 2145.800 244.110 ;
        RECT 2145.600 19.710 2145.740 243.790 ;
        RECT 2145.540 19.390 2145.800 19.710 ;
        RECT 2446.840 19.390 2447.100 19.710 ;
        RECT 2446.900 2.400 2447.040 19.390 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2159.770 243.680 2160.090 243.740 ;
        RECT 2166.210 243.680 2166.530 243.740 ;
        RECT 2159.770 243.540 2166.530 243.680 ;
        RECT 2159.770 243.480 2160.090 243.540 ;
        RECT 2166.210 243.480 2166.530 243.540 ;
        RECT 2166.210 20.640 2166.530 20.700 ;
        RECT 2464.750 20.640 2465.070 20.700 ;
        RECT 2166.210 20.500 2465.070 20.640 ;
        RECT 2166.210 20.440 2166.530 20.500 ;
        RECT 2464.750 20.440 2465.070 20.500 ;
      LAYER via ;
        RECT 2159.800 243.480 2160.060 243.740 ;
        RECT 2166.240 243.480 2166.500 243.740 ;
        RECT 2166.240 20.440 2166.500 20.700 ;
        RECT 2464.780 20.440 2465.040 20.700 ;
      LAYER met2 ;
        RECT 2159.750 260.000 2160.030 264.000 ;
        RECT 2159.860 243.770 2160.000 260.000 ;
        RECT 2159.800 243.450 2160.060 243.770 ;
        RECT 2166.240 243.450 2166.500 243.770 ;
        RECT 2166.300 20.730 2166.440 243.450 ;
        RECT 2166.240 20.410 2166.500 20.730 ;
        RECT 2464.780 20.410 2465.040 20.730 ;
        RECT 2464.840 2.400 2464.980 20.410 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 15.880 2180.330 15.940 ;
        RECT 2482.690 15.880 2483.010 15.940 ;
        RECT 2180.010 15.740 2483.010 15.880 ;
        RECT 2180.010 15.680 2180.330 15.740 ;
        RECT 2482.690 15.680 2483.010 15.740 ;
      LAYER via ;
        RECT 2180.040 15.680 2180.300 15.940 ;
        RECT 2482.720 15.680 2482.980 15.940 ;
      LAYER met2 ;
        RECT 2177.690 260.170 2177.970 264.000 ;
        RECT 2177.690 260.030 2180.240 260.170 ;
        RECT 2177.690 260.000 2177.970 260.030 ;
        RECT 2180.100 15.970 2180.240 260.030 ;
        RECT 2180.040 15.650 2180.300 15.970 ;
        RECT 2482.720 15.650 2482.980 15.970 ;
        RECT 2482.780 2.400 2482.920 15.650 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2195.650 244.020 2195.970 244.080 ;
        RECT 2200.710 244.020 2201.030 244.080 ;
        RECT 2195.650 243.880 2201.030 244.020 ;
        RECT 2195.650 243.820 2195.970 243.880 ;
        RECT 2200.710 243.820 2201.030 243.880 ;
        RECT 2200.710 16.220 2201.030 16.280 ;
        RECT 2500.630 16.220 2500.950 16.280 ;
        RECT 2200.710 16.080 2500.950 16.220 ;
        RECT 2200.710 16.020 2201.030 16.080 ;
        RECT 2500.630 16.020 2500.950 16.080 ;
      LAYER via ;
        RECT 2195.680 243.820 2195.940 244.080 ;
        RECT 2200.740 243.820 2201.000 244.080 ;
        RECT 2200.740 16.020 2201.000 16.280 ;
        RECT 2500.660 16.020 2500.920 16.280 ;
      LAYER met2 ;
        RECT 2195.630 260.000 2195.910 264.000 ;
        RECT 2195.740 244.110 2195.880 260.000 ;
        RECT 2195.680 243.790 2195.940 244.110 ;
        RECT 2200.740 243.790 2201.000 244.110 ;
        RECT 2200.800 16.310 2200.940 243.790 ;
        RECT 2200.740 15.990 2201.000 16.310 ;
        RECT 2500.660 15.990 2500.920 16.310 ;
        RECT 2500.720 2.400 2500.860 15.990 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.510 19.960 2214.830 20.020 ;
        RECT 2518.110 19.960 2518.430 20.020 ;
        RECT 2214.510 19.820 2518.430 19.960 ;
        RECT 2214.510 19.760 2214.830 19.820 ;
        RECT 2518.110 19.760 2518.430 19.820 ;
      LAYER via ;
        RECT 2214.540 19.760 2214.800 20.020 ;
        RECT 2518.140 19.760 2518.400 20.020 ;
      LAYER met2 ;
        RECT 2213.570 260.170 2213.850 264.000 ;
        RECT 2213.570 260.030 2214.740 260.170 ;
        RECT 2213.570 260.000 2213.850 260.030 ;
        RECT 2214.600 20.050 2214.740 260.030 ;
        RECT 2214.540 19.730 2214.800 20.050 ;
        RECT 2518.140 19.730 2518.400 20.050 ;
        RECT 2518.200 2.400 2518.340 19.730 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2231.070 244.020 2231.390 244.080 ;
        RECT 2235.210 244.020 2235.530 244.080 ;
        RECT 2231.070 243.880 2235.530 244.020 ;
        RECT 2231.070 243.820 2231.390 243.880 ;
        RECT 2235.210 243.820 2235.530 243.880 ;
        RECT 2235.210 15.540 2235.530 15.600 ;
        RECT 2536.050 15.540 2536.370 15.600 ;
        RECT 2235.210 15.400 2536.370 15.540 ;
        RECT 2235.210 15.340 2235.530 15.400 ;
        RECT 2536.050 15.340 2536.370 15.400 ;
      LAYER via ;
        RECT 2231.100 243.820 2231.360 244.080 ;
        RECT 2235.240 243.820 2235.500 244.080 ;
        RECT 2235.240 15.340 2235.500 15.600 ;
        RECT 2536.080 15.340 2536.340 15.600 ;
      LAYER met2 ;
        RECT 2231.050 260.000 2231.330 264.000 ;
        RECT 2231.160 244.110 2231.300 260.000 ;
        RECT 2231.100 243.790 2231.360 244.110 ;
        RECT 2235.240 243.790 2235.500 244.110 ;
        RECT 2235.300 15.630 2235.440 243.790 ;
        RECT 2235.240 15.310 2235.500 15.630 ;
        RECT 2536.080 15.310 2536.340 15.630 ;
        RECT 2536.140 2.400 2536.280 15.310 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2248.990 260.000 2249.270 264.000 ;
        RECT 2249.100 16.845 2249.240 260.000 ;
        RECT 2249.030 16.475 2249.310 16.845 ;
        RECT 2554.010 16.475 2554.290 16.845 ;
        RECT 2554.080 2.400 2554.220 16.475 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
      LAYER via2 ;
        RECT 2249.030 16.520 2249.310 16.800 ;
        RECT 2554.010 16.520 2554.290 16.800 ;
      LAYER met3 ;
        RECT 2249.005 16.810 2249.335 16.825 ;
        RECT 2553.985 16.810 2554.315 16.825 ;
        RECT 2249.005 16.510 2554.315 16.810 ;
        RECT 2249.005 16.495 2249.335 16.510 ;
        RECT 2553.985 16.495 2554.315 16.510 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 16.900 2270.030 16.960 ;
        RECT 2571.930 16.900 2572.250 16.960 ;
        RECT 2269.710 16.760 2572.250 16.900 ;
        RECT 2269.710 16.700 2270.030 16.760 ;
        RECT 2571.930 16.700 2572.250 16.760 ;
      LAYER via ;
        RECT 2269.740 16.700 2270.000 16.960 ;
        RECT 2571.960 16.700 2572.220 16.960 ;
      LAYER met2 ;
        RECT 2266.930 260.170 2267.210 264.000 ;
        RECT 2266.930 260.030 2269.940 260.170 ;
        RECT 2266.930 260.000 2267.210 260.030 ;
        RECT 2269.800 16.990 2269.940 260.030 ;
        RECT 2269.740 16.670 2270.000 16.990 ;
        RECT 2571.960 16.670 2572.220 16.990 ;
        RECT 2572.020 2.400 2572.160 16.670 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2284.890 244.020 2285.210 244.080 ;
        RECT 2290.410 244.020 2290.730 244.080 ;
        RECT 2284.890 243.880 2290.730 244.020 ;
        RECT 2284.890 243.820 2285.210 243.880 ;
        RECT 2290.410 243.820 2290.730 243.880 ;
        RECT 2290.410 16.560 2290.730 16.620 ;
        RECT 2589.410 16.560 2589.730 16.620 ;
        RECT 2290.410 16.420 2589.730 16.560 ;
        RECT 2290.410 16.360 2290.730 16.420 ;
        RECT 2589.410 16.360 2589.730 16.420 ;
      LAYER via ;
        RECT 2284.920 243.820 2285.180 244.080 ;
        RECT 2290.440 243.820 2290.700 244.080 ;
        RECT 2290.440 16.360 2290.700 16.620 ;
        RECT 2589.440 16.360 2589.700 16.620 ;
      LAYER met2 ;
        RECT 2284.870 260.000 2285.150 264.000 ;
        RECT 2284.980 244.110 2285.120 260.000 ;
        RECT 2284.920 243.790 2285.180 244.110 ;
        RECT 2290.440 243.790 2290.700 244.110 ;
        RECT 2290.500 16.650 2290.640 243.790 ;
        RECT 2290.440 16.330 2290.700 16.650 ;
        RECT 2589.440 16.330 2589.700 16.650 ;
        RECT 2589.500 2.400 2589.640 16.330 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 515.270 245.380 515.590 245.440 ;
        RECT 821.630 245.380 821.950 245.440 ;
        RECT 515.270 245.240 821.950 245.380 ;
        RECT 515.270 245.180 515.590 245.240 ;
        RECT 821.630 245.180 821.950 245.240 ;
      LAYER via ;
        RECT 515.300 245.180 515.560 245.440 ;
        RECT 821.660 245.180 821.920 245.440 ;
      LAYER met2 ;
        RECT 515.250 260.000 515.530 264.000 ;
        RECT 515.360 245.470 515.500 260.000 ;
        RECT 515.300 245.150 515.560 245.470 ;
        RECT 821.660 245.150 821.920 245.470 ;
        RECT 821.720 17.410 821.860 245.150 ;
        RECT 821.720 17.270 823.700 17.410 ;
        RECT 823.560 2.400 823.700 17.270 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2304.670 18.600 2304.990 18.660 ;
        RECT 2607.350 18.600 2607.670 18.660 ;
        RECT 2304.670 18.460 2607.670 18.600 ;
        RECT 2304.670 18.400 2304.990 18.460 ;
        RECT 2607.350 18.400 2607.670 18.460 ;
      LAYER via ;
        RECT 2304.700 18.400 2304.960 18.660 ;
        RECT 2607.380 18.400 2607.640 18.660 ;
      LAYER met2 ;
        RECT 2302.810 260.170 2303.090 264.000 ;
        RECT 2302.810 260.030 2304.440 260.170 ;
        RECT 2302.810 260.000 2303.090 260.030 ;
        RECT 2304.300 19.280 2304.440 260.030 ;
        RECT 2304.300 19.140 2304.900 19.280 ;
        RECT 2304.760 18.690 2304.900 19.140 ;
        RECT 2304.700 18.370 2304.960 18.690 ;
        RECT 2607.380 18.370 2607.640 18.690 ;
        RECT 2607.440 2.400 2607.580 18.370 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2320.770 244.020 2321.090 244.080 ;
        RECT 2324.910 244.020 2325.230 244.080 ;
        RECT 2320.770 243.880 2325.230 244.020 ;
        RECT 2320.770 243.820 2321.090 243.880 ;
        RECT 2324.910 243.820 2325.230 243.880 ;
        RECT 2324.910 20.300 2325.230 20.360 ;
        RECT 2625.290 20.300 2625.610 20.360 ;
        RECT 2324.910 20.160 2625.610 20.300 ;
        RECT 2324.910 20.100 2325.230 20.160 ;
        RECT 2625.290 20.100 2625.610 20.160 ;
      LAYER via ;
        RECT 2320.800 243.820 2321.060 244.080 ;
        RECT 2324.940 243.820 2325.200 244.080 ;
        RECT 2324.940 20.100 2325.200 20.360 ;
        RECT 2625.320 20.100 2625.580 20.360 ;
      LAYER met2 ;
        RECT 2320.750 260.000 2321.030 264.000 ;
        RECT 2320.860 244.110 2321.000 260.000 ;
        RECT 2320.800 243.790 2321.060 244.110 ;
        RECT 2324.940 243.790 2325.200 244.110 ;
        RECT 2325.000 20.390 2325.140 243.790 ;
        RECT 2324.940 20.070 2325.200 20.390 ;
        RECT 2625.320 20.070 2625.580 20.390 ;
        RECT 2625.380 2.400 2625.520 20.070 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2338.710 245.040 2339.030 245.100 ;
        RECT 2642.770 245.040 2643.090 245.100 ;
        RECT 2338.710 244.900 2643.090 245.040 ;
        RECT 2338.710 244.840 2339.030 244.900 ;
        RECT 2642.770 244.840 2643.090 244.900 ;
      LAYER via ;
        RECT 2338.740 244.840 2339.000 245.100 ;
        RECT 2642.800 244.840 2643.060 245.100 ;
      LAYER met2 ;
        RECT 2338.690 260.000 2338.970 264.000 ;
        RECT 2338.800 245.130 2338.940 260.000 ;
        RECT 2338.740 244.810 2339.000 245.130 ;
        RECT 2642.800 244.810 2643.060 245.130 ;
        RECT 2642.860 17.410 2643.000 244.810 ;
        RECT 2642.860 17.270 2643.460 17.410 ;
        RECT 2643.320 2.400 2643.460 17.270 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2642.845 16.405 2643.015 17.935 ;
      LAYER mcon ;
        RECT 2642.845 17.765 2643.015 17.935 ;
      LAYER met1 ;
        RECT 2359.410 17.920 2359.730 17.980 ;
        RECT 2642.785 17.920 2643.075 17.965 ;
        RECT 2359.410 17.780 2643.075 17.920 ;
        RECT 2359.410 17.720 2359.730 17.780 ;
        RECT 2642.785 17.735 2643.075 17.780 ;
        RECT 2642.785 16.560 2643.075 16.605 ;
        RECT 2661.170 16.560 2661.490 16.620 ;
        RECT 2642.785 16.420 2661.490 16.560 ;
        RECT 2642.785 16.375 2643.075 16.420 ;
        RECT 2661.170 16.360 2661.490 16.420 ;
      LAYER via ;
        RECT 2359.440 17.720 2359.700 17.980 ;
        RECT 2661.200 16.360 2661.460 16.620 ;
      LAYER met2 ;
        RECT 2356.630 260.170 2356.910 264.000 ;
        RECT 2356.630 260.030 2359.640 260.170 ;
        RECT 2356.630 260.000 2356.910 260.030 ;
        RECT 2359.500 18.010 2359.640 260.030 ;
        RECT 2359.440 17.690 2359.700 18.010 ;
        RECT 2661.200 16.330 2661.460 16.650 ;
        RECT 2661.260 2.400 2661.400 16.330 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2374.130 245.720 2374.450 245.780 ;
        RECT 2677.270 245.720 2677.590 245.780 ;
        RECT 2374.130 245.580 2677.590 245.720 ;
        RECT 2374.130 245.520 2374.450 245.580 ;
        RECT 2677.270 245.520 2677.590 245.580 ;
      LAYER via ;
        RECT 2374.160 245.520 2374.420 245.780 ;
        RECT 2677.300 245.520 2677.560 245.780 ;
      LAYER met2 ;
        RECT 2374.110 260.000 2374.390 264.000 ;
        RECT 2374.220 245.810 2374.360 260.000 ;
        RECT 2374.160 245.490 2374.420 245.810 ;
        RECT 2677.300 245.490 2677.560 245.810 ;
        RECT 2677.360 17.410 2677.500 245.490 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2393.910 18.940 2394.230 19.000 ;
        RECT 2696.590 18.940 2696.910 19.000 ;
        RECT 2393.910 18.800 2696.910 18.940 ;
        RECT 2393.910 18.740 2394.230 18.800 ;
        RECT 2696.590 18.740 2696.910 18.800 ;
      LAYER via ;
        RECT 2393.940 18.740 2394.200 19.000 ;
        RECT 2696.620 18.740 2696.880 19.000 ;
      LAYER met2 ;
        RECT 2392.050 260.170 2392.330 264.000 ;
        RECT 2392.050 260.030 2394.140 260.170 ;
        RECT 2392.050 260.000 2392.330 260.030 ;
        RECT 2394.000 19.030 2394.140 260.030 ;
        RECT 2393.940 18.710 2394.200 19.030 ;
        RECT 2696.620 18.710 2696.880 19.030 ;
        RECT 2696.680 2.400 2696.820 18.710 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2410.010 245.380 2410.330 245.440 ;
        RECT 2711.770 245.380 2712.090 245.440 ;
        RECT 2410.010 245.240 2712.090 245.380 ;
        RECT 2410.010 245.180 2410.330 245.240 ;
        RECT 2711.770 245.180 2712.090 245.240 ;
      LAYER via ;
        RECT 2410.040 245.180 2410.300 245.440 ;
        RECT 2711.800 245.180 2712.060 245.440 ;
      LAYER met2 ;
        RECT 2409.990 260.000 2410.270 264.000 ;
        RECT 2410.100 245.470 2410.240 260.000 ;
        RECT 2410.040 245.150 2410.300 245.470 ;
        RECT 2711.800 245.150 2712.060 245.470 ;
        RECT 2711.860 17.410 2712.000 245.150 ;
        RECT 2711.860 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2427.930 260.170 2428.210 264.000 ;
        RECT 2427.930 260.030 2428.640 260.170 ;
        RECT 2427.930 260.000 2428.210 260.030 ;
        RECT 2428.500 17.525 2428.640 260.030 ;
        RECT 2428.430 17.155 2428.710 17.525 ;
        RECT 2732.490 17.155 2732.770 17.525 ;
        RECT 2732.560 2.400 2732.700 17.155 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 2428.430 17.200 2428.710 17.480 ;
        RECT 2732.490 17.200 2732.770 17.480 ;
      LAYER met3 ;
        RECT 2428.405 17.490 2428.735 17.505 ;
        RECT 2732.465 17.490 2732.795 17.505 ;
        RECT 2428.405 17.190 2732.795 17.490 ;
        RECT 2428.405 17.175 2428.735 17.190 ;
        RECT 2732.465 17.175 2732.795 17.190 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2445.890 246.060 2446.210 246.120 ;
        RECT 2746.270 246.060 2746.590 246.120 ;
        RECT 2445.890 245.920 2746.590 246.060 ;
        RECT 2445.890 245.860 2446.210 245.920 ;
        RECT 2746.270 245.860 2746.590 245.920 ;
      LAYER via ;
        RECT 2445.920 245.860 2446.180 246.120 ;
        RECT 2746.300 245.860 2746.560 246.120 ;
      LAYER met2 ;
        RECT 2445.870 260.000 2446.150 264.000 ;
        RECT 2445.980 246.150 2446.120 260.000 ;
        RECT 2445.920 245.830 2446.180 246.150 ;
        RECT 2746.300 245.830 2746.560 246.150 ;
        RECT 2746.360 17.410 2746.500 245.830 ;
        RECT 2746.360 17.270 2750.640 17.410 ;
        RECT 2750.500 2.400 2750.640 17.270 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2463.830 244.020 2464.150 244.080 ;
        RECT 2469.810 244.020 2470.130 244.080 ;
        RECT 2463.830 243.880 2470.130 244.020 ;
        RECT 2463.830 243.820 2464.150 243.880 ;
        RECT 2469.810 243.820 2470.130 243.880 ;
        RECT 2469.810 19.280 2470.130 19.340 ;
        RECT 2767.890 19.280 2768.210 19.340 ;
        RECT 2469.810 19.140 2768.210 19.280 ;
        RECT 2469.810 19.080 2470.130 19.140 ;
        RECT 2767.890 19.080 2768.210 19.140 ;
      LAYER via ;
        RECT 2463.860 243.820 2464.120 244.080 ;
        RECT 2469.840 243.820 2470.100 244.080 ;
        RECT 2469.840 19.080 2470.100 19.340 ;
        RECT 2767.920 19.080 2768.180 19.340 ;
      LAYER met2 ;
        RECT 2463.810 260.000 2464.090 264.000 ;
        RECT 2463.920 244.110 2464.060 260.000 ;
        RECT 2463.860 243.790 2464.120 244.110 ;
        RECT 2469.840 243.790 2470.100 244.110 ;
        RECT 2469.900 19.370 2470.040 243.790 ;
        RECT 2469.840 19.050 2470.100 19.370 ;
        RECT 2767.920 19.050 2768.180 19.370 ;
        RECT 2767.980 2.400 2768.120 19.050 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 533.210 244.020 533.530 244.080 ;
        RECT 537.810 244.020 538.130 244.080 ;
        RECT 533.210 243.880 538.130 244.020 ;
        RECT 533.210 243.820 533.530 243.880 ;
        RECT 537.810 243.820 538.130 243.880 ;
        RECT 537.810 15.540 538.130 15.600 ;
        RECT 840.950 15.540 841.270 15.600 ;
        RECT 537.810 15.400 841.270 15.540 ;
        RECT 537.810 15.340 538.130 15.400 ;
        RECT 840.950 15.340 841.270 15.400 ;
      LAYER via ;
        RECT 533.240 243.820 533.500 244.080 ;
        RECT 537.840 243.820 538.100 244.080 ;
        RECT 537.840 15.340 538.100 15.600 ;
        RECT 840.980 15.340 841.240 15.600 ;
      LAYER met2 ;
        RECT 533.190 260.000 533.470 264.000 ;
        RECT 533.300 244.110 533.440 260.000 ;
        RECT 533.240 243.790 533.500 244.110 ;
        RECT 537.840 243.790 538.100 244.110 ;
        RECT 537.900 15.630 538.040 243.790 ;
        RECT 537.840 15.310 538.100 15.630 ;
        RECT 840.980 15.310 841.240 15.630 ;
        RECT 841.040 2.400 841.180 15.310 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2483.610 20.640 2483.930 20.700 ;
        RECT 2785.830 20.640 2786.150 20.700 ;
        RECT 2483.610 20.500 2786.150 20.640 ;
        RECT 2483.610 20.440 2483.930 20.500 ;
        RECT 2785.830 20.440 2786.150 20.500 ;
      LAYER via ;
        RECT 2483.640 20.440 2483.900 20.700 ;
        RECT 2785.860 20.440 2786.120 20.700 ;
      LAYER met2 ;
        RECT 2481.750 260.170 2482.030 264.000 ;
        RECT 2481.750 260.030 2483.840 260.170 ;
        RECT 2481.750 260.000 2482.030 260.030 ;
        RECT 2483.700 20.730 2483.840 260.030 ;
        RECT 2483.640 20.410 2483.900 20.730 ;
        RECT 2785.860 20.410 2786.120 20.730 ;
        RECT 2785.920 2.400 2786.060 20.410 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2499.250 244.020 2499.570 244.080 ;
        RECT 2504.310 244.020 2504.630 244.080 ;
        RECT 2499.250 243.880 2504.630 244.020 ;
        RECT 2499.250 243.820 2499.570 243.880 ;
        RECT 2504.310 243.820 2504.630 243.880 ;
        RECT 2504.310 19.620 2504.630 19.680 ;
        RECT 2803.770 19.620 2804.090 19.680 ;
        RECT 2504.310 19.480 2804.090 19.620 ;
        RECT 2504.310 19.420 2504.630 19.480 ;
        RECT 2803.770 19.420 2804.090 19.480 ;
      LAYER via ;
        RECT 2499.280 243.820 2499.540 244.080 ;
        RECT 2504.340 243.820 2504.600 244.080 ;
        RECT 2504.340 19.420 2504.600 19.680 ;
        RECT 2803.800 19.420 2804.060 19.680 ;
      LAYER met2 ;
        RECT 2499.230 260.000 2499.510 264.000 ;
        RECT 2499.340 244.110 2499.480 260.000 ;
        RECT 2499.280 243.790 2499.540 244.110 ;
        RECT 2504.340 243.790 2504.600 244.110 ;
        RECT 2504.400 19.710 2504.540 243.790 ;
        RECT 2504.340 19.390 2504.600 19.710 ;
        RECT 2803.800 19.390 2804.060 19.710 ;
        RECT 2803.860 2.400 2804.000 19.390 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2517.190 18.260 2517.510 18.320 ;
        RECT 2821.710 18.260 2822.030 18.320 ;
        RECT 2517.190 18.120 2822.030 18.260 ;
        RECT 2517.190 18.060 2517.510 18.120 ;
        RECT 2821.710 18.060 2822.030 18.120 ;
      LAYER via ;
        RECT 2517.220 18.060 2517.480 18.320 ;
        RECT 2821.740 18.060 2822.000 18.320 ;
      LAYER met2 ;
        RECT 2517.170 260.170 2517.450 264.000 ;
        RECT 2517.170 260.030 2518.340 260.170 ;
        RECT 2517.170 260.000 2517.450 260.030 ;
        RECT 2518.200 34.410 2518.340 260.030 ;
        RECT 2517.280 34.270 2518.340 34.410 ;
        RECT 2517.280 18.350 2517.420 34.270 ;
        RECT 2517.220 18.030 2517.480 18.350 ;
        RECT 2821.740 18.030 2822.000 18.350 ;
        RECT 2821.800 2.400 2821.940 18.030 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2538.810 17.580 2539.130 17.640 ;
        RECT 2839.190 17.580 2839.510 17.640 ;
        RECT 2538.810 17.440 2839.510 17.580 ;
        RECT 2538.810 17.380 2539.130 17.440 ;
        RECT 2839.190 17.380 2839.510 17.440 ;
      LAYER via ;
        RECT 2538.840 17.380 2539.100 17.640 ;
        RECT 2839.220 17.380 2839.480 17.640 ;
      LAYER met2 ;
        RECT 2535.110 260.170 2535.390 264.000 ;
        RECT 2535.110 260.030 2539.040 260.170 ;
        RECT 2535.110 260.000 2535.390 260.030 ;
        RECT 2538.900 17.670 2539.040 260.030 ;
        RECT 2538.840 17.350 2539.100 17.670 ;
        RECT 2839.220 17.350 2839.480 17.670 ;
        RECT 2839.280 2.400 2839.420 17.350 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2553.070 242.660 2553.390 242.720 ;
        RECT 2559.510 242.660 2559.830 242.720 ;
        RECT 2553.070 242.520 2559.830 242.660 ;
        RECT 2553.070 242.460 2553.390 242.520 ;
        RECT 2559.510 242.460 2559.830 242.520 ;
        RECT 2559.510 16.220 2559.830 16.280 ;
        RECT 2857.130 16.220 2857.450 16.280 ;
        RECT 2559.510 16.080 2857.450 16.220 ;
        RECT 2559.510 16.020 2559.830 16.080 ;
        RECT 2857.130 16.020 2857.450 16.080 ;
      LAYER via ;
        RECT 2553.100 242.460 2553.360 242.720 ;
        RECT 2559.540 242.460 2559.800 242.720 ;
        RECT 2559.540 16.020 2559.800 16.280 ;
        RECT 2857.160 16.020 2857.420 16.280 ;
      LAYER met2 ;
        RECT 2553.050 260.000 2553.330 264.000 ;
        RECT 2553.160 242.750 2553.300 260.000 ;
        RECT 2553.100 242.430 2553.360 242.750 ;
        RECT 2559.540 242.430 2559.800 242.750 ;
        RECT 2559.600 16.310 2559.740 242.430 ;
        RECT 2559.540 15.990 2559.800 16.310 ;
        RECT 2857.160 15.990 2857.420 16.310 ;
        RECT 2857.220 2.400 2857.360 15.990 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 19.960 2573.630 20.020 ;
        RECT 2875.070 19.960 2875.390 20.020 ;
        RECT 2573.310 19.820 2875.390 19.960 ;
        RECT 2573.310 19.760 2573.630 19.820 ;
        RECT 2875.070 19.760 2875.390 19.820 ;
      LAYER via ;
        RECT 2573.340 19.760 2573.600 20.020 ;
        RECT 2875.100 19.760 2875.360 20.020 ;
      LAYER met2 ;
        RECT 2570.990 260.170 2571.270 264.000 ;
        RECT 2570.990 260.030 2573.540 260.170 ;
        RECT 2570.990 260.000 2571.270 260.030 ;
        RECT 2573.400 20.050 2573.540 260.030 ;
        RECT 2573.340 19.730 2573.600 20.050 ;
        RECT 2875.100 19.730 2875.360 20.050 ;
        RECT 2875.160 2.400 2875.300 19.730 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2588.950 244.020 2589.270 244.080 ;
        RECT 2594.010 244.020 2594.330 244.080 ;
        RECT 2588.950 243.880 2594.330 244.020 ;
        RECT 2588.950 243.820 2589.270 243.880 ;
        RECT 2594.010 243.820 2594.330 243.880 ;
        RECT 2594.010 17.240 2594.330 17.300 ;
        RECT 2893.010 17.240 2893.330 17.300 ;
        RECT 2594.010 17.100 2893.330 17.240 ;
        RECT 2594.010 17.040 2594.330 17.100 ;
        RECT 2893.010 17.040 2893.330 17.100 ;
      LAYER via ;
        RECT 2588.980 243.820 2589.240 244.080 ;
        RECT 2594.040 243.820 2594.300 244.080 ;
        RECT 2594.040 17.040 2594.300 17.300 ;
        RECT 2893.040 17.040 2893.300 17.300 ;
      LAYER met2 ;
        RECT 2588.930 260.000 2589.210 264.000 ;
        RECT 2589.040 244.110 2589.180 260.000 ;
        RECT 2588.980 243.790 2589.240 244.110 ;
        RECT 2594.040 243.790 2594.300 244.110 ;
        RECT 2594.100 17.330 2594.240 243.790 ;
        RECT 2594.040 17.010 2594.300 17.330 ;
        RECT 2893.040 17.010 2893.300 17.330 ;
        RECT 2893.100 2.400 2893.240 17.010 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2607.810 18.600 2608.130 18.660 ;
        RECT 2910.950 18.600 2911.270 18.660 ;
        RECT 2607.810 18.460 2911.270 18.600 ;
        RECT 2607.810 18.400 2608.130 18.460 ;
        RECT 2910.950 18.400 2911.270 18.460 ;
      LAYER via ;
        RECT 2607.840 18.400 2608.100 18.660 ;
        RECT 2910.980 18.400 2911.240 18.660 ;
      LAYER met2 ;
        RECT 2606.870 260.170 2607.150 264.000 ;
        RECT 2606.870 260.030 2608.040 260.170 ;
        RECT 2606.870 260.000 2607.150 260.030 ;
        RECT 2607.900 18.690 2608.040 260.030 ;
        RECT 2607.840 18.370 2608.100 18.690 ;
        RECT 2910.980 18.370 2911.240 18.690 ;
        RECT 2911.040 2.400 2911.180 18.370 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 18.940 551.930 19.000 ;
        RECT 858.890 18.940 859.210 19.000 ;
        RECT 551.610 18.800 859.210 18.940 ;
        RECT 551.610 18.740 551.930 18.800 ;
        RECT 858.890 18.740 859.210 18.800 ;
      LAYER via ;
        RECT 551.640 18.740 551.900 19.000 ;
        RECT 858.920 18.740 859.180 19.000 ;
      LAYER met2 ;
        RECT 551.130 260.170 551.410 264.000 ;
        RECT 551.130 260.030 551.840 260.170 ;
        RECT 551.130 260.000 551.410 260.030 ;
        RECT 551.700 19.030 551.840 260.030 ;
        RECT 551.640 18.710 551.900 19.030 ;
        RECT 858.920 18.710 859.180 19.030 ;
        RECT 858.980 2.400 859.120 18.710 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 568.630 244.020 568.950 244.080 ;
        RECT 572.310 244.020 572.630 244.080 ;
        RECT 568.630 243.880 572.630 244.020 ;
        RECT 568.630 243.820 568.950 243.880 ;
        RECT 572.310 243.820 572.630 243.880 ;
        RECT 572.310 18.600 572.630 18.660 ;
        RECT 876.370 18.600 876.690 18.660 ;
        RECT 572.310 18.460 876.690 18.600 ;
        RECT 572.310 18.400 572.630 18.460 ;
        RECT 876.370 18.400 876.690 18.460 ;
      LAYER via ;
        RECT 568.660 243.820 568.920 244.080 ;
        RECT 572.340 243.820 572.600 244.080 ;
        RECT 572.340 18.400 572.600 18.660 ;
        RECT 876.400 18.400 876.660 18.660 ;
      LAYER met2 ;
        RECT 568.610 260.000 568.890 264.000 ;
        RECT 568.720 244.110 568.860 260.000 ;
        RECT 568.660 243.790 568.920 244.110 ;
        RECT 572.340 243.790 572.600 244.110 ;
        RECT 572.400 18.690 572.540 243.790 ;
        RECT 572.340 18.370 572.600 18.690 ;
        RECT 876.400 18.370 876.660 18.690 ;
        RECT 876.460 18.090 876.600 18.370 ;
        RECT 876.460 17.950 877.060 18.090 ;
        RECT 876.920 2.400 877.060 17.950 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.570 244.020 586.890 244.080 ;
        RECT 593.010 244.020 593.330 244.080 ;
        RECT 586.570 243.880 593.330 244.020 ;
        RECT 586.570 243.820 586.890 243.880 ;
        RECT 593.010 243.820 593.330 243.880 ;
        RECT 593.010 16.220 593.330 16.280 ;
        RECT 894.770 16.220 895.090 16.280 ;
        RECT 593.010 16.080 895.090 16.220 ;
        RECT 593.010 16.020 593.330 16.080 ;
        RECT 894.770 16.020 895.090 16.080 ;
      LAYER via ;
        RECT 586.600 243.820 586.860 244.080 ;
        RECT 593.040 243.820 593.300 244.080 ;
        RECT 593.040 16.020 593.300 16.280 ;
        RECT 894.800 16.020 895.060 16.280 ;
      LAYER met2 ;
        RECT 586.550 260.000 586.830 264.000 ;
        RECT 586.660 244.110 586.800 260.000 ;
        RECT 586.600 243.790 586.860 244.110 ;
        RECT 593.040 243.790 593.300 244.110 ;
        RECT 593.100 16.310 593.240 243.790 ;
        RECT 593.040 15.990 593.300 16.310 ;
        RECT 894.800 15.990 895.060 16.310 ;
        RECT 894.860 2.400 895.000 15.990 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 18.260 607.130 18.320 ;
        RECT 912.710 18.260 913.030 18.320 ;
        RECT 606.810 18.120 913.030 18.260 ;
        RECT 606.810 18.060 607.130 18.120 ;
        RECT 912.710 18.060 913.030 18.120 ;
      LAYER via ;
        RECT 606.840 18.060 607.100 18.320 ;
        RECT 912.740 18.060 913.000 18.320 ;
      LAYER met2 ;
        RECT 604.490 260.170 604.770 264.000 ;
        RECT 604.490 260.030 607.040 260.170 ;
        RECT 604.490 260.000 604.770 260.030 ;
        RECT 606.900 18.350 607.040 260.030 ;
        RECT 606.840 18.030 607.100 18.350 ;
        RECT 912.740 18.030 913.000 18.350 ;
        RECT 912.800 2.400 912.940 18.030 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 622.450 244.020 622.770 244.080 ;
        RECT 627.510 244.020 627.830 244.080 ;
        RECT 622.450 243.880 627.830 244.020 ;
        RECT 622.450 243.820 622.770 243.880 ;
        RECT 627.510 243.820 627.830 243.880 ;
        RECT 627.510 20.300 627.830 20.360 ;
        RECT 930.190 20.300 930.510 20.360 ;
        RECT 627.510 20.160 930.510 20.300 ;
        RECT 627.510 20.100 627.830 20.160 ;
        RECT 930.190 20.100 930.510 20.160 ;
      LAYER via ;
        RECT 622.480 243.820 622.740 244.080 ;
        RECT 627.540 243.820 627.800 244.080 ;
        RECT 627.540 20.100 627.800 20.360 ;
        RECT 930.220 20.100 930.480 20.360 ;
      LAYER met2 ;
        RECT 622.430 260.000 622.710 264.000 ;
        RECT 622.540 244.110 622.680 260.000 ;
        RECT 622.480 243.790 622.740 244.110 ;
        RECT 627.540 243.790 627.800 244.110 ;
        RECT 627.600 20.390 627.740 243.790 ;
        RECT 627.540 20.070 627.800 20.390 ;
        RECT 930.220 20.070 930.480 20.390 ;
        RECT 930.280 2.400 930.420 20.070 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 641.310 19.280 641.630 19.340 ;
        RECT 948.130 19.280 948.450 19.340 ;
        RECT 641.310 19.140 948.450 19.280 ;
        RECT 641.310 19.080 641.630 19.140 ;
        RECT 948.130 19.080 948.450 19.140 ;
      LAYER via ;
        RECT 641.340 19.080 641.600 19.340 ;
        RECT 948.160 19.080 948.420 19.340 ;
      LAYER met2 ;
        RECT 640.370 260.170 640.650 264.000 ;
        RECT 640.370 260.030 641.540 260.170 ;
        RECT 640.370 260.000 640.650 260.030 ;
        RECT 641.400 19.370 641.540 260.030 ;
        RECT 641.340 19.050 641.600 19.370 ;
        RECT 948.160 19.050 948.420 19.370 ;
        RECT 948.220 2.400 948.360 19.050 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.010 17.920 662.330 17.980 ;
        RECT 966.070 17.920 966.390 17.980 ;
        RECT 662.010 17.780 966.390 17.920 ;
        RECT 662.010 17.720 662.330 17.780 ;
        RECT 966.070 17.720 966.390 17.780 ;
      LAYER via ;
        RECT 662.040 17.720 662.300 17.980 ;
        RECT 966.100 17.720 966.360 17.980 ;
      LAYER met2 ;
        RECT 658.310 260.170 658.590 264.000 ;
        RECT 658.310 260.030 662.240 260.170 ;
        RECT 658.310 260.000 658.590 260.030 ;
        RECT 662.100 18.010 662.240 260.030 ;
        RECT 662.040 17.690 662.300 18.010 ;
        RECT 966.100 17.690 966.360 18.010 ;
        RECT 966.160 2.400 966.300 17.690 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 676.270 244.020 676.590 244.080 ;
        RECT 682.250 244.020 682.570 244.080 ;
        RECT 676.270 243.880 682.570 244.020 ;
        RECT 676.270 243.820 676.590 243.880 ;
        RECT 682.250 243.820 682.570 243.880 ;
        RECT 682.250 16.900 682.570 16.960 ;
        RECT 984.010 16.900 984.330 16.960 ;
        RECT 682.250 16.760 984.330 16.900 ;
        RECT 682.250 16.700 682.570 16.760 ;
        RECT 984.010 16.700 984.330 16.760 ;
      LAYER via ;
        RECT 676.300 243.820 676.560 244.080 ;
        RECT 682.280 243.820 682.540 244.080 ;
        RECT 682.280 16.700 682.540 16.960 ;
        RECT 984.040 16.700 984.300 16.960 ;
      LAYER met2 ;
        RECT 676.250 260.000 676.530 264.000 ;
        RECT 676.360 244.110 676.500 260.000 ;
        RECT 676.300 243.790 676.560 244.110 ;
        RECT 682.280 243.790 682.540 244.110 ;
        RECT 682.340 16.990 682.480 243.790 ;
        RECT 682.280 16.670 682.540 16.990 ;
        RECT 984.040 16.670 984.300 16.990 ;
        RECT 984.100 2.400 984.240 16.670 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 354.270 244.020 354.590 244.080 ;
        RECT 358.410 244.020 358.730 244.080 ;
        RECT 354.270 243.880 358.730 244.020 ;
        RECT 354.270 243.820 354.590 243.880 ;
        RECT 358.410 243.820 358.730 243.880 ;
        RECT 358.410 17.240 358.730 17.300 ;
        RECT 358.410 17.100 663.160 17.240 ;
        RECT 358.410 17.040 358.730 17.100 ;
        RECT 663.020 16.960 663.160 17.100 ;
        RECT 662.930 16.700 663.250 16.960 ;
      LAYER via ;
        RECT 354.300 243.820 354.560 244.080 ;
        RECT 358.440 243.820 358.700 244.080 ;
        RECT 358.440 17.040 358.700 17.300 ;
        RECT 662.960 16.700 663.220 16.960 ;
      LAYER met2 ;
        RECT 354.250 260.000 354.530 264.000 ;
        RECT 354.360 244.110 354.500 260.000 ;
        RECT 354.300 243.790 354.560 244.110 ;
        RECT 358.440 243.790 358.700 244.110 ;
        RECT 358.500 17.330 358.640 243.790 ;
        RECT 358.440 17.010 358.700 17.330 ;
        RECT 662.960 16.670 663.220 16.990 ;
        RECT 663.020 2.400 663.160 16.670 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.510 17.580 696.830 17.640 ;
        RECT 1001.950 17.580 1002.270 17.640 ;
        RECT 696.510 17.440 1002.270 17.580 ;
        RECT 696.510 17.380 696.830 17.440 ;
        RECT 1001.950 17.380 1002.270 17.440 ;
      LAYER via ;
        RECT 696.540 17.380 696.800 17.640 ;
        RECT 1001.980 17.380 1002.240 17.640 ;
      LAYER met2 ;
        RECT 694.190 260.170 694.470 264.000 ;
        RECT 694.190 260.030 696.740 260.170 ;
        RECT 694.190 260.000 694.470 260.030 ;
        RECT 696.600 17.670 696.740 260.030 ;
        RECT 696.540 17.350 696.800 17.670 ;
        RECT 1001.980 17.350 1002.240 17.670 ;
        RECT 1002.040 2.400 1002.180 17.350 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 711.690 244.020 712.010 244.080 ;
        RECT 717.210 244.020 717.530 244.080 ;
        RECT 711.690 243.880 717.530 244.020 ;
        RECT 711.690 243.820 712.010 243.880 ;
        RECT 717.210 243.820 717.530 243.880 ;
        RECT 717.210 20.640 717.530 20.700 ;
        RECT 1019.430 20.640 1019.750 20.700 ;
        RECT 717.210 20.500 1019.750 20.640 ;
        RECT 717.210 20.440 717.530 20.500 ;
        RECT 1019.430 20.440 1019.750 20.500 ;
      LAYER via ;
        RECT 711.720 243.820 711.980 244.080 ;
        RECT 717.240 243.820 717.500 244.080 ;
        RECT 717.240 20.440 717.500 20.700 ;
        RECT 1019.460 20.440 1019.720 20.700 ;
      LAYER met2 ;
        RECT 711.670 260.000 711.950 264.000 ;
        RECT 711.780 244.110 711.920 260.000 ;
        RECT 711.720 243.790 711.980 244.110 ;
        RECT 717.240 243.790 717.500 244.110 ;
        RECT 717.300 20.730 717.440 243.790 ;
        RECT 717.240 20.410 717.500 20.730 ;
        RECT 1019.460 20.410 1019.720 20.730 ;
        RECT 1019.520 2.400 1019.660 20.410 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 729.630 245.040 729.950 245.100 ;
        RECT 1035.530 245.040 1035.850 245.100 ;
        RECT 729.630 244.900 1035.850 245.040 ;
        RECT 729.630 244.840 729.950 244.900 ;
        RECT 1035.530 244.840 1035.850 244.900 ;
      LAYER via ;
        RECT 729.660 244.840 729.920 245.100 ;
        RECT 1035.560 244.840 1035.820 245.100 ;
      LAYER met2 ;
        RECT 729.610 260.000 729.890 264.000 ;
        RECT 729.720 245.130 729.860 260.000 ;
        RECT 729.660 244.810 729.920 245.130 ;
        RECT 1035.560 244.810 1035.820 245.130 ;
        RECT 1035.620 16.730 1035.760 244.810 ;
        RECT 1035.620 16.590 1037.600 16.730 ;
        RECT 1037.460 2.400 1037.600 16.590 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 747.570 244.020 747.890 244.080 ;
        RECT 751.710 244.020 752.030 244.080 ;
        RECT 747.570 243.880 752.030 244.020 ;
        RECT 747.570 243.820 747.890 243.880 ;
        RECT 751.710 243.820 752.030 243.880 ;
        RECT 751.710 16.560 752.030 16.620 ;
        RECT 1055.310 16.560 1055.630 16.620 ;
        RECT 751.710 16.420 1055.630 16.560 ;
        RECT 751.710 16.360 752.030 16.420 ;
        RECT 1055.310 16.360 1055.630 16.420 ;
      LAYER via ;
        RECT 747.600 243.820 747.860 244.080 ;
        RECT 751.740 243.820 752.000 244.080 ;
        RECT 751.740 16.360 752.000 16.620 ;
        RECT 1055.340 16.360 1055.600 16.620 ;
      LAYER met2 ;
        RECT 747.550 260.000 747.830 264.000 ;
        RECT 747.660 244.110 747.800 260.000 ;
        RECT 747.600 243.790 747.860 244.110 ;
        RECT 751.740 243.790 752.000 244.110 ;
        RECT 751.800 16.650 751.940 243.790 ;
        RECT 751.740 16.330 752.000 16.650 ;
        RECT 1055.340 16.330 1055.600 16.650 ;
        RECT 1055.400 2.400 1055.540 16.330 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.490 260.000 765.770 264.000 ;
        RECT 765.600 17.525 765.740 260.000 ;
        RECT 765.530 17.155 765.810 17.525 ;
        RECT 1073.270 17.155 1073.550 17.525 ;
        RECT 1073.340 2.400 1073.480 17.155 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 765.530 17.200 765.810 17.480 ;
        RECT 1073.270 17.200 1073.550 17.480 ;
      LAYER met3 ;
        RECT 765.505 17.490 765.835 17.505 ;
        RECT 1073.245 17.490 1073.575 17.505 ;
        RECT 765.505 17.190 1073.575 17.490 ;
        RECT 765.505 17.175 765.835 17.190 ;
        RECT 1073.245 17.175 1073.575 17.190 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.430 260.170 783.710 264.000 ;
        RECT 783.430 260.030 786.440 260.170 ;
        RECT 783.430 260.000 783.710 260.030 ;
        RECT 786.300 16.845 786.440 260.030 ;
        RECT 786.230 16.475 786.510 16.845 ;
        RECT 1090.750 16.475 1091.030 16.845 ;
        RECT 1090.820 2.400 1090.960 16.475 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
      LAYER via2 ;
        RECT 786.230 16.520 786.510 16.800 ;
        RECT 1090.750 16.520 1091.030 16.800 ;
      LAYER met3 ;
        RECT 786.205 16.810 786.535 16.825 ;
        RECT 1090.725 16.810 1091.055 16.825 ;
        RECT 786.205 16.510 1091.055 16.810 ;
        RECT 786.205 16.495 786.535 16.510 ;
        RECT 1090.725 16.495 1091.055 16.510 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 801.390 244.020 801.710 244.080 ;
        RECT 806.910 244.020 807.230 244.080 ;
        RECT 801.390 243.880 807.230 244.020 ;
        RECT 801.390 243.820 801.710 243.880 ;
        RECT 806.910 243.820 807.230 243.880 ;
        RECT 806.910 19.960 807.230 20.020 ;
        RECT 1108.670 19.960 1108.990 20.020 ;
        RECT 806.910 19.820 1108.990 19.960 ;
        RECT 806.910 19.760 807.230 19.820 ;
        RECT 1108.670 19.760 1108.990 19.820 ;
      LAYER via ;
        RECT 801.420 243.820 801.680 244.080 ;
        RECT 806.940 243.820 807.200 244.080 ;
        RECT 806.940 19.760 807.200 20.020 ;
        RECT 1108.700 19.760 1108.960 20.020 ;
      LAYER met2 ;
        RECT 801.370 260.000 801.650 264.000 ;
        RECT 801.480 244.110 801.620 260.000 ;
        RECT 801.420 243.790 801.680 244.110 ;
        RECT 806.940 243.790 807.200 244.110 ;
        RECT 807.000 20.050 807.140 243.790 ;
        RECT 806.940 19.730 807.200 20.050 ;
        RECT 1108.700 19.730 1108.960 20.050 ;
        RECT 1108.760 2.400 1108.900 19.730 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 820.710 17.240 821.030 17.300 ;
        RECT 1126.610 17.240 1126.930 17.300 ;
        RECT 820.710 17.100 1126.930 17.240 ;
        RECT 820.710 17.040 821.030 17.100 ;
        RECT 1126.610 17.040 1126.930 17.100 ;
      LAYER via ;
        RECT 820.740 17.040 821.000 17.300 ;
        RECT 1126.640 17.040 1126.900 17.300 ;
      LAYER met2 ;
        RECT 819.310 260.170 819.590 264.000 ;
        RECT 819.310 260.030 820.940 260.170 ;
        RECT 819.310 260.000 819.590 260.030 ;
        RECT 820.800 17.330 820.940 260.030 ;
        RECT 820.740 17.010 821.000 17.330 ;
        RECT 1126.640 17.010 1126.900 17.330 ;
        RECT 1126.700 2.400 1126.840 17.010 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 836.810 245.720 837.130 245.780 ;
        RECT 1139.490 245.720 1139.810 245.780 ;
        RECT 836.810 245.580 1139.810 245.720 ;
        RECT 836.810 245.520 837.130 245.580 ;
        RECT 1139.490 245.520 1139.810 245.580 ;
      LAYER via ;
        RECT 836.840 245.520 837.100 245.780 ;
        RECT 1139.520 245.520 1139.780 245.780 ;
      LAYER met2 ;
        RECT 836.790 260.000 837.070 264.000 ;
        RECT 836.900 245.810 837.040 260.000 ;
        RECT 836.840 245.490 837.100 245.810 ;
        RECT 1139.520 245.490 1139.780 245.810 ;
        RECT 1139.580 16.730 1139.720 245.490 ;
        RECT 1139.580 16.590 1144.780 16.730 ;
        RECT 1144.640 2.400 1144.780 16.590 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 855.210 19.620 855.530 19.680 ;
        RECT 1162.490 19.620 1162.810 19.680 ;
        RECT 855.210 19.480 1162.810 19.620 ;
        RECT 855.210 19.420 855.530 19.480 ;
        RECT 1162.490 19.420 1162.810 19.480 ;
      LAYER via ;
        RECT 855.240 19.420 855.500 19.680 ;
        RECT 1162.520 19.420 1162.780 19.680 ;
      LAYER met2 ;
        RECT 854.730 260.170 855.010 264.000 ;
        RECT 854.730 260.030 855.440 260.170 ;
        RECT 854.730 260.000 855.010 260.030 ;
        RECT 855.300 19.710 855.440 260.030 ;
        RECT 855.240 19.390 855.500 19.710 ;
        RECT 1162.520 19.390 1162.780 19.710 ;
        RECT 1162.580 2.400 1162.720 19.390 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 246.400 372.530 246.460 ;
        RECT 677.190 246.400 677.510 246.460 ;
        RECT 372.210 246.260 677.510 246.400 ;
        RECT 372.210 246.200 372.530 246.260 ;
        RECT 677.190 246.200 677.510 246.260 ;
      LAYER via ;
        RECT 372.240 246.200 372.500 246.460 ;
        RECT 677.220 246.200 677.480 246.460 ;
      LAYER met2 ;
        RECT 372.190 260.000 372.470 264.000 ;
        RECT 372.300 246.490 372.440 260.000 ;
        RECT 372.240 246.170 372.500 246.490 ;
        RECT 677.220 246.170 677.480 246.490 ;
        RECT 677.280 16.730 677.420 246.170 ;
        RECT 677.280 16.590 680.640 16.730 ;
        RECT 680.500 2.400 680.640 16.590 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 875.910 18.940 876.230 19.000 ;
        RECT 1179.970 18.940 1180.290 19.000 ;
        RECT 875.910 18.800 1180.290 18.940 ;
        RECT 875.910 18.740 876.230 18.800 ;
        RECT 1179.970 18.740 1180.290 18.800 ;
      LAYER via ;
        RECT 875.940 18.740 876.200 19.000 ;
        RECT 1180.000 18.740 1180.260 19.000 ;
      LAYER met2 ;
        RECT 872.670 260.170 872.950 264.000 ;
        RECT 872.670 260.030 876.140 260.170 ;
        RECT 872.670 260.000 872.950 260.030 ;
        RECT 876.000 19.030 876.140 260.030 ;
        RECT 875.940 18.710 876.200 19.030 ;
        RECT 1180.000 18.710 1180.260 19.030 ;
        RECT 1180.060 2.400 1180.200 18.710 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 890.630 244.020 890.950 244.080 ;
        RECT 896.610 244.020 896.930 244.080 ;
        RECT 890.630 243.880 896.930 244.020 ;
        RECT 890.630 243.820 890.950 243.880 ;
        RECT 896.610 243.820 896.930 243.880 ;
        RECT 896.610 16.220 896.930 16.280 ;
        RECT 1197.910 16.220 1198.230 16.280 ;
        RECT 896.610 16.080 1198.230 16.220 ;
        RECT 896.610 16.020 896.930 16.080 ;
        RECT 1197.910 16.020 1198.230 16.080 ;
      LAYER via ;
        RECT 890.660 243.820 890.920 244.080 ;
        RECT 896.640 243.820 896.900 244.080 ;
        RECT 896.640 16.020 896.900 16.280 ;
        RECT 1197.940 16.020 1198.200 16.280 ;
      LAYER met2 ;
        RECT 890.610 260.000 890.890 264.000 ;
        RECT 890.720 244.110 890.860 260.000 ;
        RECT 890.660 243.790 890.920 244.110 ;
        RECT 896.640 243.790 896.900 244.110 ;
        RECT 896.700 16.310 896.840 243.790 ;
        RECT 896.640 15.990 896.900 16.310 ;
        RECT 1197.940 15.990 1198.200 16.310 ;
        RECT 1198.000 2.400 1198.140 15.990 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 910.410 18.600 910.730 18.660 ;
        RECT 1215.850 18.600 1216.170 18.660 ;
        RECT 910.410 18.460 1216.170 18.600 ;
        RECT 910.410 18.400 910.730 18.460 ;
        RECT 1215.850 18.400 1216.170 18.460 ;
      LAYER via ;
        RECT 910.440 18.400 910.700 18.660 ;
        RECT 1215.880 18.400 1216.140 18.660 ;
      LAYER met2 ;
        RECT 908.550 260.170 908.830 264.000 ;
        RECT 908.550 260.030 910.640 260.170 ;
        RECT 908.550 260.000 908.830 260.030 ;
        RECT 910.500 18.690 910.640 260.030 ;
        RECT 910.440 18.370 910.700 18.690 ;
        RECT 1215.880 18.370 1216.140 18.690 ;
        RECT 1215.940 2.400 1216.080 18.370 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 926.510 244.020 926.830 244.080 ;
        RECT 931.110 244.020 931.430 244.080 ;
        RECT 926.510 243.880 931.430 244.020 ;
        RECT 926.510 243.820 926.830 243.880 ;
        RECT 931.110 243.820 931.430 243.880 ;
        RECT 931.110 15.540 931.430 15.600 ;
        RECT 1233.790 15.540 1234.110 15.600 ;
        RECT 931.110 15.400 1234.110 15.540 ;
        RECT 931.110 15.340 931.430 15.400 ;
        RECT 1233.790 15.340 1234.110 15.400 ;
      LAYER via ;
        RECT 926.540 243.820 926.800 244.080 ;
        RECT 931.140 243.820 931.400 244.080 ;
        RECT 931.140 15.340 931.400 15.600 ;
        RECT 1233.820 15.340 1234.080 15.600 ;
      LAYER met2 ;
        RECT 926.490 260.000 926.770 264.000 ;
        RECT 926.600 244.110 926.740 260.000 ;
        RECT 926.540 243.790 926.800 244.110 ;
        RECT 931.140 243.790 931.400 244.110 ;
        RECT 931.200 15.630 931.340 243.790 ;
        RECT 931.140 15.310 931.400 15.630 ;
        RECT 1233.820 15.310 1234.080 15.630 ;
        RECT 1233.880 2.400 1234.020 15.310 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 944.910 18.260 945.230 18.320 ;
        RECT 1251.730 18.260 1252.050 18.320 ;
        RECT 944.910 18.120 1252.050 18.260 ;
        RECT 944.910 18.060 945.230 18.120 ;
        RECT 1251.730 18.060 1252.050 18.120 ;
      LAYER via ;
        RECT 944.940 18.060 945.200 18.320 ;
        RECT 1251.760 18.060 1252.020 18.320 ;
      LAYER met2 ;
        RECT 944.430 260.170 944.710 264.000 ;
        RECT 944.430 260.030 945.140 260.170 ;
        RECT 944.430 260.000 944.710 260.030 ;
        RECT 945.000 18.350 945.140 260.030 ;
        RECT 944.940 18.030 945.200 18.350 ;
        RECT 1251.760 18.030 1252.020 18.350 ;
        RECT 1251.820 2.400 1251.960 18.030 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 965.610 20.300 965.930 20.360 ;
        RECT 1269.210 20.300 1269.530 20.360 ;
        RECT 965.610 20.160 1269.530 20.300 ;
        RECT 965.610 20.100 965.930 20.160 ;
        RECT 1269.210 20.100 1269.530 20.160 ;
      LAYER via ;
        RECT 965.640 20.100 965.900 20.360 ;
        RECT 1269.240 20.100 1269.500 20.360 ;
      LAYER met2 ;
        RECT 961.910 260.170 962.190 264.000 ;
        RECT 961.910 260.030 965.840 260.170 ;
        RECT 961.910 260.000 962.190 260.030 ;
        RECT 965.700 20.390 965.840 260.030 ;
        RECT 965.640 20.070 965.900 20.390 ;
        RECT 1269.240 20.070 1269.500 20.390 ;
        RECT 1269.300 2.400 1269.440 20.070 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 979.870 243.340 980.190 243.400 ;
        RECT 986.310 243.340 986.630 243.400 ;
        RECT 979.870 243.200 986.630 243.340 ;
        RECT 979.870 243.140 980.190 243.200 ;
        RECT 986.310 243.140 986.630 243.200 ;
        RECT 986.310 16.900 986.630 16.960 ;
        RECT 1287.150 16.900 1287.470 16.960 ;
        RECT 986.310 16.760 1287.470 16.900 ;
        RECT 986.310 16.700 986.630 16.760 ;
        RECT 1287.150 16.700 1287.470 16.760 ;
      LAYER via ;
        RECT 979.900 243.140 980.160 243.400 ;
        RECT 986.340 243.140 986.600 243.400 ;
        RECT 986.340 16.700 986.600 16.960 ;
        RECT 1287.180 16.700 1287.440 16.960 ;
      LAYER met2 ;
        RECT 979.850 260.000 980.130 264.000 ;
        RECT 979.960 243.430 980.100 260.000 ;
        RECT 979.900 243.110 980.160 243.430 ;
        RECT 986.340 243.110 986.600 243.430 ;
        RECT 986.400 16.990 986.540 243.110 ;
        RECT 986.340 16.670 986.600 16.990 ;
        RECT 1287.180 16.670 1287.440 16.990 ;
        RECT 1287.240 2.400 1287.380 16.670 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1000.110 17.920 1000.430 17.980 ;
        RECT 1305.090 17.920 1305.410 17.980 ;
        RECT 1000.110 17.780 1305.410 17.920 ;
        RECT 1000.110 17.720 1000.430 17.780 ;
        RECT 1305.090 17.720 1305.410 17.780 ;
      LAYER via ;
        RECT 1000.140 17.720 1000.400 17.980 ;
        RECT 1305.120 17.720 1305.380 17.980 ;
      LAYER met2 ;
        RECT 997.790 260.170 998.070 264.000 ;
        RECT 997.790 260.030 1000.340 260.170 ;
        RECT 997.790 260.000 998.070 260.030 ;
        RECT 1000.200 18.010 1000.340 260.030 ;
        RECT 1000.140 17.690 1000.400 18.010 ;
        RECT 1305.120 17.690 1305.380 18.010 ;
        RECT 1305.180 2.400 1305.320 17.690 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1015.750 244.020 1016.070 244.080 ;
        RECT 1020.810 244.020 1021.130 244.080 ;
        RECT 1015.750 243.880 1021.130 244.020 ;
        RECT 1015.750 243.820 1016.070 243.880 ;
        RECT 1020.810 243.820 1021.130 243.880 ;
        RECT 1020.810 15.880 1021.130 15.940 ;
        RECT 1323.030 15.880 1323.350 15.940 ;
        RECT 1020.810 15.740 1323.350 15.880 ;
        RECT 1020.810 15.680 1021.130 15.740 ;
        RECT 1323.030 15.680 1323.350 15.740 ;
      LAYER via ;
        RECT 1015.780 243.820 1016.040 244.080 ;
        RECT 1020.840 243.820 1021.100 244.080 ;
        RECT 1020.840 15.680 1021.100 15.940 ;
        RECT 1323.060 15.680 1323.320 15.940 ;
      LAYER met2 ;
        RECT 1015.730 260.000 1016.010 264.000 ;
        RECT 1015.840 244.110 1015.980 260.000 ;
        RECT 1015.780 243.790 1016.040 244.110 ;
        RECT 1020.840 243.790 1021.100 244.110 ;
        RECT 1020.900 15.970 1021.040 243.790 ;
        RECT 1020.840 15.650 1021.100 15.970 ;
        RECT 1323.060 15.650 1323.320 15.970 ;
        RECT 1323.120 2.400 1323.260 15.650 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1034.610 17.580 1034.930 17.640 ;
        RECT 1340.510 17.580 1340.830 17.640 ;
        RECT 1034.610 17.440 1340.830 17.580 ;
        RECT 1034.610 17.380 1034.930 17.440 ;
        RECT 1340.510 17.380 1340.830 17.440 ;
      LAYER via ;
        RECT 1034.640 17.380 1034.900 17.640 ;
        RECT 1340.540 17.380 1340.800 17.640 ;
      LAYER met2 ;
        RECT 1033.670 260.170 1033.950 264.000 ;
        RECT 1033.670 260.030 1034.840 260.170 ;
        RECT 1033.670 260.000 1033.950 260.030 ;
        RECT 1034.700 17.670 1034.840 260.030 ;
        RECT 1034.640 17.350 1034.900 17.670 ;
        RECT 1340.540 17.350 1340.800 17.670 ;
        RECT 1340.600 2.400 1340.740 17.350 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 19.960 393.230 20.020 ;
        RECT 698.350 19.960 698.670 20.020 ;
        RECT 392.910 19.820 698.670 19.960 ;
        RECT 392.910 19.760 393.230 19.820 ;
        RECT 698.350 19.760 698.670 19.820 ;
      LAYER via ;
        RECT 392.940 19.760 393.200 20.020 ;
        RECT 698.380 19.760 698.640 20.020 ;
      LAYER met2 ;
        RECT 390.130 260.170 390.410 264.000 ;
        RECT 390.130 260.030 393.140 260.170 ;
        RECT 390.130 260.000 390.410 260.030 ;
        RECT 393.000 20.050 393.140 260.030 ;
        RECT 392.940 19.730 393.200 20.050 ;
        RECT 698.380 19.730 698.640 20.050 ;
        RECT 698.440 2.400 698.580 19.730 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1051.630 246.060 1051.950 246.120 ;
        RECT 1352.470 246.060 1352.790 246.120 ;
        RECT 1051.630 245.920 1352.790 246.060 ;
        RECT 1051.630 245.860 1051.950 245.920 ;
        RECT 1352.470 245.860 1352.790 245.920 ;
        RECT 1352.470 37.640 1352.790 37.700 ;
        RECT 1358.450 37.640 1358.770 37.700 ;
        RECT 1352.470 37.500 1358.770 37.640 ;
        RECT 1352.470 37.440 1352.790 37.500 ;
        RECT 1358.450 37.440 1358.770 37.500 ;
      LAYER via ;
        RECT 1051.660 245.860 1051.920 246.120 ;
        RECT 1352.500 245.860 1352.760 246.120 ;
        RECT 1352.500 37.440 1352.760 37.700 ;
        RECT 1358.480 37.440 1358.740 37.700 ;
      LAYER met2 ;
        RECT 1051.610 260.000 1051.890 264.000 ;
        RECT 1051.720 246.150 1051.860 260.000 ;
        RECT 1051.660 245.830 1051.920 246.150 ;
        RECT 1352.500 245.830 1352.760 246.150 ;
        RECT 1352.560 37.730 1352.700 245.830 ;
        RECT 1352.500 37.410 1352.760 37.730 ;
        RECT 1358.480 37.410 1358.740 37.730 ;
        RECT 1358.540 2.400 1358.680 37.410 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1069.570 244.020 1069.890 244.080 ;
        RECT 1076.010 244.020 1076.330 244.080 ;
        RECT 1069.570 243.880 1076.330 244.020 ;
        RECT 1069.570 243.820 1069.890 243.880 ;
        RECT 1076.010 243.820 1076.330 243.880 ;
        RECT 1076.010 19.280 1076.330 19.340 ;
        RECT 1376.390 19.280 1376.710 19.340 ;
        RECT 1076.010 19.140 1376.710 19.280 ;
        RECT 1076.010 19.080 1076.330 19.140 ;
        RECT 1376.390 19.080 1376.710 19.140 ;
      LAYER via ;
        RECT 1069.600 243.820 1069.860 244.080 ;
        RECT 1076.040 243.820 1076.300 244.080 ;
        RECT 1076.040 19.080 1076.300 19.340 ;
        RECT 1376.420 19.080 1376.680 19.340 ;
      LAYER met2 ;
        RECT 1069.550 260.000 1069.830 264.000 ;
        RECT 1069.660 244.110 1069.800 260.000 ;
        RECT 1069.600 243.790 1069.860 244.110 ;
        RECT 1076.040 243.790 1076.300 244.110 ;
        RECT 1076.100 19.370 1076.240 243.790 ;
        RECT 1076.040 19.050 1076.300 19.370 ;
        RECT 1376.420 19.050 1376.680 19.370 ;
        RECT 1376.480 2.400 1376.620 19.050 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1394.865 241.485 1395.035 245.395 ;
        RECT 1394.865 48.365 1395.035 96.475 ;
      LAYER mcon ;
        RECT 1394.865 245.225 1395.035 245.395 ;
        RECT 1394.865 96.305 1395.035 96.475 ;
      LAYER met1 ;
        RECT 1087.050 245.380 1087.370 245.440 ;
        RECT 1394.805 245.380 1395.095 245.425 ;
        RECT 1087.050 245.240 1395.095 245.380 ;
        RECT 1087.050 245.180 1087.370 245.240 ;
        RECT 1394.805 245.195 1395.095 245.240 ;
        RECT 1394.790 241.640 1395.110 241.700 ;
        RECT 1394.595 241.500 1395.110 241.640 ;
        RECT 1394.790 241.440 1395.110 241.500 ;
        RECT 1394.790 96.460 1395.110 96.520 ;
        RECT 1394.595 96.320 1395.110 96.460 ;
        RECT 1394.790 96.260 1395.110 96.320 ;
        RECT 1394.790 48.520 1395.110 48.580 ;
        RECT 1394.595 48.380 1395.110 48.520 ;
        RECT 1394.790 48.320 1395.110 48.380 ;
      LAYER via ;
        RECT 1087.080 245.180 1087.340 245.440 ;
        RECT 1394.820 241.440 1395.080 241.700 ;
        RECT 1394.820 96.260 1395.080 96.520 ;
        RECT 1394.820 48.320 1395.080 48.580 ;
      LAYER met2 ;
        RECT 1087.030 260.000 1087.310 264.000 ;
        RECT 1087.140 245.470 1087.280 260.000 ;
        RECT 1087.080 245.150 1087.340 245.470 ;
        RECT 1394.820 241.410 1395.080 241.730 ;
        RECT 1394.880 96.550 1395.020 241.410 ;
        RECT 1394.820 96.230 1395.080 96.550 ;
        RECT 1394.820 48.290 1395.080 48.610 ;
        RECT 1394.880 14.690 1395.020 48.290 ;
        RECT 1394.880 14.550 1395.480 14.690 ;
        RECT 1395.340 13.330 1395.480 14.550 ;
        RECT 1394.420 13.190 1395.480 13.330 ;
        RECT 1394.420 2.400 1394.560 13.190 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1104.990 244.020 1105.310 244.080 ;
        RECT 1110.510 244.020 1110.830 244.080 ;
        RECT 1104.990 243.880 1110.830 244.020 ;
        RECT 1104.990 243.820 1105.310 243.880 ;
        RECT 1110.510 243.820 1110.830 243.880 ;
        RECT 1110.510 20.640 1110.830 20.700 ;
        RECT 1412.270 20.640 1412.590 20.700 ;
        RECT 1110.510 20.500 1412.590 20.640 ;
        RECT 1110.510 20.440 1110.830 20.500 ;
        RECT 1412.270 20.440 1412.590 20.500 ;
      LAYER via ;
        RECT 1105.020 243.820 1105.280 244.080 ;
        RECT 1110.540 243.820 1110.800 244.080 ;
        RECT 1110.540 20.440 1110.800 20.700 ;
        RECT 1412.300 20.440 1412.560 20.700 ;
      LAYER met2 ;
        RECT 1104.970 260.000 1105.250 264.000 ;
        RECT 1105.080 244.110 1105.220 260.000 ;
        RECT 1105.020 243.790 1105.280 244.110 ;
        RECT 1110.540 243.790 1110.800 244.110 ;
        RECT 1110.600 20.730 1110.740 243.790 ;
        RECT 1110.540 20.410 1110.800 20.730 ;
        RECT 1412.300 20.410 1412.560 20.730 ;
        RECT 1412.360 2.400 1412.500 20.410 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1428.905 186.405 1429.075 234.515 ;
        RECT 1428.905 48.365 1429.075 137.955 ;
      LAYER mcon ;
        RECT 1428.905 234.345 1429.075 234.515 ;
        RECT 1428.905 137.785 1429.075 137.955 ;
      LAYER met1 ;
        RECT 1122.930 245.040 1123.250 245.100 ;
        RECT 1428.830 245.040 1429.150 245.100 ;
        RECT 1122.930 244.900 1429.150 245.040 ;
        RECT 1122.930 244.840 1123.250 244.900 ;
        RECT 1428.830 244.840 1429.150 244.900 ;
        RECT 1428.830 234.500 1429.150 234.560 ;
        RECT 1428.635 234.360 1429.150 234.500 ;
        RECT 1428.830 234.300 1429.150 234.360 ;
        RECT 1428.830 186.560 1429.150 186.620 ;
        RECT 1428.635 186.420 1429.150 186.560 ;
        RECT 1428.830 186.360 1429.150 186.420 ;
        RECT 1428.830 137.940 1429.150 138.000 ;
        RECT 1428.635 137.800 1429.150 137.940 ;
        RECT 1428.830 137.740 1429.150 137.800 ;
        RECT 1428.845 48.520 1429.135 48.565 ;
        RECT 1429.750 48.520 1430.070 48.580 ;
        RECT 1428.845 48.380 1430.070 48.520 ;
        RECT 1428.845 48.335 1429.135 48.380 ;
        RECT 1429.750 48.320 1430.070 48.380 ;
      LAYER via ;
        RECT 1122.960 244.840 1123.220 245.100 ;
        RECT 1428.860 244.840 1429.120 245.100 ;
        RECT 1428.860 234.300 1429.120 234.560 ;
        RECT 1428.860 186.360 1429.120 186.620 ;
        RECT 1428.860 137.740 1429.120 138.000 ;
        RECT 1429.780 48.320 1430.040 48.580 ;
      LAYER met2 ;
        RECT 1122.910 260.000 1123.190 264.000 ;
        RECT 1123.020 245.130 1123.160 260.000 ;
        RECT 1122.960 244.810 1123.220 245.130 ;
        RECT 1428.860 244.810 1429.120 245.130 ;
        RECT 1428.920 234.590 1429.060 244.810 ;
        RECT 1428.860 234.270 1429.120 234.590 ;
        RECT 1428.860 186.330 1429.120 186.650 ;
        RECT 1428.920 138.030 1429.060 186.330 ;
        RECT 1428.860 137.710 1429.120 138.030 ;
        RECT 1429.780 48.290 1430.040 48.610 ;
        RECT 1429.840 2.400 1429.980 48.290 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1140.870 244.020 1141.190 244.080 ;
        RECT 1145.010 244.020 1145.330 244.080 ;
        RECT 1140.870 243.880 1145.330 244.020 ;
        RECT 1140.870 243.820 1141.190 243.880 ;
        RECT 1145.010 243.820 1145.330 243.880 ;
        RECT 1145.010 19.960 1145.330 20.020 ;
        RECT 1447.690 19.960 1448.010 20.020 ;
        RECT 1145.010 19.820 1448.010 19.960 ;
        RECT 1145.010 19.760 1145.330 19.820 ;
        RECT 1447.690 19.760 1448.010 19.820 ;
      LAYER via ;
        RECT 1140.900 243.820 1141.160 244.080 ;
        RECT 1145.040 243.820 1145.300 244.080 ;
        RECT 1145.040 19.760 1145.300 20.020 ;
        RECT 1447.720 19.760 1447.980 20.020 ;
      LAYER met2 ;
        RECT 1140.850 260.000 1141.130 264.000 ;
        RECT 1140.960 244.110 1141.100 260.000 ;
        RECT 1140.900 243.790 1141.160 244.110 ;
        RECT 1145.040 243.790 1145.300 244.110 ;
        RECT 1145.100 20.050 1145.240 243.790 ;
        RECT 1145.040 19.730 1145.300 20.050 ;
        RECT 1447.720 19.730 1447.980 20.050 ;
        RECT 1447.780 2.400 1447.920 19.730 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1158.790 260.000 1159.070 264.000 ;
        RECT 1158.900 16.845 1159.040 260.000 ;
        RECT 1158.830 16.475 1159.110 16.845 ;
        RECT 1465.650 16.475 1465.930 16.845 ;
        RECT 1465.720 2.400 1465.860 16.475 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
      LAYER via2 ;
        RECT 1158.830 16.520 1159.110 16.800 ;
        RECT 1465.650 16.520 1465.930 16.800 ;
      LAYER met3 ;
        RECT 1158.805 16.810 1159.135 16.825 ;
        RECT 1465.625 16.810 1465.955 16.825 ;
        RECT 1158.805 16.510 1465.955 16.810 ;
        RECT 1158.805 16.495 1159.135 16.510 ;
        RECT 1465.625 16.495 1465.955 16.510 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1176.750 244.020 1177.070 244.080 ;
        RECT 1183.190 244.020 1183.510 244.080 ;
        RECT 1176.750 243.880 1183.510 244.020 ;
        RECT 1176.750 243.820 1177.070 243.880 ;
        RECT 1183.190 243.820 1183.510 243.880 ;
        RECT 1183.190 141.680 1183.510 141.740 ;
        RECT 1483.570 141.680 1483.890 141.740 ;
        RECT 1183.190 141.540 1483.890 141.680 ;
        RECT 1183.190 141.480 1183.510 141.540 ;
        RECT 1483.570 141.480 1483.890 141.540 ;
      LAYER via ;
        RECT 1176.780 243.820 1177.040 244.080 ;
        RECT 1183.220 243.820 1183.480 244.080 ;
        RECT 1183.220 141.480 1183.480 141.740 ;
        RECT 1483.600 141.480 1483.860 141.740 ;
      LAYER met2 ;
        RECT 1176.730 260.000 1177.010 264.000 ;
        RECT 1176.840 244.110 1176.980 260.000 ;
        RECT 1176.780 243.790 1177.040 244.110 ;
        RECT 1183.220 243.790 1183.480 244.110 ;
        RECT 1183.280 141.770 1183.420 243.790 ;
        RECT 1183.220 141.450 1183.480 141.770 ;
        RECT 1483.600 141.450 1483.860 141.770 ;
        RECT 1483.660 2.400 1483.800 141.450 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.690 244.020 1195.010 244.080 ;
        RECT 1200.210 244.020 1200.530 244.080 ;
        RECT 1194.690 243.880 1200.530 244.020 ;
        RECT 1194.690 243.820 1195.010 243.880 ;
        RECT 1200.210 243.820 1200.530 243.880 ;
        RECT 1200.210 18.940 1200.530 19.000 ;
        RECT 1501.510 18.940 1501.830 19.000 ;
        RECT 1200.210 18.800 1501.830 18.940 ;
        RECT 1200.210 18.740 1200.530 18.800 ;
        RECT 1501.510 18.740 1501.830 18.800 ;
      LAYER via ;
        RECT 1194.720 243.820 1194.980 244.080 ;
        RECT 1200.240 243.820 1200.500 244.080 ;
        RECT 1200.240 18.740 1200.500 19.000 ;
        RECT 1501.540 18.740 1501.800 19.000 ;
      LAYER met2 ;
        RECT 1194.670 260.000 1194.950 264.000 ;
        RECT 1194.780 244.110 1194.920 260.000 ;
        RECT 1194.720 243.790 1194.980 244.110 ;
        RECT 1200.240 243.790 1200.500 244.110 ;
        RECT 1200.300 19.030 1200.440 243.790 ;
        RECT 1200.240 18.710 1200.500 19.030 ;
        RECT 1501.540 18.710 1501.800 19.030 ;
        RECT 1501.600 2.400 1501.740 18.710 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1212.170 237.900 1212.490 237.960 ;
        RECT 1518.070 237.900 1518.390 237.960 ;
        RECT 1212.170 237.760 1518.390 237.900 ;
        RECT 1212.170 237.700 1212.490 237.760 ;
        RECT 1518.070 237.700 1518.390 237.760 ;
      LAYER via ;
        RECT 1212.200 237.700 1212.460 237.960 ;
        RECT 1518.100 237.700 1518.360 237.960 ;
      LAYER met2 ;
        RECT 1212.150 260.000 1212.430 264.000 ;
        RECT 1212.260 237.990 1212.400 260.000 ;
        RECT 1212.200 237.670 1212.460 237.990 ;
        RECT 1518.100 237.670 1518.360 237.990 ;
        RECT 1518.160 17.410 1518.300 237.670 ;
        RECT 1518.160 17.270 1519.220 17.410 ;
        RECT 1519.080 2.400 1519.220 17.270 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 408.090 246.740 408.410 246.800 ;
        RECT 711.230 246.740 711.550 246.800 ;
        RECT 408.090 246.600 711.550 246.740 ;
        RECT 408.090 246.540 408.410 246.600 ;
        RECT 711.230 246.540 711.550 246.600 ;
      LAYER via ;
        RECT 408.120 246.540 408.380 246.800 ;
        RECT 711.260 246.540 711.520 246.800 ;
      LAYER met2 ;
        RECT 408.070 260.000 408.350 264.000 ;
        RECT 408.180 246.830 408.320 260.000 ;
        RECT 408.120 246.510 408.380 246.830 ;
        RECT 711.260 246.510 711.520 246.830 ;
        RECT 711.320 16.730 711.460 246.510 ;
        RECT 711.320 16.590 716.520 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1230.110 244.020 1230.430 244.080 ;
        RECT 1234.710 244.020 1235.030 244.080 ;
        RECT 1230.110 243.880 1235.030 244.020 ;
        RECT 1230.110 243.820 1230.430 243.880 ;
        RECT 1234.710 243.820 1235.030 243.880 ;
        RECT 1234.710 17.240 1235.030 17.300 ;
        RECT 1536.930 17.240 1537.250 17.300 ;
        RECT 1234.710 17.100 1537.250 17.240 ;
        RECT 1234.710 17.040 1235.030 17.100 ;
        RECT 1536.930 17.040 1537.250 17.100 ;
      LAYER via ;
        RECT 1230.140 243.820 1230.400 244.080 ;
        RECT 1234.740 243.820 1235.000 244.080 ;
        RECT 1234.740 17.040 1235.000 17.300 ;
        RECT 1536.960 17.040 1537.220 17.300 ;
      LAYER met2 ;
        RECT 1230.090 260.000 1230.370 264.000 ;
        RECT 1230.200 244.110 1230.340 260.000 ;
        RECT 1230.140 243.790 1230.400 244.110 ;
        RECT 1234.740 243.790 1235.000 244.110 ;
        RECT 1234.800 17.330 1234.940 243.790 ;
        RECT 1234.740 17.010 1235.000 17.330 ;
        RECT 1536.960 17.010 1537.220 17.330 ;
        RECT 1537.020 2.400 1537.160 17.010 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.510 120.940 1248.830 121.000 ;
        RECT 1552.570 120.940 1552.890 121.000 ;
        RECT 1248.510 120.800 1552.890 120.940 ;
        RECT 1248.510 120.740 1248.830 120.800 ;
        RECT 1552.570 120.740 1552.890 120.800 ;
      LAYER via ;
        RECT 1248.540 120.740 1248.800 121.000 ;
        RECT 1552.600 120.740 1552.860 121.000 ;
      LAYER met2 ;
        RECT 1248.030 260.170 1248.310 264.000 ;
        RECT 1248.030 260.030 1248.740 260.170 ;
        RECT 1248.030 260.000 1248.310 260.030 ;
        RECT 1248.600 121.030 1248.740 260.030 ;
        RECT 1248.540 120.710 1248.800 121.030 ;
        RECT 1552.600 120.710 1552.860 121.030 ;
        RECT 1552.660 16.730 1552.800 120.710 ;
        RECT 1552.660 16.590 1555.100 16.730 ;
        RECT 1554.960 2.400 1555.100 16.590 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1265.990 245.720 1266.310 245.780 ;
        RECT 1567.290 245.720 1567.610 245.780 ;
        RECT 1265.990 245.580 1567.610 245.720 ;
        RECT 1265.990 245.520 1266.310 245.580 ;
        RECT 1567.290 245.520 1567.610 245.580 ;
      LAYER via ;
        RECT 1266.020 245.520 1266.280 245.780 ;
        RECT 1567.320 245.520 1567.580 245.780 ;
      LAYER met2 ;
        RECT 1265.970 260.000 1266.250 264.000 ;
        RECT 1266.080 245.810 1266.220 260.000 ;
        RECT 1266.020 245.490 1266.280 245.810 ;
        RECT 1567.320 245.490 1567.580 245.810 ;
        RECT 1567.380 16.730 1567.520 245.490 ;
        RECT 1567.380 16.590 1573.040 16.730 ;
        RECT 1572.900 2.400 1573.040 16.590 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.930 244.020 1284.250 244.080 ;
        RECT 1289.910 244.020 1290.230 244.080 ;
        RECT 1283.930 243.880 1290.230 244.020 ;
        RECT 1283.930 243.820 1284.250 243.880 ;
        RECT 1289.910 243.820 1290.230 243.880 ;
        RECT 1289.910 45.120 1290.230 45.180 ;
        RECT 1590.290 45.120 1590.610 45.180 ;
        RECT 1289.910 44.980 1590.610 45.120 ;
        RECT 1289.910 44.920 1290.230 44.980 ;
        RECT 1590.290 44.920 1590.610 44.980 ;
      LAYER via ;
        RECT 1283.960 243.820 1284.220 244.080 ;
        RECT 1289.940 243.820 1290.200 244.080 ;
        RECT 1289.940 44.920 1290.200 45.180 ;
        RECT 1590.320 44.920 1590.580 45.180 ;
      LAYER met2 ;
        RECT 1283.910 260.000 1284.190 264.000 ;
        RECT 1284.020 244.110 1284.160 260.000 ;
        RECT 1283.960 243.790 1284.220 244.110 ;
        RECT 1289.940 243.790 1290.200 244.110 ;
        RECT 1290.000 45.210 1290.140 243.790 ;
        RECT 1289.940 44.890 1290.200 45.210 ;
        RECT 1590.320 44.890 1590.580 45.210 ;
        RECT 1590.380 2.400 1590.520 44.890 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1301.870 244.020 1302.190 244.080 ;
        RECT 1307.390 244.020 1307.710 244.080 ;
        RECT 1301.870 243.880 1307.710 244.020 ;
        RECT 1301.870 243.820 1302.190 243.880 ;
        RECT 1307.390 243.820 1307.710 243.880 ;
        RECT 1307.390 114.140 1307.710 114.200 ;
        RECT 1607.770 114.140 1608.090 114.200 ;
        RECT 1307.390 114.000 1608.090 114.140 ;
        RECT 1307.390 113.940 1307.710 114.000 ;
        RECT 1607.770 113.940 1608.090 114.000 ;
      LAYER via ;
        RECT 1301.900 243.820 1302.160 244.080 ;
        RECT 1307.420 243.820 1307.680 244.080 ;
        RECT 1307.420 113.940 1307.680 114.200 ;
        RECT 1607.800 113.940 1608.060 114.200 ;
      LAYER met2 ;
        RECT 1301.850 260.000 1302.130 264.000 ;
        RECT 1301.960 244.110 1302.100 260.000 ;
        RECT 1301.900 243.790 1302.160 244.110 ;
        RECT 1307.420 243.790 1307.680 244.110 ;
        RECT 1307.480 114.230 1307.620 243.790 ;
        RECT 1307.420 113.910 1307.680 114.230 ;
        RECT 1607.800 113.910 1608.060 114.230 ;
        RECT 1607.860 17.410 1608.000 113.910 ;
        RECT 1607.860 17.270 1608.460 17.410 ;
        RECT 1608.320 2.400 1608.460 17.270 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1319.810 243.680 1320.130 243.740 ;
        RECT 1328.090 243.680 1328.410 243.740 ;
        RECT 1319.810 243.540 1328.410 243.680 ;
        RECT 1319.810 243.480 1320.130 243.540 ;
        RECT 1328.090 243.480 1328.410 243.540 ;
        RECT 1328.090 51.920 1328.410 51.980 ;
        RECT 1621.570 51.920 1621.890 51.980 ;
        RECT 1328.090 51.780 1621.890 51.920 ;
        RECT 1328.090 51.720 1328.410 51.780 ;
        RECT 1621.570 51.720 1621.890 51.780 ;
      LAYER via ;
        RECT 1319.840 243.480 1320.100 243.740 ;
        RECT 1328.120 243.480 1328.380 243.740 ;
        RECT 1328.120 51.720 1328.380 51.980 ;
        RECT 1621.600 51.720 1621.860 51.980 ;
      LAYER met2 ;
        RECT 1319.790 260.000 1320.070 264.000 ;
        RECT 1319.900 243.770 1320.040 260.000 ;
        RECT 1319.840 243.450 1320.100 243.770 ;
        RECT 1328.120 243.450 1328.380 243.770 ;
        RECT 1328.180 52.010 1328.320 243.450 ;
        RECT 1328.120 51.690 1328.380 52.010 ;
        RECT 1621.600 51.690 1621.860 52.010 ;
        RECT 1621.660 16.730 1621.800 51.690 ;
        RECT 1621.660 16.590 1626.400 16.730 ;
        RECT 1626.260 2.400 1626.400 16.590 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1338.210 58.720 1338.530 58.780 ;
        RECT 1642.270 58.720 1642.590 58.780 ;
        RECT 1338.210 58.580 1642.590 58.720 ;
        RECT 1338.210 58.520 1338.530 58.580 ;
        RECT 1642.270 58.520 1642.590 58.580 ;
      LAYER via ;
        RECT 1338.240 58.520 1338.500 58.780 ;
        RECT 1642.300 58.520 1642.560 58.780 ;
      LAYER met2 ;
        RECT 1337.270 260.170 1337.550 264.000 ;
        RECT 1337.270 260.030 1338.440 260.170 ;
        RECT 1337.270 260.000 1337.550 260.030 ;
        RECT 1338.300 58.810 1338.440 260.030 ;
        RECT 1338.240 58.490 1338.500 58.810 ;
        RECT 1642.300 58.490 1642.560 58.810 ;
        RECT 1642.360 16.730 1642.500 58.490 ;
        RECT 1642.360 16.590 1644.340 16.730 ;
        RECT 1644.200 2.400 1644.340 16.590 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1355.230 243.680 1355.550 243.740 ;
        RECT 1362.590 243.680 1362.910 243.740 ;
        RECT 1355.230 243.540 1362.910 243.680 ;
        RECT 1355.230 243.480 1355.550 243.540 ;
        RECT 1362.590 243.480 1362.910 243.540 ;
        RECT 1362.590 66.200 1362.910 66.260 ;
        RECT 1656.070 66.200 1656.390 66.260 ;
        RECT 1362.590 66.060 1656.390 66.200 ;
        RECT 1362.590 66.000 1362.910 66.060 ;
        RECT 1656.070 66.000 1656.390 66.060 ;
        RECT 1656.070 17.580 1656.390 17.640 ;
        RECT 1662.050 17.580 1662.370 17.640 ;
        RECT 1656.070 17.440 1662.370 17.580 ;
        RECT 1656.070 17.380 1656.390 17.440 ;
        RECT 1662.050 17.380 1662.370 17.440 ;
      LAYER via ;
        RECT 1355.260 243.480 1355.520 243.740 ;
        RECT 1362.620 243.480 1362.880 243.740 ;
        RECT 1362.620 66.000 1362.880 66.260 ;
        RECT 1656.100 66.000 1656.360 66.260 ;
        RECT 1656.100 17.380 1656.360 17.640 ;
        RECT 1662.080 17.380 1662.340 17.640 ;
      LAYER met2 ;
        RECT 1355.210 260.000 1355.490 264.000 ;
        RECT 1355.320 243.770 1355.460 260.000 ;
        RECT 1355.260 243.450 1355.520 243.770 ;
        RECT 1362.620 243.450 1362.880 243.770 ;
        RECT 1362.680 66.290 1362.820 243.450 ;
        RECT 1362.620 65.970 1362.880 66.290 ;
        RECT 1656.100 65.970 1656.360 66.290 ;
        RECT 1656.160 17.670 1656.300 65.970 ;
        RECT 1656.100 17.350 1656.360 17.670 ;
        RECT 1662.080 17.350 1662.340 17.670 ;
        RECT 1662.140 2.400 1662.280 17.350 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1373.170 244.020 1373.490 244.080 ;
        RECT 1383.290 244.020 1383.610 244.080 ;
        RECT 1373.170 243.880 1383.610 244.020 ;
        RECT 1373.170 243.820 1373.490 243.880 ;
        RECT 1383.290 243.820 1383.610 243.880 ;
        RECT 1383.290 73.000 1383.610 73.060 ;
        RECT 1676.770 73.000 1677.090 73.060 ;
        RECT 1383.290 72.860 1677.090 73.000 ;
        RECT 1383.290 72.800 1383.610 72.860 ;
        RECT 1676.770 72.800 1677.090 72.860 ;
      LAYER via ;
        RECT 1373.200 243.820 1373.460 244.080 ;
        RECT 1383.320 243.820 1383.580 244.080 ;
        RECT 1383.320 72.800 1383.580 73.060 ;
        RECT 1676.800 72.800 1677.060 73.060 ;
      LAYER met2 ;
        RECT 1373.150 260.000 1373.430 264.000 ;
        RECT 1373.260 244.110 1373.400 260.000 ;
        RECT 1373.200 243.790 1373.460 244.110 ;
        RECT 1383.320 243.790 1383.580 244.110 ;
        RECT 1383.380 73.090 1383.520 243.790 ;
        RECT 1383.320 72.770 1383.580 73.090 ;
        RECT 1676.800 72.770 1677.060 73.090 ;
        RECT 1676.860 16.730 1677.000 72.770 ;
        RECT 1676.860 16.590 1679.760 16.730 ;
        RECT 1679.620 2.400 1679.760 16.590 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1391.110 243.340 1391.430 243.400 ;
        RECT 1403.990 243.340 1404.310 243.400 ;
        RECT 1391.110 243.200 1404.310 243.340 ;
        RECT 1391.110 243.140 1391.430 243.200 ;
        RECT 1403.990 243.140 1404.310 243.200 ;
        RECT 1403.990 142.020 1404.310 142.080 ;
        RECT 1697.470 142.020 1697.790 142.080 ;
        RECT 1403.990 141.880 1697.790 142.020 ;
        RECT 1403.990 141.820 1404.310 141.880 ;
        RECT 1697.470 141.820 1697.790 141.880 ;
      LAYER via ;
        RECT 1391.140 243.140 1391.400 243.400 ;
        RECT 1404.020 243.140 1404.280 243.400 ;
        RECT 1404.020 141.820 1404.280 142.080 ;
        RECT 1697.500 141.820 1697.760 142.080 ;
      LAYER met2 ;
        RECT 1391.090 260.000 1391.370 264.000 ;
        RECT 1391.200 243.430 1391.340 260.000 ;
        RECT 1391.140 243.110 1391.400 243.430 ;
        RECT 1404.020 243.110 1404.280 243.430 ;
        RECT 1404.080 142.110 1404.220 243.110 ;
        RECT 1404.020 141.790 1404.280 142.110 ;
        RECT 1697.500 141.790 1697.760 142.110 ;
        RECT 1697.560 2.400 1697.700 141.790 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 19.620 427.730 19.680 ;
        RECT 734.230 19.620 734.550 19.680 ;
        RECT 427.410 19.480 734.550 19.620 ;
        RECT 427.410 19.420 427.730 19.480 ;
        RECT 734.230 19.420 734.550 19.480 ;
      LAYER via ;
        RECT 427.440 19.420 427.700 19.680 ;
        RECT 734.260 19.420 734.520 19.680 ;
      LAYER met2 ;
        RECT 426.010 260.170 426.290 264.000 ;
        RECT 426.010 260.030 427.640 260.170 ;
        RECT 426.010 260.000 426.290 260.030 ;
        RECT 427.500 19.710 427.640 260.030 ;
        RECT 427.440 19.390 427.700 19.710 ;
        RECT 734.260 19.390 734.520 19.710 ;
        RECT 734.320 2.400 734.460 19.390 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.050 246.060 1409.370 246.120 ;
        RECT 1541.990 246.060 1542.310 246.120 ;
        RECT 1409.050 245.920 1542.310 246.060 ;
        RECT 1409.050 245.860 1409.370 245.920 ;
        RECT 1541.990 245.860 1542.310 245.920 ;
        RECT 1541.990 24.380 1542.310 24.440 ;
        RECT 1715.410 24.380 1715.730 24.440 ;
        RECT 1541.990 24.240 1715.730 24.380 ;
        RECT 1541.990 24.180 1542.310 24.240 ;
        RECT 1715.410 24.180 1715.730 24.240 ;
      LAYER via ;
        RECT 1409.080 245.860 1409.340 246.120 ;
        RECT 1542.020 245.860 1542.280 246.120 ;
        RECT 1542.020 24.180 1542.280 24.440 ;
        RECT 1715.440 24.180 1715.700 24.440 ;
      LAYER met2 ;
        RECT 1409.030 260.000 1409.310 264.000 ;
        RECT 1409.140 246.150 1409.280 260.000 ;
        RECT 1409.080 245.830 1409.340 246.150 ;
        RECT 1542.020 245.830 1542.280 246.150 ;
        RECT 1542.080 24.470 1542.220 245.830 ;
        RECT 1542.020 24.150 1542.280 24.470 ;
        RECT 1715.440 24.150 1715.700 24.470 ;
        RECT 1715.500 2.400 1715.640 24.150 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.910 79.460 1428.230 79.520 ;
        RECT 1731.970 79.460 1732.290 79.520 ;
        RECT 1427.910 79.320 1732.290 79.460 ;
        RECT 1427.910 79.260 1428.230 79.320 ;
        RECT 1731.970 79.260 1732.290 79.320 ;
      LAYER via ;
        RECT 1427.940 79.260 1428.200 79.520 ;
        RECT 1732.000 79.260 1732.260 79.520 ;
      LAYER met2 ;
        RECT 1426.970 260.170 1427.250 264.000 ;
        RECT 1426.970 260.030 1428.140 260.170 ;
        RECT 1426.970 260.000 1427.250 260.030 ;
        RECT 1428.000 79.550 1428.140 260.030 ;
        RECT 1427.940 79.230 1428.200 79.550 ;
        RECT 1732.000 79.230 1732.260 79.550 ;
        RECT 1732.060 17.410 1732.200 79.230 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.930 243.680 1445.250 243.740 ;
        RECT 1452.290 243.680 1452.610 243.740 ;
        RECT 1444.930 243.540 1452.610 243.680 ;
        RECT 1444.930 243.480 1445.250 243.540 ;
        RECT 1452.290 243.480 1452.610 243.540 ;
        RECT 1452.290 86.600 1452.610 86.660 ;
        RECT 1745.770 86.600 1746.090 86.660 ;
        RECT 1452.290 86.460 1746.090 86.600 ;
        RECT 1452.290 86.400 1452.610 86.460 ;
        RECT 1745.770 86.400 1746.090 86.460 ;
      LAYER via ;
        RECT 1444.960 243.480 1445.220 243.740 ;
        RECT 1452.320 243.480 1452.580 243.740 ;
        RECT 1452.320 86.400 1452.580 86.660 ;
        RECT 1745.800 86.400 1746.060 86.660 ;
      LAYER met2 ;
        RECT 1444.910 260.000 1445.190 264.000 ;
        RECT 1445.020 243.770 1445.160 260.000 ;
        RECT 1444.960 243.450 1445.220 243.770 ;
        RECT 1452.320 243.450 1452.580 243.770 ;
        RECT 1452.380 86.690 1452.520 243.450 ;
        RECT 1452.320 86.370 1452.580 86.690 ;
        RECT 1745.800 86.370 1746.060 86.690 ;
        RECT 1745.860 17.410 1746.000 86.370 ;
        RECT 1745.860 17.270 1751.520 17.410 ;
        RECT 1751.380 2.400 1751.520 17.270 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.870 243.340 1463.190 243.400 ;
        RECT 1469.310 243.340 1469.630 243.400 ;
        RECT 1462.870 243.200 1469.630 243.340 ;
        RECT 1462.870 243.140 1463.190 243.200 ;
        RECT 1469.310 243.140 1469.630 243.200 ;
        RECT 1469.310 38.660 1469.630 38.720 ;
        RECT 1768.770 38.660 1769.090 38.720 ;
        RECT 1469.310 38.520 1769.090 38.660 ;
        RECT 1469.310 38.460 1469.630 38.520 ;
        RECT 1768.770 38.460 1769.090 38.520 ;
      LAYER via ;
        RECT 1462.900 243.140 1463.160 243.400 ;
        RECT 1469.340 243.140 1469.600 243.400 ;
        RECT 1469.340 38.460 1469.600 38.720 ;
        RECT 1768.800 38.460 1769.060 38.720 ;
      LAYER met2 ;
        RECT 1462.850 260.000 1463.130 264.000 ;
        RECT 1462.960 243.430 1463.100 260.000 ;
        RECT 1462.900 243.110 1463.160 243.430 ;
        RECT 1469.340 243.110 1469.600 243.430 ;
        RECT 1469.400 38.750 1469.540 243.110 ;
        RECT 1469.340 38.430 1469.600 38.750 ;
        RECT 1768.800 38.430 1769.060 38.750 ;
        RECT 1768.860 2.400 1769.000 38.430 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1480.350 245.380 1480.670 245.440 ;
        RECT 1666.190 245.380 1666.510 245.440 ;
        RECT 1480.350 245.240 1666.510 245.380 ;
        RECT 1480.350 245.180 1480.670 245.240 ;
        RECT 1666.190 245.180 1666.510 245.240 ;
        RECT 1666.190 24.040 1666.510 24.100 ;
        RECT 1786.250 24.040 1786.570 24.100 ;
        RECT 1666.190 23.900 1786.570 24.040 ;
        RECT 1666.190 23.840 1666.510 23.900 ;
        RECT 1786.250 23.840 1786.570 23.900 ;
      LAYER via ;
        RECT 1480.380 245.180 1480.640 245.440 ;
        RECT 1666.220 245.180 1666.480 245.440 ;
        RECT 1666.220 23.840 1666.480 24.100 ;
        RECT 1786.280 23.840 1786.540 24.100 ;
      LAYER met2 ;
        RECT 1480.330 260.000 1480.610 264.000 ;
        RECT 1480.440 245.470 1480.580 260.000 ;
        RECT 1480.380 245.150 1480.640 245.470 ;
        RECT 1666.220 245.150 1666.480 245.470 ;
        RECT 1666.280 24.130 1666.420 245.150 ;
        RECT 1666.220 23.810 1666.480 24.130 ;
        RECT 1786.280 23.810 1786.540 24.130 ;
        RECT 1786.340 19.450 1786.480 23.810 ;
        RECT 1786.340 19.310 1786.940 19.450 ;
        RECT 1786.800 2.400 1786.940 19.310 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1498.290 244.020 1498.610 244.080 ;
        RECT 1507.490 244.020 1507.810 244.080 ;
        RECT 1498.290 243.880 1507.810 244.020 ;
        RECT 1498.290 243.820 1498.610 243.880 ;
        RECT 1507.490 243.820 1507.810 243.880 ;
        RECT 1507.490 31.520 1507.810 31.580 ;
        RECT 1804.650 31.520 1804.970 31.580 ;
        RECT 1507.490 31.380 1804.970 31.520 ;
        RECT 1507.490 31.320 1507.810 31.380 ;
        RECT 1804.650 31.320 1804.970 31.380 ;
      LAYER via ;
        RECT 1498.320 243.820 1498.580 244.080 ;
        RECT 1507.520 243.820 1507.780 244.080 ;
        RECT 1507.520 31.320 1507.780 31.580 ;
        RECT 1804.680 31.320 1804.940 31.580 ;
      LAYER met2 ;
        RECT 1498.270 260.000 1498.550 264.000 ;
        RECT 1498.380 244.110 1498.520 260.000 ;
        RECT 1498.320 243.790 1498.580 244.110 ;
        RECT 1507.520 243.790 1507.780 244.110 ;
        RECT 1507.580 31.610 1507.720 243.790 ;
        RECT 1507.520 31.290 1507.780 31.610 ;
        RECT 1804.680 31.290 1804.940 31.610 ;
        RECT 1804.740 2.400 1804.880 31.290 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.610 93.060 1517.930 93.120 ;
        RECT 1821.670 93.060 1821.990 93.120 ;
        RECT 1517.610 92.920 1821.990 93.060 ;
        RECT 1517.610 92.860 1517.930 92.920 ;
        RECT 1821.670 92.860 1821.990 92.920 ;
      LAYER via ;
        RECT 1517.640 92.860 1517.900 93.120 ;
        RECT 1821.700 92.860 1821.960 93.120 ;
      LAYER met2 ;
        RECT 1516.210 260.170 1516.490 264.000 ;
        RECT 1516.210 260.030 1517.840 260.170 ;
        RECT 1516.210 260.000 1516.490 260.030 ;
        RECT 1517.700 93.150 1517.840 260.030 ;
        RECT 1517.640 92.830 1517.900 93.150 ;
        RECT 1821.700 92.830 1821.960 93.150 ;
        RECT 1821.760 16.730 1821.900 92.830 ;
        RECT 1821.760 16.590 1822.820 16.730 ;
        RECT 1822.680 2.400 1822.820 16.590 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1534.170 243.680 1534.490 243.740 ;
        RECT 1562.690 243.680 1563.010 243.740 ;
        RECT 1534.170 243.540 1563.010 243.680 ;
        RECT 1534.170 243.480 1534.490 243.540 ;
        RECT 1562.690 243.480 1563.010 243.540 ;
        RECT 1562.690 100.200 1563.010 100.260 ;
        RECT 1835.470 100.200 1835.790 100.260 ;
        RECT 1562.690 100.060 1835.790 100.200 ;
        RECT 1562.690 100.000 1563.010 100.060 ;
        RECT 1835.470 100.000 1835.790 100.060 ;
      LAYER via ;
        RECT 1534.200 243.480 1534.460 243.740 ;
        RECT 1562.720 243.480 1562.980 243.740 ;
        RECT 1562.720 100.000 1562.980 100.260 ;
        RECT 1835.500 100.000 1835.760 100.260 ;
      LAYER met2 ;
        RECT 1534.150 260.000 1534.430 264.000 ;
        RECT 1534.260 243.770 1534.400 260.000 ;
        RECT 1534.200 243.450 1534.460 243.770 ;
        RECT 1562.720 243.450 1562.980 243.770 ;
        RECT 1562.780 100.290 1562.920 243.450 ;
        RECT 1562.720 99.970 1562.980 100.290 ;
        RECT 1835.500 99.970 1835.760 100.290 ;
        RECT 1835.560 16.730 1835.700 99.970 ;
        RECT 1835.560 16.590 1840.300 16.730 ;
        RECT 1840.160 2.400 1840.300 16.590 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1552.110 44.780 1552.430 44.840 ;
        RECT 1858.010 44.780 1858.330 44.840 ;
        RECT 1552.110 44.640 1858.330 44.780 ;
        RECT 1552.110 44.580 1552.430 44.640 ;
        RECT 1858.010 44.580 1858.330 44.640 ;
      LAYER via ;
        RECT 1552.140 44.580 1552.400 44.840 ;
        RECT 1858.040 44.580 1858.300 44.840 ;
      LAYER met2 ;
        RECT 1552.090 260.000 1552.370 264.000 ;
        RECT 1552.200 44.870 1552.340 260.000 ;
        RECT 1552.140 44.550 1552.400 44.870 ;
        RECT 1858.040 44.550 1858.300 44.870 ;
        RECT 1858.100 2.400 1858.240 44.550 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 17.240 1573.130 17.300 ;
        RECT 1572.810 17.100 1573.500 17.240 ;
        RECT 1572.810 17.040 1573.130 17.100 ;
        RECT 1573.360 16.560 1573.500 17.100 ;
        RECT 1875.950 16.560 1876.270 16.620 ;
        RECT 1573.360 16.420 1876.270 16.560 ;
        RECT 1875.950 16.360 1876.270 16.420 ;
      LAYER via ;
        RECT 1572.840 17.040 1573.100 17.300 ;
        RECT 1875.980 16.360 1876.240 16.620 ;
      LAYER met2 ;
        RECT 1570.030 260.170 1570.310 264.000 ;
        RECT 1570.030 260.030 1573.040 260.170 ;
        RECT 1570.030 260.000 1570.310 260.030 ;
        RECT 1572.900 17.330 1573.040 260.030 ;
        RECT 1572.840 17.010 1573.100 17.330 ;
        RECT 1875.980 16.330 1876.240 16.650 ;
        RECT 1876.040 2.400 1876.180 16.330 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 443.510 246.060 443.830 246.120 ;
        RECT 753.090 246.060 753.410 246.120 ;
        RECT 443.510 245.920 753.410 246.060 ;
        RECT 443.510 245.860 443.830 245.920 ;
        RECT 753.090 245.860 753.410 245.920 ;
      LAYER via ;
        RECT 443.540 245.860 443.800 246.120 ;
        RECT 753.120 245.860 753.380 246.120 ;
      LAYER met2 ;
        RECT 443.490 260.000 443.770 264.000 ;
        RECT 443.600 246.150 443.740 260.000 ;
        RECT 443.540 245.830 443.800 246.150 ;
        RECT 753.120 245.830 753.380 246.150 ;
        RECT 753.180 17.410 753.320 245.830 ;
        RECT 752.260 17.270 753.320 17.410 ;
        RECT 752.260 2.400 752.400 17.270 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.990 241.640 1588.310 241.700 ;
        RECT 1593.510 241.640 1593.830 241.700 ;
        RECT 1587.990 241.500 1593.830 241.640 ;
        RECT 1587.990 241.440 1588.310 241.500 ;
        RECT 1593.510 241.440 1593.830 241.500 ;
        RECT 1893.890 17.920 1894.210 17.980 ;
        RECT 1614.760 17.780 1894.210 17.920 ;
        RECT 1593.510 17.580 1593.830 17.640 ;
        RECT 1614.760 17.580 1614.900 17.780 ;
        RECT 1893.890 17.720 1894.210 17.780 ;
        RECT 1593.510 17.440 1614.900 17.580 ;
        RECT 1593.510 17.380 1593.830 17.440 ;
      LAYER via ;
        RECT 1588.020 241.440 1588.280 241.700 ;
        RECT 1593.540 241.440 1593.800 241.700 ;
        RECT 1593.540 17.380 1593.800 17.640 ;
        RECT 1893.920 17.720 1894.180 17.980 ;
      LAYER met2 ;
        RECT 1587.970 260.000 1588.250 264.000 ;
        RECT 1588.080 241.730 1588.220 260.000 ;
        RECT 1588.020 241.410 1588.280 241.730 ;
        RECT 1593.540 241.410 1593.800 241.730 ;
        RECT 1593.600 17.670 1593.740 241.410 ;
        RECT 1893.920 17.690 1894.180 18.010 ;
        RECT 1593.540 17.350 1593.800 17.670 ;
        RECT 1893.980 2.400 1894.120 17.690 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1607.310 18.260 1607.630 18.320 ;
        RECT 1911.370 18.260 1911.690 18.320 ;
        RECT 1607.310 18.120 1911.690 18.260 ;
        RECT 1607.310 18.060 1607.630 18.120 ;
        RECT 1911.370 18.060 1911.690 18.120 ;
      LAYER via ;
        RECT 1607.340 18.060 1607.600 18.320 ;
        RECT 1911.400 18.060 1911.660 18.320 ;
      LAYER met2 ;
        RECT 1605.450 260.170 1605.730 264.000 ;
        RECT 1605.450 260.030 1607.540 260.170 ;
        RECT 1605.450 260.000 1605.730 260.030 ;
        RECT 1607.400 18.350 1607.540 260.030 ;
        RECT 1607.340 18.030 1607.600 18.350 ;
        RECT 1911.400 18.030 1911.660 18.350 ;
        RECT 1911.460 17.410 1911.600 18.030 ;
        RECT 1911.460 17.270 1912.060 17.410 ;
        RECT 1911.920 2.400 1912.060 17.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1623.410 244.020 1623.730 244.080 ;
        RECT 1628.010 244.020 1628.330 244.080 ;
        RECT 1623.410 243.880 1628.330 244.020 ;
        RECT 1623.410 243.820 1623.730 243.880 ;
        RECT 1628.010 243.820 1628.330 243.880 ;
        RECT 1628.010 15.880 1628.330 15.940 ;
        RECT 1929.310 15.880 1929.630 15.940 ;
        RECT 1628.010 15.740 1929.630 15.880 ;
        RECT 1628.010 15.680 1628.330 15.740 ;
        RECT 1929.310 15.680 1929.630 15.740 ;
      LAYER via ;
        RECT 1623.440 243.820 1623.700 244.080 ;
        RECT 1628.040 243.820 1628.300 244.080 ;
        RECT 1628.040 15.680 1628.300 15.940 ;
        RECT 1929.340 15.680 1929.600 15.940 ;
      LAYER met2 ;
        RECT 1623.390 260.000 1623.670 264.000 ;
        RECT 1623.500 244.110 1623.640 260.000 ;
        RECT 1623.440 243.790 1623.700 244.110 ;
        RECT 1628.040 243.790 1628.300 244.110 ;
        RECT 1628.100 15.970 1628.240 243.790 ;
        RECT 1628.040 15.650 1628.300 15.970 ;
        RECT 1929.340 15.650 1929.600 15.970 ;
        RECT 1929.400 2.400 1929.540 15.650 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1641.810 18.600 1642.130 18.660 ;
        RECT 1947.250 18.600 1947.570 18.660 ;
        RECT 1641.810 18.460 1947.570 18.600 ;
        RECT 1641.810 18.400 1642.130 18.460 ;
        RECT 1947.250 18.400 1947.570 18.460 ;
      LAYER via ;
        RECT 1641.840 18.400 1642.100 18.660 ;
        RECT 1947.280 18.400 1947.540 18.660 ;
      LAYER met2 ;
        RECT 1641.330 260.170 1641.610 264.000 ;
        RECT 1641.330 260.030 1642.040 260.170 ;
        RECT 1641.330 260.000 1641.610 260.030 ;
        RECT 1641.900 18.690 1642.040 260.030 ;
        RECT 1641.840 18.370 1642.100 18.690 ;
        RECT 1947.280 18.370 1947.540 18.690 ;
        RECT 1947.340 2.400 1947.480 18.370 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.510 19.280 1662.830 19.340 ;
        RECT 1965.190 19.280 1965.510 19.340 ;
        RECT 1662.510 19.140 1965.510 19.280 ;
        RECT 1662.510 19.080 1662.830 19.140 ;
        RECT 1965.190 19.080 1965.510 19.140 ;
      LAYER via ;
        RECT 1662.540 19.080 1662.800 19.340 ;
        RECT 1965.220 19.080 1965.480 19.340 ;
      LAYER met2 ;
        RECT 1659.270 260.170 1659.550 264.000 ;
        RECT 1659.270 260.030 1662.740 260.170 ;
        RECT 1659.270 260.000 1659.550 260.030 ;
        RECT 1662.600 19.370 1662.740 260.030 ;
        RECT 1662.540 19.050 1662.800 19.370 ;
        RECT 1965.220 19.050 1965.480 19.370 ;
        RECT 1965.280 2.400 1965.420 19.050 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1677.230 244.020 1677.550 244.080 ;
        RECT 1683.210 244.020 1683.530 244.080 ;
        RECT 1677.230 243.880 1683.530 244.020 ;
        RECT 1677.230 243.820 1677.550 243.880 ;
        RECT 1683.210 243.820 1683.530 243.880 ;
        RECT 1683.210 20.640 1683.530 20.700 ;
        RECT 1983.130 20.640 1983.450 20.700 ;
        RECT 1683.210 20.500 1983.450 20.640 ;
        RECT 1683.210 20.440 1683.530 20.500 ;
        RECT 1983.130 20.440 1983.450 20.500 ;
      LAYER via ;
        RECT 1677.260 243.820 1677.520 244.080 ;
        RECT 1683.240 243.820 1683.500 244.080 ;
        RECT 1683.240 20.440 1683.500 20.700 ;
        RECT 1983.160 20.440 1983.420 20.700 ;
      LAYER met2 ;
        RECT 1677.210 260.000 1677.490 264.000 ;
        RECT 1677.320 244.110 1677.460 260.000 ;
        RECT 1677.260 243.790 1677.520 244.110 ;
        RECT 1683.240 243.790 1683.500 244.110 ;
        RECT 1683.300 20.730 1683.440 243.790 ;
        RECT 1683.240 20.410 1683.500 20.730 ;
        RECT 1983.160 20.410 1983.420 20.730 ;
        RECT 1983.220 2.400 1983.360 20.410 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1752.285 17.085 1753.375 17.255 ;
      LAYER mcon ;
        RECT 1753.205 17.085 1753.375 17.255 ;
      LAYER met1 ;
        RECT 1697.010 17.240 1697.330 17.300 ;
        RECT 1752.225 17.240 1752.515 17.285 ;
        RECT 1697.010 17.100 1752.515 17.240 ;
        RECT 1697.010 17.040 1697.330 17.100 ;
        RECT 1752.225 17.055 1752.515 17.100 ;
        RECT 1753.145 17.240 1753.435 17.285 ;
        RECT 2001.070 17.240 2001.390 17.300 ;
        RECT 1753.145 17.100 2001.390 17.240 ;
        RECT 1753.145 17.055 1753.435 17.100 ;
        RECT 2001.070 17.040 2001.390 17.100 ;
      LAYER via ;
        RECT 1697.040 17.040 1697.300 17.300 ;
        RECT 2001.100 17.040 2001.360 17.300 ;
      LAYER met2 ;
        RECT 1695.150 260.170 1695.430 264.000 ;
        RECT 1695.150 260.030 1697.240 260.170 ;
        RECT 1695.150 260.000 1695.430 260.030 ;
        RECT 1697.100 17.330 1697.240 260.030 ;
        RECT 1697.040 17.010 1697.300 17.330 ;
        RECT 2001.100 17.010 2001.360 17.330 ;
        RECT 2001.160 2.400 2001.300 17.010 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1713.110 242.660 1713.430 242.720 ;
        RECT 1717.710 242.660 1718.030 242.720 ;
        RECT 1713.110 242.520 1718.030 242.660 ;
        RECT 1713.110 242.460 1713.430 242.520 ;
        RECT 1717.710 242.460 1718.030 242.520 ;
        RECT 1717.710 19.960 1718.030 20.020 ;
        RECT 2018.550 19.960 2018.870 20.020 ;
        RECT 1717.710 19.820 2018.870 19.960 ;
        RECT 1717.710 19.760 1718.030 19.820 ;
        RECT 2018.550 19.760 2018.870 19.820 ;
      LAYER via ;
        RECT 1713.140 242.460 1713.400 242.720 ;
        RECT 1717.740 242.460 1718.000 242.720 ;
        RECT 1717.740 19.760 1718.000 20.020 ;
        RECT 2018.580 19.760 2018.840 20.020 ;
      LAYER met2 ;
        RECT 1713.090 260.000 1713.370 264.000 ;
        RECT 1713.200 242.750 1713.340 260.000 ;
        RECT 1713.140 242.430 1713.400 242.750 ;
        RECT 1717.740 242.430 1718.000 242.750 ;
        RECT 1717.800 20.050 1717.940 242.430 ;
        RECT 1717.740 19.730 1718.000 20.050 ;
        RECT 2018.580 19.730 2018.840 20.050 ;
        RECT 2018.640 2.400 2018.780 19.730 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2036.490 17.580 2036.810 17.640 ;
        RECT 1752.760 17.440 2036.810 17.580 ;
        RECT 1731.510 16.900 1731.830 16.960 ;
        RECT 1752.760 16.900 1752.900 17.440 ;
        RECT 2036.490 17.380 2036.810 17.440 ;
        RECT 1731.510 16.760 1752.900 16.900 ;
        RECT 1731.510 16.700 1731.830 16.760 ;
      LAYER via ;
        RECT 1731.540 16.700 1731.800 16.960 ;
        RECT 2036.520 17.380 2036.780 17.640 ;
      LAYER met2 ;
        RECT 1730.570 260.170 1730.850 264.000 ;
        RECT 1730.570 260.030 1731.740 260.170 ;
        RECT 1730.570 260.000 1730.850 260.030 ;
        RECT 1731.600 16.990 1731.740 260.030 ;
        RECT 2036.520 17.350 2036.780 17.670 ;
        RECT 1731.540 16.670 1731.800 16.990 ;
        RECT 2036.580 2.400 2036.720 17.350 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1752.210 18.940 1752.530 19.000 ;
        RECT 2054.430 18.940 2054.750 19.000 ;
        RECT 1752.210 18.800 2054.750 18.940 ;
        RECT 1752.210 18.740 1752.530 18.800 ;
        RECT 2054.430 18.740 2054.750 18.800 ;
      LAYER via ;
        RECT 1752.240 18.740 1752.500 19.000 ;
        RECT 2054.460 18.740 2054.720 19.000 ;
      LAYER met2 ;
        RECT 1748.510 260.170 1748.790 264.000 ;
        RECT 1748.510 260.030 1752.440 260.170 ;
        RECT 1748.510 260.000 1748.790 260.030 ;
        RECT 1752.300 19.030 1752.440 260.030 ;
        RECT 1752.240 18.710 1752.500 19.030 ;
        RECT 2054.460 18.710 2054.720 19.030 ;
        RECT 2054.520 2.400 2054.660 18.710 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.430 260.170 461.710 264.000 ;
        RECT 461.430 260.030 462.140 260.170 ;
        RECT 461.430 260.000 461.710 260.030 ;
        RECT 462.000 16.845 462.140 260.030 ;
        RECT 461.930 16.475 462.210 16.845 ;
        RECT 769.670 16.475 769.950 16.845 ;
        RECT 769.740 2.400 769.880 16.475 ;
        RECT 769.530 -4.800 770.090 2.400 ;
      LAYER via2 ;
        RECT 461.930 16.520 462.210 16.800 ;
        RECT 769.670 16.520 769.950 16.800 ;
      LAYER met3 ;
        RECT 461.905 16.810 462.235 16.825 ;
        RECT 769.645 16.810 769.975 16.825 ;
        RECT 461.905 16.510 769.975 16.810 ;
        RECT 461.905 16.495 462.235 16.510 ;
        RECT 769.645 16.495 769.975 16.510 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.470 244.020 1766.790 244.080 ;
        RECT 1772.910 244.020 1773.230 244.080 ;
        RECT 1766.470 243.880 1773.230 244.020 ;
        RECT 1766.470 243.820 1766.790 243.880 ;
        RECT 1772.910 243.820 1773.230 243.880 ;
        RECT 1772.910 16.900 1773.230 16.960 ;
        RECT 2072.370 16.900 2072.690 16.960 ;
        RECT 1772.910 16.760 2072.690 16.900 ;
        RECT 1772.910 16.700 1773.230 16.760 ;
        RECT 2072.370 16.700 2072.690 16.760 ;
      LAYER via ;
        RECT 1766.500 243.820 1766.760 244.080 ;
        RECT 1772.940 243.820 1773.200 244.080 ;
        RECT 1772.940 16.700 1773.200 16.960 ;
        RECT 2072.400 16.700 2072.660 16.960 ;
      LAYER met2 ;
        RECT 1766.450 260.000 1766.730 264.000 ;
        RECT 1766.560 244.110 1766.700 260.000 ;
        RECT 1766.500 243.790 1766.760 244.110 ;
        RECT 1772.940 243.790 1773.200 244.110 ;
        RECT 1773.000 16.990 1773.140 243.790 ;
        RECT 1772.940 16.670 1773.200 16.990 ;
        RECT 2072.400 16.670 2072.660 16.990 ;
        RECT 2072.460 2.400 2072.600 16.670 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 20.300 1787.030 20.360 ;
        RECT 2089.850 20.300 2090.170 20.360 ;
        RECT 1786.710 20.160 2090.170 20.300 ;
        RECT 1786.710 20.100 1787.030 20.160 ;
        RECT 2089.850 20.100 2090.170 20.160 ;
      LAYER via ;
        RECT 1786.740 20.100 1787.000 20.360 ;
        RECT 2089.880 20.100 2090.140 20.360 ;
      LAYER met2 ;
        RECT 1784.390 260.170 1784.670 264.000 ;
        RECT 1784.390 260.030 1786.940 260.170 ;
        RECT 1784.390 260.000 1784.670 260.030 ;
        RECT 1786.800 20.390 1786.940 260.030 ;
        RECT 1786.740 20.070 1787.000 20.390 ;
        RECT 2089.880 20.070 2090.140 20.390 ;
        RECT 2089.940 2.400 2090.080 20.070 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1802.350 243.680 1802.670 243.740 ;
        RECT 1807.410 243.680 1807.730 243.740 ;
        RECT 1802.350 243.540 1807.730 243.680 ;
        RECT 1802.350 243.480 1802.670 243.540 ;
        RECT 1807.410 243.480 1807.730 243.540 ;
        RECT 1807.410 19.620 1807.730 19.680 ;
        RECT 2107.790 19.620 2108.110 19.680 ;
        RECT 1807.410 19.480 2108.110 19.620 ;
        RECT 1807.410 19.420 1807.730 19.480 ;
        RECT 2107.790 19.420 2108.110 19.480 ;
      LAYER via ;
        RECT 1802.380 243.480 1802.640 243.740 ;
        RECT 1807.440 243.480 1807.700 243.740 ;
        RECT 1807.440 19.420 1807.700 19.680 ;
        RECT 2107.820 19.420 2108.080 19.680 ;
      LAYER met2 ;
        RECT 1802.330 260.000 1802.610 264.000 ;
        RECT 1802.440 243.770 1802.580 260.000 ;
        RECT 1802.380 243.450 1802.640 243.770 ;
        RECT 1807.440 243.450 1807.700 243.770 ;
        RECT 1807.500 19.710 1807.640 243.450 ;
        RECT 1807.440 19.390 1807.700 19.710 ;
        RECT 2107.820 19.390 2108.080 19.710 ;
        RECT 2107.880 2.400 2108.020 19.390 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1820.270 260.170 1820.550 264.000 ;
        RECT 1820.270 260.030 1821.440 260.170 ;
        RECT 1820.270 260.000 1820.550 260.030 ;
        RECT 1821.300 16.845 1821.440 260.030 ;
        RECT 1821.230 16.475 1821.510 16.845 ;
        RECT 2125.750 16.475 2126.030 16.845 ;
        RECT 2125.820 2.400 2125.960 16.475 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
      LAYER via2 ;
        RECT 1821.230 16.520 1821.510 16.800 ;
        RECT 2125.750 16.520 2126.030 16.800 ;
      LAYER met3 ;
        RECT 1821.205 16.810 1821.535 16.825 ;
        RECT 2125.725 16.810 2126.055 16.825 ;
        RECT 1821.205 16.510 2126.055 16.810 ;
        RECT 1821.205 16.495 1821.535 16.510 ;
        RECT 2125.725 16.495 2126.055 16.510 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2139.605 241.485 2139.775 245.735 ;
        RECT 2139.605 144.925 2139.775 193.035 ;
        RECT 2139.605 48.365 2139.775 96.475 ;
      LAYER mcon ;
        RECT 2139.605 245.565 2139.775 245.735 ;
        RECT 2139.605 192.865 2139.775 193.035 ;
        RECT 2139.605 96.305 2139.775 96.475 ;
      LAYER met1 ;
        RECT 1838.230 245.720 1838.550 245.780 ;
        RECT 2139.545 245.720 2139.835 245.765 ;
        RECT 1838.230 245.580 2139.835 245.720 ;
        RECT 1838.230 245.520 1838.550 245.580 ;
        RECT 2139.545 245.535 2139.835 245.580 ;
        RECT 2139.530 241.640 2139.850 241.700 ;
        RECT 2139.335 241.500 2139.850 241.640 ;
        RECT 2139.530 241.440 2139.850 241.500 ;
        RECT 2139.530 193.020 2139.850 193.080 ;
        RECT 2139.335 192.880 2139.850 193.020 ;
        RECT 2139.530 192.820 2139.850 192.880 ;
        RECT 2139.530 145.080 2139.850 145.140 ;
        RECT 2139.335 144.940 2139.850 145.080 ;
        RECT 2139.530 144.880 2139.850 144.940 ;
        RECT 2139.530 96.460 2139.850 96.520 ;
        RECT 2139.335 96.320 2139.850 96.460 ;
        RECT 2139.530 96.260 2139.850 96.320 ;
        RECT 2139.530 48.520 2139.850 48.580 ;
        RECT 2139.335 48.380 2139.850 48.520 ;
        RECT 2139.530 48.320 2139.850 48.380 ;
        RECT 2139.530 14.180 2139.850 14.240 ;
        RECT 2139.530 14.040 2143.900 14.180 ;
        RECT 2139.530 13.980 2139.850 14.040 ;
        RECT 2143.760 13.900 2143.900 14.040 ;
        RECT 2143.670 13.640 2143.990 13.900 ;
      LAYER via ;
        RECT 1838.260 245.520 1838.520 245.780 ;
        RECT 2139.560 241.440 2139.820 241.700 ;
        RECT 2139.560 192.820 2139.820 193.080 ;
        RECT 2139.560 144.880 2139.820 145.140 ;
        RECT 2139.560 96.260 2139.820 96.520 ;
        RECT 2139.560 48.320 2139.820 48.580 ;
        RECT 2139.560 13.980 2139.820 14.240 ;
        RECT 2143.700 13.640 2143.960 13.900 ;
      LAYER met2 ;
        RECT 1838.210 260.000 1838.490 264.000 ;
        RECT 1838.320 245.810 1838.460 260.000 ;
        RECT 1838.260 245.490 1838.520 245.810 ;
        RECT 2139.560 241.410 2139.820 241.730 ;
        RECT 2139.620 193.110 2139.760 241.410 ;
        RECT 2139.560 192.790 2139.820 193.110 ;
        RECT 2139.560 144.850 2139.820 145.170 ;
        RECT 2139.620 96.550 2139.760 144.850 ;
        RECT 2139.560 96.230 2139.820 96.550 ;
        RECT 2139.560 48.290 2139.820 48.610 ;
        RECT 2139.620 14.270 2139.760 48.290 ;
        RECT 2139.560 13.950 2139.820 14.270 ;
        RECT 2143.700 13.610 2143.960 13.930 ;
        RECT 2143.760 2.400 2143.900 13.610 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1855.690 260.000 1855.970 264.000 ;
        RECT 1855.800 18.205 1855.940 260.000 ;
        RECT 1855.730 17.835 1856.010 18.205 ;
        RECT 2161.630 17.835 2161.910 18.205 ;
        RECT 2161.700 2.400 2161.840 17.835 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 1855.730 17.880 1856.010 18.160 ;
        RECT 2161.630 17.880 2161.910 18.160 ;
      LAYER met3 ;
        RECT 1855.705 18.170 1856.035 18.185 ;
        RECT 2161.605 18.170 2161.935 18.185 ;
        RECT 1855.705 17.870 2161.935 18.170 ;
        RECT 1855.705 17.855 1856.035 17.870 ;
        RECT 2161.605 17.855 2161.935 17.870 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2174.105 241.485 2174.275 245.395 ;
        RECT 2174.105 144.925 2174.275 193.035 ;
        RECT 2174.105 48.365 2174.275 96.475 ;
      LAYER mcon ;
        RECT 2174.105 245.225 2174.275 245.395 ;
        RECT 2174.105 192.865 2174.275 193.035 ;
        RECT 2174.105 96.305 2174.275 96.475 ;
      LAYER met1 ;
        RECT 1873.650 245.380 1873.970 245.440 ;
        RECT 2174.045 245.380 2174.335 245.425 ;
        RECT 1873.650 245.240 2174.335 245.380 ;
        RECT 1873.650 245.180 1873.970 245.240 ;
        RECT 2174.045 245.195 2174.335 245.240 ;
        RECT 2174.030 241.640 2174.350 241.700 ;
        RECT 2173.835 241.500 2174.350 241.640 ;
        RECT 2174.030 241.440 2174.350 241.500 ;
        RECT 2174.030 193.020 2174.350 193.080 ;
        RECT 2173.835 192.880 2174.350 193.020 ;
        RECT 2174.030 192.820 2174.350 192.880 ;
        RECT 2174.030 145.080 2174.350 145.140 ;
        RECT 2173.835 144.940 2174.350 145.080 ;
        RECT 2174.030 144.880 2174.350 144.940 ;
        RECT 2174.030 96.460 2174.350 96.520 ;
        RECT 2173.835 96.320 2174.350 96.460 ;
        RECT 2174.030 96.260 2174.350 96.320 ;
        RECT 2174.030 48.520 2174.350 48.580 ;
        RECT 2173.835 48.380 2174.350 48.520 ;
        RECT 2174.030 48.320 2174.350 48.380 ;
        RECT 2174.030 14.180 2174.350 14.240 ;
        RECT 2174.030 14.040 2179.320 14.180 ;
        RECT 2174.030 13.980 2174.350 14.040 ;
        RECT 2179.180 13.900 2179.320 14.040 ;
        RECT 2179.090 13.640 2179.410 13.900 ;
      LAYER via ;
        RECT 1873.680 245.180 1873.940 245.440 ;
        RECT 2174.060 241.440 2174.320 241.700 ;
        RECT 2174.060 192.820 2174.320 193.080 ;
        RECT 2174.060 144.880 2174.320 145.140 ;
        RECT 2174.060 96.260 2174.320 96.520 ;
        RECT 2174.060 48.320 2174.320 48.580 ;
        RECT 2174.060 13.980 2174.320 14.240 ;
        RECT 2179.120 13.640 2179.380 13.900 ;
      LAYER met2 ;
        RECT 1873.630 260.000 1873.910 264.000 ;
        RECT 1873.740 245.470 1873.880 260.000 ;
        RECT 1873.680 245.150 1873.940 245.470 ;
        RECT 2174.060 241.410 2174.320 241.730 ;
        RECT 2174.120 193.110 2174.260 241.410 ;
        RECT 2174.060 192.790 2174.320 193.110 ;
        RECT 2174.060 144.850 2174.320 145.170 ;
        RECT 2174.120 96.550 2174.260 144.850 ;
        RECT 2174.060 96.230 2174.320 96.550 ;
        RECT 2174.060 48.290 2174.320 48.610 ;
        RECT 2174.120 14.270 2174.260 48.290 ;
        RECT 2174.060 13.950 2174.320 14.270 ;
        RECT 2179.120 13.610 2179.380 13.930 ;
        RECT 2179.180 2.400 2179.320 13.610 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.590 244.020 1891.910 244.080 ;
        RECT 1897.110 244.020 1897.430 244.080 ;
        RECT 1891.590 243.880 1897.430 244.020 ;
        RECT 1891.590 243.820 1891.910 243.880 ;
        RECT 1897.110 243.820 1897.430 243.880 ;
        RECT 1897.110 16.220 1897.430 16.280 ;
        RECT 2197.030 16.220 2197.350 16.280 ;
        RECT 1897.110 16.080 2197.350 16.220 ;
        RECT 1897.110 16.020 1897.430 16.080 ;
        RECT 2197.030 16.020 2197.350 16.080 ;
      LAYER via ;
        RECT 1891.620 243.820 1891.880 244.080 ;
        RECT 1897.140 243.820 1897.400 244.080 ;
        RECT 1897.140 16.020 1897.400 16.280 ;
        RECT 2197.060 16.020 2197.320 16.280 ;
      LAYER met2 ;
        RECT 1891.570 260.000 1891.850 264.000 ;
        RECT 1891.680 244.110 1891.820 260.000 ;
        RECT 1891.620 243.790 1891.880 244.110 ;
        RECT 1897.140 243.790 1897.400 244.110 ;
        RECT 1897.200 16.310 1897.340 243.790 ;
        RECT 1897.140 15.990 1897.400 16.310 ;
        RECT 2197.060 15.990 2197.320 16.310 ;
        RECT 2197.120 2.400 2197.260 15.990 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1910.910 17.920 1911.230 17.980 ;
        RECT 2214.970 17.920 2215.290 17.980 ;
        RECT 1910.910 17.780 2215.290 17.920 ;
        RECT 1910.910 17.720 1911.230 17.780 ;
        RECT 2214.970 17.720 2215.290 17.780 ;
      LAYER via ;
        RECT 1910.940 17.720 1911.200 17.980 ;
        RECT 2215.000 17.720 2215.260 17.980 ;
      LAYER met2 ;
        RECT 1909.510 260.170 1909.790 264.000 ;
        RECT 1909.510 260.030 1911.140 260.170 ;
        RECT 1909.510 260.000 1909.790 260.030 ;
        RECT 1911.000 18.010 1911.140 260.030 ;
        RECT 1910.940 17.690 1911.200 18.010 ;
        RECT 2215.000 17.690 2215.260 18.010 ;
        RECT 2215.060 2.400 2215.200 17.690 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1927.470 244.020 1927.790 244.080 ;
        RECT 1931.610 244.020 1931.930 244.080 ;
        RECT 1927.470 243.880 1931.930 244.020 ;
        RECT 1927.470 243.820 1927.790 243.880 ;
        RECT 1931.610 243.820 1931.930 243.880 ;
        RECT 1931.610 16.560 1931.930 16.620 ;
        RECT 2232.910 16.560 2233.230 16.620 ;
        RECT 1931.610 16.420 2233.230 16.560 ;
        RECT 1931.610 16.360 1931.930 16.420 ;
        RECT 2232.910 16.360 2233.230 16.420 ;
      LAYER via ;
        RECT 1927.500 243.820 1927.760 244.080 ;
        RECT 1931.640 243.820 1931.900 244.080 ;
        RECT 1931.640 16.360 1931.900 16.620 ;
        RECT 2232.940 16.360 2233.200 16.620 ;
      LAYER met2 ;
        RECT 1927.450 260.000 1927.730 264.000 ;
        RECT 1927.560 244.110 1927.700 260.000 ;
        RECT 1927.500 243.790 1927.760 244.110 ;
        RECT 1931.640 243.790 1931.900 244.110 ;
        RECT 1931.700 16.650 1931.840 243.790 ;
        RECT 1931.640 16.330 1931.900 16.650 ;
        RECT 2232.940 16.330 2233.200 16.650 ;
        RECT 2233.000 2.400 2233.140 16.330 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 479.390 245.720 479.710 245.780 ;
        RECT 787.130 245.720 787.450 245.780 ;
        RECT 479.390 245.580 787.450 245.720 ;
        RECT 479.390 245.520 479.710 245.580 ;
        RECT 787.130 245.520 787.450 245.580 ;
      LAYER via ;
        RECT 479.420 245.520 479.680 245.780 ;
        RECT 787.160 245.520 787.420 245.780 ;
      LAYER met2 ;
        RECT 479.370 260.000 479.650 264.000 ;
        RECT 479.480 245.810 479.620 260.000 ;
        RECT 479.420 245.490 479.680 245.810 ;
        RECT 787.160 245.490 787.420 245.810 ;
        RECT 787.220 7.890 787.360 245.490 ;
        RECT 787.220 7.750 787.820 7.890 ;
        RECT 787.680 2.400 787.820 7.750 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1945.410 245.040 1945.730 245.100 ;
        RECT 2249.470 245.040 2249.790 245.100 ;
        RECT 1945.410 244.900 2249.790 245.040 ;
        RECT 1945.410 244.840 1945.730 244.900 ;
        RECT 2249.470 244.840 2249.790 244.900 ;
      LAYER via ;
        RECT 1945.440 244.840 1945.700 245.100 ;
        RECT 2249.500 244.840 2249.760 245.100 ;
      LAYER met2 ;
        RECT 1945.390 260.000 1945.670 264.000 ;
        RECT 1945.500 245.130 1945.640 260.000 ;
        RECT 1945.440 244.810 1945.700 245.130 ;
        RECT 2249.500 244.810 2249.760 245.130 ;
        RECT 2249.560 16.730 2249.700 244.810 ;
        RECT 2249.560 16.590 2251.080 16.730 ;
        RECT 2250.940 2.400 2251.080 16.590 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 19.280 1966.430 19.340 ;
        RECT 2268.330 19.280 2268.650 19.340 ;
        RECT 1966.110 19.140 2268.650 19.280 ;
        RECT 1966.110 19.080 1966.430 19.140 ;
        RECT 2268.330 19.080 2268.650 19.140 ;
      LAYER via ;
        RECT 1966.140 19.080 1966.400 19.340 ;
        RECT 2268.360 19.080 2268.620 19.340 ;
      LAYER met2 ;
        RECT 1963.330 260.170 1963.610 264.000 ;
        RECT 1963.330 260.030 1966.340 260.170 ;
        RECT 1963.330 260.000 1963.610 260.030 ;
        RECT 1966.200 19.370 1966.340 260.030 ;
        RECT 1966.140 19.050 1966.400 19.370 ;
        RECT 2268.360 19.050 2268.620 19.370 ;
        RECT 2268.420 2.400 2268.560 19.050 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1980.830 246.400 1981.150 246.460 ;
        RECT 2284.430 246.400 2284.750 246.460 ;
        RECT 1980.830 246.260 2284.750 246.400 ;
        RECT 1980.830 246.200 1981.150 246.260 ;
        RECT 2284.430 246.200 2284.750 246.260 ;
      LAYER via ;
        RECT 1980.860 246.200 1981.120 246.460 ;
        RECT 2284.460 246.200 2284.720 246.460 ;
      LAYER met2 ;
        RECT 1980.810 260.000 1981.090 264.000 ;
        RECT 1980.920 246.490 1981.060 260.000 ;
        RECT 1980.860 246.170 1981.120 246.490 ;
        RECT 2284.460 246.170 2284.720 246.490 ;
        RECT 2284.520 3.130 2284.660 246.170 ;
        RECT 2284.520 2.990 2286.040 3.130 ;
        RECT 2285.900 2.960 2286.040 2.990 ;
        RECT 2285.900 2.820 2286.500 2.960 ;
        RECT 2286.360 2.400 2286.500 2.820 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2000.610 18.600 2000.930 18.660 ;
        RECT 2304.210 18.600 2304.530 18.660 ;
        RECT 2000.610 18.460 2304.530 18.600 ;
        RECT 2000.610 18.400 2000.930 18.460 ;
        RECT 2304.210 18.400 2304.530 18.460 ;
      LAYER via ;
        RECT 2000.640 18.400 2000.900 18.660 ;
        RECT 2304.240 18.400 2304.500 18.660 ;
      LAYER met2 ;
        RECT 1998.750 260.170 1999.030 264.000 ;
        RECT 1998.750 260.030 2000.840 260.170 ;
        RECT 1998.750 260.000 1999.030 260.030 ;
        RECT 2000.700 18.690 2000.840 260.030 ;
        RECT 2000.640 18.370 2000.900 18.690 ;
        RECT 2304.240 18.370 2304.500 18.690 ;
        RECT 2304.300 2.400 2304.440 18.370 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2016.710 246.060 2017.030 246.120 ;
        RECT 2318.930 246.060 2319.250 246.120 ;
        RECT 2016.710 245.920 2319.250 246.060 ;
        RECT 2016.710 245.860 2017.030 245.920 ;
        RECT 2318.930 245.860 2319.250 245.920 ;
        RECT 2318.930 2.960 2319.250 3.020 ;
        RECT 2322.150 2.960 2322.470 3.020 ;
        RECT 2318.930 2.820 2322.470 2.960 ;
        RECT 2318.930 2.760 2319.250 2.820 ;
        RECT 2322.150 2.760 2322.470 2.820 ;
      LAYER via ;
        RECT 2016.740 245.860 2017.000 246.120 ;
        RECT 2318.960 245.860 2319.220 246.120 ;
        RECT 2318.960 2.760 2319.220 3.020 ;
        RECT 2322.180 2.760 2322.440 3.020 ;
      LAYER met2 ;
        RECT 2016.690 260.000 2016.970 264.000 ;
        RECT 2016.800 246.150 2016.940 260.000 ;
        RECT 2016.740 245.830 2017.000 246.150 ;
        RECT 2318.960 245.830 2319.220 246.150 ;
        RECT 2319.020 3.050 2319.160 245.830 ;
        RECT 2318.960 2.730 2319.220 3.050 ;
        RECT 2322.180 2.730 2322.440 3.050 ;
        RECT 2322.240 2.400 2322.380 2.730 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2034.630 260.170 2034.910 264.000 ;
        RECT 2034.630 260.030 2035.340 260.170 ;
        RECT 2034.630 260.000 2034.910 260.030 ;
        RECT 2035.200 17.525 2035.340 260.030 ;
        RECT 2035.130 17.155 2035.410 17.525 ;
        RECT 2339.650 17.155 2339.930 17.525 ;
        RECT 2339.720 2.400 2339.860 17.155 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
      LAYER via2 ;
        RECT 2035.130 17.200 2035.410 17.480 ;
        RECT 2339.650 17.200 2339.930 17.480 ;
      LAYER met3 ;
        RECT 2035.105 17.490 2035.435 17.505 ;
        RECT 2339.625 17.490 2339.955 17.505 ;
        RECT 2035.105 17.190 2339.955 17.490 ;
        RECT 2035.105 17.175 2035.435 17.190 ;
        RECT 2339.625 17.175 2339.955 17.190 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 18.940 2056.130 19.000 ;
        RECT 2357.570 18.940 2357.890 19.000 ;
        RECT 2055.810 18.800 2357.890 18.940 ;
        RECT 2055.810 18.740 2056.130 18.800 ;
        RECT 2357.570 18.740 2357.890 18.800 ;
      LAYER via ;
        RECT 2055.840 18.740 2056.100 19.000 ;
        RECT 2357.600 18.740 2357.860 19.000 ;
      LAYER met2 ;
        RECT 2052.570 260.170 2052.850 264.000 ;
        RECT 2052.570 260.030 2056.040 260.170 ;
        RECT 2052.570 260.000 2052.850 260.030 ;
        RECT 2055.900 19.030 2056.040 260.030 ;
        RECT 2055.840 18.710 2056.100 19.030 ;
        RECT 2357.600 18.710 2357.860 19.030 ;
        RECT 2357.660 2.400 2357.800 18.710 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2070.530 244.020 2070.850 244.080 ;
        RECT 2076.510 244.020 2076.830 244.080 ;
        RECT 2070.530 243.880 2076.830 244.020 ;
        RECT 2070.530 243.820 2070.850 243.880 ;
        RECT 2076.510 243.820 2076.830 243.880 ;
        RECT 2076.510 17.580 2076.830 17.640 ;
        RECT 2375.510 17.580 2375.830 17.640 ;
        RECT 2076.510 17.440 2375.830 17.580 ;
        RECT 2076.510 17.380 2076.830 17.440 ;
        RECT 2375.510 17.380 2375.830 17.440 ;
      LAYER via ;
        RECT 2070.560 243.820 2070.820 244.080 ;
        RECT 2076.540 243.820 2076.800 244.080 ;
        RECT 2076.540 17.380 2076.800 17.640 ;
        RECT 2375.540 17.380 2375.800 17.640 ;
      LAYER met2 ;
        RECT 2070.510 260.000 2070.790 264.000 ;
        RECT 2070.620 244.110 2070.760 260.000 ;
        RECT 2070.560 243.790 2070.820 244.110 ;
        RECT 2076.540 243.790 2076.800 244.110 ;
        RECT 2076.600 17.670 2076.740 243.790 ;
        RECT 2076.540 17.350 2076.800 17.670 ;
        RECT 2375.540 17.350 2375.800 17.670 ;
        RECT 2375.600 2.400 2375.740 17.350 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 18.260 2090.630 18.320 ;
        RECT 2393.450 18.260 2393.770 18.320 ;
        RECT 2090.310 18.120 2393.770 18.260 ;
        RECT 2090.310 18.060 2090.630 18.120 ;
        RECT 2393.450 18.060 2393.770 18.120 ;
      LAYER via ;
        RECT 2090.340 18.060 2090.600 18.320 ;
        RECT 2393.480 18.060 2393.740 18.320 ;
      LAYER met2 ;
        RECT 2088.450 260.170 2088.730 264.000 ;
        RECT 2088.450 260.030 2090.540 260.170 ;
        RECT 2088.450 260.000 2088.730 260.030 ;
        RECT 2090.400 18.350 2090.540 260.030 ;
        RECT 2090.340 18.030 2090.600 18.350 ;
        RECT 2393.480 18.030 2393.740 18.350 ;
        RECT 2393.540 2.400 2393.680 18.030 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2105.950 244.020 2106.270 244.080 ;
        RECT 2111.010 244.020 2111.330 244.080 ;
        RECT 2105.950 243.880 2111.330 244.020 ;
        RECT 2105.950 243.820 2106.270 243.880 ;
        RECT 2111.010 243.820 2111.330 243.880 ;
        RECT 2111.010 17.240 2111.330 17.300 ;
        RECT 2411.390 17.240 2411.710 17.300 ;
        RECT 2111.010 17.100 2411.710 17.240 ;
        RECT 2111.010 17.040 2111.330 17.100 ;
        RECT 2411.390 17.040 2411.710 17.100 ;
      LAYER via ;
        RECT 2105.980 243.820 2106.240 244.080 ;
        RECT 2111.040 243.820 2111.300 244.080 ;
        RECT 2111.040 17.040 2111.300 17.300 ;
        RECT 2411.420 17.040 2411.680 17.300 ;
      LAYER met2 ;
        RECT 2105.930 260.000 2106.210 264.000 ;
        RECT 2106.040 244.110 2106.180 260.000 ;
        RECT 2105.980 243.790 2106.240 244.110 ;
        RECT 2111.040 243.790 2111.300 244.110 ;
        RECT 2111.100 17.330 2111.240 243.790 ;
        RECT 2111.040 17.010 2111.300 17.330 ;
        RECT 2411.420 17.010 2411.680 17.330 ;
        RECT 2411.480 2.400 2411.620 17.010 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 497.330 244.020 497.650 244.080 ;
        RECT 503.310 244.020 503.630 244.080 ;
        RECT 497.330 243.880 503.630 244.020 ;
        RECT 497.330 243.820 497.650 243.880 ;
        RECT 503.310 243.820 503.630 243.880 ;
        RECT 503.310 15.880 503.630 15.940 ;
        RECT 805.530 15.880 805.850 15.940 ;
        RECT 503.310 15.740 805.850 15.880 ;
        RECT 503.310 15.680 503.630 15.740 ;
        RECT 805.530 15.680 805.850 15.740 ;
      LAYER via ;
        RECT 497.360 243.820 497.620 244.080 ;
        RECT 503.340 243.820 503.600 244.080 ;
        RECT 503.340 15.680 503.600 15.940 ;
        RECT 805.560 15.680 805.820 15.940 ;
      LAYER met2 ;
        RECT 497.310 260.000 497.590 264.000 ;
        RECT 497.420 244.110 497.560 260.000 ;
        RECT 497.360 243.790 497.620 244.110 ;
        RECT 503.340 243.790 503.600 244.110 ;
        RECT 503.400 15.970 503.540 243.790 ;
        RECT 503.340 15.650 503.600 15.970 ;
        RECT 805.560 15.650 805.820 15.970 ;
        RECT 805.620 2.400 805.760 15.650 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 310.570 17.240 310.890 17.300 ;
        RECT 2.830 17.100 310.890 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 310.570 17.040 310.890 17.100 ;
      LAYER via ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 310.600 17.040 310.860 17.300 ;
      LAYER met2 ;
        RECT 312.850 260.170 313.130 264.000 ;
        RECT 310.660 260.030 313.130 260.170 ;
        RECT 310.660 17.330 310.800 260.030 ;
        RECT 312.850 260.000 313.130 260.030 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 310.600 17.010 310.860 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 317.470 17.580 317.790 17.640 ;
        RECT 8.350 17.440 317.790 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 317.470 17.380 317.790 17.440 ;
      LAYER via ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 317.500 17.380 317.760 17.640 ;
      LAYER met2 ;
        RECT 318.370 260.170 318.650 264.000 ;
        RECT 317.560 260.030 318.650 260.170 ;
        RECT 317.560 17.670 317.700 260.030 ;
        RECT 318.370 260.000 318.650 260.030 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 317.500 17.350 317.760 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 3260.000 367.020 3528.900 ;
        RECT 544.020 3260.000 547.020 3528.900 ;
        RECT 724.020 3260.000 727.020 3528.900 ;
        RECT 904.020 3260.000 907.020 3528.900 ;
        RECT 1084.020 3260.000 1087.020 3528.900 ;
        RECT 1264.020 3260.000 1267.020 3528.900 ;
        RECT 1444.020 3260.000 1447.020 3528.900 ;
        RECT 1624.020 3260.000 1627.020 3528.900 ;
        RECT 1804.020 3260.000 1807.020 3528.900 ;
        RECT 1984.020 3260.000 1987.020 3528.900 ;
        RECT 2164.020 3260.000 2167.020 3528.900 ;
        RECT 2344.020 3260.000 2347.020 3528.900 ;
        RECT 2524.020 3260.000 2527.020 3528.900 ;
        RECT 364.020 -9.220 367.020 260.000 ;
        RECT 544.020 -9.220 547.020 260.000 ;
        RECT 724.020 -9.220 727.020 260.000 ;
        RECT 904.020 -9.220 907.020 260.000 ;
        RECT 1084.020 -9.220 1087.020 260.000 ;
        RECT 1264.020 -9.220 1267.020 260.000 ;
        RECT 1444.020 -9.220 1447.020 260.000 ;
        RECT 1624.020 -9.220 1627.020 260.000 ;
        RECT 1804.020 -9.220 1807.020 260.000 ;
        RECT 1984.020 -9.220 1987.020 260.000 ;
        RECT 2164.020 -9.220 2167.020 260.000 ;
        RECT 2344.020 -9.220 2347.020 260.000 ;
        RECT 2524.020 -9.220 2527.020 260.000 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 3260.000 457.020 3528.900 ;
        RECT 634.020 3260.000 637.020 3528.900 ;
        RECT 814.020 3260.000 817.020 3528.900 ;
        RECT 994.020 3260.000 997.020 3528.900 ;
        RECT 1174.020 3260.000 1177.020 3528.900 ;
        RECT 1354.020 3260.000 1357.020 3528.900 ;
        RECT 1534.020 3260.000 1537.020 3528.900 ;
        RECT 1714.020 3260.000 1717.020 3528.900 ;
        RECT 1894.020 3260.000 1897.020 3528.900 ;
        RECT 2074.020 3260.000 2077.020 3528.900 ;
        RECT 2254.020 3260.000 2257.020 3528.900 ;
        RECT 2434.020 3260.000 2437.020 3528.900 ;
        RECT 454.020 -9.220 457.020 260.000 ;
        RECT 634.020 -9.220 637.020 260.000 ;
        RECT 814.020 -9.220 817.020 260.000 ;
        RECT 994.020 -9.220 997.020 260.000 ;
        RECT 1174.020 -9.220 1177.020 260.000 ;
        RECT 1354.020 -9.220 1357.020 260.000 ;
        RECT 1534.020 -9.220 1537.020 260.000 ;
        RECT 1714.020 -9.220 1717.020 260.000 ;
        RECT 1894.020 -9.220 1897.020 260.000 ;
        RECT 2074.020 -9.220 2077.020 260.000 ;
        RECT 2254.020 -9.220 2257.020 260.000 ;
        RECT 2434.020 -9.220 2437.020 260.000 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 3260.000 385.020 3538.100 ;
        RECT 562.020 3260.000 565.020 3538.100 ;
        RECT 742.020 3260.000 745.020 3538.100 ;
        RECT 922.020 3260.000 925.020 3538.100 ;
        RECT 1102.020 3260.000 1105.020 3538.100 ;
        RECT 1282.020 3260.000 1285.020 3538.100 ;
        RECT 1462.020 3260.000 1465.020 3538.100 ;
        RECT 1642.020 3260.000 1645.020 3538.100 ;
        RECT 1822.020 3260.000 1825.020 3538.100 ;
        RECT 2002.020 3260.000 2005.020 3538.100 ;
        RECT 2182.020 3260.000 2185.020 3538.100 ;
        RECT 2362.020 3260.000 2365.020 3538.100 ;
        RECT 2542.020 3260.000 2545.020 3538.100 ;
        RECT 382.020 -18.420 385.020 260.000 ;
        RECT 562.020 -18.420 565.020 260.000 ;
        RECT 742.020 -18.420 745.020 260.000 ;
        RECT 922.020 -18.420 925.020 260.000 ;
        RECT 1102.020 -18.420 1105.020 260.000 ;
        RECT 1282.020 -18.420 1285.020 260.000 ;
        RECT 1462.020 -18.420 1465.020 260.000 ;
        RECT 1642.020 -18.420 1645.020 260.000 ;
        RECT 1822.020 -18.420 1825.020 260.000 ;
        RECT 2002.020 -18.420 2005.020 260.000 ;
        RECT 2182.020 -18.420 2185.020 260.000 ;
        RECT 2362.020 -18.420 2365.020 260.000 ;
        RECT 2542.020 -18.420 2545.020 260.000 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 3260.000 475.020 3538.100 ;
        RECT 652.020 3260.000 655.020 3538.100 ;
        RECT 832.020 3260.000 835.020 3538.100 ;
        RECT 1012.020 3260.000 1015.020 3538.100 ;
        RECT 1192.020 3260.000 1195.020 3538.100 ;
        RECT 1372.020 3260.000 1375.020 3538.100 ;
        RECT 1552.020 3260.000 1555.020 3538.100 ;
        RECT 1732.020 3260.000 1735.020 3538.100 ;
        RECT 1912.020 3260.000 1915.020 3538.100 ;
        RECT 2092.020 3260.000 2095.020 3538.100 ;
        RECT 2272.020 3260.000 2275.020 3538.100 ;
        RECT 2452.020 3260.000 2455.020 3538.100 ;
        RECT 472.020 -18.420 475.020 260.000 ;
        RECT 652.020 -18.420 655.020 260.000 ;
        RECT 832.020 -18.420 835.020 260.000 ;
        RECT 1012.020 -18.420 1015.020 260.000 ;
        RECT 1192.020 -18.420 1195.020 260.000 ;
        RECT 1372.020 -18.420 1375.020 260.000 ;
        RECT 1552.020 -18.420 1555.020 260.000 ;
        RECT 1732.020 -18.420 1735.020 260.000 ;
        RECT 1912.020 -18.420 1915.020 260.000 ;
        RECT 2092.020 -18.420 2095.020 260.000 ;
        RECT 2272.020 -18.420 2275.020 260.000 ;
        RECT 2452.020 -18.420 2455.020 260.000 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 3260.000 403.020 3547.300 ;
        RECT 580.020 3260.000 583.020 3547.300 ;
        RECT 760.020 3260.000 763.020 3547.300 ;
        RECT 940.020 3260.000 943.020 3547.300 ;
        RECT 1120.020 3260.000 1123.020 3547.300 ;
        RECT 1300.020 3260.000 1303.020 3547.300 ;
        RECT 1480.020 3260.000 1483.020 3547.300 ;
        RECT 1660.020 3260.000 1663.020 3547.300 ;
        RECT 1840.020 3260.000 1843.020 3547.300 ;
        RECT 2020.020 3260.000 2023.020 3547.300 ;
        RECT 2200.020 3260.000 2203.020 3547.300 ;
        RECT 2380.020 3260.000 2383.020 3547.300 ;
        RECT 2560.020 3260.000 2563.020 3547.300 ;
        RECT 400.020 -27.620 403.020 260.000 ;
        RECT 580.020 -27.620 583.020 260.000 ;
        RECT 760.020 -27.620 763.020 260.000 ;
        RECT 940.020 -27.620 943.020 260.000 ;
        RECT 1120.020 -27.620 1123.020 260.000 ;
        RECT 1300.020 -27.620 1303.020 260.000 ;
        RECT 1480.020 -27.620 1483.020 260.000 ;
        RECT 1660.020 -27.620 1663.020 260.000 ;
        RECT 1840.020 -27.620 1843.020 260.000 ;
        RECT 2020.020 -27.620 2023.020 260.000 ;
        RECT 2200.020 -27.620 2203.020 260.000 ;
        RECT 2380.020 -27.620 2383.020 260.000 ;
        RECT 2560.020 -27.620 2563.020 260.000 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 3260.000 313.020 3547.300 ;
        RECT 490.020 3260.000 493.020 3547.300 ;
        RECT 670.020 3260.000 673.020 3547.300 ;
        RECT 850.020 3260.000 853.020 3547.300 ;
        RECT 1030.020 3260.000 1033.020 3547.300 ;
        RECT 1210.020 3260.000 1213.020 3547.300 ;
        RECT 1390.020 3260.000 1393.020 3547.300 ;
        RECT 1570.020 3260.000 1573.020 3547.300 ;
        RECT 1750.020 3260.000 1753.020 3547.300 ;
        RECT 1930.020 3260.000 1933.020 3547.300 ;
        RECT 2110.020 3260.000 2113.020 3547.300 ;
        RECT 2290.020 3260.000 2293.020 3547.300 ;
        RECT 2470.020 3260.000 2473.020 3547.300 ;
        RECT 310.020 -27.620 313.020 260.000 ;
        RECT 490.020 -27.620 493.020 260.000 ;
        RECT 670.020 -27.620 673.020 260.000 ;
        RECT 850.020 -27.620 853.020 260.000 ;
        RECT 1030.020 -27.620 1033.020 260.000 ;
        RECT 1210.020 -27.620 1213.020 260.000 ;
        RECT 1390.020 -27.620 1393.020 260.000 ;
        RECT 1570.020 -27.620 1573.020 260.000 ;
        RECT 1750.020 -27.620 1753.020 260.000 ;
        RECT 1930.020 -27.620 1933.020 260.000 ;
        RECT 2110.020 -27.620 2113.020 260.000 ;
        RECT 2290.020 -27.620 2293.020 260.000 ;
        RECT 2470.020 -27.620 2473.020 260.000 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 3260.000 421.020 3556.500 ;
        RECT 598.020 3260.000 601.020 3556.500 ;
        RECT 778.020 3260.000 781.020 3556.500 ;
        RECT 958.020 3260.000 961.020 3556.500 ;
        RECT 1138.020 3260.000 1141.020 3556.500 ;
        RECT 1318.020 3260.000 1321.020 3556.500 ;
        RECT 1498.020 3260.000 1501.020 3556.500 ;
        RECT 1678.020 3260.000 1681.020 3556.500 ;
        RECT 1858.020 3260.000 1861.020 3556.500 ;
        RECT 2038.020 3260.000 2041.020 3556.500 ;
        RECT 2218.020 3260.000 2221.020 3556.500 ;
        RECT 2398.020 3260.000 2401.020 3556.500 ;
        RECT 2578.020 3260.000 2581.020 3556.500 ;
        RECT 418.020 -36.820 421.020 260.000 ;
        RECT 598.020 -36.820 601.020 260.000 ;
        RECT 778.020 -36.820 781.020 260.000 ;
        RECT 958.020 -36.820 961.020 260.000 ;
        RECT 1138.020 -36.820 1141.020 260.000 ;
        RECT 1318.020 -36.820 1321.020 260.000 ;
        RECT 1498.020 -36.820 1501.020 260.000 ;
        RECT 1678.020 -36.820 1681.020 260.000 ;
        RECT 1858.020 -36.820 1861.020 260.000 ;
        RECT 2038.020 -36.820 2041.020 260.000 ;
        RECT 2218.020 -36.820 2221.020 260.000 ;
        RECT 2398.020 -36.820 2401.020 260.000 ;
        RECT 2578.020 -36.820 2581.020 260.000 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 3260.000 331.020 3556.500 ;
        RECT 508.020 3260.000 511.020 3556.500 ;
        RECT 688.020 3260.000 691.020 3556.500 ;
        RECT 868.020 3260.000 871.020 3556.500 ;
        RECT 1048.020 3260.000 1051.020 3556.500 ;
        RECT 1228.020 3260.000 1231.020 3556.500 ;
        RECT 1408.020 3260.000 1411.020 3556.500 ;
        RECT 1588.020 3260.000 1591.020 3556.500 ;
        RECT 1768.020 3260.000 1771.020 3556.500 ;
        RECT 1948.020 3260.000 1951.020 3556.500 ;
        RECT 2128.020 3260.000 2131.020 3556.500 ;
        RECT 2308.020 3260.000 2311.020 3556.500 ;
        RECT 2488.020 3260.000 2491.020 3556.500 ;
        RECT 328.020 -36.820 331.020 260.000 ;
        RECT 508.020 -36.820 511.020 260.000 ;
        RECT 688.020 -36.820 691.020 260.000 ;
        RECT 868.020 -36.820 871.020 260.000 ;
        RECT 1048.020 -36.820 1051.020 260.000 ;
        RECT 1228.020 -36.820 1231.020 260.000 ;
        RECT 1408.020 -36.820 1411.020 260.000 ;
        RECT 1588.020 -36.820 1591.020 260.000 ;
        RECT 1768.020 -36.820 1771.020 260.000 ;
        RECT 1948.020 -36.820 1951.020 260.000 ;
        RECT 2128.020 -36.820 2131.020 260.000 ;
        RECT 2308.020 -36.820 2311.020 260.000 ;
        RECT 2488.020 -36.820 2491.020 260.000 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 315.520 270.795 2605.715 3246.645 ;
      LAYER met1 ;
        RECT 312.830 264.460 2605.775 3246.800 ;
      LAYER met2 ;
        RECT 312.860 3255.720 352.130 3256.000 ;
        RECT 352.970 3255.720 437.230 3256.000 ;
        RECT 438.070 3255.720 522.330 3256.000 ;
        RECT 523.170 3255.720 607.430 3256.000 ;
        RECT 608.270 3255.720 692.530 3256.000 ;
        RECT 693.370 3255.720 777.630 3256.000 ;
        RECT 778.470 3255.720 863.190 3256.000 ;
        RECT 864.030 3255.720 948.290 3256.000 ;
        RECT 949.130 3255.720 1033.390 3256.000 ;
        RECT 1034.230 3255.720 1118.490 3256.000 ;
        RECT 1119.330 3255.720 1203.590 3256.000 ;
        RECT 1204.430 3255.720 1289.150 3256.000 ;
        RECT 1289.990 3255.720 1374.250 3256.000 ;
        RECT 1375.090 3255.720 1459.350 3256.000 ;
        RECT 1460.190 3255.720 1544.450 3256.000 ;
        RECT 1545.290 3255.720 1629.550 3256.000 ;
        RECT 1630.390 3255.720 1714.650 3256.000 ;
        RECT 1715.490 3255.720 1800.210 3256.000 ;
        RECT 1801.050 3255.720 1885.310 3256.000 ;
        RECT 1886.150 3255.720 1970.410 3256.000 ;
        RECT 1971.250 3255.720 2055.510 3256.000 ;
        RECT 2056.350 3255.720 2140.610 3256.000 ;
        RECT 2141.450 3255.720 2226.170 3256.000 ;
        RECT 2227.010 3255.720 2311.270 3256.000 ;
        RECT 2312.110 3255.720 2396.370 3256.000 ;
        RECT 2397.210 3255.720 2481.470 3256.000 ;
        RECT 2482.310 3255.720 2566.570 3256.000 ;
        RECT 2567.410 3255.720 2602.080 3256.000 ;
        RECT 312.860 264.280 2602.080 3255.720 ;
        RECT 313.410 264.000 318.090 264.280 ;
        RECT 318.930 264.000 324.070 264.280 ;
        RECT 324.910 264.000 330.050 264.280 ;
        RECT 330.890 264.000 336.030 264.280 ;
        RECT 336.870 264.000 342.010 264.280 ;
        RECT 342.850 264.000 347.990 264.280 ;
        RECT 348.830 264.000 353.970 264.280 ;
        RECT 354.810 264.000 359.950 264.280 ;
        RECT 360.790 264.000 365.930 264.280 ;
        RECT 366.770 264.000 371.910 264.280 ;
        RECT 372.750 264.000 377.890 264.280 ;
        RECT 378.730 264.000 383.870 264.280 ;
        RECT 384.710 264.000 389.850 264.280 ;
        RECT 390.690 264.000 395.830 264.280 ;
        RECT 396.670 264.000 401.810 264.280 ;
        RECT 402.650 264.000 407.790 264.280 ;
        RECT 408.630 264.000 413.770 264.280 ;
        RECT 414.610 264.000 419.750 264.280 ;
        RECT 420.590 264.000 425.730 264.280 ;
        RECT 426.570 264.000 431.710 264.280 ;
        RECT 432.550 264.000 437.690 264.280 ;
        RECT 438.530 264.000 443.210 264.280 ;
        RECT 444.050 264.000 449.190 264.280 ;
        RECT 450.030 264.000 455.170 264.280 ;
        RECT 456.010 264.000 461.150 264.280 ;
        RECT 461.990 264.000 467.130 264.280 ;
        RECT 467.970 264.000 473.110 264.280 ;
        RECT 473.950 264.000 479.090 264.280 ;
        RECT 479.930 264.000 485.070 264.280 ;
        RECT 485.910 264.000 491.050 264.280 ;
        RECT 491.890 264.000 497.030 264.280 ;
        RECT 497.870 264.000 503.010 264.280 ;
        RECT 503.850 264.000 508.990 264.280 ;
        RECT 509.830 264.000 514.970 264.280 ;
        RECT 515.810 264.000 520.950 264.280 ;
        RECT 521.790 264.000 526.930 264.280 ;
        RECT 527.770 264.000 532.910 264.280 ;
        RECT 533.750 264.000 538.890 264.280 ;
        RECT 539.730 264.000 544.870 264.280 ;
        RECT 545.710 264.000 550.850 264.280 ;
        RECT 551.690 264.000 556.830 264.280 ;
        RECT 557.670 264.000 562.810 264.280 ;
        RECT 563.650 264.000 568.330 264.280 ;
        RECT 569.170 264.000 574.310 264.280 ;
        RECT 575.150 264.000 580.290 264.280 ;
        RECT 581.130 264.000 586.270 264.280 ;
        RECT 587.110 264.000 592.250 264.280 ;
        RECT 593.090 264.000 598.230 264.280 ;
        RECT 599.070 264.000 604.210 264.280 ;
        RECT 605.050 264.000 610.190 264.280 ;
        RECT 611.030 264.000 616.170 264.280 ;
        RECT 617.010 264.000 622.150 264.280 ;
        RECT 622.990 264.000 628.130 264.280 ;
        RECT 628.970 264.000 634.110 264.280 ;
        RECT 634.950 264.000 640.090 264.280 ;
        RECT 640.930 264.000 646.070 264.280 ;
        RECT 646.910 264.000 652.050 264.280 ;
        RECT 652.890 264.000 658.030 264.280 ;
        RECT 658.870 264.000 664.010 264.280 ;
        RECT 664.850 264.000 669.990 264.280 ;
        RECT 670.830 264.000 675.970 264.280 ;
        RECT 676.810 264.000 681.950 264.280 ;
        RECT 682.790 264.000 687.930 264.280 ;
        RECT 688.770 264.000 693.910 264.280 ;
        RECT 694.750 264.000 699.430 264.280 ;
        RECT 700.270 264.000 705.410 264.280 ;
        RECT 706.250 264.000 711.390 264.280 ;
        RECT 712.230 264.000 717.370 264.280 ;
        RECT 718.210 264.000 723.350 264.280 ;
        RECT 724.190 264.000 729.330 264.280 ;
        RECT 730.170 264.000 735.310 264.280 ;
        RECT 736.150 264.000 741.290 264.280 ;
        RECT 742.130 264.000 747.270 264.280 ;
        RECT 748.110 264.000 753.250 264.280 ;
        RECT 754.090 264.000 759.230 264.280 ;
        RECT 760.070 264.000 765.210 264.280 ;
        RECT 766.050 264.000 771.190 264.280 ;
        RECT 772.030 264.000 777.170 264.280 ;
        RECT 778.010 264.000 783.150 264.280 ;
        RECT 783.990 264.000 789.130 264.280 ;
        RECT 789.970 264.000 795.110 264.280 ;
        RECT 795.950 264.000 801.090 264.280 ;
        RECT 801.930 264.000 807.070 264.280 ;
        RECT 807.910 264.000 813.050 264.280 ;
        RECT 813.890 264.000 819.030 264.280 ;
        RECT 819.870 264.000 824.550 264.280 ;
        RECT 825.390 264.000 830.530 264.280 ;
        RECT 831.370 264.000 836.510 264.280 ;
        RECT 837.350 264.000 842.490 264.280 ;
        RECT 843.330 264.000 848.470 264.280 ;
        RECT 849.310 264.000 854.450 264.280 ;
        RECT 855.290 264.000 860.430 264.280 ;
        RECT 861.270 264.000 866.410 264.280 ;
        RECT 867.250 264.000 872.390 264.280 ;
        RECT 873.230 264.000 878.370 264.280 ;
        RECT 879.210 264.000 884.350 264.280 ;
        RECT 885.190 264.000 890.330 264.280 ;
        RECT 891.170 264.000 896.310 264.280 ;
        RECT 897.150 264.000 902.290 264.280 ;
        RECT 903.130 264.000 908.270 264.280 ;
        RECT 909.110 264.000 914.250 264.280 ;
        RECT 915.090 264.000 920.230 264.280 ;
        RECT 921.070 264.000 926.210 264.280 ;
        RECT 927.050 264.000 932.190 264.280 ;
        RECT 933.030 264.000 938.170 264.280 ;
        RECT 939.010 264.000 944.150 264.280 ;
        RECT 944.990 264.000 950.130 264.280 ;
        RECT 950.970 264.000 955.650 264.280 ;
        RECT 956.490 264.000 961.630 264.280 ;
        RECT 962.470 264.000 967.610 264.280 ;
        RECT 968.450 264.000 973.590 264.280 ;
        RECT 974.430 264.000 979.570 264.280 ;
        RECT 980.410 264.000 985.550 264.280 ;
        RECT 986.390 264.000 991.530 264.280 ;
        RECT 992.370 264.000 997.510 264.280 ;
        RECT 998.350 264.000 1003.490 264.280 ;
        RECT 1004.330 264.000 1009.470 264.280 ;
        RECT 1010.310 264.000 1015.450 264.280 ;
        RECT 1016.290 264.000 1021.430 264.280 ;
        RECT 1022.270 264.000 1027.410 264.280 ;
        RECT 1028.250 264.000 1033.390 264.280 ;
        RECT 1034.230 264.000 1039.370 264.280 ;
        RECT 1040.210 264.000 1045.350 264.280 ;
        RECT 1046.190 264.000 1051.330 264.280 ;
        RECT 1052.170 264.000 1057.310 264.280 ;
        RECT 1058.150 264.000 1063.290 264.280 ;
        RECT 1064.130 264.000 1069.270 264.280 ;
        RECT 1070.110 264.000 1075.250 264.280 ;
        RECT 1076.090 264.000 1080.770 264.280 ;
        RECT 1081.610 264.000 1086.750 264.280 ;
        RECT 1087.590 264.000 1092.730 264.280 ;
        RECT 1093.570 264.000 1098.710 264.280 ;
        RECT 1099.550 264.000 1104.690 264.280 ;
        RECT 1105.530 264.000 1110.670 264.280 ;
        RECT 1111.510 264.000 1116.650 264.280 ;
        RECT 1117.490 264.000 1122.630 264.280 ;
        RECT 1123.470 264.000 1128.610 264.280 ;
        RECT 1129.450 264.000 1134.590 264.280 ;
        RECT 1135.430 264.000 1140.570 264.280 ;
        RECT 1141.410 264.000 1146.550 264.280 ;
        RECT 1147.390 264.000 1152.530 264.280 ;
        RECT 1153.370 264.000 1158.510 264.280 ;
        RECT 1159.350 264.000 1164.490 264.280 ;
        RECT 1165.330 264.000 1170.470 264.280 ;
        RECT 1171.310 264.000 1176.450 264.280 ;
        RECT 1177.290 264.000 1182.430 264.280 ;
        RECT 1183.270 264.000 1188.410 264.280 ;
        RECT 1189.250 264.000 1194.390 264.280 ;
        RECT 1195.230 264.000 1200.370 264.280 ;
        RECT 1201.210 264.000 1206.350 264.280 ;
        RECT 1207.190 264.000 1211.870 264.280 ;
        RECT 1212.710 264.000 1217.850 264.280 ;
        RECT 1218.690 264.000 1223.830 264.280 ;
        RECT 1224.670 264.000 1229.810 264.280 ;
        RECT 1230.650 264.000 1235.790 264.280 ;
        RECT 1236.630 264.000 1241.770 264.280 ;
        RECT 1242.610 264.000 1247.750 264.280 ;
        RECT 1248.590 264.000 1253.730 264.280 ;
        RECT 1254.570 264.000 1259.710 264.280 ;
        RECT 1260.550 264.000 1265.690 264.280 ;
        RECT 1266.530 264.000 1271.670 264.280 ;
        RECT 1272.510 264.000 1277.650 264.280 ;
        RECT 1278.490 264.000 1283.630 264.280 ;
        RECT 1284.470 264.000 1289.610 264.280 ;
        RECT 1290.450 264.000 1295.590 264.280 ;
        RECT 1296.430 264.000 1301.570 264.280 ;
        RECT 1302.410 264.000 1307.550 264.280 ;
        RECT 1308.390 264.000 1313.530 264.280 ;
        RECT 1314.370 264.000 1319.510 264.280 ;
        RECT 1320.350 264.000 1325.490 264.280 ;
        RECT 1326.330 264.000 1331.470 264.280 ;
        RECT 1332.310 264.000 1336.990 264.280 ;
        RECT 1337.830 264.000 1342.970 264.280 ;
        RECT 1343.810 264.000 1348.950 264.280 ;
        RECT 1349.790 264.000 1354.930 264.280 ;
        RECT 1355.770 264.000 1360.910 264.280 ;
        RECT 1361.750 264.000 1366.890 264.280 ;
        RECT 1367.730 264.000 1372.870 264.280 ;
        RECT 1373.710 264.000 1378.850 264.280 ;
        RECT 1379.690 264.000 1384.830 264.280 ;
        RECT 1385.670 264.000 1390.810 264.280 ;
        RECT 1391.650 264.000 1396.790 264.280 ;
        RECT 1397.630 264.000 1402.770 264.280 ;
        RECT 1403.610 264.000 1408.750 264.280 ;
        RECT 1409.590 264.000 1414.730 264.280 ;
        RECT 1415.570 264.000 1420.710 264.280 ;
        RECT 1421.550 264.000 1426.690 264.280 ;
        RECT 1427.530 264.000 1432.670 264.280 ;
        RECT 1433.510 264.000 1438.650 264.280 ;
        RECT 1439.490 264.000 1444.630 264.280 ;
        RECT 1445.470 264.000 1450.610 264.280 ;
        RECT 1451.450 264.000 1456.590 264.280 ;
        RECT 1457.430 264.000 1462.570 264.280 ;
        RECT 1463.410 264.000 1468.090 264.280 ;
        RECT 1468.930 264.000 1474.070 264.280 ;
        RECT 1474.910 264.000 1480.050 264.280 ;
        RECT 1480.890 264.000 1486.030 264.280 ;
        RECT 1486.870 264.000 1492.010 264.280 ;
        RECT 1492.850 264.000 1497.990 264.280 ;
        RECT 1498.830 264.000 1503.970 264.280 ;
        RECT 1504.810 264.000 1509.950 264.280 ;
        RECT 1510.790 264.000 1515.930 264.280 ;
        RECT 1516.770 264.000 1521.910 264.280 ;
        RECT 1522.750 264.000 1527.890 264.280 ;
        RECT 1528.730 264.000 1533.870 264.280 ;
        RECT 1534.710 264.000 1539.850 264.280 ;
        RECT 1540.690 264.000 1545.830 264.280 ;
        RECT 1546.670 264.000 1551.810 264.280 ;
        RECT 1552.650 264.000 1557.790 264.280 ;
        RECT 1558.630 264.000 1563.770 264.280 ;
        RECT 1564.610 264.000 1569.750 264.280 ;
        RECT 1570.590 264.000 1575.730 264.280 ;
        RECT 1576.570 264.000 1581.710 264.280 ;
        RECT 1582.550 264.000 1587.690 264.280 ;
        RECT 1588.530 264.000 1593.210 264.280 ;
        RECT 1594.050 264.000 1599.190 264.280 ;
        RECT 1600.030 264.000 1605.170 264.280 ;
        RECT 1606.010 264.000 1611.150 264.280 ;
        RECT 1611.990 264.000 1617.130 264.280 ;
        RECT 1617.970 264.000 1623.110 264.280 ;
        RECT 1623.950 264.000 1629.090 264.280 ;
        RECT 1629.930 264.000 1635.070 264.280 ;
        RECT 1635.910 264.000 1641.050 264.280 ;
        RECT 1641.890 264.000 1647.030 264.280 ;
        RECT 1647.870 264.000 1653.010 264.280 ;
        RECT 1653.850 264.000 1658.990 264.280 ;
        RECT 1659.830 264.000 1664.970 264.280 ;
        RECT 1665.810 264.000 1670.950 264.280 ;
        RECT 1671.790 264.000 1676.930 264.280 ;
        RECT 1677.770 264.000 1682.910 264.280 ;
        RECT 1683.750 264.000 1688.890 264.280 ;
        RECT 1689.730 264.000 1694.870 264.280 ;
        RECT 1695.710 264.000 1700.850 264.280 ;
        RECT 1701.690 264.000 1706.830 264.280 ;
        RECT 1707.670 264.000 1712.810 264.280 ;
        RECT 1713.650 264.000 1718.330 264.280 ;
        RECT 1719.170 264.000 1724.310 264.280 ;
        RECT 1725.150 264.000 1730.290 264.280 ;
        RECT 1731.130 264.000 1736.270 264.280 ;
        RECT 1737.110 264.000 1742.250 264.280 ;
        RECT 1743.090 264.000 1748.230 264.280 ;
        RECT 1749.070 264.000 1754.210 264.280 ;
        RECT 1755.050 264.000 1760.190 264.280 ;
        RECT 1761.030 264.000 1766.170 264.280 ;
        RECT 1767.010 264.000 1772.150 264.280 ;
        RECT 1772.990 264.000 1778.130 264.280 ;
        RECT 1778.970 264.000 1784.110 264.280 ;
        RECT 1784.950 264.000 1790.090 264.280 ;
        RECT 1790.930 264.000 1796.070 264.280 ;
        RECT 1796.910 264.000 1802.050 264.280 ;
        RECT 1802.890 264.000 1808.030 264.280 ;
        RECT 1808.870 264.000 1814.010 264.280 ;
        RECT 1814.850 264.000 1819.990 264.280 ;
        RECT 1820.830 264.000 1825.970 264.280 ;
        RECT 1826.810 264.000 1831.950 264.280 ;
        RECT 1832.790 264.000 1837.930 264.280 ;
        RECT 1838.770 264.000 1843.910 264.280 ;
        RECT 1844.750 264.000 1849.430 264.280 ;
        RECT 1850.270 264.000 1855.410 264.280 ;
        RECT 1856.250 264.000 1861.390 264.280 ;
        RECT 1862.230 264.000 1867.370 264.280 ;
        RECT 1868.210 264.000 1873.350 264.280 ;
        RECT 1874.190 264.000 1879.330 264.280 ;
        RECT 1880.170 264.000 1885.310 264.280 ;
        RECT 1886.150 264.000 1891.290 264.280 ;
        RECT 1892.130 264.000 1897.270 264.280 ;
        RECT 1898.110 264.000 1903.250 264.280 ;
        RECT 1904.090 264.000 1909.230 264.280 ;
        RECT 1910.070 264.000 1915.210 264.280 ;
        RECT 1916.050 264.000 1921.190 264.280 ;
        RECT 1922.030 264.000 1927.170 264.280 ;
        RECT 1928.010 264.000 1933.150 264.280 ;
        RECT 1933.990 264.000 1939.130 264.280 ;
        RECT 1939.970 264.000 1945.110 264.280 ;
        RECT 1945.950 264.000 1951.090 264.280 ;
        RECT 1951.930 264.000 1957.070 264.280 ;
        RECT 1957.910 264.000 1963.050 264.280 ;
        RECT 1963.890 264.000 1969.030 264.280 ;
        RECT 1969.870 264.000 1974.550 264.280 ;
        RECT 1975.390 264.000 1980.530 264.280 ;
        RECT 1981.370 264.000 1986.510 264.280 ;
        RECT 1987.350 264.000 1992.490 264.280 ;
        RECT 1993.330 264.000 1998.470 264.280 ;
        RECT 1999.310 264.000 2004.450 264.280 ;
        RECT 2005.290 264.000 2010.430 264.280 ;
        RECT 2011.270 264.000 2016.410 264.280 ;
        RECT 2017.250 264.000 2022.390 264.280 ;
        RECT 2023.230 264.000 2028.370 264.280 ;
        RECT 2029.210 264.000 2034.350 264.280 ;
        RECT 2035.190 264.000 2040.330 264.280 ;
        RECT 2041.170 264.000 2046.310 264.280 ;
        RECT 2047.150 264.000 2052.290 264.280 ;
        RECT 2053.130 264.000 2058.270 264.280 ;
        RECT 2059.110 264.000 2064.250 264.280 ;
        RECT 2065.090 264.000 2070.230 264.280 ;
        RECT 2071.070 264.000 2076.210 264.280 ;
        RECT 2077.050 264.000 2082.190 264.280 ;
        RECT 2083.030 264.000 2088.170 264.280 ;
        RECT 2089.010 264.000 2094.150 264.280 ;
        RECT 2094.990 264.000 2100.130 264.280 ;
        RECT 2100.970 264.000 2105.650 264.280 ;
        RECT 2106.490 264.000 2111.630 264.280 ;
        RECT 2112.470 264.000 2117.610 264.280 ;
        RECT 2118.450 264.000 2123.590 264.280 ;
        RECT 2124.430 264.000 2129.570 264.280 ;
        RECT 2130.410 264.000 2135.550 264.280 ;
        RECT 2136.390 264.000 2141.530 264.280 ;
        RECT 2142.370 264.000 2147.510 264.280 ;
        RECT 2148.350 264.000 2153.490 264.280 ;
        RECT 2154.330 264.000 2159.470 264.280 ;
        RECT 2160.310 264.000 2165.450 264.280 ;
        RECT 2166.290 264.000 2171.430 264.280 ;
        RECT 2172.270 264.000 2177.410 264.280 ;
        RECT 2178.250 264.000 2183.390 264.280 ;
        RECT 2184.230 264.000 2189.370 264.280 ;
        RECT 2190.210 264.000 2195.350 264.280 ;
        RECT 2196.190 264.000 2201.330 264.280 ;
        RECT 2202.170 264.000 2207.310 264.280 ;
        RECT 2208.150 264.000 2213.290 264.280 ;
        RECT 2214.130 264.000 2219.270 264.280 ;
        RECT 2220.110 264.000 2225.250 264.280 ;
        RECT 2226.090 264.000 2230.770 264.280 ;
        RECT 2231.610 264.000 2236.750 264.280 ;
        RECT 2237.590 264.000 2242.730 264.280 ;
        RECT 2243.570 264.000 2248.710 264.280 ;
        RECT 2249.550 264.000 2254.690 264.280 ;
        RECT 2255.530 264.000 2260.670 264.280 ;
        RECT 2261.510 264.000 2266.650 264.280 ;
        RECT 2267.490 264.000 2272.630 264.280 ;
        RECT 2273.470 264.000 2278.610 264.280 ;
        RECT 2279.450 264.000 2284.590 264.280 ;
        RECT 2285.430 264.000 2290.570 264.280 ;
        RECT 2291.410 264.000 2296.550 264.280 ;
        RECT 2297.390 264.000 2302.530 264.280 ;
        RECT 2303.370 264.000 2308.510 264.280 ;
        RECT 2309.350 264.000 2314.490 264.280 ;
        RECT 2315.330 264.000 2320.470 264.280 ;
        RECT 2321.310 264.000 2326.450 264.280 ;
        RECT 2327.290 264.000 2332.430 264.280 ;
        RECT 2333.270 264.000 2338.410 264.280 ;
        RECT 2339.250 264.000 2344.390 264.280 ;
        RECT 2345.230 264.000 2350.370 264.280 ;
        RECT 2351.210 264.000 2356.350 264.280 ;
        RECT 2357.190 264.000 2361.870 264.280 ;
        RECT 2362.710 264.000 2367.850 264.280 ;
        RECT 2368.690 264.000 2373.830 264.280 ;
        RECT 2374.670 264.000 2379.810 264.280 ;
        RECT 2380.650 264.000 2385.790 264.280 ;
        RECT 2386.630 264.000 2391.770 264.280 ;
        RECT 2392.610 264.000 2397.750 264.280 ;
        RECT 2398.590 264.000 2403.730 264.280 ;
        RECT 2404.570 264.000 2409.710 264.280 ;
        RECT 2410.550 264.000 2415.690 264.280 ;
        RECT 2416.530 264.000 2421.670 264.280 ;
        RECT 2422.510 264.000 2427.650 264.280 ;
        RECT 2428.490 264.000 2433.630 264.280 ;
        RECT 2434.470 264.000 2439.610 264.280 ;
        RECT 2440.450 264.000 2445.590 264.280 ;
        RECT 2446.430 264.000 2451.570 264.280 ;
        RECT 2452.410 264.000 2457.550 264.280 ;
        RECT 2458.390 264.000 2463.530 264.280 ;
        RECT 2464.370 264.000 2469.510 264.280 ;
        RECT 2470.350 264.000 2475.490 264.280 ;
        RECT 2476.330 264.000 2481.470 264.280 ;
        RECT 2482.310 264.000 2486.990 264.280 ;
        RECT 2487.830 264.000 2492.970 264.280 ;
        RECT 2493.810 264.000 2498.950 264.280 ;
        RECT 2499.790 264.000 2504.930 264.280 ;
        RECT 2505.770 264.000 2510.910 264.280 ;
        RECT 2511.750 264.000 2516.890 264.280 ;
        RECT 2517.730 264.000 2522.870 264.280 ;
        RECT 2523.710 264.000 2528.850 264.280 ;
        RECT 2529.690 264.000 2534.830 264.280 ;
        RECT 2535.670 264.000 2540.810 264.280 ;
        RECT 2541.650 264.000 2546.790 264.280 ;
        RECT 2547.630 264.000 2552.770 264.280 ;
        RECT 2553.610 264.000 2558.750 264.280 ;
        RECT 2559.590 264.000 2564.730 264.280 ;
        RECT 2565.570 264.000 2570.710 264.280 ;
        RECT 2571.550 264.000 2576.690 264.280 ;
        RECT 2577.530 264.000 2582.670 264.280 ;
        RECT 2583.510 264.000 2588.650 264.280 ;
        RECT 2589.490 264.000 2594.630 264.280 ;
        RECT 2595.470 264.000 2600.610 264.280 ;
        RECT 2601.450 264.000 2602.080 264.280 ;
      LAYER met3 ;
        RECT 314.000 3227.200 2606.000 3246.725 ;
        RECT 314.000 3225.800 2605.600 3227.200 ;
        RECT 314.000 3224.480 2606.000 3225.800 ;
        RECT 314.400 3223.080 2606.000 3224.480 ;
        RECT 314.000 3160.560 2606.000 3223.080 ;
        RECT 314.000 3159.160 2605.600 3160.560 ;
        RECT 314.000 3153.080 2606.000 3159.160 ;
        RECT 314.400 3151.680 2606.000 3153.080 ;
        RECT 314.000 3093.920 2606.000 3151.680 ;
        RECT 314.000 3092.520 2605.600 3093.920 ;
        RECT 314.000 3081.680 2606.000 3092.520 ;
        RECT 314.400 3080.280 2606.000 3081.680 ;
        RECT 314.000 3027.280 2606.000 3080.280 ;
        RECT 314.000 3025.880 2605.600 3027.280 ;
        RECT 314.000 3010.280 2606.000 3025.880 ;
        RECT 314.400 3008.880 2606.000 3010.280 ;
        RECT 314.000 2960.640 2606.000 3008.880 ;
        RECT 314.000 2959.240 2605.600 2960.640 ;
        RECT 314.000 2938.880 2606.000 2959.240 ;
        RECT 314.400 2937.480 2606.000 2938.880 ;
        RECT 314.000 2894.000 2606.000 2937.480 ;
        RECT 314.000 2892.600 2605.600 2894.000 ;
        RECT 314.000 2867.480 2606.000 2892.600 ;
        RECT 314.400 2866.080 2606.000 2867.480 ;
        RECT 314.000 2827.360 2606.000 2866.080 ;
        RECT 314.000 2825.960 2605.600 2827.360 ;
        RECT 314.000 2796.080 2606.000 2825.960 ;
        RECT 314.400 2794.680 2606.000 2796.080 ;
        RECT 314.000 2760.720 2606.000 2794.680 ;
        RECT 314.000 2759.320 2605.600 2760.720 ;
        RECT 314.000 2724.680 2606.000 2759.320 ;
        RECT 314.400 2723.280 2606.000 2724.680 ;
        RECT 314.000 2694.080 2606.000 2723.280 ;
        RECT 314.000 2692.680 2605.600 2694.080 ;
        RECT 314.000 2653.280 2606.000 2692.680 ;
        RECT 314.400 2651.880 2606.000 2653.280 ;
        RECT 314.000 2627.440 2606.000 2651.880 ;
        RECT 314.000 2626.040 2605.600 2627.440 ;
        RECT 314.000 2581.880 2606.000 2626.040 ;
        RECT 314.400 2580.480 2606.000 2581.880 ;
        RECT 314.000 2560.800 2606.000 2580.480 ;
        RECT 314.000 2559.400 2605.600 2560.800 ;
        RECT 314.000 2510.480 2606.000 2559.400 ;
        RECT 314.400 2509.080 2606.000 2510.480 ;
        RECT 314.000 2494.160 2606.000 2509.080 ;
        RECT 314.000 2492.760 2605.600 2494.160 ;
        RECT 314.000 2439.080 2606.000 2492.760 ;
        RECT 314.400 2437.680 2606.000 2439.080 ;
        RECT 314.000 2427.520 2606.000 2437.680 ;
        RECT 314.000 2426.120 2605.600 2427.520 ;
        RECT 314.000 2367.680 2606.000 2426.120 ;
        RECT 314.400 2366.280 2606.000 2367.680 ;
        RECT 314.000 2360.880 2606.000 2366.280 ;
        RECT 314.000 2359.480 2605.600 2360.880 ;
        RECT 314.000 2296.280 2606.000 2359.480 ;
        RECT 314.400 2294.880 2606.000 2296.280 ;
        RECT 314.000 2294.240 2606.000 2294.880 ;
        RECT 314.000 2292.840 2605.600 2294.240 ;
        RECT 314.000 2227.600 2606.000 2292.840 ;
        RECT 314.000 2226.200 2605.600 2227.600 ;
        RECT 314.000 2224.880 2606.000 2226.200 ;
        RECT 314.400 2223.480 2606.000 2224.880 ;
        RECT 314.000 2160.960 2606.000 2223.480 ;
        RECT 314.000 2159.560 2605.600 2160.960 ;
        RECT 314.000 2153.480 2606.000 2159.560 ;
        RECT 314.400 2152.080 2606.000 2153.480 ;
        RECT 314.000 2094.320 2606.000 2152.080 ;
        RECT 314.000 2092.920 2605.600 2094.320 ;
        RECT 314.000 2082.080 2606.000 2092.920 ;
        RECT 314.400 2080.680 2606.000 2082.080 ;
        RECT 314.000 2027.680 2606.000 2080.680 ;
        RECT 314.000 2026.280 2605.600 2027.680 ;
        RECT 314.000 2010.680 2606.000 2026.280 ;
        RECT 314.400 2009.280 2606.000 2010.680 ;
        RECT 314.000 1961.040 2606.000 2009.280 ;
        RECT 314.000 1959.640 2605.600 1961.040 ;
        RECT 314.000 1939.280 2606.000 1959.640 ;
        RECT 314.400 1937.880 2606.000 1939.280 ;
        RECT 314.000 1894.400 2606.000 1937.880 ;
        RECT 314.000 1893.000 2605.600 1894.400 ;
        RECT 314.000 1867.880 2606.000 1893.000 ;
        RECT 314.400 1866.480 2606.000 1867.880 ;
        RECT 314.000 1827.760 2606.000 1866.480 ;
        RECT 314.000 1826.360 2605.600 1827.760 ;
        RECT 314.000 1796.480 2606.000 1826.360 ;
        RECT 314.400 1795.080 2606.000 1796.480 ;
        RECT 314.000 1760.440 2606.000 1795.080 ;
        RECT 314.000 1759.040 2605.600 1760.440 ;
        RECT 314.000 1724.400 2606.000 1759.040 ;
        RECT 314.400 1723.000 2606.000 1724.400 ;
        RECT 314.000 1693.800 2606.000 1723.000 ;
        RECT 314.000 1692.400 2605.600 1693.800 ;
        RECT 314.000 1653.000 2606.000 1692.400 ;
        RECT 314.400 1651.600 2606.000 1653.000 ;
        RECT 314.000 1627.160 2606.000 1651.600 ;
        RECT 314.000 1625.760 2605.600 1627.160 ;
        RECT 314.000 1581.600 2606.000 1625.760 ;
        RECT 314.400 1580.200 2606.000 1581.600 ;
        RECT 314.000 1560.520 2606.000 1580.200 ;
        RECT 314.000 1559.120 2605.600 1560.520 ;
        RECT 314.000 1510.200 2606.000 1559.120 ;
        RECT 314.400 1508.800 2606.000 1510.200 ;
        RECT 314.000 1493.880 2606.000 1508.800 ;
        RECT 314.000 1492.480 2605.600 1493.880 ;
        RECT 314.000 1438.800 2606.000 1492.480 ;
        RECT 314.400 1437.400 2606.000 1438.800 ;
        RECT 314.000 1427.240 2606.000 1437.400 ;
        RECT 314.000 1425.840 2605.600 1427.240 ;
        RECT 314.000 1367.400 2606.000 1425.840 ;
        RECT 314.400 1366.000 2606.000 1367.400 ;
        RECT 314.000 1360.600 2606.000 1366.000 ;
        RECT 314.000 1359.200 2605.600 1360.600 ;
        RECT 314.000 1296.000 2606.000 1359.200 ;
        RECT 314.400 1294.600 2606.000 1296.000 ;
        RECT 314.000 1293.960 2606.000 1294.600 ;
        RECT 314.000 1292.560 2605.600 1293.960 ;
        RECT 314.000 1227.320 2606.000 1292.560 ;
        RECT 314.000 1225.920 2605.600 1227.320 ;
        RECT 314.000 1224.600 2606.000 1225.920 ;
        RECT 314.400 1223.200 2606.000 1224.600 ;
        RECT 314.000 1160.680 2606.000 1223.200 ;
        RECT 314.000 1159.280 2605.600 1160.680 ;
        RECT 314.000 1153.200 2606.000 1159.280 ;
        RECT 314.400 1151.800 2606.000 1153.200 ;
        RECT 314.000 1094.040 2606.000 1151.800 ;
        RECT 314.000 1092.640 2605.600 1094.040 ;
        RECT 314.000 1081.800 2606.000 1092.640 ;
        RECT 314.400 1080.400 2606.000 1081.800 ;
        RECT 314.000 1027.400 2606.000 1080.400 ;
        RECT 314.000 1026.000 2605.600 1027.400 ;
        RECT 314.000 1010.400 2606.000 1026.000 ;
        RECT 314.400 1009.000 2606.000 1010.400 ;
        RECT 314.000 960.760 2606.000 1009.000 ;
        RECT 314.000 959.360 2605.600 960.760 ;
        RECT 314.000 939.000 2606.000 959.360 ;
        RECT 314.400 937.600 2606.000 939.000 ;
        RECT 314.000 894.120 2606.000 937.600 ;
        RECT 314.000 892.720 2605.600 894.120 ;
        RECT 314.000 867.600 2606.000 892.720 ;
        RECT 314.400 866.200 2606.000 867.600 ;
        RECT 314.000 827.480 2606.000 866.200 ;
        RECT 314.000 826.080 2605.600 827.480 ;
        RECT 314.000 796.200 2606.000 826.080 ;
        RECT 314.400 794.800 2606.000 796.200 ;
        RECT 314.000 760.840 2606.000 794.800 ;
        RECT 314.000 759.440 2605.600 760.840 ;
        RECT 314.000 724.800 2606.000 759.440 ;
        RECT 314.400 723.400 2606.000 724.800 ;
        RECT 314.000 694.200 2606.000 723.400 ;
        RECT 314.000 692.800 2605.600 694.200 ;
        RECT 314.000 653.400 2606.000 692.800 ;
        RECT 314.400 652.000 2606.000 653.400 ;
        RECT 314.000 627.560 2606.000 652.000 ;
        RECT 314.000 626.160 2605.600 627.560 ;
        RECT 314.000 582.000 2606.000 626.160 ;
        RECT 314.400 580.600 2606.000 582.000 ;
        RECT 314.000 560.920 2606.000 580.600 ;
        RECT 314.000 559.520 2605.600 560.920 ;
        RECT 314.000 510.600 2606.000 559.520 ;
        RECT 314.400 509.200 2606.000 510.600 ;
        RECT 314.000 494.280 2606.000 509.200 ;
        RECT 314.000 492.880 2605.600 494.280 ;
        RECT 314.000 439.200 2606.000 492.880 ;
        RECT 314.400 437.800 2606.000 439.200 ;
        RECT 314.000 427.640 2606.000 437.800 ;
        RECT 314.000 426.240 2605.600 427.640 ;
        RECT 314.000 367.800 2606.000 426.240 ;
        RECT 314.400 366.400 2606.000 367.800 ;
        RECT 314.000 361.000 2606.000 366.400 ;
        RECT 314.000 359.600 2605.600 361.000 ;
        RECT 314.000 296.400 2606.000 359.600 ;
        RECT 314.400 295.000 2606.000 296.400 ;
        RECT 314.000 294.360 2606.000 295.000 ;
        RECT 314.000 292.960 2605.600 294.360 ;
        RECT 314.000 270.715 2606.000 292.960 ;
      LAYER met4 ;
        RECT 325.015 270.640 330.640 3246.800 ;
      LAYER met4 ;
        RECT 331.040 270.640 332.640 3246.800 ;
      LAYER met4 ;
        RECT 333.040 270.640 407.440 3246.800 ;
      LAYER met4 ;
        RECT 407.840 270.640 409.440 3246.800 ;
      LAYER met4 ;
        RECT 409.840 270.640 2591.305 3246.800 ;
  END
END user_project_wrapper
END LIBRARY

