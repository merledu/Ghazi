VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ghazi_top_dffram_csv
  CLASS BLOCK ;
  FOREIGN ghazi_top_dffram_csv ;
  ORIGIN 0.000 0.000 ;
  SIZE 2300.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2899.560 4.000 2900.160 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1368.200 2300.000 1368.800 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1696.570 2996.000 1696.850 3000.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1904.490 0.000 1904.770 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1440.280 4.000 1440.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 2996.000 80.410 3000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.410 2996.000 1238.690 3000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2276.170 0.000 2276.450 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 838.210 2996.000 838.490 3000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 945.240 2300.000 945.840 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1653.330 2996.000 1653.610 3000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 267.960 2300.000 268.560 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1103.000 4.000 1103.600 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2445.320 2300.000 2445.920 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2560.920 4.000 2561.520 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.930 0.000 2233.210 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.410 2996.000 824.690 3000.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.490 2996.000 938.770 3000.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 766.450 2996.000 766.730 3000.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2509.240 2300.000 2509.840 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2168.530 2996.000 2168.810 3000.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1853.720 2300.000 1854.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2296.410 2996.000 2296.690 3000.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1196.090 2996.000 1196.370 3000.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 2996.000 23.370 3000.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.730 2996.000 338.010 3000.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1833.320 2300.000 1833.920 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2741.800 2300.000 2742.400 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1536.840 2300.000 1537.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 366.250 2996.000 366.530 3000.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 586.200 2300.000 586.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1494.680 2300.000 1495.280 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1847.450 0.000 1847.730 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.530 2996.000 466.810 3000.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2699.640 2300.000 2700.240 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1553.050 2996.000 1553.330 3000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1472.920 2300.000 1473.520 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1918.290 0.000 1918.570 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1532.810 0.000 1533.090 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2267.890 2996.000 2268.170 3000.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2011.210 2996.000 2011.490 3000.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 15.000 2300.000 15.600 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1139.050 2996.000 1139.330 3000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1389.290 0.000 1389.570 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.290 2996.000 9.570 3000.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2687.400 4.000 2688.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 4.000 1251.840 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2835.640 4.000 2836.240 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1938.040 2300.000 1938.640 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2125.290 2996.000 2125.570 3000.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 552.090 2996.000 552.370 3000.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2239.370 2996.000 2239.650 3000.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1782.130 2996.000 1782.410 3000.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.490 2996.000 409.770 3000.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.490 2996.000 294.770 3000.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1775.690 0.000 1775.970 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1861.250 0.000 1861.530 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1769.400 2300.000 1770.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2805.720 2300.000 2806.320 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2307.960 4.000 2308.560 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1295.450 2996.000 1295.730 3000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1432.530 0.000 1432.810 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2075.610 0.000 2075.890 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2001.960 2300.000 2002.560 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1969.320 4.000 1969.920 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 2996.000 423.570 3000.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2910.440 2300.000 2911.040 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.970 2996.000 910.250 3000.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 797.000 2300.000 797.600 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1353.410 2996.000 1353.690 3000.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 809.690 2996.000 809.970 3000.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 223.650 2996.000 223.930 3000.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 923.480 2300.000 924.080 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1546.360 4.000 1546.960 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2868.280 2300.000 2868.880 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1395.730 2996.000 1396.010 3000.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1262.120 2300.000 1262.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.880 4.000 1420.480 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1839.170 2996.000 1839.450 3000.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1417.810 0.000 1418.090 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 2996.000 95.130 3000.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1231.970 0.000 1232.250 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 733.080 2300.000 733.680 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 331.880 2300.000 332.480 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.810 2996.000 567.090 3000.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1967.970 2996.000 1968.250 3000.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1438.970 2996.000 1439.250 3000.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1990.050 0.000 1990.330 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.080 4.000 1039.680 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1093.480 2300.000 1094.080 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2110.570 2996.000 2110.850 3000.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1905.400 4.000 1906.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2118.850 0.000 2119.130 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2261.450 0.000 2261.730 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 595.330 2996.000 595.610 3000.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 912.600 4.000 913.200 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1624.810 2996.000 1625.090 3000.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.170 0.000 1632.450 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2709.160 4.000 2709.760 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2159.720 4.000 2160.320 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2053.640 4.000 2054.240 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1430.760 2300.000 1431.360 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 225.800 2300.000 226.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2424.920 2300.000 2425.520 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2815.240 4.000 2815.840 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2254.090 2996.000 2254.370 3000.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.650 2996.000 752.930 3000.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2540.520 4.000 2541.120 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.970 2996.000 381.250 3000.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 35.400 2300.000 36.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1825.370 2996.000 1825.650 3000.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 903.080 2300.000 903.680 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1660.690 0.000 1660.970 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2826.120 2300.000 2826.720 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1705.480 2300.000 1706.080 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2128.440 2300.000 2129.040 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 623.850 2996.000 624.130 3000.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1588.520 4.000 1589.120 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 881.320 2300.000 881.920 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.570 2996.000 523.850 3000.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1800.680 4.000 1801.280 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2890.040 2300.000 2890.640 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1452.520 2300.000 1453.120 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2382.760 2300.000 2383.360 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1510.730 2996.000 1511.010 3000.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2137.960 4.000 2138.560 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2498.360 4.000 2498.960 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2573.160 2300.000 2573.760 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2254.920 2300.000 2255.520 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2201.880 4.000 2202.480 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.170 2996.000 1310.450 3000.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2454.840 4.000 2455.440 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 818.760 2300.000 819.360 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1338.690 2996.000 1338.970 3000.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2667.000 4.000 2667.600 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.570 0.000 2018.850 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1539.250 2996.000 1539.530 3000.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2318.840 2300.000 2319.440 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1663.320 2300.000 1663.920 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1610.090 2996.000 1610.370 3000.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2140.010 2996.000 2140.290 3000.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2763.560 2300.000 2764.160 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2847.880 2300.000 2848.480 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2175.890 0.000 2176.170 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 163.240 2300.000 163.840 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1818.010 0.000 1818.290 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1668.050 2996.000 1668.330 3000.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 416.200 2300.000 416.800 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1610.280 4.000 1610.880 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.290 2996.000 1596.570 3000.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1618.370 0.000 1618.650 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1388.600 2300.000 1389.200 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2518.760 4.000 2519.360 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2011.480 4.000 2012.080 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2952.600 2300.000 2953.200 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1324.890 2996.000 1325.170 3000.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2033.290 0.000 2033.570 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2941.720 4.000 2942.320 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.970 2996.000 266.250 3000.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 974.370 0.000 974.650 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1219.960 2300.000 1220.560 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 564.440 2300.000 565.040 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 806.520 4.000 807.120 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2247.650 0.000 2247.930 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1917.640 2300.000 1918.240 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2004.770 0.000 2005.050 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 247.560 2300.000 248.160 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2783.960 2300.000 2784.560 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 923.770 2996.000 924.050 3000.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1461.050 0.000 1461.330 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2328.360 4.000 2328.960 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1975.330 0.000 1975.610 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 394.770 2996.000 395.050 3000.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 121.080 2300.000 121.680 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.410 2996.000 709.690 3000.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1896.210 2996.000 1896.490 3000.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.120 4.000 1398.720 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.810 0.000 1004.090 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 2996.000 252.450 3000.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 860.920 2300.000 861.520 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2117.560 4.000 2118.160 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1747.170 0.000 1747.450 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1980.200 2300.000 1980.800 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1504.200 4.000 1504.800 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1203.450 0.000 1203.730 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2289.970 0.000 2290.250 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 374.040 2300.000 374.640 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1600.760 2300.000 1601.360 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2350.120 4.000 2350.720 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2265.800 4.000 2266.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2180.120 4.000 2180.720 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.250 2996.000 2068.530 3000.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1303.730 0.000 1304.010 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2751.320 4.000 2751.920 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1518.090 0.000 1518.370 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1630.680 4.000 1631.280 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1953.250 2996.000 1953.530 3000.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2932.200 2300.000 2932.800 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1240.360 2300.000 1240.960 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1579.000 2300.000 1579.600 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1821.080 4.000 1821.680 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 2996.000 738.210 3000.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 2996.000 137.450 3000.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1482.210 2996.000 1482.490 3000.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 839.160 2300.000 839.760 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2132.650 0.000 2132.930 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.890 2996.000 1210.170 3000.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1424.250 2996.000 1424.530 3000.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.090 0.000 989.370 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 57.160 2300.000 57.760 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 451.810 2996.000 452.090 3000.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1832.730 0.000 1833.010 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2361.000 2300.000 2361.600 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.050 2996.000 1024.330 3000.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2615.320 2300.000 2615.920 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 481.250 2996.000 481.530 3000.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1736.760 4.000 1737.360 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1135.640 2300.000 1136.240 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1229.480 4.000 1230.080 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2720.040 2300.000 2720.640 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1875.480 2300.000 1876.080 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1758.520 4.000 1759.120 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1346.440 2300.000 1347.040 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1326.040 2300.000 1326.640 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1778.920 4.000 1779.520 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1639.530 2996.000 1639.810 3000.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 311.480 2300.000 312.080 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 965.640 2300.000 966.240 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 670.520 2300.000 671.120 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1289.010 0.000 1289.290 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2212.760 2300.000 2213.360 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 2996.000 66.610 3000.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2645.240 4.000 2645.840 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1725.090 2996.000 1725.370 3000.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1567.770 2996.000 1568.050 3000.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1895.880 2300.000 1896.480 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 652.370 2996.000 652.650 3000.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1038.770 2996.000 1039.050 3000.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2210.850 2996.000 2211.130 3000.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.610 2996.000 166.890 3000.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2412.680 4.000 2413.280 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2551.400 2300.000 2552.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1853.890 2996.000 1854.170 3000.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1381.930 2996.000 1382.210 3000.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1177.800 2300.000 1178.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2403.160 2300.000 2403.760 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 99.320 2300.000 99.920 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1266.930 2996.000 1267.210 3000.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1642.920 2300.000 1643.520 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 702.970 0.000 703.250 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1681.850 2996.000 1682.130 3000.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1675.410 0.000 1675.690 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1718.650 0.000 1718.930 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1946.810 0.000 1947.090 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 981.730 2996.000 982.010 3000.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1685.080 2300.000 1685.680 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.610 0.000 2190.890 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 437.960 2300.000 438.560 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 78.920 2300.000 79.520 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 609.130 2996.000 609.410 3000.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2153.810 2996.000 2154.090 3000.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1060.850 0.000 1061.130 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2047.090 0.000 2047.370 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1007.800 2300.000 1008.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1575.130 0.000 1575.410 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1767.410 2996.000 1767.690 3000.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.960 4.000 1356.560 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1747.640 2300.000 1748.240 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1603.650 0.000 1603.930 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2075.400 4.000 2076.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1789.490 0.000 1789.770 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.000 4.000 1715.600 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2476.600 4.000 2477.200 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2603.080 4.000 2603.680 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1558.600 2300.000 1559.200 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 667.090 2996.000 667.370 3000.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1515.080 2300.000 1515.680 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 141.480 2300.000 142.080 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.890 2996.000 152.170 3000.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2082.050 2996.000 2082.330 3000.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1996.490 2996.000 1996.770 3000.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2773.080 4.000 2773.680 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2033.240 4.000 2033.840 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2340.600 2300.000 2341.200 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.250 2996.000 1010.530 3000.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 960.570 0.000 960.850 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1811.560 2300.000 1812.160 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1410.360 2300.000 1410.960 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1103.170 0.000 1103.450 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2467.080 2300.000 2467.680 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.450 2996.000 881.730 3000.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2044.120 2300.000 2044.720 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 895.250 2996.000 895.530 3000.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.530 2996.000 1524.810 3000.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1690.130 0.000 1690.410 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 0.000 1160.490 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2434.440 4.000 2435.040 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.610 2996.000 580.890 3000.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1124.330 2996.000 1124.610 3000.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1029.560 2300.000 1030.160 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.010 2996.000 438.290 3000.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1452.770 2996.000 1453.050 3000.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 480.120 2300.000 480.720 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1095.810 2996.000 1096.090 3000.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 205.400 2300.000 206.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2974.360 2300.000 2974.960 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 690.920 2300.000 691.520 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 4.000 975.760 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1795.930 2996.000 1796.210 3000.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2090.330 0.000 2090.610 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1051.320 2300.000 1051.920 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1156.040 2300.000 1156.640 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2298.440 2300.000 2299.040 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1224.610 2996.000 1224.890 3000.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1525.960 4.000 1526.560 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1117.890 0.000 1118.170 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1727.240 2300.000 1727.840 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1181.370 2996.000 1181.650 3000.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 775.240 2300.000 775.840 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1991.080 4.000 1991.680 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2192.360 2300.000 2192.960 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1089.370 0.000 1089.650 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 395.800 2300.000 396.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1317.530 0.000 1317.810 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 628.360 2300.000 628.960 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1332.250 0.000 1332.530 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1760.970 0.000 1761.250 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2204.410 0.000 2204.690 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 289.720 2300.000 290.320 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 2996.000 324.210 3000.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 2996.000 123.650 3000.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2793.480 4.000 2794.080 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1885.000 4.000 1885.600 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1313.800 4.000 1314.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2234.520 2300.000 2235.120 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2635.720 2300.000 2636.320 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1939.450 2996.000 1939.730 3000.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2276.680 2300.000 2277.280 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2582.680 4.000 2583.280 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 522.280 2300.000 522.880 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1867.690 2996.000 1867.970 3000.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2108.040 2300.000 2108.640 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1198.200 2300.000 1198.800 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1081.090 2996.000 1081.370 3000.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1253.130 2996.000 1253.410 3000.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.890 2996.000 681.170 3000.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.650 2996.000 1810.930 3000.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1189.650 0.000 1189.930 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1959.800 2300.000 1960.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.450 2996.000 237.730 3000.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2182.330 2996.000 2182.610 3000.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.130 2996.000 195.410 3000.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1581.570 2996.000 1581.850 3000.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2223.640 4.000 2224.240 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1123.400 4.000 1124.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2531.000 2300.000 2531.600 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.690 2996.000 280.970 3000.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2244.040 4.000 2244.640 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.010 2996.000 967.290 3000.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1375.490 0.000 1375.770 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1304.280 2300.000 1304.880 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1933.010 0.000 1933.290 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1982.690 2996.000 1982.970 3000.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1483.800 4.000 1484.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2677.880 2300.000 2678.480 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2286.200 4.000 2286.800 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1496.010 2996.000 1496.290 3000.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1910.930 2996.000 1911.210 3000.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2392.280 4.000 2392.880 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1071.720 2300.000 1072.320 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1074.650 0.000 1074.930 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.450 2996.000 352.730 3000.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1067.290 2996.000 1067.570 3000.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2086.280 2300.000 2086.880 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.410 2996.000 180.690 3000.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2370.520 4.000 2371.120 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2857.400 4.000 2858.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 754.840 2300.000 755.440 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1281.650 2996.000 1281.930 3000.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1113.880 2300.000 1114.480 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2487.480 2300.000 2488.080 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2197.050 2996.000 2197.330 3000.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 544.040 2300.000 544.640 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1842.840 4.000 1843.440 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 458.360 2300.000 458.960 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.170 2996.000 781.450 3000.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 648.760 2300.000 649.360 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1187.320 4.000 1187.920 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1738.890 2996.000 1739.170 3000.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2162.090 0.000 2162.370 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1410.450 2996.000 1410.730 3000.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2104.130 0.000 2104.410 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 353.640 2300.000 354.240 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1694.600 4.000 1695.200 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.930 0.000 1704.210 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2624.840 4.000 2625.440 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 794.970 2996.000 795.250 3000.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2657.480 2300.000 2658.080 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1446.330 0.000 1446.610 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1546.610 0.000 1546.890 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 2996.000 38.090 3000.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2730.920 4.000 2731.520 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.610 2996.000 1109.890 3000.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2919.960 4.000 2920.560 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2025.010 2996.000 2025.290 3000.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1467.490 2996.000 1467.770 3000.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 987.400 2300.000 988.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1165.560 4.000 1166.160 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.530 2996.000 995.810 3000.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2096.770 2996.000 2097.050 3000.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1568.120 4.000 1568.720 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 500.520 2300.000 501.120 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2170.600 2300.000 2171.200 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 952.290 2996.000 952.570 3000.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.770 2996.000 510.050 3000.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2150.200 2300.000 2150.800 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.210 0.000 1804.490 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.570 2996.000 1052.850 3000.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2061.810 0.000 2062.090 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1283.880 2300.000 1284.480 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.730 2996.000 867.010 3000.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.970 0.000 1347.250 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1561.330 0.000 1561.610 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1889.770 0.000 1890.050 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 2996.000 108.930 3000.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.690 0.000 1131.970 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.720 4.000 1378.320 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2053.530 2996.000 2053.810 3000.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2039.730 2996.000 2040.010 3000.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2282.610 2996.000 2282.890 3000.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1753.610 2996.000 1753.890 3000.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.330 0.000 917.610 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 2996.000 51.890 3000.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2095.800 4.000 2096.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.850 2996.000 1153.130 3000.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2023.720 2300.000 2024.320 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2065.880 2300.000 2066.480 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2963.480 4.000 2964.080 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 606.600 2300.000 607.200 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 712.680 2300.000 713.280 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1961.530 0.000 1961.810 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1791.160 2300.000 1791.760 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.330 0.000 1032.610 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.570 0.000 1489.850 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1947.560 4.000 1948.160 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2147.370 0.000 2147.650 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1167.570 2996.000 1167.850 3000.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.130 2996.000 724.410 3000.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1882.410 2996.000 1882.690 3000.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1672.840 4.000 1673.440 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.930 2996.000 853.210 3000.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2219.130 0.000 2219.410 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1335.560 4.000 1336.160 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 183.640 2300.000 184.240 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1260.490 0.000 1260.770 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2983.880 4.000 2984.480 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2225.570 2996.000 2225.850 3000.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1924.730 2996.000 1925.010 3000.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.210 2996.000 309.490 3000.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.570 2996.000 638.850 3000.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1621.160 2300.000 1621.760 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1646.890 0.000 1647.170 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1875.970 0.000 1876.250 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1863.240 4.000 1863.840 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 495.050 2996.000 495.330 3000.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.160 4.000 1927.760 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2593.560 2300.000 2594.160 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 695.610 2996.000 695.890 3000.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2877.800 4.000 2878.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.290 2996.000 538.570 3000.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1710.370 2996.000 1710.650 3000.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1367.210 2996.000 1367.490 3000.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 2996.000 209.210 3000.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1504.290 0.000 1504.570 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2294.480 2986.645 ;
      LAYER met1 ;
        RECT 5.520 4.460 2294.480 2992.300 ;
      LAYER met2 ;
        RECT 6.080 2995.720 9.010 2996.000 ;
        RECT 9.850 2995.720 22.810 2996.000 ;
        RECT 23.650 2995.720 37.530 2996.000 ;
        RECT 38.370 2995.720 51.330 2996.000 ;
        RECT 52.170 2995.720 66.050 2996.000 ;
        RECT 66.890 2995.720 79.850 2996.000 ;
        RECT 80.690 2995.720 94.570 2996.000 ;
        RECT 95.410 2995.720 108.370 2996.000 ;
        RECT 109.210 2995.720 123.090 2996.000 ;
        RECT 123.930 2995.720 136.890 2996.000 ;
        RECT 137.730 2995.720 151.610 2996.000 ;
        RECT 152.450 2995.720 166.330 2996.000 ;
        RECT 167.170 2995.720 180.130 2996.000 ;
        RECT 180.970 2995.720 194.850 2996.000 ;
        RECT 195.690 2995.720 208.650 2996.000 ;
        RECT 209.490 2995.720 223.370 2996.000 ;
        RECT 224.210 2995.720 237.170 2996.000 ;
        RECT 238.010 2995.720 251.890 2996.000 ;
        RECT 252.730 2995.720 265.690 2996.000 ;
        RECT 266.530 2995.720 280.410 2996.000 ;
        RECT 281.250 2995.720 294.210 2996.000 ;
        RECT 295.050 2995.720 308.930 2996.000 ;
        RECT 309.770 2995.720 323.650 2996.000 ;
        RECT 324.490 2995.720 337.450 2996.000 ;
        RECT 338.290 2995.720 352.170 2996.000 ;
        RECT 353.010 2995.720 365.970 2996.000 ;
        RECT 366.810 2995.720 380.690 2996.000 ;
        RECT 381.530 2995.720 394.490 2996.000 ;
        RECT 395.330 2995.720 409.210 2996.000 ;
        RECT 410.050 2995.720 423.010 2996.000 ;
        RECT 423.850 2995.720 437.730 2996.000 ;
        RECT 438.570 2995.720 451.530 2996.000 ;
        RECT 452.370 2995.720 466.250 2996.000 ;
        RECT 467.090 2995.720 480.970 2996.000 ;
        RECT 481.810 2995.720 494.770 2996.000 ;
        RECT 495.610 2995.720 509.490 2996.000 ;
        RECT 510.330 2995.720 523.290 2996.000 ;
        RECT 524.130 2995.720 538.010 2996.000 ;
        RECT 538.850 2995.720 551.810 2996.000 ;
        RECT 552.650 2995.720 566.530 2996.000 ;
        RECT 567.370 2995.720 580.330 2996.000 ;
        RECT 581.170 2995.720 595.050 2996.000 ;
        RECT 595.890 2995.720 608.850 2996.000 ;
        RECT 609.690 2995.720 623.570 2996.000 ;
        RECT 624.410 2995.720 638.290 2996.000 ;
        RECT 639.130 2995.720 652.090 2996.000 ;
        RECT 652.930 2995.720 666.810 2996.000 ;
        RECT 667.650 2995.720 680.610 2996.000 ;
        RECT 681.450 2995.720 695.330 2996.000 ;
        RECT 696.170 2995.720 709.130 2996.000 ;
        RECT 709.970 2995.720 723.850 2996.000 ;
        RECT 724.690 2995.720 737.650 2996.000 ;
        RECT 738.490 2995.720 752.370 2996.000 ;
        RECT 753.210 2995.720 766.170 2996.000 ;
        RECT 767.010 2995.720 780.890 2996.000 ;
        RECT 781.730 2995.720 794.690 2996.000 ;
        RECT 795.530 2995.720 809.410 2996.000 ;
        RECT 810.250 2995.720 824.130 2996.000 ;
        RECT 824.970 2995.720 837.930 2996.000 ;
        RECT 838.770 2995.720 852.650 2996.000 ;
        RECT 853.490 2995.720 866.450 2996.000 ;
        RECT 867.290 2995.720 881.170 2996.000 ;
        RECT 882.010 2995.720 894.970 2996.000 ;
        RECT 895.810 2995.720 909.690 2996.000 ;
        RECT 910.530 2995.720 923.490 2996.000 ;
        RECT 924.330 2995.720 938.210 2996.000 ;
        RECT 939.050 2995.720 952.010 2996.000 ;
        RECT 952.850 2995.720 966.730 2996.000 ;
        RECT 967.570 2995.720 981.450 2996.000 ;
        RECT 982.290 2995.720 995.250 2996.000 ;
        RECT 996.090 2995.720 1009.970 2996.000 ;
        RECT 1010.810 2995.720 1023.770 2996.000 ;
        RECT 1024.610 2995.720 1038.490 2996.000 ;
        RECT 1039.330 2995.720 1052.290 2996.000 ;
        RECT 1053.130 2995.720 1067.010 2996.000 ;
        RECT 1067.850 2995.720 1080.810 2996.000 ;
        RECT 1081.650 2995.720 1095.530 2996.000 ;
        RECT 1096.370 2995.720 1109.330 2996.000 ;
        RECT 1110.170 2995.720 1124.050 2996.000 ;
        RECT 1124.890 2995.720 1138.770 2996.000 ;
        RECT 1139.610 2995.720 1152.570 2996.000 ;
        RECT 1153.410 2995.720 1167.290 2996.000 ;
        RECT 1168.130 2995.720 1181.090 2996.000 ;
        RECT 1181.930 2995.720 1195.810 2996.000 ;
        RECT 1196.650 2995.720 1209.610 2996.000 ;
        RECT 1210.450 2995.720 1224.330 2996.000 ;
        RECT 1225.170 2995.720 1238.130 2996.000 ;
        RECT 1238.970 2995.720 1252.850 2996.000 ;
        RECT 1253.690 2995.720 1266.650 2996.000 ;
        RECT 1267.490 2995.720 1281.370 2996.000 ;
        RECT 1282.210 2995.720 1295.170 2996.000 ;
        RECT 1296.010 2995.720 1309.890 2996.000 ;
        RECT 1310.730 2995.720 1324.610 2996.000 ;
        RECT 1325.450 2995.720 1338.410 2996.000 ;
        RECT 1339.250 2995.720 1353.130 2996.000 ;
        RECT 1353.970 2995.720 1366.930 2996.000 ;
        RECT 1367.770 2995.720 1381.650 2996.000 ;
        RECT 1382.490 2995.720 1395.450 2996.000 ;
        RECT 1396.290 2995.720 1410.170 2996.000 ;
        RECT 1411.010 2995.720 1423.970 2996.000 ;
        RECT 1424.810 2995.720 1438.690 2996.000 ;
        RECT 1439.530 2995.720 1452.490 2996.000 ;
        RECT 1453.330 2995.720 1467.210 2996.000 ;
        RECT 1468.050 2995.720 1481.930 2996.000 ;
        RECT 1482.770 2995.720 1495.730 2996.000 ;
        RECT 1496.570 2995.720 1510.450 2996.000 ;
        RECT 1511.290 2995.720 1524.250 2996.000 ;
        RECT 1525.090 2995.720 1538.970 2996.000 ;
        RECT 1539.810 2995.720 1552.770 2996.000 ;
        RECT 1553.610 2995.720 1567.490 2996.000 ;
        RECT 1568.330 2995.720 1581.290 2996.000 ;
        RECT 1582.130 2995.720 1596.010 2996.000 ;
        RECT 1596.850 2995.720 1609.810 2996.000 ;
        RECT 1610.650 2995.720 1624.530 2996.000 ;
        RECT 1625.370 2995.720 1639.250 2996.000 ;
        RECT 1640.090 2995.720 1653.050 2996.000 ;
        RECT 1653.890 2995.720 1667.770 2996.000 ;
        RECT 1668.610 2995.720 1681.570 2996.000 ;
        RECT 1682.410 2995.720 1696.290 2996.000 ;
        RECT 1697.130 2995.720 1710.090 2996.000 ;
        RECT 1710.930 2995.720 1724.810 2996.000 ;
        RECT 1725.650 2995.720 1738.610 2996.000 ;
        RECT 1739.450 2995.720 1753.330 2996.000 ;
        RECT 1754.170 2995.720 1767.130 2996.000 ;
        RECT 1767.970 2995.720 1781.850 2996.000 ;
        RECT 1782.690 2995.720 1795.650 2996.000 ;
        RECT 1796.490 2995.720 1810.370 2996.000 ;
        RECT 1811.210 2995.720 1825.090 2996.000 ;
        RECT 1825.930 2995.720 1838.890 2996.000 ;
        RECT 1839.730 2995.720 1853.610 2996.000 ;
        RECT 1854.450 2995.720 1867.410 2996.000 ;
        RECT 1868.250 2995.720 1882.130 2996.000 ;
        RECT 1882.970 2995.720 1895.930 2996.000 ;
        RECT 1896.770 2995.720 1910.650 2996.000 ;
        RECT 1911.490 2995.720 1924.450 2996.000 ;
        RECT 1925.290 2995.720 1939.170 2996.000 ;
        RECT 1940.010 2995.720 1952.970 2996.000 ;
        RECT 1953.810 2995.720 1967.690 2996.000 ;
        RECT 1968.530 2995.720 1982.410 2996.000 ;
        RECT 1983.250 2995.720 1996.210 2996.000 ;
        RECT 1997.050 2995.720 2010.930 2996.000 ;
        RECT 2011.770 2995.720 2024.730 2996.000 ;
        RECT 2025.570 2995.720 2039.450 2996.000 ;
        RECT 2040.290 2995.720 2053.250 2996.000 ;
        RECT 2054.090 2995.720 2067.970 2996.000 ;
        RECT 2068.810 2995.720 2081.770 2996.000 ;
        RECT 2082.610 2995.720 2096.490 2996.000 ;
        RECT 2097.330 2995.720 2110.290 2996.000 ;
        RECT 2111.130 2995.720 2125.010 2996.000 ;
        RECT 2125.850 2995.720 2139.730 2996.000 ;
        RECT 2140.570 2995.720 2153.530 2996.000 ;
        RECT 2154.370 2995.720 2168.250 2996.000 ;
        RECT 2169.090 2995.720 2182.050 2996.000 ;
        RECT 2182.890 2995.720 2196.770 2996.000 ;
        RECT 2197.610 2995.720 2210.570 2996.000 ;
        RECT 2211.410 2995.720 2225.290 2996.000 ;
        RECT 2226.130 2995.720 2239.090 2996.000 ;
        RECT 2239.930 2995.720 2253.810 2996.000 ;
        RECT 2254.650 2995.720 2267.610 2996.000 ;
        RECT 2268.450 2995.720 2282.330 2996.000 ;
        RECT 2283.170 2995.720 2296.130 2996.000 ;
        RECT 6.080 4.280 2296.620 2995.720 ;
        RECT 6.080 4.000 16.370 4.280 ;
        RECT 17.210 4.000 31.090 4.280 ;
        RECT 31.930 4.000 44.890 4.280 ;
        RECT 45.730 4.000 59.610 4.280 ;
        RECT 60.450 4.000 73.410 4.280 ;
        RECT 74.250 4.000 88.130 4.280 ;
        RECT 88.970 4.000 101.930 4.280 ;
        RECT 102.770 4.000 116.650 4.280 ;
        RECT 117.490 4.000 130.450 4.280 ;
        RECT 131.290 4.000 145.170 4.280 ;
        RECT 146.010 4.000 158.970 4.280 ;
        RECT 159.810 4.000 173.690 4.280 ;
        RECT 174.530 4.000 188.410 4.280 ;
        RECT 189.250 4.000 202.210 4.280 ;
        RECT 203.050 4.000 216.930 4.280 ;
        RECT 217.770 4.000 230.730 4.280 ;
        RECT 231.570 4.000 245.450 4.280 ;
        RECT 246.290 4.000 259.250 4.280 ;
        RECT 260.090 4.000 273.970 4.280 ;
        RECT 274.810 4.000 287.770 4.280 ;
        RECT 288.610 4.000 302.490 4.280 ;
        RECT 303.330 4.000 316.290 4.280 ;
        RECT 317.130 4.000 331.010 4.280 ;
        RECT 331.850 4.000 345.730 4.280 ;
        RECT 346.570 4.000 359.530 4.280 ;
        RECT 360.370 4.000 374.250 4.280 ;
        RECT 375.090 4.000 388.050 4.280 ;
        RECT 388.890 4.000 402.770 4.280 ;
        RECT 403.610 4.000 416.570 4.280 ;
        RECT 417.410 4.000 431.290 4.280 ;
        RECT 432.130 4.000 445.090 4.280 ;
        RECT 445.930 4.000 459.810 4.280 ;
        RECT 460.650 4.000 473.610 4.280 ;
        RECT 474.450 4.000 488.330 4.280 ;
        RECT 489.170 4.000 503.050 4.280 ;
        RECT 503.890 4.000 516.850 4.280 ;
        RECT 517.690 4.000 531.570 4.280 ;
        RECT 532.410 4.000 545.370 4.280 ;
        RECT 546.210 4.000 560.090 4.280 ;
        RECT 560.930 4.000 573.890 4.280 ;
        RECT 574.730 4.000 588.610 4.280 ;
        RECT 589.450 4.000 602.410 4.280 ;
        RECT 603.250 4.000 617.130 4.280 ;
        RECT 617.970 4.000 630.930 4.280 ;
        RECT 631.770 4.000 645.650 4.280 ;
        RECT 646.490 4.000 659.450 4.280 ;
        RECT 660.290 4.000 674.170 4.280 ;
        RECT 675.010 4.000 688.890 4.280 ;
        RECT 689.730 4.000 702.690 4.280 ;
        RECT 703.530 4.000 717.410 4.280 ;
        RECT 718.250 4.000 731.210 4.280 ;
        RECT 732.050 4.000 745.930 4.280 ;
        RECT 746.770 4.000 759.730 4.280 ;
        RECT 760.570 4.000 774.450 4.280 ;
        RECT 775.290 4.000 788.250 4.280 ;
        RECT 789.090 4.000 802.970 4.280 ;
        RECT 803.810 4.000 816.770 4.280 ;
        RECT 817.610 4.000 831.490 4.280 ;
        RECT 832.330 4.000 846.210 4.280 ;
        RECT 847.050 4.000 860.010 4.280 ;
        RECT 860.850 4.000 874.730 4.280 ;
        RECT 875.570 4.000 888.530 4.280 ;
        RECT 889.370 4.000 903.250 4.280 ;
        RECT 904.090 4.000 917.050 4.280 ;
        RECT 917.890 4.000 931.770 4.280 ;
        RECT 932.610 4.000 945.570 4.280 ;
        RECT 946.410 4.000 960.290 4.280 ;
        RECT 961.130 4.000 974.090 4.280 ;
        RECT 974.930 4.000 988.810 4.280 ;
        RECT 989.650 4.000 1003.530 4.280 ;
        RECT 1004.370 4.000 1017.330 4.280 ;
        RECT 1018.170 4.000 1032.050 4.280 ;
        RECT 1032.890 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1060.570 4.280 ;
        RECT 1061.410 4.000 1074.370 4.280 ;
        RECT 1075.210 4.000 1089.090 4.280 ;
        RECT 1089.930 4.000 1102.890 4.280 ;
        RECT 1103.730 4.000 1117.610 4.280 ;
        RECT 1118.450 4.000 1131.410 4.280 ;
        RECT 1132.250 4.000 1146.130 4.280 ;
        RECT 1146.970 4.000 1159.930 4.280 ;
        RECT 1160.770 4.000 1174.650 4.280 ;
        RECT 1175.490 4.000 1189.370 4.280 ;
        RECT 1190.210 4.000 1203.170 4.280 ;
        RECT 1204.010 4.000 1217.890 4.280 ;
        RECT 1218.730 4.000 1231.690 4.280 ;
        RECT 1232.530 4.000 1246.410 4.280 ;
        RECT 1247.250 4.000 1260.210 4.280 ;
        RECT 1261.050 4.000 1274.930 4.280 ;
        RECT 1275.770 4.000 1288.730 4.280 ;
        RECT 1289.570 4.000 1303.450 4.280 ;
        RECT 1304.290 4.000 1317.250 4.280 ;
        RECT 1318.090 4.000 1331.970 4.280 ;
        RECT 1332.810 4.000 1346.690 4.280 ;
        RECT 1347.530 4.000 1360.490 4.280 ;
        RECT 1361.330 4.000 1375.210 4.280 ;
        RECT 1376.050 4.000 1389.010 4.280 ;
        RECT 1389.850 4.000 1403.730 4.280 ;
        RECT 1404.570 4.000 1417.530 4.280 ;
        RECT 1418.370 4.000 1432.250 4.280 ;
        RECT 1433.090 4.000 1446.050 4.280 ;
        RECT 1446.890 4.000 1460.770 4.280 ;
        RECT 1461.610 4.000 1474.570 4.280 ;
        RECT 1475.410 4.000 1489.290 4.280 ;
        RECT 1490.130 4.000 1504.010 4.280 ;
        RECT 1504.850 4.000 1517.810 4.280 ;
        RECT 1518.650 4.000 1532.530 4.280 ;
        RECT 1533.370 4.000 1546.330 4.280 ;
        RECT 1547.170 4.000 1561.050 4.280 ;
        RECT 1561.890 4.000 1574.850 4.280 ;
        RECT 1575.690 4.000 1589.570 4.280 ;
        RECT 1590.410 4.000 1603.370 4.280 ;
        RECT 1604.210 4.000 1618.090 4.280 ;
        RECT 1618.930 4.000 1631.890 4.280 ;
        RECT 1632.730 4.000 1646.610 4.280 ;
        RECT 1647.450 4.000 1660.410 4.280 ;
        RECT 1661.250 4.000 1675.130 4.280 ;
        RECT 1675.970 4.000 1689.850 4.280 ;
        RECT 1690.690 4.000 1703.650 4.280 ;
        RECT 1704.490 4.000 1718.370 4.280 ;
        RECT 1719.210 4.000 1732.170 4.280 ;
        RECT 1733.010 4.000 1746.890 4.280 ;
        RECT 1747.730 4.000 1760.690 4.280 ;
        RECT 1761.530 4.000 1775.410 4.280 ;
        RECT 1776.250 4.000 1789.210 4.280 ;
        RECT 1790.050 4.000 1803.930 4.280 ;
        RECT 1804.770 4.000 1817.730 4.280 ;
        RECT 1818.570 4.000 1832.450 4.280 ;
        RECT 1833.290 4.000 1847.170 4.280 ;
        RECT 1848.010 4.000 1860.970 4.280 ;
        RECT 1861.810 4.000 1875.690 4.280 ;
        RECT 1876.530 4.000 1889.490 4.280 ;
        RECT 1890.330 4.000 1904.210 4.280 ;
        RECT 1905.050 4.000 1918.010 4.280 ;
        RECT 1918.850 4.000 1932.730 4.280 ;
        RECT 1933.570 4.000 1946.530 4.280 ;
        RECT 1947.370 4.000 1961.250 4.280 ;
        RECT 1962.090 4.000 1975.050 4.280 ;
        RECT 1975.890 4.000 1989.770 4.280 ;
        RECT 1990.610 4.000 2004.490 4.280 ;
        RECT 2005.330 4.000 2018.290 4.280 ;
        RECT 2019.130 4.000 2033.010 4.280 ;
        RECT 2033.850 4.000 2046.810 4.280 ;
        RECT 2047.650 4.000 2061.530 4.280 ;
        RECT 2062.370 4.000 2075.330 4.280 ;
        RECT 2076.170 4.000 2090.050 4.280 ;
        RECT 2090.890 4.000 2103.850 4.280 ;
        RECT 2104.690 4.000 2118.570 4.280 ;
        RECT 2119.410 4.000 2132.370 4.280 ;
        RECT 2133.210 4.000 2147.090 4.280 ;
        RECT 2147.930 4.000 2161.810 4.280 ;
        RECT 2162.650 4.000 2175.610 4.280 ;
        RECT 2176.450 4.000 2190.330 4.280 ;
        RECT 2191.170 4.000 2204.130 4.280 ;
        RECT 2204.970 4.000 2218.850 4.280 ;
        RECT 2219.690 4.000 2232.650 4.280 ;
        RECT 2233.490 4.000 2247.370 4.280 ;
        RECT 2248.210 4.000 2261.170 4.280 ;
        RECT 2262.010 4.000 2275.890 4.280 ;
        RECT 2276.730 4.000 2289.690 4.280 ;
        RECT 2290.530 4.000 2296.620 4.280 ;
      LAYER met3 ;
        RECT 4.000 2984.880 2296.000 2987.745 ;
        RECT 4.400 2983.480 2296.000 2984.880 ;
        RECT 4.000 2975.360 2296.000 2983.480 ;
        RECT 4.000 2973.960 2295.600 2975.360 ;
        RECT 4.000 2964.480 2296.000 2973.960 ;
        RECT 4.400 2963.080 2296.000 2964.480 ;
        RECT 4.000 2953.600 2296.000 2963.080 ;
        RECT 4.000 2952.200 2295.600 2953.600 ;
        RECT 4.000 2942.720 2296.000 2952.200 ;
        RECT 4.400 2941.320 2296.000 2942.720 ;
        RECT 4.000 2933.200 2296.000 2941.320 ;
        RECT 4.000 2931.800 2295.600 2933.200 ;
        RECT 4.000 2920.960 2296.000 2931.800 ;
        RECT 4.400 2919.560 2296.000 2920.960 ;
        RECT 4.000 2911.440 2296.000 2919.560 ;
        RECT 4.000 2910.040 2295.600 2911.440 ;
        RECT 4.000 2900.560 2296.000 2910.040 ;
        RECT 4.400 2899.160 2296.000 2900.560 ;
        RECT 4.000 2891.040 2296.000 2899.160 ;
        RECT 4.000 2889.640 2295.600 2891.040 ;
        RECT 4.000 2878.800 2296.000 2889.640 ;
        RECT 4.400 2877.400 2296.000 2878.800 ;
        RECT 4.000 2869.280 2296.000 2877.400 ;
        RECT 4.000 2867.880 2295.600 2869.280 ;
        RECT 4.000 2858.400 2296.000 2867.880 ;
        RECT 4.400 2857.000 2296.000 2858.400 ;
        RECT 4.000 2848.880 2296.000 2857.000 ;
        RECT 4.000 2847.480 2295.600 2848.880 ;
        RECT 4.000 2836.640 2296.000 2847.480 ;
        RECT 4.400 2835.240 2296.000 2836.640 ;
        RECT 4.000 2827.120 2296.000 2835.240 ;
        RECT 4.000 2825.720 2295.600 2827.120 ;
        RECT 4.000 2816.240 2296.000 2825.720 ;
        RECT 4.400 2814.840 2296.000 2816.240 ;
        RECT 4.000 2806.720 2296.000 2814.840 ;
        RECT 4.000 2805.320 2295.600 2806.720 ;
        RECT 4.000 2794.480 2296.000 2805.320 ;
        RECT 4.400 2793.080 2296.000 2794.480 ;
        RECT 4.000 2784.960 2296.000 2793.080 ;
        RECT 4.000 2783.560 2295.600 2784.960 ;
        RECT 4.000 2774.080 2296.000 2783.560 ;
        RECT 4.400 2772.680 2296.000 2774.080 ;
        RECT 4.000 2764.560 2296.000 2772.680 ;
        RECT 4.000 2763.160 2295.600 2764.560 ;
        RECT 4.000 2752.320 2296.000 2763.160 ;
        RECT 4.400 2750.920 2296.000 2752.320 ;
        RECT 4.000 2742.800 2296.000 2750.920 ;
        RECT 4.000 2741.400 2295.600 2742.800 ;
        RECT 4.000 2731.920 2296.000 2741.400 ;
        RECT 4.400 2730.520 2296.000 2731.920 ;
        RECT 4.000 2721.040 2296.000 2730.520 ;
        RECT 4.000 2719.640 2295.600 2721.040 ;
        RECT 4.000 2710.160 2296.000 2719.640 ;
        RECT 4.400 2708.760 2296.000 2710.160 ;
        RECT 4.000 2700.640 2296.000 2708.760 ;
        RECT 4.000 2699.240 2295.600 2700.640 ;
        RECT 4.000 2688.400 2296.000 2699.240 ;
        RECT 4.400 2687.000 2296.000 2688.400 ;
        RECT 4.000 2678.880 2296.000 2687.000 ;
        RECT 4.000 2677.480 2295.600 2678.880 ;
        RECT 4.000 2668.000 2296.000 2677.480 ;
        RECT 4.400 2666.600 2296.000 2668.000 ;
        RECT 4.000 2658.480 2296.000 2666.600 ;
        RECT 4.000 2657.080 2295.600 2658.480 ;
        RECT 4.000 2646.240 2296.000 2657.080 ;
        RECT 4.400 2644.840 2296.000 2646.240 ;
        RECT 4.000 2636.720 2296.000 2644.840 ;
        RECT 4.000 2635.320 2295.600 2636.720 ;
        RECT 4.000 2625.840 2296.000 2635.320 ;
        RECT 4.400 2624.440 2296.000 2625.840 ;
        RECT 4.000 2616.320 2296.000 2624.440 ;
        RECT 4.000 2614.920 2295.600 2616.320 ;
        RECT 4.000 2604.080 2296.000 2614.920 ;
        RECT 4.400 2602.680 2296.000 2604.080 ;
        RECT 4.000 2594.560 2296.000 2602.680 ;
        RECT 4.000 2593.160 2295.600 2594.560 ;
        RECT 4.000 2583.680 2296.000 2593.160 ;
        RECT 4.400 2582.280 2296.000 2583.680 ;
        RECT 4.000 2574.160 2296.000 2582.280 ;
        RECT 4.000 2572.760 2295.600 2574.160 ;
        RECT 4.000 2561.920 2296.000 2572.760 ;
        RECT 4.400 2560.520 2296.000 2561.920 ;
        RECT 4.000 2552.400 2296.000 2560.520 ;
        RECT 4.000 2551.000 2295.600 2552.400 ;
        RECT 4.000 2541.520 2296.000 2551.000 ;
        RECT 4.400 2540.120 2296.000 2541.520 ;
        RECT 4.000 2532.000 2296.000 2540.120 ;
        RECT 4.000 2530.600 2295.600 2532.000 ;
        RECT 4.000 2519.760 2296.000 2530.600 ;
        RECT 4.400 2518.360 2296.000 2519.760 ;
        RECT 4.000 2510.240 2296.000 2518.360 ;
        RECT 4.000 2508.840 2295.600 2510.240 ;
        RECT 4.000 2499.360 2296.000 2508.840 ;
        RECT 4.400 2497.960 2296.000 2499.360 ;
        RECT 4.000 2488.480 2296.000 2497.960 ;
        RECT 4.000 2487.080 2295.600 2488.480 ;
        RECT 4.000 2477.600 2296.000 2487.080 ;
        RECT 4.400 2476.200 2296.000 2477.600 ;
        RECT 4.000 2468.080 2296.000 2476.200 ;
        RECT 4.000 2466.680 2295.600 2468.080 ;
        RECT 4.000 2455.840 2296.000 2466.680 ;
        RECT 4.400 2454.440 2296.000 2455.840 ;
        RECT 4.000 2446.320 2296.000 2454.440 ;
        RECT 4.000 2444.920 2295.600 2446.320 ;
        RECT 4.000 2435.440 2296.000 2444.920 ;
        RECT 4.400 2434.040 2296.000 2435.440 ;
        RECT 4.000 2425.920 2296.000 2434.040 ;
        RECT 4.000 2424.520 2295.600 2425.920 ;
        RECT 4.000 2413.680 2296.000 2424.520 ;
        RECT 4.400 2412.280 2296.000 2413.680 ;
        RECT 4.000 2404.160 2296.000 2412.280 ;
        RECT 4.000 2402.760 2295.600 2404.160 ;
        RECT 4.000 2393.280 2296.000 2402.760 ;
        RECT 4.400 2391.880 2296.000 2393.280 ;
        RECT 4.000 2383.760 2296.000 2391.880 ;
        RECT 4.000 2382.360 2295.600 2383.760 ;
        RECT 4.000 2371.520 2296.000 2382.360 ;
        RECT 4.400 2370.120 2296.000 2371.520 ;
        RECT 4.000 2362.000 2296.000 2370.120 ;
        RECT 4.000 2360.600 2295.600 2362.000 ;
        RECT 4.000 2351.120 2296.000 2360.600 ;
        RECT 4.400 2349.720 2296.000 2351.120 ;
        RECT 4.000 2341.600 2296.000 2349.720 ;
        RECT 4.000 2340.200 2295.600 2341.600 ;
        RECT 4.000 2329.360 2296.000 2340.200 ;
        RECT 4.400 2327.960 2296.000 2329.360 ;
        RECT 4.000 2319.840 2296.000 2327.960 ;
        RECT 4.000 2318.440 2295.600 2319.840 ;
        RECT 4.000 2308.960 2296.000 2318.440 ;
        RECT 4.400 2307.560 2296.000 2308.960 ;
        RECT 4.000 2299.440 2296.000 2307.560 ;
        RECT 4.000 2298.040 2295.600 2299.440 ;
        RECT 4.000 2287.200 2296.000 2298.040 ;
        RECT 4.400 2285.800 2296.000 2287.200 ;
        RECT 4.000 2277.680 2296.000 2285.800 ;
        RECT 4.000 2276.280 2295.600 2277.680 ;
        RECT 4.000 2266.800 2296.000 2276.280 ;
        RECT 4.400 2265.400 2296.000 2266.800 ;
        RECT 4.000 2255.920 2296.000 2265.400 ;
        RECT 4.000 2254.520 2295.600 2255.920 ;
        RECT 4.000 2245.040 2296.000 2254.520 ;
        RECT 4.400 2243.640 2296.000 2245.040 ;
        RECT 4.000 2235.520 2296.000 2243.640 ;
        RECT 4.000 2234.120 2295.600 2235.520 ;
        RECT 4.000 2224.640 2296.000 2234.120 ;
        RECT 4.400 2223.240 2296.000 2224.640 ;
        RECT 4.000 2213.760 2296.000 2223.240 ;
        RECT 4.000 2212.360 2295.600 2213.760 ;
        RECT 4.000 2202.880 2296.000 2212.360 ;
        RECT 4.400 2201.480 2296.000 2202.880 ;
        RECT 4.000 2193.360 2296.000 2201.480 ;
        RECT 4.000 2191.960 2295.600 2193.360 ;
        RECT 4.000 2181.120 2296.000 2191.960 ;
        RECT 4.400 2179.720 2296.000 2181.120 ;
        RECT 4.000 2171.600 2296.000 2179.720 ;
        RECT 4.000 2170.200 2295.600 2171.600 ;
        RECT 4.000 2160.720 2296.000 2170.200 ;
        RECT 4.400 2159.320 2296.000 2160.720 ;
        RECT 4.000 2151.200 2296.000 2159.320 ;
        RECT 4.000 2149.800 2295.600 2151.200 ;
        RECT 4.000 2138.960 2296.000 2149.800 ;
        RECT 4.400 2137.560 2296.000 2138.960 ;
        RECT 4.000 2129.440 2296.000 2137.560 ;
        RECT 4.000 2128.040 2295.600 2129.440 ;
        RECT 4.000 2118.560 2296.000 2128.040 ;
        RECT 4.400 2117.160 2296.000 2118.560 ;
        RECT 4.000 2109.040 2296.000 2117.160 ;
        RECT 4.000 2107.640 2295.600 2109.040 ;
        RECT 4.000 2096.800 2296.000 2107.640 ;
        RECT 4.400 2095.400 2296.000 2096.800 ;
        RECT 4.000 2087.280 2296.000 2095.400 ;
        RECT 4.000 2085.880 2295.600 2087.280 ;
        RECT 4.000 2076.400 2296.000 2085.880 ;
        RECT 4.400 2075.000 2296.000 2076.400 ;
        RECT 4.000 2066.880 2296.000 2075.000 ;
        RECT 4.000 2065.480 2295.600 2066.880 ;
        RECT 4.000 2054.640 2296.000 2065.480 ;
        RECT 4.400 2053.240 2296.000 2054.640 ;
        RECT 4.000 2045.120 2296.000 2053.240 ;
        RECT 4.000 2043.720 2295.600 2045.120 ;
        RECT 4.000 2034.240 2296.000 2043.720 ;
        RECT 4.400 2032.840 2296.000 2034.240 ;
        RECT 4.000 2024.720 2296.000 2032.840 ;
        RECT 4.000 2023.320 2295.600 2024.720 ;
        RECT 4.000 2012.480 2296.000 2023.320 ;
        RECT 4.400 2011.080 2296.000 2012.480 ;
        RECT 4.000 2002.960 2296.000 2011.080 ;
        RECT 4.000 2001.560 2295.600 2002.960 ;
        RECT 4.000 1992.080 2296.000 2001.560 ;
        RECT 4.400 1990.680 2296.000 1992.080 ;
        RECT 4.000 1981.200 2296.000 1990.680 ;
        RECT 4.000 1979.800 2295.600 1981.200 ;
        RECT 4.000 1970.320 2296.000 1979.800 ;
        RECT 4.400 1968.920 2296.000 1970.320 ;
        RECT 4.000 1960.800 2296.000 1968.920 ;
        RECT 4.000 1959.400 2295.600 1960.800 ;
        RECT 4.000 1948.560 2296.000 1959.400 ;
        RECT 4.400 1947.160 2296.000 1948.560 ;
        RECT 4.000 1939.040 2296.000 1947.160 ;
        RECT 4.000 1937.640 2295.600 1939.040 ;
        RECT 4.000 1928.160 2296.000 1937.640 ;
        RECT 4.400 1926.760 2296.000 1928.160 ;
        RECT 4.000 1918.640 2296.000 1926.760 ;
        RECT 4.000 1917.240 2295.600 1918.640 ;
        RECT 4.000 1906.400 2296.000 1917.240 ;
        RECT 4.400 1905.000 2296.000 1906.400 ;
        RECT 4.000 1896.880 2296.000 1905.000 ;
        RECT 4.000 1895.480 2295.600 1896.880 ;
        RECT 4.000 1886.000 2296.000 1895.480 ;
        RECT 4.400 1884.600 2296.000 1886.000 ;
        RECT 4.000 1876.480 2296.000 1884.600 ;
        RECT 4.000 1875.080 2295.600 1876.480 ;
        RECT 4.000 1864.240 2296.000 1875.080 ;
        RECT 4.400 1862.840 2296.000 1864.240 ;
        RECT 4.000 1854.720 2296.000 1862.840 ;
        RECT 4.000 1853.320 2295.600 1854.720 ;
        RECT 4.000 1843.840 2296.000 1853.320 ;
        RECT 4.400 1842.440 2296.000 1843.840 ;
        RECT 4.000 1834.320 2296.000 1842.440 ;
        RECT 4.000 1832.920 2295.600 1834.320 ;
        RECT 4.000 1822.080 2296.000 1832.920 ;
        RECT 4.400 1820.680 2296.000 1822.080 ;
        RECT 4.000 1812.560 2296.000 1820.680 ;
        RECT 4.000 1811.160 2295.600 1812.560 ;
        RECT 4.000 1801.680 2296.000 1811.160 ;
        RECT 4.400 1800.280 2296.000 1801.680 ;
        RECT 4.000 1792.160 2296.000 1800.280 ;
        RECT 4.000 1790.760 2295.600 1792.160 ;
        RECT 4.000 1779.920 2296.000 1790.760 ;
        RECT 4.400 1778.520 2296.000 1779.920 ;
        RECT 4.000 1770.400 2296.000 1778.520 ;
        RECT 4.000 1769.000 2295.600 1770.400 ;
        RECT 4.000 1759.520 2296.000 1769.000 ;
        RECT 4.400 1758.120 2296.000 1759.520 ;
        RECT 4.000 1748.640 2296.000 1758.120 ;
        RECT 4.000 1747.240 2295.600 1748.640 ;
        RECT 4.000 1737.760 2296.000 1747.240 ;
        RECT 4.400 1736.360 2296.000 1737.760 ;
        RECT 4.000 1728.240 2296.000 1736.360 ;
        RECT 4.000 1726.840 2295.600 1728.240 ;
        RECT 4.000 1716.000 2296.000 1726.840 ;
        RECT 4.400 1714.600 2296.000 1716.000 ;
        RECT 4.000 1706.480 2296.000 1714.600 ;
        RECT 4.000 1705.080 2295.600 1706.480 ;
        RECT 4.000 1695.600 2296.000 1705.080 ;
        RECT 4.400 1694.200 2296.000 1695.600 ;
        RECT 4.000 1686.080 2296.000 1694.200 ;
        RECT 4.000 1684.680 2295.600 1686.080 ;
        RECT 4.000 1673.840 2296.000 1684.680 ;
        RECT 4.400 1672.440 2296.000 1673.840 ;
        RECT 4.000 1664.320 2296.000 1672.440 ;
        RECT 4.000 1662.920 2295.600 1664.320 ;
        RECT 4.000 1653.440 2296.000 1662.920 ;
        RECT 4.400 1652.040 2296.000 1653.440 ;
        RECT 4.000 1643.920 2296.000 1652.040 ;
        RECT 4.000 1642.520 2295.600 1643.920 ;
        RECT 4.000 1631.680 2296.000 1642.520 ;
        RECT 4.400 1630.280 2296.000 1631.680 ;
        RECT 4.000 1622.160 2296.000 1630.280 ;
        RECT 4.000 1620.760 2295.600 1622.160 ;
        RECT 4.000 1611.280 2296.000 1620.760 ;
        RECT 4.400 1609.880 2296.000 1611.280 ;
        RECT 4.000 1601.760 2296.000 1609.880 ;
        RECT 4.000 1600.360 2295.600 1601.760 ;
        RECT 4.000 1589.520 2296.000 1600.360 ;
        RECT 4.400 1588.120 2296.000 1589.520 ;
        RECT 4.000 1580.000 2296.000 1588.120 ;
        RECT 4.000 1578.600 2295.600 1580.000 ;
        RECT 4.000 1569.120 2296.000 1578.600 ;
        RECT 4.400 1567.720 2296.000 1569.120 ;
        RECT 4.000 1559.600 2296.000 1567.720 ;
        RECT 4.000 1558.200 2295.600 1559.600 ;
        RECT 4.000 1547.360 2296.000 1558.200 ;
        RECT 4.400 1545.960 2296.000 1547.360 ;
        RECT 4.000 1537.840 2296.000 1545.960 ;
        RECT 4.000 1536.440 2295.600 1537.840 ;
        RECT 4.000 1526.960 2296.000 1536.440 ;
        RECT 4.400 1525.560 2296.000 1526.960 ;
        RECT 4.000 1516.080 2296.000 1525.560 ;
        RECT 4.000 1514.680 2295.600 1516.080 ;
        RECT 4.000 1505.200 2296.000 1514.680 ;
        RECT 4.400 1503.800 2296.000 1505.200 ;
        RECT 4.000 1495.680 2296.000 1503.800 ;
        RECT 4.000 1494.280 2295.600 1495.680 ;
        RECT 4.000 1484.800 2296.000 1494.280 ;
        RECT 4.400 1483.400 2296.000 1484.800 ;
        RECT 4.000 1473.920 2296.000 1483.400 ;
        RECT 4.000 1472.520 2295.600 1473.920 ;
        RECT 4.000 1463.040 2296.000 1472.520 ;
        RECT 4.400 1461.640 2296.000 1463.040 ;
        RECT 4.000 1453.520 2296.000 1461.640 ;
        RECT 4.000 1452.120 2295.600 1453.520 ;
        RECT 4.000 1441.280 2296.000 1452.120 ;
        RECT 4.400 1439.880 2296.000 1441.280 ;
        RECT 4.000 1431.760 2296.000 1439.880 ;
        RECT 4.000 1430.360 2295.600 1431.760 ;
        RECT 4.000 1420.880 2296.000 1430.360 ;
        RECT 4.400 1419.480 2296.000 1420.880 ;
        RECT 4.000 1411.360 2296.000 1419.480 ;
        RECT 4.000 1409.960 2295.600 1411.360 ;
        RECT 4.000 1399.120 2296.000 1409.960 ;
        RECT 4.400 1397.720 2296.000 1399.120 ;
        RECT 4.000 1389.600 2296.000 1397.720 ;
        RECT 4.000 1388.200 2295.600 1389.600 ;
        RECT 4.000 1378.720 2296.000 1388.200 ;
        RECT 4.400 1377.320 2296.000 1378.720 ;
        RECT 4.000 1369.200 2296.000 1377.320 ;
        RECT 4.000 1367.800 2295.600 1369.200 ;
        RECT 4.000 1356.960 2296.000 1367.800 ;
        RECT 4.400 1355.560 2296.000 1356.960 ;
        RECT 4.000 1347.440 2296.000 1355.560 ;
        RECT 4.000 1346.040 2295.600 1347.440 ;
        RECT 4.000 1336.560 2296.000 1346.040 ;
        RECT 4.400 1335.160 2296.000 1336.560 ;
        RECT 4.000 1327.040 2296.000 1335.160 ;
        RECT 4.000 1325.640 2295.600 1327.040 ;
        RECT 4.000 1314.800 2296.000 1325.640 ;
        RECT 4.400 1313.400 2296.000 1314.800 ;
        RECT 4.000 1305.280 2296.000 1313.400 ;
        RECT 4.000 1303.880 2295.600 1305.280 ;
        RECT 4.000 1294.400 2296.000 1303.880 ;
        RECT 4.400 1293.000 2296.000 1294.400 ;
        RECT 4.000 1284.880 2296.000 1293.000 ;
        RECT 4.000 1283.480 2295.600 1284.880 ;
        RECT 4.000 1272.640 2296.000 1283.480 ;
        RECT 4.400 1271.240 2296.000 1272.640 ;
        RECT 4.000 1263.120 2296.000 1271.240 ;
        RECT 4.000 1261.720 2295.600 1263.120 ;
        RECT 4.000 1252.240 2296.000 1261.720 ;
        RECT 4.400 1250.840 2296.000 1252.240 ;
        RECT 4.000 1241.360 2296.000 1250.840 ;
        RECT 4.000 1239.960 2295.600 1241.360 ;
        RECT 4.000 1230.480 2296.000 1239.960 ;
        RECT 4.400 1229.080 2296.000 1230.480 ;
        RECT 4.000 1220.960 2296.000 1229.080 ;
        RECT 4.000 1219.560 2295.600 1220.960 ;
        RECT 4.000 1208.720 2296.000 1219.560 ;
        RECT 4.400 1207.320 2296.000 1208.720 ;
        RECT 4.000 1199.200 2296.000 1207.320 ;
        RECT 4.000 1197.800 2295.600 1199.200 ;
        RECT 4.000 1188.320 2296.000 1197.800 ;
        RECT 4.400 1186.920 2296.000 1188.320 ;
        RECT 4.000 1178.800 2296.000 1186.920 ;
        RECT 4.000 1177.400 2295.600 1178.800 ;
        RECT 4.000 1166.560 2296.000 1177.400 ;
        RECT 4.400 1165.160 2296.000 1166.560 ;
        RECT 4.000 1157.040 2296.000 1165.160 ;
        RECT 4.000 1155.640 2295.600 1157.040 ;
        RECT 4.000 1146.160 2296.000 1155.640 ;
        RECT 4.400 1144.760 2296.000 1146.160 ;
        RECT 4.000 1136.640 2296.000 1144.760 ;
        RECT 4.000 1135.240 2295.600 1136.640 ;
        RECT 4.000 1124.400 2296.000 1135.240 ;
        RECT 4.400 1123.000 2296.000 1124.400 ;
        RECT 4.000 1114.880 2296.000 1123.000 ;
        RECT 4.000 1113.480 2295.600 1114.880 ;
        RECT 4.000 1104.000 2296.000 1113.480 ;
        RECT 4.400 1102.600 2296.000 1104.000 ;
        RECT 4.000 1094.480 2296.000 1102.600 ;
        RECT 4.000 1093.080 2295.600 1094.480 ;
        RECT 4.000 1082.240 2296.000 1093.080 ;
        RECT 4.400 1080.840 2296.000 1082.240 ;
        RECT 4.000 1072.720 2296.000 1080.840 ;
        RECT 4.000 1071.320 2295.600 1072.720 ;
        RECT 4.000 1061.840 2296.000 1071.320 ;
        RECT 4.400 1060.440 2296.000 1061.840 ;
        RECT 4.000 1052.320 2296.000 1060.440 ;
        RECT 4.000 1050.920 2295.600 1052.320 ;
        RECT 4.000 1040.080 2296.000 1050.920 ;
        RECT 4.400 1038.680 2296.000 1040.080 ;
        RECT 4.000 1030.560 2296.000 1038.680 ;
        RECT 4.000 1029.160 2295.600 1030.560 ;
        RECT 4.000 1019.680 2296.000 1029.160 ;
        RECT 4.400 1018.280 2296.000 1019.680 ;
        RECT 4.000 1008.800 2296.000 1018.280 ;
        RECT 4.000 1007.400 2295.600 1008.800 ;
        RECT 4.000 997.920 2296.000 1007.400 ;
        RECT 4.400 996.520 2296.000 997.920 ;
        RECT 4.000 988.400 2296.000 996.520 ;
        RECT 4.000 987.000 2295.600 988.400 ;
        RECT 4.000 976.160 2296.000 987.000 ;
        RECT 4.400 974.760 2296.000 976.160 ;
        RECT 4.000 966.640 2296.000 974.760 ;
        RECT 4.000 965.240 2295.600 966.640 ;
        RECT 4.000 955.760 2296.000 965.240 ;
        RECT 4.400 954.360 2296.000 955.760 ;
        RECT 4.000 946.240 2296.000 954.360 ;
        RECT 4.000 944.840 2295.600 946.240 ;
        RECT 4.000 934.000 2296.000 944.840 ;
        RECT 4.400 932.600 2296.000 934.000 ;
        RECT 4.000 924.480 2296.000 932.600 ;
        RECT 4.000 923.080 2295.600 924.480 ;
        RECT 4.000 913.600 2296.000 923.080 ;
        RECT 4.400 912.200 2296.000 913.600 ;
        RECT 4.000 904.080 2296.000 912.200 ;
        RECT 4.000 902.680 2295.600 904.080 ;
        RECT 4.000 891.840 2296.000 902.680 ;
        RECT 4.400 890.440 2296.000 891.840 ;
        RECT 4.000 882.320 2296.000 890.440 ;
        RECT 4.000 880.920 2295.600 882.320 ;
        RECT 4.000 871.440 2296.000 880.920 ;
        RECT 4.400 870.040 2296.000 871.440 ;
        RECT 4.000 861.920 2296.000 870.040 ;
        RECT 4.000 860.520 2295.600 861.920 ;
        RECT 4.000 849.680 2296.000 860.520 ;
        RECT 4.400 848.280 2296.000 849.680 ;
        RECT 4.000 840.160 2296.000 848.280 ;
        RECT 4.000 838.760 2295.600 840.160 ;
        RECT 4.000 829.280 2296.000 838.760 ;
        RECT 4.400 827.880 2296.000 829.280 ;
        RECT 4.000 819.760 2296.000 827.880 ;
        RECT 4.000 818.360 2295.600 819.760 ;
        RECT 4.000 807.520 2296.000 818.360 ;
        RECT 4.400 806.120 2296.000 807.520 ;
        RECT 4.000 798.000 2296.000 806.120 ;
        RECT 4.000 796.600 2295.600 798.000 ;
        RECT 4.000 787.120 2296.000 796.600 ;
        RECT 4.400 785.720 2296.000 787.120 ;
        RECT 4.000 776.240 2296.000 785.720 ;
        RECT 4.000 774.840 2295.600 776.240 ;
        RECT 4.000 765.360 2296.000 774.840 ;
        RECT 4.400 763.960 2296.000 765.360 ;
        RECT 4.000 755.840 2296.000 763.960 ;
        RECT 4.000 754.440 2295.600 755.840 ;
        RECT 4.000 744.960 2296.000 754.440 ;
        RECT 4.400 743.560 2296.000 744.960 ;
        RECT 4.000 734.080 2296.000 743.560 ;
        RECT 4.000 732.680 2295.600 734.080 ;
        RECT 4.000 723.200 2296.000 732.680 ;
        RECT 4.400 721.800 2296.000 723.200 ;
        RECT 4.000 713.680 2296.000 721.800 ;
        RECT 4.000 712.280 2295.600 713.680 ;
        RECT 4.000 701.440 2296.000 712.280 ;
        RECT 4.400 700.040 2296.000 701.440 ;
        RECT 4.000 691.920 2296.000 700.040 ;
        RECT 4.000 690.520 2295.600 691.920 ;
        RECT 4.000 681.040 2296.000 690.520 ;
        RECT 4.400 679.640 2296.000 681.040 ;
        RECT 4.000 671.520 2296.000 679.640 ;
        RECT 4.000 670.120 2295.600 671.520 ;
        RECT 4.000 659.280 2296.000 670.120 ;
        RECT 4.400 657.880 2296.000 659.280 ;
        RECT 4.000 649.760 2296.000 657.880 ;
        RECT 4.000 648.360 2295.600 649.760 ;
        RECT 4.000 638.880 2296.000 648.360 ;
        RECT 4.400 637.480 2296.000 638.880 ;
        RECT 4.000 629.360 2296.000 637.480 ;
        RECT 4.000 627.960 2295.600 629.360 ;
        RECT 4.000 617.120 2296.000 627.960 ;
        RECT 4.400 615.720 2296.000 617.120 ;
        RECT 4.000 607.600 2296.000 615.720 ;
        RECT 4.000 606.200 2295.600 607.600 ;
        RECT 4.000 596.720 2296.000 606.200 ;
        RECT 4.400 595.320 2296.000 596.720 ;
        RECT 4.000 587.200 2296.000 595.320 ;
        RECT 4.000 585.800 2295.600 587.200 ;
        RECT 4.000 574.960 2296.000 585.800 ;
        RECT 4.400 573.560 2296.000 574.960 ;
        RECT 4.000 565.440 2296.000 573.560 ;
        RECT 4.000 564.040 2295.600 565.440 ;
        RECT 4.000 554.560 2296.000 564.040 ;
        RECT 4.400 553.160 2296.000 554.560 ;
        RECT 4.000 545.040 2296.000 553.160 ;
        RECT 4.000 543.640 2295.600 545.040 ;
        RECT 4.000 532.800 2296.000 543.640 ;
        RECT 4.400 531.400 2296.000 532.800 ;
        RECT 4.000 523.280 2296.000 531.400 ;
        RECT 4.000 521.880 2295.600 523.280 ;
        RECT 4.000 512.400 2296.000 521.880 ;
        RECT 4.400 511.000 2296.000 512.400 ;
        RECT 4.000 501.520 2296.000 511.000 ;
        RECT 4.000 500.120 2295.600 501.520 ;
        RECT 4.000 490.640 2296.000 500.120 ;
        RECT 4.400 489.240 2296.000 490.640 ;
        RECT 4.000 481.120 2296.000 489.240 ;
        RECT 4.000 479.720 2295.600 481.120 ;
        RECT 4.000 468.880 2296.000 479.720 ;
        RECT 4.400 467.480 2296.000 468.880 ;
        RECT 4.000 459.360 2296.000 467.480 ;
        RECT 4.000 457.960 2295.600 459.360 ;
        RECT 4.000 448.480 2296.000 457.960 ;
        RECT 4.400 447.080 2296.000 448.480 ;
        RECT 4.000 438.960 2296.000 447.080 ;
        RECT 4.000 437.560 2295.600 438.960 ;
        RECT 4.000 426.720 2296.000 437.560 ;
        RECT 4.400 425.320 2296.000 426.720 ;
        RECT 4.000 417.200 2296.000 425.320 ;
        RECT 4.000 415.800 2295.600 417.200 ;
        RECT 4.000 406.320 2296.000 415.800 ;
        RECT 4.400 404.920 2296.000 406.320 ;
        RECT 4.000 396.800 2296.000 404.920 ;
        RECT 4.000 395.400 2295.600 396.800 ;
        RECT 4.000 384.560 2296.000 395.400 ;
        RECT 4.400 383.160 2296.000 384.560 ;
        RECT 4.000 375.040 2296.000 383.160 ;
        RECT 4.000 373.640 2295.600 375.040 ;
        RECT 4.000 364.160 2296.000 373.640 ;
        RECT 4.400 362.760 2296.000 364.160 ;
        RECT 4.000 354.640 2296.000 362.760 ;
        RECT 4.000 353.240 2295.600 354.640 ;
        RECT 4.000 342.400 2296.000 353.240 ;
        RECT 4.400 341.000 2296.000 342.400 ;
        RECT 4.000 332.880 2296.000 341.000 ;
        RECT 4.000 331.480 2295.600 332.880 ;
        RECT 4.000 322.000 2296.000 331.480 ;
        RECT 4.400 320.600 2296.000 322.000 ;
        RECT 4.000 312.480 2296.000 320.600 ;
        RECT 4.000 311.080 2295.600 312.480 ;
        RECT 4.000 300.240 2296.000 311.080 ;
        RECT 4.400 298.840 2296.000 300.240 ;
        RECT 4.000 290.720 2296.000 298.840 ;
        RECT 4.000 289.320 2295.600 290.720 ;
        RECT 4.000 279.840 2296.000 289.320 ;
        RECT 4.400 278.440 2296.000 279.840 ;
        RECT 4.000 268.960 2296.000 278.440 ;
        RECT 4.000 267.560 2295.600 268.960 ;
        RECT 4.000 258.080 2296.000 267.560 ;
        RECT 4.400 256.680 2296.000 258.080 ;
        RECT 4.000 248.560 2296.000 256.680 ;
        RECT 4.000 247.160 2295.600 248.560 ;
        RECT 4.000 236.320 2296.000 247.160 ;
        RECT 4.400 234.920 2296.000 236.320 ;
        RECT 4.000 226.800 2296.000 234.920 ;
        RECT 4.000 225.400 2295.600 226.800 ;
        RECT 4.000 215.920 2296.000 225.400 ;
        RECT 4.400 214.520 2296.000 215.920 ;
        RECT 4.000 206.400 2296.000 214.520 ;
        RECT 4.000 205.000 2295.600 206.400 ;
        RECT 4.000 194.160 2296.000 205.000 ;
        RECT 4.400 192.760 2296.000 194.160 ;
        RECT 4.000 184.640 2296.000 192.760 ;
        RECT 4.000 183.240 2295.600 184.640 ;
        RECT 4.000 173.760 2296.000 183.240 ;
        RECT 4.400 172.360 2296.000 173.760 ;
        RECT 4.000 164.240 2296.000 172.360 ;
        RECT 4.000 162.840 2295.600 164.240 ;
        RECT 4.000 152.000 2296.000 162.840 ;
        RECT 4.400 150.600 2296.000 152.000 ;
        RECT 4.000 142.480 2296.000 150.600 ;
        RECT 4.000 141.080 2295.600 142.480 ;
        RECT 4.000 131.600 2296.000 141.080 ;
        RECT 4.400 130.200 2296.000 131.600 ;
        RECT 4.000 122.080 2296.000 130.200 ;
        RECT 4.000 120.680 2295.600 122.080 ;
        RECT 4.000 109.840 2296.000 120.680 ;
        RECT 4.400 108.440 2296.000 109.840 ;
        RECT 4.000 100.320 2296.000 108.440 ;
        RECT 4.000 98.920 2295.600 100.320 ;
        RECT 4.000 89.440 2296.000 98.920 ;
        RECT 4.400 88.040 2296.000 89.440 ;
        RECT 4.000 79.920 2296.000 88.040 ;
        RECT 4.000 78.520 2295.600 79.920 ;
        RECT 4.000 67.680 2296.000 78.520 ;
        RECT 4.400 66.280 2296.000 67.680 ;
        RECT 4.000 58.160 2296.000 66.280 ;
        RECT 4.000 56.760 2295.600 58.160 ;
        RECT 4.000 47.280 2296.000 56.760 ;
        RECT 4.400 45.880 2296.000 47.280 ;
        RECT 4.000 36.400 2296.000 45.880 ;
        RECT 4.000 35.000 2295.600 36.400 ;
        RECT 4.000 25.520 2296.000 35.000 ;
        RECT 4.400 24.120 2296.000 25.520 ;
        RECT 4.000 16.000 2296.000 24.120 ;
        RECT 4.000 14.600 2295.600 16.000 ;
        RECT 4.000 4.255 2296.000 14.600 ;
      LAYER met4 ;
        RECT 7.655 10.640 20.640 2986.800 ;
        RECT 23.040 10.640 97.440 2986.800 ;
        RECT 99.840 10.640 2280.385 2986.800 ;
  END
END ghazi_top_dffram_csv
END LIBRARY

