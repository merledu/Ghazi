VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 41.380 2618.710 41.440 ;
        RECT 2900.830 41.380 2901.150 41.440 ;
        RECT 2618.390 41.240 2901.150 41.380 ;
        RECT 2618.390 41.180 2618.710 41.240 ;
        RECT 2900.830 41.180 2901.150 41.240 ;
      LAYER via ;
        RECT 2618.420 41.180 2618.680 41.440 ;
        RECT 2900.860 41.180 2901.120 41.440 ;
      LAYER met2 ;
        RECT 2618.410 293.235 2618.690 293.605 ;
        RECT 2618.480 41.470 2618.620 293.235 ;
        RECT 2618.420 41.150 2618.680 41.470 ;
        RECT 2900.860 41.150 2901.120 41.470 ;
        RECT 2900.920 39.285 2901.060 41.150 ;
        RECT 2900.850 38.915 2901.130 39.285 ;
      LAYER via2 ;
        RECT 2618.410 293.280 2618.690 293.560 ;
        RECT 2900.850 38.960 2901.130 39.240 ;
      LAYER met3 ;
        RECT 2606.000 293.570 2610.000 293.960 ;
        RECT 2618.385 293.570 2618.715 293.585 ;
        RECT 2606.000 293.360 2618.715 293.570 ;
        RECT 2609.580 293.270 2618.715 293.360 ;
        RECT 2618.385 293.255 2618.715 293.270 ;
        RECT 2900.825 39.250 2901.155 39.265 ;
        RECT 2917.600 39.250 2924.800 39.700 ;
        RECT 2900.825 38.950 2924.800 39.250 ;
        RECT 2900.825 38.935 2901.155 38.950 ;
        RECT 2917.600 38.500 2924.800 38.950 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2380.580 2618.710 2380.640 ;
        RECT 2900.830 2380.580 2901.150 2380.640 ;
        RECT 2618.390 2380.440 2901.150 2380.580 ;
        RECT 2618.390 2380.380 2618.710 2380.440 ;
        RECT 2900.830 2380.380 2901.150 2380.440 ;
      LAYER via ;
        RECT 2618.420 2380.380 2618.680 2380.640 ;
        RECT 2900.860 2380.380 2901.120 2380.640 ;
      LAYER met2 ;
        RECT 2900.850 2384.915 2901.130 2385.285 ;
        RECT 2900.920 2380.670 2901.060 2384.915 ;
        RECT 2618.420 2380.350 2618.680 2380.670 ;
        RECT 2900.860 2380.350 2901.120 2380.670 ;
        RECT 2618.480 2293.485 2618.620 2380.350 ;
        RECT 2618.410 2293.115 2618.690 2293.485 ;
      LAYER via2 ;
        RECT 2900.850 2384.960 2901.130 2385.240 ;
        RECT 2618.410 2293.160 2618.690 2293.440 ;
      LAYER met3 ;
        RECT 2900.825 2385.250 2901.155 2385.265 ;
        RECT 2917.600 2385.250 2924.800 2385.700 ;
        RECT 2900.825 2384.950 2924.800 2385.250 ;
        RECT 2900.825 2384.935 2901.155 2384.950 ;
        RECT 2917.600 2384.500 2924.800 2384.950 ;
        RECT 2606.000 2293.450 2610.000 2293.840 ;
        RECT 2618.385 2293.450 2618.715 2293.465 ;
        RECT 2606.000 2293.240 2618.715 2293.450 ;
        RECT 2609.580 2293.150 2618.715 2293.240 ;
        RECT 2618.385 2293.135 2618.715 2293.150 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2615.180 2619.170 2615.240 ;
        RECT 2900.830 2615.180 2901.150 2615.240 ;
        RECT 2618.850 2615.040 2901.150 2615.180 ;
        RECT 2618.850 2614.980 2619.170 2615.040 ;
        RECT 2900.830 2614.980 2901.150 2615.040 ;
      LAYER via ;
        RECT 2618.880 2614.980 2619.140 2615.240 ;
        RECT 2900.860 2614.980 2901.120 2615.240 ;
      LAYER met2 ;
        RECT 2900.850 2619.515 2901.130 2619.885 ;
        RECT 2900.920 2615.270 2901.060 2619.515 ;
        RECT 2618.880 2614.950 2619.140 2615.270 ;
        RECT 2900.860 2614.950 2901.120 2615.270 ;
        RECT 2618.940 2493.405 2619.080 2614.950 ;
        RECT 2618.870 2493.035 2619.150 2493.405 ;
      LAYER via2 ;
        RECT 2900.850 2619.560 2901.130 2619.840 ;
        RECT 2618.870 2493.080 2619.150 2493.360 ;
      LAYER met3 ;
        RECT 2900.825 2619.850 2901.155 2619.865 ;
        RECT 2917.600 2619.850 2924.800 2620.300 ;
        RECT 2900.825 2619.550 2924.800 2619.850 ;
        RECT 2900.825 2619.535 2901.155 2619.550 ;
        RECT 2917.600 2619.100 2924.800 2619.550 ;
        RECT 2606.000 2493.370 2610.000 2493.760 ;
        RECT 2618.845 2493.370 2619.175 2493.385 ;
        RECT 2606.000 2493.160 2619.175 2493.370 ;
        RECT 2609.580 2493.070 2619.175 2493.160 ;
        RECT 2618.845 2493.055 2619.175 2493.070 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2697.800 2618.710 2697.860 ;
        RECT 2901.290 2697.800 2901.610 2697.860 ;
        RECT 2618.390 2697.660 2901.610 2697.800 ;
        RECT 2618.390 2697.600 2618.710 2697.660 ;
        RECT 2901.290 2697.600 2901.610 2697.660 ;
      LAYER via ;
        RECT 2618.420 2697.600 2618.680 2697.860 ;
        RECT 2901.320 2697.600 2901.580 2697.860 ;
      LAYER met2 ;
        RECT 2901.310 2854.115 2901.590 2854.485 ;
        RECT 2901.380 2697.890 2901.520 2854.115 ;
        RECT 2618.420 2697.570 2618.680 2697.890 ;
        RECT 2901.320 2697.570 2901.580 2697.890 ;
        RECT 2618.480 2693.325 2618.620 2697.570 ;
        RECT 2618.410 2692.955 2618.690 2693.325 ;
      LAYER via2 ;
        RECT 2901.310 2854.160 2901.590 2854.440 ;
        RECT 2618.410 2693.000 2618.690 2693.280 ;
      LAYER met3 ;
        RECT 2901.285 2854.450 2901.615 2854.465 ;
        RECT 2917.600 2854.450 2924.800 2854.900 ;
        RECT 2901.285 2854.150 2924.800 2854.450 ;
        RECT 2901.285 2854.135 2901.615 2854.150 ;
        RECT 2917.600 2853.700 2924.800 2854.150 ;
        RECT 2606.000 2693.290 2610.000 2693.680 ;
        RECT 2618.385 2693.290 2618.715 2693.305 ;
        RECT 2606.000 2693.080 2618.715 2693.290 ;
        RECT 2609.580 2692.990 2618.715 2693.080 ;
        RECT 2618.385 2692.975 2618.715 2692.990 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 2898.060 2621.930 2898.120 ;
        RECT 2901.290 2898.060 2901.610 2898.120 ;
        RECT 2621.610 2897.920 2901.610 2898.060 ;
        RECT 2621.610 2897.860 2621.930 2897.920 ;
        RECT 2901.290 2897.860 2901.610 2897.920 ;
      LAYER via ;
        RECT 2621.640 2897.860 2621.900 2898.120 ;
        RECT 2901.320 2897.860 2901.580 2898.120 ;
      LAYER met2 ;
        RECT 2901.310 3088.715 2901.590 3089.085 ;
        RECT 2901.380 2898.150 2901.520 3088.715 ;
        RECT 2621.640 2897.830 2621.900 2898.150 ;
        RECT 2901.320 2897.830 2901.580 2898.150 ;
        RECT 2621.700 2893.245 2621.840 2897.830 ;
        RECT 2621.630 2892.875 2621.910 2893.245 ;
      LAYER via2 ;
        RECT 2901.310 3088.760 2901.590 3089.040 ;
        RECT 2621.630 2892.920 2621.910 2893.200 ;
      LAYER met3 ;
        RECT 2901.285 3089.050 2901.615 3089.065 ;
        RECT 2917.600 3089.050 2924.800 3089.500 ;
        RECT 2901.285 3088.750 2924.800 3089.050 ;
        RECT 2901.285 3088.735 2901.615 3088.750 ;
        RECT 2917.600 3088.300 2924.800 3088.750 ;
        RECT 2606.000 2893.210 2610.000 2893.600 ;
        RECT 2621.605 2893.210 2621.935 2893.225 ;
        RECT 2606.000 2893.000 2621.935 2893.210 ;
        RECT 2609.580 2892.910 2621.935 2893.000 ;
        RECT 2621.605 2892.895 2621.935 2892.910 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 3097.980 2621.930 3098.040 ;
        RECT 2901.290 3097.980 2901.610 3098.040 ;
        RECT 2621.610 3097.840 2901.610 3097.980 ;
        RECT 2621.610 3097.780 2621.930 3097.840 ;
        RECT 2901.290 3097.780 2901.610 3097.840 ;
      LAYER via ;
        RECT 2621.640 3097.780 2621.900 3098.040 ;
        RECT 2901.320 3097.780 2901.580 3098.040 ;
      LAYER met2 ;
        RECT 2901.310 3323.315 2901.590 3323.685 ;
        RECT 2901.380 3098.070 2901.520 3323.315 ;
        RECT 2621.640 3097.750 2621.900 3098.070 ;
        RECT 2901.320 3097.750 2901.580 3098.070 ;
        RECT 2621.700 3093.165 2621.840 3097.750 ;
        RECT 2621.630 3092.795 2621.910 3093.165 ;
      LAYER via2 ;
        RECT 2901.310 3323.360 2901.590 3323.640 ;
        RECT 2621.630 3092.840 2621.910 3093.120 ;
      LAYER met3 ;
        RECT 2901.285 3323.650 2901.615 3323.665 ;
        RECT 2917.600 3323.650 2924.800 3324.100 ;
        RECT 2901.285 3323.350 2924.800 3323.650 ;
        RECT 2901.285 3323.335 2901.615 3323.350 ;
        RECT 2917.600 3322.900 2924.800 3323.350 ;
        RECT 2606.000 3093.130 2610.000 3093.520 ;
        RECT 2621.605 3093.130 2621.935 3093.145 ;
        RECT 2606.000 3092.920 2621.935 3093.130 ;
        RECT 2609.580 3092.830 2621.935 3092.920 ;
        RECT 2621.605 3092.815 2621.935 3092.830 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 3501.560 2573.630 3501.620 ;
        RECT 2865.410 3501.560 2865.730 3501.620 ;
        RECT 2573.310 3501.420 2865.730 3501.560 ;
        RECT 2573.310 3501.360 2573.630 3501.420 ;
        RECT 2865.410 3501.360 2865.730 3501.420 ;
        RECT 2566.870 3276.480 2567.190 3276.540 ;
        RECT 2573.310 3276.480 2573.630 3276.540 ;
        RECT 2566.870 3276.340 2573.630 3276.480 ;
        RECT 2566.870 3276.280 2567.190 3276.340 ;
        RECT 2573.310 3276.280 2573.630 3276.340 ;
      LAYER via ;
        RECT 2573.340 3501.360 2573.600 3501.620 ;
        RECT 2865.440 3501.360 2865.700 3501.620 ;
        RECT 2566.900 3276.280 2567.160 3276.540 ;
        RECT 2573.340 3276.280 2573.600 3276.540 ;
      LAYER met2 ;
        RECT 2865.290 3517.600 2865.850 3524.800 ;
        RECT 2865.500 3501.650 2865.640 3517.600 ;
        RECT 2573.340 3501.330 2573.600 3501.650 ;
        RECT 2865.440 3501.330 2865.700 3501.650 ;
        RECT 2573.400 3276.570 2573.540 3501.330 ;
        RECT 2566.900 3276.250 2567.160 3276.570 ;
        RECT 2573.340 3276.250 2573.600 3276.570 ;
        RECT 2566.960 3260.000 2567.100 3276.250 ;
        RECT 2566.850 3256.000 2567.130 3260.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2318.010 3501.560 2318.330 3501.620 ;
        RECT 2541.110 3501.560 2541.430 3501.620 ;
        RECT 2318.010 3501.420 2541.430 3501.560 ;
        RECT 2318.010 3501.360 2318.330 3501.420 ;
        RECT 2541.110 3501.360 2541.430 3501.420 ;
        RECT 2311.570 3277.500 2311.890 3277.560 ;
        RECT 2318.010 3277.500 2318.330 3277.560 ;
        RECT 2311.570 3277.360 2318.330 3277.500 ;
        RECT 2311.570 3277.300 2311.890 3277.360 ;
        RECT 2318.010 3277.300 2318.330 3277.360 ;
      LAYER via ;
        RECT 2318.040 3501.360 2318.300 3501.620 ;
        RECT 2541.140 3501.360 2541.400 3501.620 ;
        RECT 2311.600 3277.300 2311.860 3277.560 ;
        RECT 2318.040 3277.300 2318.300 3277.560 ;
      LAYER met2 ;
        RECT 2540.990 3517.600 2541.550 3524.800 ;
        RECT 2541.200 3501.650 2541.340 3517.600 ;
        RECT 2318.040 3501.330 2318.300 3501.650 ;
        RECT 2541.140 3501.330 2541.400 3501.650 ;
        RECT 2318.100 3277.590 2318.240 3501.330 ;
        RECT 2311.600 3277.270 2311.860 3277.590 ;
        RECT 2318.040 3277.270 2318.300 3277.590 ;
        RECT 2311.660 3260.000 2311.800 3277.270 ;
        RECT 2311.550 3256.000 2311.830 3260.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 3501.560 2056.130 3501.620 ;
        RECT 2216.810 3501.560 2217.130 3501.620 ;
        RECT 2055.810 3501.420 2217.130 3501.560 ;
        RECT 2055.810 3501.360 2056.130 3501.420 ;
        RECT 2216.810 3501.360 2217.130 3501.420 ;
      LAYER via ;
        RECT 2055.840 3501.360 2056.100 3501.620 ;
        RECT 2216.840 3501.360 2217.100 3501.620 ;
      LAYER met2 ;
        RECT 2216.690 3517.600 2217.250 3524.800 ;
        RECT 2216.900 3501.650 2217.040 3517.600 ;
        RECT 2055.840 3501.330 2056.100 3501.650 ;
        RECT 2216.840 3501.330 2217.100 3501.650 ;
        RECT 2055.900 3260.000 2056.040 3501.330 ;
        RECT 2055.790 3256.000 2056.070 3260.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.510 3501.900 1800.830 3501.960 ;
        RECT 1892.050 3501.900 1892.370 3501.960 ;
        RECT 1800.510 3501.760 1892.370 3501.900 ;
        RECT 1800.510 3501.700 1800.830 3501.760 ;
        RECT 1892.050 3501.700 1892.370 3501.760 ;
      LAYER via ;
        RECT 1800.540 3501.700 1800.800 3501.960 ;
        RECT 1892.080 3501.700 1892.340 3501.960 ;
      LAYER met2 ;
        RECT 1891.930 3517.600 1892.490 3524.800 ;
        RECT 1892.140 3501.990 1892.280 3517.600 ;
        RECT 1800.540 3501.670 1800.800 3501.990 ;
        RECT 1892.080 3501.670 1892.340 3501.990 ;
        RECT 1800.600 3260.000 1800.740 3501.670 ;
        RECT 1800.490 3256.000 1800.770 3260.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 3498.500 1545.530 3498.560 ;
        RECT 1567.750 3498.500 1568.070 3498.560 ;
        RECT 1545.210 3498.360 1568.070 3498.500 ;
        RECT 1545.210 3498.300 1545.530 3498.360 ;
        RECT 1567.750 3498.300 1568.070 3498.360 ;
      LAYER via ;
        RECT 1545.240 3498.300 1545.500 3498.560 ;
        RECT 1567.780 3498.300 1568.040 3498.560 ;
      LAYER met2 ;
        RECT 1567.630 3517.600 1568.190 3524.800 ;
        RECT 1567.840 3498.590 1567.980 3517.600 ;
        RECT 1545.240 3498.270 1545.500 3498.590 ;
        RECT 1567.780 3498.270 1568.040 3498.590 ;
        RECT 1544.730 3259.650 1545.010 3260.000 ;
        RECT 1545.300 3259.650 1545.440 3498.270 ;
        RECT 1544.730 3259.510 1545.440 3259.650 ;
        RECT 1544.730 3256.000 1545.010 3259.510 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.770 275.980 2620.090 276.040 ;
        RECT 2900.830 275.980 2901.150 276.040 ;
        RECT 2619.770 275.840 2901.150 275.980 ;
        RECT 2619.770 275.780 2620.090 275.840 ;
        RECT 2900.830 275.780 2901.150 275.840 ;
      LAYER via ;
        RECT 2619.800 275.780 2620.060 276.040 ;
        RECT 2900.860 275.780 2901.120 276.040 ;
      LAYER met2 ;
        RECT 2619.790 493.155 2620.070 493.525 ;
        RECT 2619.860 276.070 2620.000 493.155 ;
        RECT 2619.800 275.750 2620.060 276.070 ;
        RECT 2900.860 275.750 2901.120 276.070 ;
        RECT 2900.920 273.885 2901.060 275.750 ;
        RECT 2900.850 273.515 2901.130 273.885 ;
      LAYER via2 ;
        RECT 2619.790 493.200 2620.070 493.480 ;
        RECT 2900.850 273.560 2901.130 273.840 ;
      LAYER met3 ;
        RECT 2606.000 493.490 2610.000 493.880 ;
        RECT 2619.765 493.490 2620.095 493.505 ;
        RECT 2606.000 493.280 2620.095 493.490 ;
        RECT 2609.580 493.190 2620.095 493.280 ;
        RECT 2619.765 493.175 2620.095 493.190 ;
        RECT 2900.825 273.850 2901.155 273.865 ;
        RECT 2917.600 273.850 2924.800 274.300 ;
        RECT 2900.825 273.550 2924.800 273.850 ;
        RECT 2900.825 273.535 2901.155 273.550 ;
        RECT 2917.600 273.100 2924.800 273.550 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1243.450 3498.500 1243.770 3498.560 ;
        RECT 1248.510 3498.500 1248.830 3498.560 ;
        RECT 1243.450 3498.360 1248.830 3498.500 ;
        RECT 1243.450 3498.300 1243.770 3498.360 ;
        RECT 1248.510 3498.300 1248.830 3498.360 ;
        RECT 1248.510 3277.500 1248.830 3277.560 ;
        RECT 1289.450 3277.500 1289.770 3277.560 ;
        RECT 1248.510 3277.360 1289.770 3277.500 ;
        RECT 1248.510 3277.300 1248.830 3277.360 ;
        RECT 1289.450 3277.300 1289.770 3277.360 ;
      LAYER via ;
        RECT 1243.480 3498.300 1243.740 3498.560 ;
        RECT 1248.540 3498.300 1248.800 3498.560 ;
        RECT 1248.540 3277.300 1248.800 3277.560 ;
        RECT 1289.480 3277.300 1289.740 3277.560 ;
      LAYER met2 ;
        RECT 1243.330 3517.600 1243.890 3524.800 ;
        RECT 1243.540 3498.590 1243.680 3517.600 ;
        RECT 1243.480 3498.270 1243.740 3498.590 ;
        RECT 1248.540 3498.270 1248.800 3498.590 ;
        RECT 1248.600 3277.590 1248.740 3498.270 ;
        RECT 1248.540 3277.270 1248.800 3277.590 ;
        RECT 1289.480 3277.270 1289.740 3277.590 ;
        RECT 1289.540 3260.000 1289.680 3277.270 ;
        RECT 1289.430 3256.000 1289.710 3260.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 918.690 3500.880 919.010 3500.940 ;
        RECT 924.210 3500.880 924.530 3500.940 ;
        RECT 918.690 3500.740 924.530 3500.880 ;
        RECT 918.690 3500.680 919.010 3500.740 ;
        RECT 924.210 3500.680 924.530 3500.740 ;
        RECT 924.210 3274.100 924.530 3274.160 ;
        RECT 1033.690 3274.100 1034.010 3274.160 ;
        RECT 924.210 3273.960 1034.010 3274.100 ;
        RECT 924.210 3273.900 924.530 3273.960 ;
        RECT 1033.690 3273.900 1034.010 3273.960 ;
      LAYER via ;
        RECT 918.720 3500.680 918.980 3500.940 ;
        RECT 924.240 3500.680 924.500 3500.940 ;
        RECT 924.240 3273.900 924.500 3274.160 ;
        RECT 1033.720 3273.900 1033.980 3274.160 ;
      LAYER met2 ;
        RECT 918.570 3517.600 919.130 3524.800 ;
        RECT 918.780 3500.970 918.920 3517.600 ;
        RECT 918.720 3500.650 918.980 3500.970 ;
        RECT 924.240 3500.650 924.500 3500.970 ;
        RECT 924.300 3274.190 924.440 3500.650 ;
        RECT 924.240 3273.870 924.500 3274.190 ;
        RECT 1033.720 3273.870 1033.980 3274.190 ;
        RECT 1033.780 3260.000 1033.920 3273.870 ;
        RECT 1033.670 3256.000 1033.950 3260.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 594.390 3498.500 594.710 3498.560 ;
        RECT 599.910 3498.500 600.230 3498.560 ;
        RECT 594.390 3498.360 600.230 3498.500 ;
        RECT 594.390 3498.300 594.710 3498.360 ;
        RECT 599.910 3498.300 600.230 3498.360 ;
        RECT 599.910 3274.780 600.230 3274.840 ;
        RECT 777.930 3274.780 778.250 3274.840 ;
        RECT 599.910 3274.640 778.250 3274.780 ;
        RECT 599.910 3274.580 600.230 3274.640 ;
        RECT 777.930 3274.580 778.250 3274.640 ;
      LAYER via ;
        RECT 594.420 3498.300 594.680 3498.560 ;
        RECT 599.940 3498.300 600.200 3498.560 ;
        RECT 599.940 3274.580 600.200 3274.840 ;
        RECT 777.960 3274.580 778.220 3274.840 ;
      LAYER met2 ;
        RECT 594.270 3517.600 594.830 3524.800 ;
        RECT 594.480 3498.590 594.620 3517.600 ;
        RECT 594.420 3498.270 594.680 3498.590 ;
        RECT 599.940 3498.270 600.200 3498.590 ;
        RECT 600.000 3274.870 600.140 3498.270 ;
        RECT 599.940 3274.550 600.200 3274.870 ;
        RECT 777.960 3274.550 778.220 3274.870 ;
        RECT 778.020 3260.000 778.160 3274.550 ;
        RECT 777.910 3256.000 778.190 3260.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 270.090 3504.280 270.410 3504.340 ;
        RECT 275.610 3504.280 275.930 3504.340 ;
        RECT 270.090 3504.140 275.930 3504.280 ;
        RECT 270.090 3504.080 270.410 3504.140 ;
        RECT 275.610 3504.080 275.930 3504.140 ;
        RECT 275.610 3274.780 275.930 3274.840 ;
        RECT 522.630 3274.780 522.950 3274.840 ;
        RECT 275.610 3274.640 522.950 3274.780 ;
        RECT 275.610 3274.580 275.930 3274.640 ;
        RECT 522.630 3274.580 522.950 3274.640 ;
      LAYER via ;
        RECT 270.120 3504.080 270.380 3504.340 ;
        RECT 275.640 3504.080 275.900 3504.340 ;
        RECT 275.640 3274.580 275.900 3274.840 ;
        RECT 522.660 3274.580 522.920 3274.840 ;
      LAYER met2 ;
        RECT 269.970 3517.600 270.530 3524.800 ;
        RECT 270.180 3504.370 270.320 3517.600 ;
        RECT 270.120 3504.050 270.380 3504.370 ;
        RECT 275.640 3504.050 275.900 3504.370 ;
        RECT 275.700 3274.870 275.840 3504.050 ;
        RECT 275.640 3274.550 275.900 3274.870 ;
        RECT 522.660 3274.550 522.920 3274.870 ;
        RECT 522.720 3260.000 522.860 3274.550 ;
        RECT 522.610 3256.000 522.890 3260.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3229.220 17.410 3229.280 ;
        RECT 296.770 3229.220 297.090 3229.280 ;
        RECT 17.090 3229.080 297.090 3229.220 ;
        RECT 17.090 3229.020 17.410 3229.080 ;
        RECT 296.770 3229.020 297.090 3229.080 ;
      LAYER via ;
        RECT 17.120 3229.020 17.380 3229.280 ;
        RECT 296.800 3229.020 297.060 3229.280 ;
      LAYER met2 ;
        RECT 17.110 3476.995 17.390 3477.365 ;
        RECT 17.180 3229.310 17.320 3476.995 ;
        RECT 17.120 3228.990 17.380 3229.310 ;
        RECT 296.800 3228.990 297.060 3229.310 ;
        RECT 296.860 3223.725 297.000 3228.990 ;
        RECT 296.790 3223.355 297.070 3223.725 ;
      LAYER via2 ;
        RECT 17.110 3477.040 17.390 3477.320 ;
        RECT 296.790 3223.400 297.070 3223.680 ;
      LAYER met3 ;
        RECT -4.800 3477.330 2.400 3477.780 ;
        RECT 17.085 3477.330 17.415 3477.345 ;
        RECT -4.800 3477.030 17.415 3477.330 ;
        RECT -4.800 3476.580 2.400 3477.030 ;
        RECT 17.085 3477.015 17.415 3477.030 ;
        RECT 296.765 3223.690 297.095 3223.705 ;
        RECT 310.000 3223.690 314.000 3224.080 ;
        RECT 296.765 3223.480 314.000 3223.690 ;
        RECT 296.765 3223.390 310.500 3223.480 ;
        RECT 296.765 3223.375 297.095 3223.390 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.470 3015.360 18.790 3015.420 ;
        RECT 296.770 3015.360 297.090 3015.420 ;
        RECT 18.470 3015.220 297.090 3015.360 ;
        RECT 18.470 3015.160 18.790 3015.220 ;
        RECT 296.770 3015.160 297.090 3015.220 ;
      LAYER via ;
        RECT 18.500 3015.160 18.760 3015.420 ;
        RECT 296.800 3015.160 297.060 3015.420 ;
      LAYER met2 ;
        RECT 18.490 3226.075 18.770 3226.445 ;
        RECT 18.560 3015.450 18.700 3226.075 ;
        RECT 18.500 3015.130 18.760 3015.450 ;
        RECT 296.800 3015.130 297.060 3015.450 ;
        RECT 296.860 3009.525 297.000 3015.130 ;
        RECT 296.790 3009.155 297.070 3009.525 ;
      LAYER via2 ;
        RECT 18.490 3226.120 18.770 3226.400 ;
        RECT 296.790 3009.200 297.070 3009.480 ;
      LAYER met3 ;
        RECT -4.800 3226.410 2.400 3226.860 ;
        RECT 18.465 3226.410 18.795 3226.425 ;
        RECT -4.800 3226.110 18.795 3226.410 ;
        RECT -4.800 3225.660 2.400 3226.110 ;
        RECT 18.465 3226.095 18.795 3226.110 ;
        RECT 296.765 3009.490 297.095 3009.505 ;
        RECT 310.000 3009.490 314.000 3009.880 ;
        RECT 296.765 3009.280 314.000 3009.490 ;
        RECT 296.765 3009.190 310.500 3009.280 ;
        RECT 296.765 3009.175 297.095 3009.190 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 2801.160 18.330 2801.220 ;
        RECT 296.770 2801.160 297.090 2801.220 ;
        RECT 18.010 2801.020 297.090 2801.160 ;
        RECT 18.010 2800.960 18.330 2801.020 ;
        RECT 296.770 2800.960 297.090 2801.020 ;
      LAYER via ;
        RECT 18.040 2800.960 18.300 2801.220 ;
        RECT 296.800 2800.960 297.060 2801.220 ;
      LAYER met2 ;
        RECT 18.030 2974.475 18.310 2974.845 ;
        RECT 18.100 2801.250 18.240 2974.475 ;
        RECT 18.040 2800.930 18.300 2801.250 ;
        RECT 296.800 2800.930 297.060 2801.250 ;
        RECT 296.860 2795.325 297.000 2800.930 ;
        RECT 296.790 2794.955 297.070 2795.325 ;
      LAYER via2 ;
        RECT 18.030 2974.520 18.310 2974.800 ;
        RECT 296.790 2795.000 297.070 2795.280 ;
      LAYER met3 ;
        RECT -4.800 2974.810 2.400 2975.260 ;
        RECT 18.005 2974.810 18.335 2974.825 ;
        RECT -4.800 2974.510 18.335 2974.810 ;
        RECT -4.800 2974.060 2.400 2974.510 ;
        RECT 18.005 2974.495 18.335 2974.510 ;
        RECT 296.765 2795.290 297.095 2795.305 ;
        RECT 310.000 2795.290 314.000 2795.680 ;
        RECT 296.765 2795.080 314.000 2795.290 ;
        RECT 296.765 2794.990 310.500 2795.080 ;
        RECT 296.765 2794.975 297.095 2794.990 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 2587.300 18.330 2587.360 ;
        RECT 296.770 2587.300 297.090 2587.360 ;
        RECT 18.010 2587.160 297.090 2587.300 ;
        RECT 18.010 2587.100 18.330 2587.160 ;
        RECT 296.770 2587.100 297.090 2587.160 ;
      LAYER via ;
        RECT 18.040 2587.100 18.300 2587.360 ;
        RECT 296.800 2587.100 297.060 2587.360 ;
      LAYER met2 ;
        RECT 18.030 2722.875 18.310 2723.245 ;
        RECT 18.100 2587.390 18.240 2722.875 ;
        RECT 18.040 2587.070 18.300 2587.390 ;
        RECT 296.800 2587.070 297.060 2587.390 ;
        RECT 296.860 2581.125 297.000 2587.070 ;
        RECT 296.790 2580.755 297.070 2581.125 ;
      LAYER via2 ;
        RECT 18.030 2722.920 18.310 2723.200 ;
        RECT 296.790 2580.800 297.070 2581.080 ;
      LAYER met3 ;
        RECT -4.800 2723.210 2.400 2723.660 ;
        RECT 18.005 2723.210 18.335 2723.225 ;
        RECT -4.800 2722.910 18.335 2723.210 ;
        RECT -4.800 2722.460 2.400 2722.910 ;
        RECT 18.005 2722.895 18.335 2722.910 ;
        RECT 296.765 2581.090 297.095 2581.105 ;
        RECT 310.000 2581.090 314.000 2581.480 ;
        RECT 296.765 2580.880 314.000 2581.090 ;
        RECT 296.765 2580.790 310.500 2580.880 ;
        RECT 296.765 2580.775 297.095 2580.790 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2373.440 17.410 2373.500 ;
        RECT 296.770 2373.440 297.090 2373.500 ;
        RECT 17.090 2373.300 297.090 2373.440 ;
        RECT 17.090 2373.240 17.410 2373.300 ;
        RECT 296.770 2373.240 297.090 2373.300 ;
      LAYER via ;
        RECT 17.120 2373.240 17.380 2373.500 ;
        RECT 296.800 2373.240 297.060 2373.500 ;
      LAYER met2 ;
        RECT 17.110 2471.275 17.390 2471.645 ;
        RECT 17.180 2373.530 17.320 2471.275 ;
        RECT 17.120 2373.210 17.380 2373.530 ;
        RECT 296.800 2373.210 297.060 2373.530 ;
        RECT 296.860 2366.925 297.000 2373.210 ;
        RECT 296.790 2366.555 297.070 2366.925 ;
      LAYER via2 ;
        RECT 17.110 2471.320 17.390 2471.600 ;
        RECT 296.790 2366.600 297.070 2366.880 ;
      LAYER met3 ;
        RECT -4.800 2471.610 2.400 2472.060 ;
        RECT 17.085 2471.610 17.415 2471.625 ;
        RECT -4.800 2471.310 17.415 2471.610 ;
        RECT -4.800 2470.860 2.400 2471.310 ;
        RECT 17.085 2471.295 17.415 2471.310 ;
        RECT 296.765 2366.890 297.095 2366.905 ;
        RECT 310.000 2366.890 314.000 2367.280 ;
        RECT 296.765 2366.680 314.000 2366.890 ;
        RECT 296.765 2366.590 310.500 2366.680 ;
        RECT 296.765 2366.575 297.095 2366.590 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2152.780 17.410 2152.840 ;
        RECT 296.770 2152.780 297.090 2152.840 ;
        RECT 17.090 2152.640 297.090 2152.780 ;
        RECT 17.090 2152.580 17.410 2152.640 ;
        RECT 296.770 2152.580 297.090 2152.640 ;
      LAYER via ;
        RECT 17.120 2152.580 17.380 2152.840 ;
        RECT 296.800 2152.580 297.060 2152.840 ;
      LAYER met2 ;
        RECT 17.110 2220.355 17.390 2220.725 ;
        RECT 17.180 2152.870 17.320 2220.355 ;
        RECT 17.120 2152.550 17.380 2152.870 ;
        RECT 296.800 2152.725 297.060 2152.870 ;
        RECT 296.790 2152.355 297.070 2152.725 ;
      LAYER via2 ;
        RECT 17.110 2220.400 17.390 2220.680 ;
        RECT 296.790 2152.400 297.070 2152.680 ;
      LAYER met3 ;
        RECT -4.800 2220.690 2.400 2221.140 ;
        RECT 17.085 2220.690 17.415 2220.705 ;
        RECT -4.800 2220.390 17.415 2220.690 ;
        RECT -4.800 2219.940 2.400 2220.390 ;
        RECT 17.085 2220.375 17.415 2220.390 ;
        RECT 296.765 2152.690 297.095 2152.705 ;
        RECT 310.000 2152.690 314.000 2153.080 ;
        RECT 296.765 2152.480 314.000 2152.690 ;
        RECT 296.765 2152.390 310.500 2152.480 ;
        RECT 296.765 2152.375 297.095 2152.390 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 510.580 2619.630 510.640 ;
        RECT 2900.830 510.580 2901.150 510.640 ;
        RECT 2619.310 510.440 2901.150 510.580 ;
        RECT 2619.310 510.380 2619.630 510.440 ;
        RECT 2900.830 510.380 2901.150 510.440 ;
      LAYER via ;
        RECT 2619.340 510.380 2619.600 510.640 ;
        RECT 2900.860 510.380 2901.120 510.640 ;
      LAYER met2 ;
        RECT 2619.330 693.075 2619.610 693.445 ;
        RECT 2619.400 510.670 2619.540 693.075 ;
        RECT 2619.340 510.350 2619.600 510.670 ;
        RECT 2900.860 510.350 2901.120 510.670 ;
        RECT 2900.920 508.485 2901.060 510.350 ;
        RECT 2900.850 508.115 2901.130 508.485 ;
      LAYER via2 ;
        RECT 2619.330 693.120 2619.610 693.400 ;
        RECT 2900.850 508.160 2901.130 508.440 ;
      LAYER met3 ;
        RECT 2606.000 693.410 2610.000 693.800 ;
        RECT 2619.305 693.410 2619.635 693.425 ;
        RECT 2606.000 693.200 2619.635 693.410 ;
        RECT 2609.580 693.110 2619.635 693.200 ;
        RECT 2619.305 693.095 2619.635 693.110 ;
        RECT 2900.825 508.450 2901.155 508.465 ;
        RECT 2917.600 508.450 2924.800 508.900 ;
        RECT 2900.825 508.150 2924.800 508.450 ;
        RECT 2900.825 508.135 2901.155 508.150 ;
        RECT 2917.600 507.700 2924.800 508.150 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 1938.920 19.710 1938.980 ;
        RECT 296.770 1938.920 297.090 1938.980 ;
        RECT 19.390 1938.780 297.090 1938.920 ;
        RECT 19.390 1938.720 19.710 1938.780 ;
        RECT 296.770 1938.720 297.090 1938.780 ;
      LAYER via ;
        RECT 19.420 1938.720 19.680 1938.980 ;
        RECT 296.800 1938.720 297.060 1938.980 ;
      LAYER met2 ;
        RECT 19.410 1968.755 19.690 1969.125 ;
        RECT 19.480 1939.010 19.620 1968.755 ;
        RECT 19.420 1938.690 19.680 1939.010 ;
        RECT 296.800 1938.690 297.060 1939.010 ;
        RECT 296.860 1938.525 297.000 1938.690 ;
        RECT 296.790 1938.155 297.070 1938.525 ;
      LAYER via2 ;
        RECT 19.410 1968.800 19.690 1969.080 ;
        RECT 296.790 1938.200 297.070 1938.480 ;
      LAYER met3 ;
        RECT -4.800 1969.090 2.400 1969.540 ;
        RECT 19.385 1969.090 19.715 1969.105 ;
        RECT -4.800 1968.790 19.715 1969.090 ;
        RECT -4.800 1968.340 2.400 1968.790 ;
        RECT 19.385 1968.775 19.715 1968.790 ;
        RECT 296.765 1938.490 297.095 1938.505 ;
        RECT 310.000 1938.490 314.000 1938.880 ;
        RECT 296.765 1938.280 314.000 1938.490 ;
        RECT 296.765 1938.190 310.500 1938.280 ;
        RECT 296.765 1938.175 297.095 1938.190 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1717.920 17.410 1717.980 ;
        RECT 296.770 1717.920 297.090 1717.980 ;
        RECT 17.090 1717.780 297.090 1717.920 ;
        RECT 17.090 1717.720 17.410 1717.780 ;
        RECT 296.770 1717.720 297.090 1717.780 ;
      LAYER via ;
        RECT 17.120 1717.720 17.380 1717.980 ;
        RECT 296.800 1717.720 297.060 1717.980 ;
      LAYER met2 ;
        RECT 296.790 1723.275 297.070 1723.645 ;
        RECT 296.860 1718.010 297.000 1723.275 ;
        RECT 17.120 1717.690 17.380 1718.010 ;
        RECT 296.800 1717.690 297.060 1718.010 ;
        RECT 17.180 1717.525 17.320 1717.690 ;
        RECT 17.110 1717.155 17.390 1717.525 ;
      LAYER via2 ;
        RECT 296.790 1723.320 297.070 1723.600 ;
        RECT 17.110 1717.200 17.390 1717.480 ;
      LAYER met3 ;
        RECT 296.765 1723.610 297.095 1723.625 ;
        RECT 310.000 1723.610 314.000 1724.000 ;
        RECT 296.765 1723.400 314.000 1723.610 ;
        RECT 296.765 1723.310 310.500 1723.400 ;
        RECT 296.765 1723.295 297.095 1723.310 ;
        RECT -4.800 1717.490 2.400 1717.940 ;
        RECT 17.085 1717.490 17.415 1717.505 ;
        RECT -4.800 1717.190 17.415 1717.490 ;
        RECT -4.800 1716.740 2.400 1717.190 ;
        RECT 17.085 1717.175 17.415 1717.190 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1469.720 16.030 1469.780 ;
        RECT 299.990 1469.720 300.310 1469.780 ;
        RECT 15.710 1469.580 300.310 1469.720 ;
        RECT 15.710 1469.520 16.030 1469.580 ;
        RECT 299.990 1469.520 300.310 1469.580 ;
      LAYER via ;
        RECT 15.740 1469.520 16.000 1469.780 ;
        RECT 300.020 1469.520 300.280 1469.780 ;
      LAYER met2 ;
        RECT 300.010 1509.075 300.290 1509.445 ;
        RECT 300.080 1469.810 300.220 1509.075 ;
        RECT 15.740 1469.490 16.000 1469.810 ;
        RECT 300.020 1469.490 300.280 1469.810 ;
        RECT 15.800 1466.605 15.940 1469.490 ;
        RECT 15.730 1466.235 16.010 1466.605 ;
      LAYER via2 ;
        RECT 300.010 1509.120 300.290 1509.400 ;
        RECT 15.730 1466.280 16.010 1466.560 ;
      LAYER met3 ;
        RECT 299.985 1509.410 300.315 1509.425 ;
        RECT 310.000 1509.410 314.000 1509.800 ;
        RECT 299.985 1509.200 314.000 1509.410 ;
        RECT 299.985 1509.110 310.500 1509.200 ;
        RECT 299.985 1509.095 300.315 1509.110 ;
        RECT -4.800 1466.570 2.400 1467.020 ;
        RECT 15.705 1466.570 16.035 1466.585 ;
        RECT -4.800 1466.270 16.035 1466.570 ;
        RECT -4.800 1465.820 2.400 1466.270 ;
        RECT 15.705 1466.255 16.035 1466.270 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1221.180 17.410 1221.240 ;
        RECT 299.990 1221.180 300.310 1221.240 ;
        RECT 17.090 1221.040 300.310 1221.180 ;
        RECT 17.090 1220.980 17.410 1221.040 ;
        RECT 299.990 1220.980 300.310 1221.040 ;
      LAYER via ;
        RECT 17.120 1220.980 17.380 1221.240 ;
        RECT 300.020 1220.980 300.280 1221.240 ;
      LAYER met2 ;
        RECT 300.010 1294.875 300.290 1295.245 ;
        RECT 300.080 1221.270 300.220 1294.875 ;
        RECT 17.120 1220.950 17.380 1221.270 ;
        RECT 300.020 1220.950 300.280 1221.270 ;
        RECT 17.180 1215.005 17.320 1220.950 ;
        RECT 17.110 1214.635 17.390 1215.005 ;
      LAYER via2 ;
        RECT 300.010 1294.920 300.290 1295.200 ;
        RECT 17.110 1214.680 17.390 1214.960 ;
      LAYER met3 ;
        RECT 299.985 1295.210 300.315 1295.225 ;
        RECT 310.000 1295.210 314.000 1295.600 ;
        RECT 299.985 1295.000 314.000 1295.210 ;
        RECT 299.985 1294.910 310.500 1295.000 ;
        RECT 299.985 1294.895 300.315 1294.910 ;
        RECT -4.800 1214.970 2.400 1215.420 ;
        RECT 17.085 1214.970 17.415 1214.985 ;
        RECT -4.800 1214.670 17.415 1214.970 ;
        RECT -4.800 1214.220 2.400 1214.670 ;
        RECT 17.085 1214.655 17.415 1214.670 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 965.840 17.870 965.900 ;
        RECT 300.450 965.840 300.770 965.900 ;
        RECT 17.550 965.700 300.770 965.840 ;
        RECT 17.550 965.640 17.870 965.700 ;
        RECT 300.450 965.640 300.770 965.700 ;
      LAYER via ;
        RECT 17.580 965.640 17.840 965.900 ;
        RECT 300.480 965.640 300.740 965.900 ;
      LAYER met2 ;
        RECT 300.470 1080.675 300.750 1081.045 ;
        RECT 300.540 965.930 300.680 1080.675 ;
        RECT 17.580 965.610 17.840 965.930 ;
        RECT 300.480 965.610 300.740 965.930 ;
        RECT 17.640 963.405 17.780 965.610 ;
        RECT 17.570 963.035 17.850 963.405 ;
      LAYER via2 ;
        RECT 300.470 1080.720 300.750 1081.000 ;
        RECT 17.570 963.080 17.850 963.360 ;
      LAYER met3 ;
        RECT 300.445 1081.010 300.775 1081.025 ;
        RECT 310.000 1081.010 314.000 1081.400 ;
        RECT 300.445 1080.800 314.000 1081.010 ;
        RECT 300.445 1080.710 310.500 1080.800 ;
        RECT 300.445 1080.695 300.775 1080.710 ;
        RECT -4.800 963.370 2.400 963.820 ;
        RECT 17.545 963.370 17.875 963.385 ;
        RECT -4.800 963.070 17.875 963.370 ;
        RECT -4.800 962.620 2.400 963.070 ;
        RECT 17.545 963.055 17.875 963.070 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 717.640 16.490 717.700 ;
        RECT 300.450 717.640 300.770 717.700 ;
        RECT 16.170 717.500 300.770 717.640 ;
        RECT 16.170 717.440 16.490 717.500 ;
        RECT 300.450 717.440 300.770 717.500 ;
      LAYER via ;
        RECT 16.200 717.440 16.460 717.700 ;
        RECT 300.480 717.440 300.740 717.700 ;
      LAYER met2 ;
        RECT 300.470 866.475 300.750 866.845 ;
        RECT 300.540 717.730 300.680 866.475 ;
        RECT 16.200 717.410 16.460 717.730 ;
        RECT 300.480 717.410 300.740 717.730 ;
        RECT 16.260 711.805 16.400 717.410 ;
        RECT 16.190 711.435 16.470 711.805 ;
      LAYER via2 ;
        RECT 300.470 866.520 300.750 866.800 ;
        RECT 16.190 711.480 16.470 711.760 ;
      LAYER met3 ;
        RECT 300.445 866.810 300.775 866.825 ;
        RECT 310.000 866.810 314.000 867.200 ;
        RECT 300.445 866.600 314.000 866.810 ;
        RECT 300.445 866.510 310.500 866.600 ;
        RECT 300.445 866.495 300.775 866.510 ;
        RECT -4.800 711.770 2.400 712.220 ;
        RECT 16.165 711.770 16.495 711.785 ;
        RECT -4.800 711.470 16.495 711.770 ;
        RECT -4.800 711.020 2.400 711.470 ;
        RECT 16.165 711.455 16.495 711.470 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 462.300 16.950 462.360 ;
        RECT 300.450 462.300 300.770 462.360 ;
        RECT 16.630 462.160 300.770 462.300 ;
        RECT 16.630 462.100 16.950 462.160 ;
        RECT 300.450 462.100 300.770 462.160 ;
      LAYER via ;
        RECT 16.660 462.100 16.920 462.360 ;
        RECT 300.480 462.100 300.740 462.360 ;
      LAYER met2 ;
        RECT 300.470 652.275 300.750 652.645 ;
        RECT 300.540 462.390 300.680 652.275 ;
        RECT 16.660 462.070 16.920 462.390 ;
        RECT 300.480 462.070 300.740 462.390 ;
        RECT 16.720 460.885 16.860 462.070 ;
        RECT 16.650 460.515 16.930 460.885 ;
      LAYER via2 ;
        RECT 300.470 652.320 300.750 652.600 ;
        RECT 16.650 460.560 16.930 460.840 ;
      LAYER met3 ;
        RECT 300.445 652.610 300.775 652.625 ;
        RECT 310.000 652.610 314.000 653.000 ;
        RECT 300.445 652.400 314.000 652.610 ;
        RECT 300.445 652.310 310.500 652.400 ;
        RECT 300.445 652.295 300.775 652.310 ;
        RECT -4.800 460.850 2.400 461.300 ;
        RECT 16.625 460.850 16.955 460.865 ;
        RECT -4.800 460.550 16.955 460.850 ;
        RECT -4.800 460.100 2.400 460.550 ;
        RECT 16.625 460.535 16.955 460.550 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 213.760 17.410 213.820 ;
        RECT 300.910 213.760 301.230 213.820 ;
        RECT 17.090 213.620 301.230 213.760 ;
        RECT 17.090 213.560 17.410 213.620 ;
        RECT 300.910 213.560 301.230 213.620 ;
      LAYER via ;
        RECT 17.120 213.560 17.380 213.820 ;
        RECT 300.940 213.560 301.200 213.820 ;
      LAYER met2 ;
        RECT 300.930 438.075 301.210 438.445 ;
        RECT 301.000 213.850 301.140 438.075 ;
        RECT 17.120 213.530 17.380 213.850 ;
        RECT 300.940 213.530 301.200 213.850 ;
        RECT 17.180 209.285 17.320 213.530 ;
        RECT 17.110 208.915 17.390 209.285 ;
      LAYER via2 ;
        RECT 300.930 438.120 301.210 438.400 ;
        RECT 17.110 208.960 17.390 209.240 ;
      LAYER met3 ;
        RECT 300.905 438.410 301.235 438.425 ;
        RECT 310.000 438.410 314.000 438.800 ;
        RECT 300.905 438.200 314.000 438.410 ;
        RECT 300.905 438.110 310.500 438.200 ;
        RECT 300.905 438.095 301.235 438.110 ;
        RECT -4.800 209.250 2.400 209.700 ;
        RECT 17.085 209.250 17.415 209.265 ;
        RECT -4.800 208.950 17.415 209.250 ;
        RECT -4.800 208.500 2.400 208.950 ;
        RECT 17.085 208.935 17.415 208.950 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 745.180 2619.630 745.240 ;
        RECT 2900.830 745.180 2901.150 745.240 ;
        RECT 2619.310 745.040 2901.150 745.180 ;
        RECT 2619.310 744.980 2619.630 745.040 ;
        RECT 2900.830 744.980 2901.150 745.040 ;
      LAYER via ;
        RECT 2619.340 744.980 2619.600 745.240 ;
        RECT 2900.860 744.980 2901.120 745.240 ;
      LAYER met2 ;
        RECT 2619.330 892.995 2619.610 893.365 ;
        RECT 2619.400 745.270 2619.540 892.995 ;
        RECT 2619.340 744.950 2619.600 745.270 ;
        RECT 2900.860 744.950 2901.120 745.270 ;
        RECT 2900.920 743.085 2901.060 744.950 ;
        RECT 2900.850 742.715 2901.130 743.085 ;
      LAYER via2 ;
        RECT 2619.330 893.040 2619.610 893.320 ;
        RECT 2900.850 742.760 2901.130 743.040 ;
      LAYER met3 ;
        RECT 2606.000 893.330 2610.000 893.720 ;
        RECT 2619.305 893.330 2619.635 893.345 ;
        RECT 2606.000 893.120 2619.635 893.330 ;
        RECT 2609.580 893.030 2619.635 893.120 ;
        RECT 2619.305 893.015 2619.635 893.030 ;
        RECT 2900.825 743.050 2901.155 743.065 ;
        RECT 2917.600 743.050 2924.800 743.500 ;
        RECT 2900.825 742.750 2924.800 743.050 ;
        RECT 2900.825 742.735 2901.155 742.750 ;
        RECT 2917.600 742.300 2924.800 742.750 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 979.780 2618.710 979.840 ;
        RECT 2900.830 979.780 2901.150 979.840 ;
        RECT 2618.390 979.640 2901.150 979.780 ;
        RECT 2618.390 979.580 2618.710 979.640 ;
        RECT 2900.830 979.580 2901.150 979.640 ;
      LAYER via ;
        RECT 2618.420 979.580 2618.680 979.840 ;
        RECT 2900.860 979.580 2901.120 979.840 ;
      LAYER met2 ;
        RECT 2618.410 1092.915 2618.690 1093.285 ;
        RECT 2618.480 979.870 2618.620 1092.915 ;
        RECT 2618.420 979.550 2618.680 979.870 ;
        RECT 2900.860 979.550 2901.120 979.870 ;
        RECT 2900.920 977.685 2901.060 979.550 ;
        RECT 2900.850 977.315 2901.130 977.685 ;
      LAYER via2 ;
        RECT 2618.410 1092.960 2618.690 1093.240 ;
        RECT 2900.850 977.360 2901.130 977.640 ;
      LAYER met3 ;
        RECT 2606.000 1093.250 2610.000 1093.640 ;
        RECT 2618.385 1093.250 2618.715 1093.265 ;
        RECT 2606.000 1093.040 2618.715 1093.250 ;
        RECT 2609.580 1092.950 2618.715 1093.040 ;
        RECT 2618.385 1092.935 2618.715 1092.950 ;
        RECT 2900.825 977.650 2901.155 977.665 ;
        RECT 2917.600 977.650 2924.800 978.100 ;
        RECT 2900.825 977.350 2924.800 977.650 ;
        RECT 2900.825 977.335 2901.155 977.350 ;
        RECT 2917.600 976.900 2924.800 977.350 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1214.380 2619.170 1214.440 ;
        RECT 2900.830 1214.380 2901.150 1214.440 ;
        RECT 2618.850 1214.240 2901.150 1214.380 ;
        RECT 2618.850 1214.180 2619.170 1214.240 ;
        RECT 2900.830 1214.180 2901.150 1214.240 ;
      LAYER via ;
        RECT 2618.880 1214.180 2619.140 1214.440 ;
        RECT 2900.860 1214.180 2901.120 1214.440 ;
      LAYER met2 ;
        RECT 2618.870 1292.835 2619.150 1293.205 ;
        RECT 2618.940 1214.470 2619.080 1292.835 ;
        RECT 2618.880 1214.150 2619.140 1214.470 ;
        RECT 2900.860 1214.150 2901.120 1214.470 ;
        RECT 2900.920 1212.285 2901.060 1214.150 ;
        RECT 2900.850 1211.915 2901.130 1212.285 ;
      LAYER via2 ;
        RECT 2618.870 1292.880 2619.150 1293.160 ;
        RECT 2900.850 1211.960 2901.130 1212.240 ;
      LAYER met3 ;
        RECT 2606.000 1293.170 2610.000 1293.560 ;
        RECT 2618.845 1293.170 2619.175 1293.185 ;
        RECT 2606.000 1292.960 2619.175 1293.170 ;
        RECT 2609.580 1292.870 2619.175 1292.960 ;
        RECT 2618.845 1292.855 2619.175 1292.870 ;
        RECT 2900.825 1212.250 2901.155 1212.265 ;
        RECT 2917.600 1212.250 2924.800 1212.700 ;
        RECT 2900.825 1211.950 2924.800 1212.250 ;
        RECT 2900.825 1211.935 2901.155 1211.950 ;
        RECT 2917.600 1211.500 2924.800 1211.950 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1448.980 2618.710 1449.040 ;
        RECT 2900.830 1448.980 2901.150 1449.040 ;
        RECT 2618.390 1448.840 2901.150 1448.980 ;
        RECT 2618.390 1448.780 2618.710 1448.840 ;
        RECT 2900.830 1448.780 2901.150 1448.840 ;
      LAYER via ;
        RECT 2618.420 1448.780 2618.680 1449.040 ;
        RECT 2900.860 1448.780 2901.120 1449.040 ;
      LAYER met2 ;
        RECT 2618.410 1492.755 2618.690 1493.125 ;
        RECT 2618.480 1449.070 2618.620 1492.755 ;
        RECT 2618.420 1448.750 2618.680 1449.070 ;
        RECT 2900.860 1448.750 2901.120 1449.070 ;
        RECT 2900.920 1446.885 2901.060 1448.750 ;
        RECT 2900.850 1446.515 2901.130 1446.885 ;
      LAYER via2 ;
        RECT 2618.410 1492.800 2618.690 1493.080 ;
        RECT 2900.850 1446.560 2901.130 1446.840 ;
      LAYER met3 ;
        RECT 2606.000 1493.090 2610.000 1493.480 ;
        RECT 2618.385 1493.090 2618.715 1493.105 ;
        RECT 2606.000 1492.880 2618.715 1493.090 ;
        RECT 2609.580 1492.790 2618.715 1492.880 ;
        RECT 2618.385 1492.775 2618.715 1492.790 ;
        RECT 2900.825 1446.850 2901.155 1446.865 ;
        RECT 2917.600 1446.850 2924.800 1447.300 ;
        RECT 2900.825 1446.550 2924.800 1446.850 ;
        RECT 2900.825 1446.535 2901.155 1446.550 ;
        RECT 2917.600 1446.100 2924.800 1446.550 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2617.010 1683.580 2617.330 1683.640 ;
        RECT 2900.830 1683.580 2901.150 1683.640 ;
        RECT 2617.010 1683.440 2901.150 1683.580 ;
        RECT 2617.010 1683.380 2617.330 1683.440 ;
        RECT 2900.830 1683.380 2901.150 1683.440 ;
      LAYER via ;
        RECT 2617.040 1683.380 2617.300 1683.640 ;
        RECT 2900.860 1683.380 2901.120 1683.640 ;
      LAYER met2 ;
        RECT 2617.030 1692.675 2617.310 1693.045 ;
        RECT 2617.100 1683.670 2617.240 1692.675 ;
        RECT 2617.040 1683.350 2617.300 1683.670 ;
        RECT 2900.860 1683.350 2901.120 1683.670 ;
        RECT 2900.920 1681.485 2901.060 1683.350 ;
        RECT 2900.850 1681.115 2901.130 1681.485 ;
      LAYER via2 ;
        RECT 2617.030 1692.720 2617.310 1693.000 ;
        RECT 2900.850 1681.160 2901.130 1681.440 ;
      LAYER met3 ;
        RECT 2606.000 1693.010 2610.000 1693.400 ;
        RECT 2617.005 1693.010 2617.335 1693.025 ;
        RECT 2606.000 1692.800 2617.335 1693.010 ;
        RECT 2609.580 1692.710 2617.335 1692.800 ;
        RECT 2617.005 1692.695 2617.335 1692.710 ;
        RECT 2900.825 1681.450 2901.155 1681.465 ;
        RECT 2917.600 1681.450 2924.800 1681.900 ;
        RECT 2900.825 1681.150 2924.800 1681.450 ;
        RECT 2900.825 1681.135 2901.155 1681.150 ;
        RECT 2917.600 1680.700 2924.800 1681.150 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.630 1911.380 2615.950 1911.440 ;
        RECT 2900.830 1911.380 2901.150 1911.440 ;
        RECT 2615.630 1911.240 2901.150 1911.380 ;
        RECT 2615.630 1911.180 2615.950 1911.240 ;
        RECT 2900.830 1911.180 2901.150 1911.240 ;
      LAYER via ;
        RECT 2615.660 1911.180 2615.920 1911.440 ;
        RECT 2900.860 1911.180 2901.120 1911.440 ;
      LAYER met2 ;
        RECT 2900.850 1915.715 2901.130 1916.085 ;
        RECT 2900.920 1911.470 2901.060 1915.715 ;
        RECT 2615.660 1911.150 2615.920 1911.470 ;
        RECT 2900.860 1911.150 2901.120 1911.470 ;
        RECT 2615.720 1893.645 2615.860 1911.150 ;
        RECT 2615.650 1893.275 2615.930 1893.645 ;
      LAYER via2 ;
        RECT 2900.850 1915.760 2901.130 1916.040 ;
        RECT 2615.650 1893.320 2615.930 1893.600 ;
      LAYER met3 ;
        RECT 2900.825 1916.050 2901.155 1916.065 ;
        RECT 2917.600 1916.050 2924.800 1916.500 ;
        RECT 2900.825 1915.750 2924.800 1916.050 ;
        RECT 2900.825 1915.735 2901.155 1915.750 ;
        RECT 2917.600 1915.300 2924.800 1915.750 ;
        RECT 2606.000 1893.610 2610.000 1894.000 ;
        RECT 2615.625 1893.610 2615.955 1893.625 ;
        RECT 2606.000 1893.400 2615.955 1893.610 ;
        RECT 2609.580 1893.310 2615.955 1893.400 ;
        RECT 2615.625 1893.295 2615.955 1893.310 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2145.980 2618.710 2146.040 ;
        RECT 2900.830 2145.980 2901.150 2146.040 ;
        RECT 2618.390 2145.840 2901.150 2145.980 ;
        RECT 2618.390 2145.780 2618.710 2145.840 ;
        RECT 2900.830 2145.780 2901.150 2145.840 ;
      LAYER via ;
        RECT 2618.420 2145.780 2618.680 2146.040 ;
        RECT 2900.860 2145.780 2901.120 2146.040 ;
      LAYER met2 ;
        RECT 2900.850 2150.315 2901.130 2150.685 ;
        RECT 2900.920 2146.070 2901.060 2150.315 ;
        RECT 2618.420 2145.750 2618.680 2146.070 ;
        RECT 2900.860 2145.750 2901.120 2146.070 ;
        RECT 2618.480 2093.565 2618.620 2145.750 ;
        RECT 2618.410 2093.195 2618.690 2093.565 ;
      LAYER via2 ;
        RECT 2900.850 2150.360 2901.130 2150.640 ;
        RECT 2618.410 2093.240 2618.690 2093.520 ;
      LAYER met3 ;
        RECT 2900.825 2150.650 2901.155 2150.665 ;
        RECT 2917.600 2150.650 2924.800 2151.100 ;
        RECT 2900.825 2150.350 2924.800 2150.650 ;
        RECT 2900.825 2150.335 2901.155 2150.350 ;
        RECT 2917.600 2149.900 2924.800 2150.350 ;
        RECT 2606.000 2093.530 2610.000 2093.920 ;
        RECT 2618.385 2093.530 2618.715 2093.545 ;
        RECT 2606.000 2093.320 2618.715 2093.530 ;
        RECT 2609.580 2093.230 2618.715 2093.320 ;
        RECT 2618.385 2093.215 2618.715 2093.230 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.310 200.160 2619.630 200.220 ;
        RECT 2900.830 200.160 2901.150 200.220 ;
        RECT 2619.310 200.020 2901.150 200.160 ;
        RECT 2619.310 199.960 2619.630 200.020 ;
        RECT 2900.830 199.960 2901.150 200.020 ;
      LAYER via ;
        RECT 2619.340 199.960 2619.600 200.220 ;
        RECT 2900.860 199.960 2901.120 200.220 ;
      LAYER met2 ;
        RECT 2619.330 426.515 2619.610 426.885 ;
        RECT 2619.400 200.250 2619.540 426.515 ;
        RECT 2619.340 199.930 2619.600 200.250 ;
        RECT 2900.860 199.930 2901.120 200.250 ;
        RECT 2900.920 195.685 2901.060 199.930 ;
        RECT 2900.850 195.315 2901.130 195.685 ;
      LAYER via2 ;
        RECT 2619.330 426.560 2619.610 426.840 ;
        RECT 2900.850 195.360 2901.130 195.640 ;
      LAYER met3 ;
        RECT 2606.000 426.850 2610.000 427.240 ;
        RECT 2619.305 426.850 2619.635 426.865 ;
        RECT 2606.000 426.640 2619.635 426.850 ;
        RECT 2609.580 426.550 2619.635 426.640 ;
        RECT 2619.305 426.535 2619.635 426.550 ;
        RECT 2900.825 195.650 2901.155 195.665 ;
        RECT 2917.600 195.650 2924.800 196.100 ;
        RECT 2900.825 195.350 2924.800 195.650 ;
        RECT 2900.825 195.335 2901.155 195.350 ;
        RECT 2917.600 194.900 2924.800 195.350 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2539.360 2618.710 2539.420 ;
        RECT 2900.830 2539.360 2901.150 2539.420 ;
        RECT 2618.390 2539.220 2901.150 2539.360 ;
        RECT 2618.390 2539.160 2618.710 2539.220 ;
        RECT 2900.830 2539.160 2901.150 2539.220 ;
      LAYER via ;
        RECT 2618.420 2539.160 2618.680 2539.420 ;
        RECT 2900.860 2539.160 2901.120 2539.420 ;
      LAYER met2 ;
        RECT 2900.850 2541.315 2901.130 2541.685 ;
        RECT 2900.920 2539.450 2901.060 2541.315 ;
        RECT 2618.420 2539.130 2618.680 2539.450 ;
        RECT 2900.860 2539.130 2901.120 2539.450 ;
        RECT 2618.480 2426.765 2618.620 2539.130 ;
        RECT 2618.410 2426.395 2618.690 2426.765 ;
      LAYER via2 ;
        RECT 2900.850 2541.360 2901.130 2541.640 ;
        RECT 2618.410 2426.440 2618.690 2426.720 ;
      LAYER met3 ;
        RECT 2900.825 2541.650 2901.155 2541.665 ;
        RECT 2917.600 2541.650 2924.800 2542.100 ;
        RECT 2900.825 2541.350 2924.800 2541.650 ;
        RECT 2900.825 2541.335 2901.155 2541.350 ;
        RECT 2917.600 2540.900 2924.800 2541.350 ;
        RECT 2606.000 2426.730 2610.000 2427.120 ;
        RECT 2618.385 2426.730 2618.715 2426.745 ;
        RECT 2606.000 2426.520 2618.715 2426.730 ;
        RECT 2609.580 2426.430 2618.715 2426.520 ;
        RECT 2618.385 2426.415 2618.715 2426.430 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2773.960 2619.170 2774.020 ;
        RECT 2900.830 2773.960 2901.150 2774.020 ;
        RECT 2618.850 2773.820 2901.150 2773.960 ;
        RECT 2618.850 2773.760 2619.170 2773.820 ;
        RECT 2900.830 2773.760 2901.150 2773.820 ;
      LAYER via ;
        RECT 2618.880 2773.760 2619.140 2774.020 ;
        RECT 2900.860 2773.760 2901.120 2774.020 ;
      LAYER met2 ;
        RECT 2900.850 2775.915 2901.130 2776.285 ;
        RECT 2900.920 2774.050 2901.060 2775.915 ;
        RECT 2618.880 2773.730 2619.140 2774.050 ;
        RECT 2900.860 2773.730 2901.120 2774.050 ;
        RECT 2618.940 2626.685 2619.080 2773.730 ;
        RECT 2618.870 2626.315 2619.150 2626.685 ;
      LAYER via2 ;
        RECT 2900.850 2775.960 2901.130 2776.240 ;
        RECT 2618.870 2626.360 2619.150 2626.640 ;
      LAYER met3 ;
        RECT 2900.825 2776.250 2901.155 2776.265 ;
        RECT 2917.600 2776.250 2924.800 2776.700 ;
        RECT 2900.825 2775.950 2924.800 2776.250 ;
        RECT 2900.825 2775.935 2901.155 2775.950 ;
        RECT 2917.600 2775.500 2924.800 2775.950 ;
        RECT 2606.000 2626.650 2610.000 2627.040 ;
        RECT 2618.845 2626.650 2619.175 2626.665 ;
        RECT 2606.000 2626.440 2619.175 2626.650 ;
        RECT 2609.580 2626.350 2619.175 2626.440 ;
        RECT 2618.845 2626.335 2619.175 2626.350 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3008.560 2619.170 3008.620 ;
        RECT 2900.830 3008.560 2901.150 3008.620 ;
        RECT 2618.850 3008.420 2901.150 3008.560 ;
        RECT 2618.850 3008.360 2619.170 3008.420 ;
        RECT 2900.830 3008.360 2901.150 3008.420 ;
      LAYER via ;
        RECT 2618.880 3008.360 2619.140 3008.620 ;
        RECT 2900.860 3008.360 2901.120 3008.620 ;
      LAYER met2 ;
        RECT 2900.850 3010.515 2901.130 3010.885 ;
        RECT 2900.920 3008.650 2901.060 3010.515 ;
        RECT 2618.880 3008.330 2619.140 3008.650 ;
        RECT 2900.860 3008.330 2901.120 3008.650 ;
        RECT 2618.940 2826.605 2619.080 3008.330 ;
        RECT 2618.870 2826.235 2619.150 2826.605 ;
      LAYER via2 ;
        RECT 2900.850 3010.560 2901.130 3010.840 ;
        RECT 2618.870 2826.280 2619.150 2826.560 ;
      LAYER met3 ;
        RECT 2900.825 3010.850 2901.155 3010.865 ;
        RECT 2917.600 3010.850 2924.800 3011.300 ;
        RECT 2900.825 3010.550 2924.800 3010.850 ;
        RECT 2900.825 3010.535 2901.155 3010.550 ;
        RECT 2917.600 3010.100 2924.800 3010.550 ;
        RECT 2606.000 2826.570 2610.000 2826.960 ;
        RECT 2618.845 2826.570 2619.175 2826.585 ;
        RECT 2606.000 2826.360 2619.175 2826.570 ;
        RECT 2609.580 2826.270 2619.175 2826.360 ;
        RECT 2618.845 2826.255 2619.175 2826.270 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.630 3028.960 2615.950 3029.020 ;
        RECT 2901.750 3028.960 2902.070 3029.020 ;
        RECT 2615.630 3028.820 2902.070 3028.960 ;
        RECT 2615.630 3028.760 2615.950 3028.820 ;
        RECT 2901.750 3028.760 2902.070 3028.820 ;
      LAYER via ;
        RECT 2615.660 3028.760 2615.920 3029.020 ;
        RECT 2901.780 3028.760 2902.040 3029.020 ;
      LAYER met2 ;
        RECT 2901.770 3245.115 2902.050 3245.485 ;
        RECT 2901.840 3029.050 2901.980 3245.115 ;
        RECT 2615.660 3028.730 2615.920 3029.050 ;
        RECT 2901.780 3028.730 2902.040 3029.050 ;
        RECT 2615.720 3026.525 2615.860 3028.730 ;
        RECT 2615.650 3026.155 2615.930 3026.525 ;
      LAYER via2 ;
        RECT 2901.770 3245.160 2902.050 3245.440 ;
        RECT 2615.650 3026.200 2615.930 3026.480 ;
      LAYER met3 ;
        RECT 2901.745 3245.450 2902.075 3245.465 ;
        RECT 2917.600 3245.450 2924.800 3245.900 ;
        RECT 2901.745 3245.150 2924.800 3245.450 ;
        RECT 2901.745 3245.135 2902.075 3245.150 ;
        RECT 2917.600 3244.700 2924.800 3245.150 ;
        RECT 2606.000 3026.490 2610.000 3026.880 ;
        RECT 2615.625 3026.490 2615.955 3026.505 ;
        RECT 2606.000 3026.280 2615.955 3026.490 ;
        RECT 2609.580 3026.190 2615.955 3026.280 ;
        RECT 2615.625 3026.175 2615.955 3026.190 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 3477.760 2618.710 3477.820 ;
        RECT 2900.830 3477.760 2901.150 3477.820 ;
        RECT 2618.390 3477.620 2901.150 3477.760 ;
        RECT 2618.390 3477.560 2618.710 3477.620 ;
        RECT 2900.830 3477.560 2901.150 3477.620 ;
      LAYER via ;
        RECT 2618.420 3477.560 2618.680 3477.820 ;
        RECT 2900.860 3477.560 2901.120 3477.820 ;
      LAYER met2 ;
        RECT 2900.850 3479.715 2901.130 3480.085 ;
        RECT 2900.920 3477.850 2901.060 3479.715 ;
        RECT 2618.420 3477.530 2618.680 3477.850 ;
        RECT 2900.860 3477.530 2901.120 3477.850 ;
        RECT 2618.480 3226.445 2618.620 3477.530 ;
        RECT 2618.410 3226.075 2618.690 3226.445 ;
      LAYER via2 ;
        RECT 2900.850 3479.760 2901.130 3480.040 ;
        RECT 2618.410 3226.120 2618.690 3226.400 ;
      LAYER met3 ;
        RECT 2900.825 3480.050 2901.155 3480.065 ;
        RECT 2917.600 3480.050 2924.800 3480.500 ;
        RECT 2900.825 3479.750 2924.800 3480.050 ;
        RECT 2900.825 3479.735 2901.155 3479.750 ;
        RECT 2917.600 3479.300 2924.800 3479.750 ;
        RECT 2606.000 3226.410 2610.000 3226.800 ;
        RECT 2618.385 3226.410 2618.715 3226.425 ;
        RECT 2606.000 3226.200 2618.715 3226.410 ;
        RECT 2609.580 3226.110 2618.715 3226.200 ;
        RECT 2618.385 3226.095 2618.715 3226.110 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2400.810 3502.240 2401.130 3502.300 ;
        RECT 2649.210 3502.240 2649.530 3502.300 ;
        RECT 2400.810 3502.100 2649.530 3502.240 ;
        RECT 2400.810 3502.040 2401.130 3502.100 ;
        RECT 2649.210 3502.040 2649.530 3502.100 ;
        RECT 2396.670 3277.500 2396.990 3277.560 ;
        RECT 2400.810 3277.500 2401.130 3277.560 ;
        RECT 2396.670 3277.360 2401.130 3277.500 ;
        RECT 2396.670 3277.300 2396.990 3277.360 ;
        RECT 2400.810 3277.300 2401.130 3277.360 ;
      LAYER via ;
        RECT 2400.840 3502.040 2401.100 3502.300 ;
        RECT 2649.240 3502.040 2649.500 3502.300 ;
        RECT 2396.700 3277.300 2396.960 3277.560 ;
        RECT 2400.840 3277.300 2401.100 3277.560 ;
      LAYER met2 ;
        RECT 2649.090 3517.600 2649.650 3524.800 ;
        RECT 2649.300 3502.330 2649.440 3517.600 ;
        RECT 2400.840 3502.010 2401.100 3502.330 ;
        RECT 2649.240 3502.010 2649.500 3502.330 ;
        RECT 2400.900 3277.590 2401.040 3502.010 ;
        RECT 2396.700 3277.270 2396.960 3277.590 ;
        RECT 2400.840 3277.270 2401.100 3277.590 ;
        RECT 2396.760 3260.000 2396.900 3277.270 ;
        RECT 2396.650 3256.000 2396.930 3260.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2145.510 3502.240 2145.830 3502.300 ;
        RECT 2324.910 3502.240 2325.230 3502.300 ;
        RECT 2145.510 3502.100 2325.230 3502.240 ;
        RECT 2145.510 3502.040 2145.830 3502.100 ;
        RECT 2324.910 3502.040 2325.230 3502.100 ;
        RECT 2140.910 3277.500 2141.230 3277.560 ;
        RECT 2145.510 3277.500 2145.830 3277.560 ;
        RECT 2140.910 3277.360 2145.830 3277.500 ;
        RECT 2140.910 3277.300 2141.230 3277.360 ;
        RECT 2145.510 3277.300 2145.830 3277.360 ;
      LAYER via ;
        RECT 2145.540 3502.040 2145.800 3502.300 ;
        RECT 2324.940 3502.040 2325.200 3502.300 ;
        RECT 2140.940 3277.300 2141.200 3277.560 ;
        RECT 2145.540 3277.300 2145.800 3277.560 ;
      LAYER met2 ;
        RECT 2324.790 3517.600 2325.350 3524.800 ;
        RECT 2325.000 3502.330 2325.140 3517.600 ;
        RECT 2145.540 3502.010 2145.800 3502.330 ;
        RECT 2324.940 3502.010 2325.200 3502.330 ;
        RECT 2145.600 3277.590 2145.740 3502.010 ;
        RECT 2140.940 3277.270 2141.200 3277.590 ;
        RECT 2145.540 3277.270 2145.800 3277.590 ;
        RECT 2141.000 3260.000 2141.140 3277.270 ;
        RECT 2140.890 3256.000 2141.170 3260.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1890.210 3501.560 1890.530 3501.620 ;
        RECT 2000.610 3501.560 2000.930 3501.620 ;
        RECT 1890.210 3501.420 2000.930 3501.560 ;
        RECT 1890.210 3501.360 1890.530 3501.420 ;
        RECT 2000.610 3501.360 2000.930 3501.420 ;
        RECT 1885.610 3277.500 1885.930 3277.560 ;
        RECT 1890.210 3277.500 1890.530 3277.560 ;
        RECT 1885.610 3277.360 1890.530 3277.500 ;
        RECT 1885.610 3277.300 1885.930 3277.360 ;
        RECT 1890.210 3277.300 1890.530 3277.360 ;
      LAYER via ;
        RECT 1890.240 3501.360 1890.500 3501.620 ;
        RECT 2000.640 3501.360 2000.900 3501.620 ;
        RECT 1885.640 3277.300 1885.900 3277.560 ;
        RECT 1890.240 3277.300 1890.500 3277.560 ;
      LAYER met2 ;
        RECT 2000.490 3517.600 2001.050 3524.800 ;
        RECT 2000.700 3501.650 2000.840 3517.600 ;
        RECT 1890.240 3501.330 1890.500 3501.650 ;
        RECT 2000.640 3501.330 2000.900 3501.650 ;
        RECT 1890.300 3277.590 1890.440 3501.330 ;
        RECT 1885.640 3277.270 1885.900 3277.590 ;
        RECT 1890.240 3277.270 1890.500 3277.590 ;
        RECT 1885.700 3260.000 1885.840 3277.270 ;
        RECT 1885.590 3256.000 1885.870 3260.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1634.910 3498.500 1635.230 3498.560 ;
        RECT 1675.850 3498.500 1676.170 3498.560 ;
        RECT 1634.910 3498.360 1676.170 3498.500 ;
        RECT 1634.910 3498.300 1635.230 3498.360 ;
        RECT 1675.850 3498.300 1676.170 3498.360 ;
        RECT 1629.850 3275.800 1630.170 3275.860 ;
        RECT 1634.910 3275.800 1635.230 3275.860 ;
        RECT 1629.850 3275.660 1635.230 3275.800 ;
        RECT 1629.850 3275.600 1630.170 3275.660 ;
        RECT 1634.910 3275.600 1635.230 3275.660 ;
      LAYER via ;
        RECT 1634.940 3498.300 1635.200 3498.560 ;
        RECT 1675.880 3498.300 1676.140 3498.560 ;
        RECT 1629.880 3275.600 1630.140 3275.860 ;
        RECT 1634.940 3275.600 1635.200 3275.860 ;
      LAYER met2 ;
        RECT 1675.730 3517.600 1676.290 3524.800 ;
        RECT 1675.940 3498.590 1676.080 3517.600 ;
        RECT 1634.940 3498.270 1635.200 3498.590 ;
        RECT 1675.880 3498.270 1676.140 3498.590 ;
        RECT 1635.000 3275.890 1635.140 3498.270 ;
        RECT 1629.880 3275.570 1630.140 3275.890 ;
        RECT 1634.940 3275.570 1635.200 3275.890 ;
        RECT 1629.940 3260.000 1630.080 3275.570 ;
        RECT 1629.830 3256.000 1630.110 3260.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1351.625 3429.325 1351.795 3477.435 ;
      LAYER mcon ;
        RECT 1351.625 3477.265 1351.795 3477.435 ;
      LAYER met1 ;
        RECT 1351.565 3477.420 1351.855 3477.465 ;
        RECT 1352.010 3477.420 1352.330 3477.480 ;
        RECT 1351.565 3477.280 1352.330 3477.420 ;
        RECT 1351.565 3477.235 1351.855 3477.280 ;
        RECT 1352.010 3477.220 1352.330 3477.280 ;
        RECT 1351.550 3429.480 1351.870 3429.540 ;
        RECT 1351.355 3429.340 1351.870 3429.480 ;
        RECT 1351.550 3429.280 1351.870 3429.340 ;
        RECT 1351.550 3395.140 1351.870 3395.200 ;
        RECT 1351.180 3395.000 1351.870 3395.140 ;
        RECT 1351.180 3394.860 1351.320 3395.000 ;
        RECT 1351.550 3394.940 1351.870 3395.000 ;
        RECT 1351.090 3394.600 1351.410 3394.860 ;
        RECT 1351.090 3367.600 1351.410 3367.660 ;
        RECT 1352.010 3367.600 1352.330 3367.660 ;
        RECT 1351.090 3367.460 1352.330 3367.600 ;
        RECT 1351.090 3367.400 1351.410 3367.460 ;
        RECT 1352.010 3367.400 1352.330 3367.460 ;
        RECT 1351.090 3277.500 1351.410 3277.560 ;
        RECT 1374.550 3277.500 1374.870 3277.560 ;
        RECT 1351.090 3277.360 1374.870 3277.500 ;
        RECT 1351.090 3277.300 1351.410 3277.360 ;
        RECT 1374.550 3277.300 1374.870 3277.360 ;
      LAYER via ;
        RECT 1352.040 3477.220 1352.300 3477.480 ;
        RECT 1351.580 3429.280 1351.840 3429.540 ;
        RECT 1351.580 3394.940 1351.840 3395.200 ;
        RECT 1351.120 3394.600 1351.380 3394.860 ;
        RECT 1351.120 3367.400 1351.380 3367.660 ;
        RECT 1352.040 3367.400 1352.300 3367.660 ;
        RECT 1351.120 3277.300 1351.380 3277.560 ;
        RECT 1374.580 3277.300 1374.840 3277.560 ;
      LAYER met2 ;
        RECT 1351.430 3517.600 1351.990 3524.800 ;
        RECT 1351.640 3517.370 1351.780 3517.600 ;
        RECT 1351.640 3517.230 1352.240 3517.370 ;
        RECT 1352.100 3477.510 1352.240 3517.230 ;
        RECT 1352.040 3477.190 1352.300 3477.510 ;
        RECT 1351.580 3429.250 1351.840 3429.570 ;
        RECT 1351.640 3395.230 1351.780 3429.250 ;
        RECT 1351.580 3394.910 1351.840 3395.230 ;
        RECT 1351.120 3394.570 1351.380 3394.890 ;
        RECT 1351.180 3367.690 1351.320 3394.570 ;
        RECT 1351.120 3367.370 1351.380 3367.690 ;
        RECT 1352.040 3367.370 1352.300 3367.690 ;
        RECT 1352.100 3318.810 1352.240 3367.370 ;
        RECT 1351.180 3318.670 1352.240 3318.810 ;
        RECT 1351.180 3277.590 1351.320 3318.670 ;
        RECT 1351.120 3277.270 1351.380 3277.590 ;
        RECT 1374.580 3277.270 1374.840 3277.590 ;
        RECT 1374.640 3260.000 1374.780 3277.270 ;
        RECT 1374.530 3256.000 1374.810 3260.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 434.760 2619.170 434.820 ;
        RECT 2900.830 434.760 2901.150 434.820 ;
        RECT 2618.850 434.620 2901.150 434.760 ;
        RECT 2618.850 434.560 2619.170 434.620 ;
        RECT 2900.830 434.560 2901.150 434.620 ;
      LAYER via ;
        RECT 2618.880 434.560 2619.140 434.820 ;
        RECT 2900.860 434.560 2901.120 434.820 ;
      LAYER met2 ;
        RECT 2618.870 626.435 2619.150 626.805 ;
        RECT 2618.940 434.850 2619.080 626.435 ;
        RECT 2618.880 434.530 2619.140 434.850 ;
        RECT 2900.860 434.530 2901.120 434.850 ;
        RECT 2900.920 430.285 2901.060 434.530 ;
        RECT 2900.850 429.915 2901.130 430.285 ;
      LAYER via2 ;
        RECT 2618.870 626.480 2619.150 626.760 ;
        RECT 2900.850 429.960 2901.130 430.240 ;
      LAYER met3 ;
        RECT 2606.000 626.770 2610.000 627.160 ;
        RECT 2618.845 626.770 2619.175 626.785 ;
        RECT 2606.000 626.560 2619.175 626.770 ;
        RECT 2609.580 626.470 2619.175 626.560 ;
        RECT 2618.845 626.455 2619.175 626.470 ;
        RECT 2900.825 430.250 2901.155 430.265 ;
        RECT 2917.600 430.250 2924.800 430.700 ;
        RECT 2900.825 429.950 2924.800 430.250 ;
        RECT 2900.825 429.935 2901.155 429.950 ;
        RECT 2917.600 429.500 2924.800 429.950 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1027.785 3422.525 1027.955 3470.635 ;
      LAYER mcon ;
        RECT 1027.785 3470.465 1027.955 3470.635 ;
      LAYER met1 ;
        RECT 1027.725 3470.620 1028.015 3470.665 ;
        RECT 1028.170 3470.620 1028.490 3470.680 ;
        RECT 1027.725 3470.480 1028.490 3470.620 ;
        RECT 1027.725 3470.435 1028.015 3470.480 ;
        RECT 1028.170 3470.420 1028.490 3470.480 ;
        RECT 1027.710 3422.680 1028.030 3422.740 ;
        RECT 1027.515 3422.540 1028.030 3422.680 ;
        RECT 1027.710 3422.480 1028.030 3422.540 ;
        RECT 1027.710 3395.140 1028.030 3395.200 ;
        RECT 1027.340 3395.000 1028.030 3395.140 ;
        RECT 1027.340 3394.860 1027.480 3395.000 ;
        RECT 1027.710 3394.940 1028.030 3395.000 ;
        RECT 1027.250 3394.600 1027.570 3394.860 ;
        RECT 1027.250 3346.860 1027.570 3346.920 ;
        RECT 1026.880 3346.720 1027.570 3346.860 ;
        RECT 1026.880 3346.580 1027.020 3346.720 ;
        RECT 1027.250 3346.660 1027.570 3346.720 ;
        RECT 1026.790 3346.320 1027.110 3346.580 ;
        RECT 1026.790 3298.580 1027.110 3298.640 ;
        RECT 1026.420 3298.440 1027.110 3298.580 ;
        RECT 1026.420 3298.300 1026.560 3298.440 ;
        RECT 1026.790 3298.380 1027.110 3298.440 ;
        RECT 1026.330 3298.040 1026.650 3298.300 ;
        RECT 1026.330 3274.440 1026.650 3274.500 ;
        RECT 1118.790 3274.440 1119.110 3274.500 ;
        RECT 1026.330 3274.300 1119.110 3274.440 ;
        RECT 1026.330 3274.240 1026.650 3274.300 ;
        RECT 1118.790 3274.240 1119.110 3274.300 ;
      LAYER via ;
        RECT 1028.200 3470.420 1028.460 3470.680 ;
        RECT 1027.740 3422.480 1028.000 3422.740 ;
        RECT 1027.740 3394.940 1028.000 3395.200 ;
        RECT 1027.280 3394.600 1027.540 3394.860 ;
        RECT 1027.280 3346.660 1027.540 3346.920 ;
        RECT 1026.820 3346.320 1027.080 3346.580 ;
        RECT 1026.820 3298.380 1027.080 3298.640 ;
        RECT 1026.360 3298.040 1026.620 3298.300 ;
        RECT 1026.360 3274.240 1026.620 3274.500 ;
        RECT 1118.820 3274.240 1119.080 3274.500 ;
      LAYER met2 ;
        RECT 1027.130 3517.600 1027.690 3524.800 ;
        RECT 1027.340 3492.210 1027.480 3517.600 ;
        RECT 1027.340 3492.070 1028.400 3492.210 ;
        RECT 1028.260 3470.710 1028.400 3492.070 ;
        RECT 1028.200 3470.390 1028.460 3470.710 ;
        RECT 1027.740 3422.450 1028.000 3422.770 ;
        RECT 1027.800 3395.230 1027.940 3422.450 ;
        RECT 1027.740 3394.910 1028.000 3395.230 ;
        RECT 1027.280 3394.570 1027.540 3394.890 ;
        RECT 1027.340 3346.950 1027.480 3394.570 ;
        RECT 1027.280 3346.630 1027.540 3346.950 ;
        RECT 1026.820 3346.290 1027.080 3346.610 ;
        RECT 1026.880 3298.670 1027.020 3346.290 ;
        RECT 1026.820 3298.350 1027.080 3298.670 ;
        RECT 1026.360 3298.010 1026.620 3298.330 ;
        RECT 1026.420 3274.530 1026.560 3298.010 ;
        RECT 1026.360 3274.210 1026.620 3274.530 ;
        RECT 1118.820 3274.210 1119.080 3274.530 ;
        RECT 1118.880 3260.000 1119.020 3274.210 ;
        RECT 1118.770 3256.000 1119.050 3260.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 702.565 3381.045 702.735 3429.155 ;
      LAYER mcon ;
        RECT 702.565 3428.985 702.735 3429.155 ;
      LAYER met1 ;
        RECT 702.030 3477.760 702.350 3477.820 ;
        RECT 702.490 3477.760 702.810 3477.820 ;
        RECT 702.030 3477.620 702.810 3477.760 ;
        RECT 702.030 3477.560 702.350 3477.620 ;
        RECT 702.490 3477.560 702.810 3477.620 ;
        RECT 702.030 3443.080 702.350 3443.140 ;
        RECT 702.950 3443.080 703.270 3443.140 ;
        RECT 702.030 3442.940 703.270 3443.080 ;
        RECT 702.030 3442.880 702.350 3442.940 ;
        RECT 702.950 3442.880 703.270 3442.940 ;
        RECT 702.505 3429.140 702.795 3429.185 ;
        RECT 702.950 3429.140 703.270 3429.200 ;
        RECT 702.505 3429.000 703.270 3429.140 ;
        RECT 702.505 3428.955 702.795 3429.000 ;
        RECT 702.950 3428.940 703.270 3429.000 ;
        RECT 702.490 3381.200 702.810 3381.260 ;
        RECT 702.295 3381.060 702.810 3381.200 ;
        RECT 702.490 3381.000 702.810 3381.060 ;
        RECT 702.490 3367.600 702.810 3367.660 ;
        RECT 703.410 3367.600 703.730 3367.660 ;
        RECT 702.490 3367.460 703.730 3367.600 ;
        RECT 702.490 3367.400 702.810 3367.460 ;
        RECT 703.410 3367.400 703.730 3367.460 ;
        RECT 702.490 3274.100 702.810 3274.160 ;
        RECT 863.490 3274.100 863.810 3274.160 ;
        RECT 702.490 3273.960 863.810 3274.100 ;
        RECT 702.490 3273.900 702.810 3273.960 ;
        RECT 863.490 3273.900 863.810 3273.960 ;
      LAYER via ;
        RECT 702.060 3477.560 702.320 3477.820 ;
        RECT 702.520 3477.560 702.780 3477.820 ;
        RECT 702.060 3442.880 702.320 3443.140 ;
        RECT 702.980 3442.880 703.240 3443.140 ;
        RECT 702.980 3428.940 703.240 3429.200 ;
        RECT 702.520 3381.000 702.780 3381.260 ;
        RECT 702.520 3367.400 702.780 3367.660 ;
        RECT 703.440 3367.400 703.700 3367.660 ;
        RECT 702.520 3273.900 702.780 3274.160 ;
        RECT 863.520 3273.900 863.780 3274.160 ;
      LAYER met2 ;
        RECT 702.370 3517.600 702.930 3524.800 ;
        RECT 702.580 3477.850 702.720 3517.600 ;
        RECT 702.060 3477.530 702.320 3477.850 ;
        RECT 702.520 3477.530 702.780 3477.850 ;
        RECT 702.120 3443.170 702.260 3477.530 ;
        RECT 702.060 3442.850 702.320 3443.170 ;
        RECT 702.980 3442.850 703.240 3443.170 ;
        RECT 703.040 3429.230 703.180 3442.850 ;
        RECT 702.980 3428.910 703.240 3429.230 ;
        RECT 702.520 3380.970 702.780 3381.290 ;
        RECT 702.580 3367.690 702.720 3380.970 ;
        RECT 702.520 3367.370 702.780 3367.690 ;
        RECT 703.440 3367.370 703.700 3367.690 ;
        RECT 703.500 3318.810 703.640 3367.370 ;
        RECT 702.580 3318.670 703.640 3318.810 ;
        RECT 702.580 3274.190 702.720 3318.670 ;
        RECT 702.520 3273.870 702.780 3274.190 ;
        RECT 863.520 3273.870 863.780 3274.190 ;
        RECT 863.580 3260.000 863.720 3273.870 ;
        RECT 863.470 3256.000 863.750 3260.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 378.265 3470.805 378.435 3491.715 ;
        RECT 377.805 3284.485 377.975 3332.595 ;
      LAYER mcon ;
        RECT 378.265 3491.545 378.435 3491.715 ;
        RECT 377.805 3332.425 377.975 3332.595 ;
      LAYER met1 ;
        RECT 378.190 3491.700 378.510 3491.760 ;
        RECT 377.995 3491.560 378.510 3491.700 ;
        RECT 378.190 3491.500 378.510 3491.560 ;
        RECT 378.190 3470.960 378.510 3471.020 ;
        RECT 377.995 3470.820 378.510 3470.960 ;
        RECT 378.190 3470.760 378.510 3470.820 ;
        RECT 378.190 3443.420 378.510 3443.480 ;
        RECT 377.820 3443.280 378.510 3443.420 ;
        RECT 377.820 3443.140 377.960 3443.280 ;
        RECT 378.190 3443.220 378.510 3443.280 ;
        RECT 377.730 3442.880 378.050 3443.140 ;
        RECT 377.730 3395.140 378.050 3395.200 ;
        RECT 377.360 3395.000 378.050 3395.140 ;
        RECT 377.360 3394.860 377.500 3395.000 ;
        RECT 377.730 3394.940 378.050 3395.000 ;
        RECT 377.270 3394.600 377.590 3394.860 ;
        RECT 377.270 3346.520 377.590 3346.580 ;
        RECT 378.190 3346.520 378.510 3346.580 ;
        RECT 377.270 3346.380 378.510 3346.520 ;
        RECT 377.270 3346.320 377.590 3346.380 ;
        RECT 378.190 3346.320 378.510 3346.380 ;
        RECT 377.745 3332.580 378.035 3332.625 ;
        RECT 378.190 3332.580 378.510 3332.640 ;
        RECT 377.745 3332.440 378.510 3332.580 ;
        RECT 377.745 3332.395 378.035 3332.440 ;
        RECT 378.190 3332.380 378.510 3332.440 ;
        RECT 377.730 3284.640 378.050 3284.700 ;
        RECT 377.535 3284.500 378.050 3284.640 ;
        RECT 377.730 3284.440 378.050 3284.500 ;
        RECT 377.730 3274.100 378.050 3274.160 ;
        RECT 607.730 3274.100 608.050 3274.160 ;
        RECT 377.730 3273.960 608.050 3274.100 ;
        RECT 377.730 3273.900 378.050 3273.960 ;
        RECT 607.730 3273.900 608.050 3273.960 ;
      LAYER via ;
        RECT 378.220 3491.500 378.480 3491.760 ;
        RECT 378.220 3470.760 378.480 3471.020 ;
        RECT 378.220 3443.220 378.480 3443.480 ;
        RECT 377.760 3442.880 378.020 3443.140 ;
        RECT 377.760 3394.940 378.020 3395.200 ;
        RECT 377.300 3394.600 377.560 3394.860 ;
        RECT 377.300 3346.320 377.560 3346.580 ;
        RECT 378.220 3346.320 378.480 3346.580 ;
        RECT 378.220 3332.380 378.480 3332.640 ;
        RECT 377.760 3284.440 378.020 3284.700 ;
        RECT 377.760 3273.900 378.020 3274.160 ;
        RECT 607.760 3273.900 608.020 3274.160 ;
      LAYER met2 ;
        RECT 378.070 3517.600 378.630 3524.800 ;
        RECT 378.280 3491.790 378.420 3517.600 ;
        RECT 378.220 3491.470 378.480 3491.790 ;
        RECT 378.220 3470.730 378.480 3471.050 ;
        RECT 378.280 3443.510 378.420 3470.730 ;
        RECT 378.220 3443.190 378.480 3443.510 ;
        RECT 377.760 3442.850 378.020 3443.170 ;
        RECT 377.820 3395.230 377.960 3442.850 ;
        RECT 377.760 3394.910 378.020 3395.230 ;
        RECT 377.300 3394.570 377.560 3394.890 ;
        RECT 377.360 3346.610 377.500 3394.570 ;
        RECT 377.300 3346.290 377.560 3346.610 ;
        RECT 378.220 3346.290 378.480 3346.610 ;
        RECT 378.280 3332.670 378.420 3346.290 ;
        RECT 378.220 3332.350 378.480 3332.670 ;
        RECT 377.760 3284.410 378.020 3284.730 ;
        RECT 377.820 3274.190 377.960 3284.410 ;
        RECT 377.760 3273.870 378.020 3274.190 ;
        RECT 607.760 3273.870 608.020 3274.190 ;
        RECT 607.820 3260.000 607.960 3273.870 ;
        RECT 607.710 3256.000 607.990 3260.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 53.965 3381.045 54.135 3429.155 ;
      LAYER mcon ;
        RECT 53.965 3428.985 54.135 3429.155 ;
      LAYER met1 ;
        RECT 53.430 3477.760 53.750 3477.820 ;
        RECT 53.890 3477.760 54.210 3477.820 ;
        RECT 53.430 3477.620 54.210 3477.760 ;
        RECT 53.430 3477.560 53.750 3477.620 ;
        RECT 53.890 3477.560 54.210 3477.620 ;
        RECT 53.430 3443.080 53.750 3443.140 ;
        RECT 54.350 3443.080 54.670 3443.140 ;
        RECT 53.430 3442.940 54.670 3443.080 ;
        RECT 53.430 3442.880 53.750 3442.940 ;
        RECT 54.350 3442.880 54.670 3442.940 ;
        RECT 53.905 3429.140 54.195 3429.185 ;
        RECT 54.350 3429.140 54.670 3429.200 ;
        RECT 53.905 3429.000 54.670 3429.140 ;
        RECT 53.905 3428.955 54.195 3429.000 ;
        RECT 54.350 3428.940 54.670 3429.000 ;
        RECT 53.890 3381.200 54.210 3381.260 ;
        RECT 53.695 3381.060 54.210 3381.200 ;
        RECT 53.890 3381.000 54.210 3381.060 ;
        RECT 53.890 3367.600 54.210 3367.660 ;
        RECT 54.810 3367.600 55.130 3367.660 ;
        RECT 53.890 3367.460 55.130 3367.600 ;
        RECT 53.890 3367.400 54.210 3367.460 ;
        RECT 54.810 3367.400 55.130 3367.460 ;
        RECT 53.890 3274.100 54.210 3274.160 ;
        RECT 352.430 3274.100 352.750 3274.160 ;
        RECT 53.890 3273.960 352.750 3274.100 ;
        RECT 53.890 3273.900 54.210 3273.960 ;
        RECT 352.430 3273.900 352.750 3273.960 ;
      LAYER via ;
        RECT 53.460 3477.560 53.720 3477.820 ;
        RECT 53.920 3477.560 54.180 3477.820 ;
        RECT 53.460 3442.880 53.720 3443.140 ;
        RECT 54.380 3442.880 54.640 3443.140 ;
        RECT 54.380 3428.940 54.640 3429.200 ;
        RECT 53.920 3381.000 54.180 3381.260 ;
        RECT 53.920 3367.400 54.180 3367.660 ;
        RECT 54.840 3367.400 55.100 3367.660 ;
        RECT 53.920 3273.900 54.180 3274.160 ;
        RECT 352.460 3273.900 352.720 3274.160 ;
      LAYER met2 ;
        RECT 53.770 3517.600 54.330 3524.800 ;
        RECT 53.980 3477.850 54.120 3517.600 ;
        RECT 53.460 3477.530 53.720 3477.850 ;
        RECT 53.920 3477.530 54.180 3477.850 ;
        RECT 53.520 3443.170 53.660 3477.530 ;
        RECT 53.460 3442.850 53.720 3443.170 ;
        RECT 54.380 3442.850 54.640 3443.170 ;
        RECT 54.440 3429.230 54.580 3442.850 ;
        RECT 54.380 3428.910 54.640 3429.230 ;
        RECT 53.920 3380.970 54.180 3381.290 ;
        RECT 53.980 3367.690 54.120 3380.970 ;
        RECT 53.920 3367.370 54.180 3367.690 ;
        RECT 54.840 3367.370 55.100 3367.690 ;
        RECT 54.900 3318.810 55.040 3367.370 ;
        RECT 53.980 3318.670 55.040 3318.810 ;
        RECT 53.980 3274.190 54.120 3318.670 ;
        RECT 53.920 3273.870 54.180 3274.190 ;
        RECT 352.460 3273.870 352.720 3274.190 ;
        RECT 352.520 3260.000 352.660 3273.870 ;
        RECT 352.410 3256.000 352.690 3260.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 3084.040 18.330 3084.100 ;
        RECT 296.770 3084.040 297.090 3084.100 ;
        RECT 18.010 3083.900 297.090 3084.040 ;
        RECT 18.010 3083.840 18.330 3083.900 ;
        RECT 296.770 3083.840 297.090 3083.900 ;
      LAYER via ;
        RECT 18.040 3083.840 18.300 3084.100 ;
        RECT 296.800 3083.840 297.060 3084.100 ;
      LAYER met2 ;
        RECT 18.030 3309.715 18.310 3310.085 ;
        RECT 18.100 3084.130 18.240 3309.715 ;
        RECT 18.040 3083.810 18.300 3084.130 ;
        RECT 296.800 3083.810 297.060 3084.130 ;
        RECT 296.860 3080.925 297.000 3083.810 ;
        RECT 296.790 3080.555 297.070 3080.925 ;
      LAYER via2 ;
        RECT 18.030 3309.760 18.310 3310.040 ;
        RECT 296.790 3080.600 297.070 3080.880 ;
      LAYER met3 ;
        RECT -4.800 3310.050 2.400 3310.500 ;
        RECT 18.005 3310.050 18.335 3310.065 ;
        RECT -4.800 3309.750 18.335 3310.050 ;
        RECT -4.800 3309.300 2.400 3309.750 ;
        RECT 18.005 3309.735 18.335 3309.750 ;
        RECT 296.765 3080.890 297.095 3080.905 ;
        RECT 310.000 3080.890 314.000 3081.280 ;
        RECT 296.765 3080.680 314.000 3080.890 ;
        RECT 296.765 3080.590 310.500 3080.680 ;
        RECT 296.765 3080.575 297.095 3080.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2870.180 17.870 2870.240 ;
        RECT 296.770 2870.180 297.090 2870.240 ;
        RECT 17.550 2870.040 297.090 2870.180 ;
        RECT 17.550 2869.980 17.870 2870.040 ;
        RECT 296.770 2869.980 297.090 2870.040 ;
      LAYER via ;
        RECT 17.580 2869.980 17.840 2870.240 ;
        RECT 296.800 2869.980 297.060 2870.240 ;
      LAYER met2 ;
        RECT 17.570 3058.115 17.850 3058.485 ;
        RECT 17.640 2870.270 17.780 3058.115 ;
        RECT 17.580 2869.950 17.840 2870.270 ;
        RECT 296.800 2869.950 297.060 2870.270 ;
        RECT 296.860 2866.725 297.000 2869.950 ;
        RECT 296.790 2866.355 297.070 2866.725 ;
      LAYER via2 ;
        RECT 17.570 3058.160 17.850 3058.440 ;
        RECT 296.790 2866.400 297.070 2866.680 ;
      LAYER met3 ;
        RECT -4.800 3058.450 2.400 3058.900 ;
        RECT 17.545 3058.450 17.875 3058.465 ;
        RECT -4.800 3058.150 17.875 3058.450 ;
        RECT -4.800 3057.700 2.400 3058.150 ;
        RECT 17.545 3058.135 17.875 3058.150 ;
        RECT 296.765 2866.690 297.095 2866.705 ;
        RECT 310.000 2866.690 314.000 2867.080 ;
        RECT 296.765 2866.480 314.000 2866.690 ;
        RECT 296.765 2866.390 310.500 2866.480 ;
        RECT 296.765 2866.375 297.095 2866.390 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2656.320 17.870 2656.380 ;
        RECT 296.770 2656.320 297.090 2656.380 ;
        RECT 17.550 2656.180 297.090 2656.320 ;
        RECT 17.550 2656.120 17.870 2656.180 ;
        RECT 296.770 2656.120 297.090 2656.180 ;
      LAYER via ;
        RECT 17.580 2656.120 17.840 2656.380 ;
        RECT 296.800 2656.120 297.060 2656.380 ;
      LAYER met2 ;
        RECT 17.570 2806.515 17.850 2806.885 ;
        RECT 17.640 2656.410 17.780 2806.515 ;
        RECT 17.580 2656.090 17.840 2656.410 ;
        RECT 296.800 2656.090 297.060 2656.410 ;
        RECT 296.860 2652.525 297.000 2656.090 ;
        RECT 296.790 2652.155 297.070 2652.525 ;
      LAYER via2 ;
        RECT 17.570 2806.560 17.850 2806.840 ;
        RECT 296.790 2652.200 297.070 2652.480 ;
      LAYER met3 ;
        RECT -4.800 2806.850 2.400 2807.300 ;
        RECT 17.545 2806.850 17.875 2806.865 ;
        RECT -4.800 2806.550 17.875 2806.850 ;
        RECT -4.800 2806.100 2.400 2806.550 ;
        RECT 17.545 2806.535 17.875 2806.550 ;
        RECT 296.765 2652.490 297.095 2652.505 ;
        RECT 310.000 2652.490 314.000 2652.880 ;
        RECT 296.765 2652.280 314.000 2652.490 ;
        RECT 296.765 2652.190 310.500 2652.280 ;
        RECT 296.765 2652.175 297.095 2652.190 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2442.460 17.870 2442.520 ;
        RECT 296.770 2442.460 297.090 2442.520 ;
        RECT 17.550 2442.320 297.090 2442.460 ;
        RECT 17.550 2442.260 17.870 2442.320 ;
        RECT 296.770 2442.260 297.090 2442.320 ;
      LAYER via ;
        RECT 17.580 2442.260 17.840 2442.520 ;
        RECT 296.800 2442.260 297.060 2442.520 ;
      LAYER met2 ;
        RECT 17.570 2555.595 17.850 2555.965 ;
        RECT 17.640 2442.550 17.780 2555.595 ;
        RECT 17.580 2442.230 17.840 2442.550 ;
        RECT 296.800 2442.230 297.060 2442.550 ;
        RECT 296.860 2438.325 297.000 2442.230 ;
        RECT 296.790 2437.955 297.070 2438.325 ;
      LAYER via2 ;
        RECT 17.570 2555.640 17.850 2555.920 ;
        RECT 296.790 2438.000 297.070 2438.280 ;
      LAYER met3 ;
        RECT -4.800 2555.930 2.400 2556.380 ;
        RECT 17.545 2555.930 17.875 2555.945 ;
        RECT -4.800 2555.630 17.875 2555.930 ;
        RECT -4.800 2555.180 2.400 2555.630 ;
        RECT 17.545 2555.615 17.875 2555.630 ;
        RECT 296.765 2438.290 297.095 2438.305 ;
        RECT 310.000 2438.290 314.000 2438.680 ;
        RECT 296.765 2438.080 314.000 2438.290 ;
        RECT 296.765 2437.990 310.500 2438.080 ;
        RECT 296.765 2437.975 297.095 2437.990 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2228.600 17.410 2228.660 ;
        RECT 296.770 2228.600 297.090 2228.660 ;
        RECT 17.090 2228.460 297.090 2228.600 ;
        RECT 17.090 2228.400 17.410 2228.460 ;
        RECT 296.770 2228.400 297.090 2228.460 ;
      LAYER via ;
        RECT 17.120 2228.400 17.380 2228.660 ;
        RECT 296.800 2228.400 297.060 2228.660 ;
      LAYER met2 ;
        RECT 17.110 2303.995 17.390 2304.365 ;
        RECT 17.180 2228.690 17.320 2303.995 ;
        RECT 17.120 2228.370 17.380 2228.690 ;
        RECT 296.800 2228.370 297.060 2228.690 ;
        RECT 296.860 2224.125 297.000 2228.370 ;
        RECT 296.790 2223.755 297.070 2224.125 ;
      LAYER via2 ;
        RECT 17.110 2304.040 17.390 2304.320 ;
        RECT 296.790 2223.800 297.070 2224.080 ;
      LAYER met3 ;
        RECT -4.800 2304.330 2.400 2304.780 ;
        RECT 17.085 2304.330 17.415 2304.345 ;
        RECT -4.800 2304.030 17.415 2304.330 ;
        RECT -4.800 2303.580 2.400 2304.030 ;
        RECT 17.085 2304.015 17.415 2304.030 ;
        RECT 296.765 2224.090 297.095 2224.105 ;
        RECT 310.000 2224.090 314.000 2224.480 ;
        RECT 296.765 2223.880 314.000 2224.090 ;
        RECT 296.765 2223.790 310.500 2223.880 ;
        RECT 296.765 2223.775 297.095 2223.790 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2014.740 17.410 2014.800 ;
        RECT 296.770 2014.740 297.090 2014.800 ;
        RECT 17.090 2014.600 297.090 2014.740 ;
        RECT 17.090 2014.540 17.410 2014.600 ;
        RECT 296.770 2014.540 297.090 2014.600 ;
      LAYER via ;
        RECT 17.120 2014.540 17.380 2014.800 ;
        RECT 296.800 2014.540 297.060 2014.800 ;
      LAYER met2 ;
        RECT 17.110 2052.395 17.390 2052.765 ;
        RECT 17.180 2014.830 17.320 2052.395 ;
        RECT 17.120 2014.510 17.380 2014.830 ;
        RECT 296.800 2014.510 297.060 2014.830 ;
        RECT 296.860 2009.925 297.000 2014.510 ;
        RECT 296.790 2009.555 297.070 2009.925 ;
      LAYER via2 ;
        RECT 17.110 2052.440 17.390 2052.720 ;
        RECT 296.790 2009.600 297.070 2009.880 ;
      LAYER met3 ;
        RECT -4.800 2052.730 2.400 2053.180 ;
        RECT 17.085 2052.730 17.415 2052.745 ;
        RECT -4.800 2052.430 17.415 2052.730 ;
        RECT -4.800 2051.980 2.400 2052.430 ;
        RECT 17.085 2052.415 17.415 2052.430 ;
        RECT 296.765 2009.890 297.095 2009.905 ;
        RECT 310.000 2009.890 314.000 2010.280 ;
        RECT 296.765 2009.680 314.000 2009.890 ;
        RECT 296.765 2009.590 310.500 2009.680 ;
        RECT 296.765 2009.575 297.095 2009.590 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 669.360 2619.170 669.420 ;
        RECT 2900.830 669.360 2901.150 669.420 ;
        RECT 2618.850 669.220 2901.150 669.360 ;
        RECT 2618.850 669.160 2619.170 669.220 ;
        RECT 2900.830 669.160 2901.150 669.220 ;
      LAYER via ;
        RECT 2618.880 669.160 2619.140 669.420 ;
        RECT 2900.860 669.160 2901.120 669.420 ;
      LAYER met2 ;
        RECT 2618.870 826.355 2619.150 826.725 ;
        RECT 2618.940 669.450 2619.080 826.355 ;
        RECT 2618.880 669.130 2619.140 669.450 ;
        RECT 2900.860 669.130 2901.120 669.450 ;
        RECT 2900.920 664.885 2901.060 669.130 ;
        RECT 2900.850 664.515 2901.130 664.885 ;
      LAYER via2 ;
        RECT 2618.870 826.400 2619.150 826.680 ;
        RECT 2900.850 664.560 2901.130 664.840 ;
      LAYER met3 ;
        RECT 2606.000 826.690 2610.000 827.080 ;
        RECT 2618.845 826.690 2619.175 826.705 ;
        RECT 2606.000 826.480 2619.175 826.690 ;
        RECT 2609.580 826.390 2619.175 826.480 ;
        RECT 2618.845 826.375 2619.175 826.390 ;
        RECT 2900.825 664.850 2901.155 664.865 ;
        RECT 2917.600 664.850 2924.800 665.300 ;
        RECT 2900.825 664.550 2924.800 664.850 ;
        RECT 2900.825 664.535 2901.155 664.550 ;
        RECT 2917.600 664.100 2924.800 664.550 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1800.880 17.410 1800.940 ;
        RECT 296.770 1800.880 297.090 1800.940 ;
        RECT 17.090 1800.740 297.090 1800.880 ;
        RECT 17.090 1800.680 17.410 1800.740 ;
        RECT 296.770 1800.680 297.090 1800.740 ;
      LAYER via ;
        RECT 17.120 1800.680 17.380 1800.940 ;
        RECT 296.800 1800.680 297.060 1800.940 ;
      LAYER met2 ;
        RECT 17.110 1801.475 17.390 1801.845 ;
        RECT 17.180 1800.970 17.320 1801.475 ;
        RECT 17.120 1800.650 17.380 1800.970 ;
        RECT 296.800 1800.650 297.060 1800.970 ;
        RECT 296.860 1795.725 297.000 1800.650 ;
        RECT 296.790 1795.355 297.070 1795.725 ;
      LAYER via2 ;
        RECT 17.110 1801.520 17.390 1801.800 ;
        RECT 296.790 1795.400 297.070 1795.680 ;
      LAYER met3 ;
        RECT -4.800 1801.810 2.400 1802.260 ;
        RECT 17.085 1801.810 17.415 1801.825 ;
        RECT -4.800 1801.510 17.415 1801.810 ;
        RECT -4.800 1801.060 2.400 1801.510 ;
        RECT 17.085 1801.495 17.415 1801.510 ;
        RECT 296.765 1795.690 297.095 1795.705 ;
        RECT 310.000 1795.690 314.000 1796.080 ;
        RECT 296.765 1795.480 314.000 1795.690 ;
        RECT 296.765 1795.390 310.500 1795.480 ;
        RECT 296.765 1795.375 297.095 1795.390 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1552.340 17.410 1552.400 ;
        RECT 299.990 1552.340 300.310 1552.400 ;
        RECT 17.090 1552.200 300.310 1552.340 ;
        RECT 17.090 1552.140 17.410 1552.200 ;
        RECT 299.990 1552.140 300.310 1552.200 ;
      LAYER via ;
        RECT 17.120 1552.140 17.380 1552.400 ;
        RECT 300.020 1552.140 300.280 1552.400 ;
      LAYER met2 ;
        RECT 300.010 1580.475 300.290 1580.845 ;
        RECT 300.080 1552.430 300.220 1580.475 ;
        RECT 17.120 1552.110 17.380 1552.430 ;
        RECT 300.020 1552.110 300.280 1552.430 ;
        RECT 17.180 1550.245 17.320 1552.110 ;
        RECT 17.110 1549.875 17.390 1550.245 ;
      LAYER via2 ;
        RECT 300.010 1580.520 300.290 1580.800 ;
        RECT 17.110 1549.920 17.390 1550.200 ;
      LAYER met3 ;
        RECT 299.985 1580.810 300.315 1580.825 ;
        RECT 310.000 1580.810 314.000 1581.200 ;
        RECT 299.985 1580.600 314.000 1580.810 ;
        RECT 299.985 1580.510 310.500 1580.600 ;
        RECT 299.985 1580.495 300.315 1580.510 ;
        RECT -4.800 1550.210 2.400 1550.660 ;
        RECT 17.085 1550.210 17.415 1550.225 ;
        RECT -4.800 1549.910 17.415 1550.210 ;
        RECT -4.800 1549.460 2.400 1549.910 ;
        RECT 17.085 1549.895 17.415 1549.910 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1304.140 17.410 1304.200 ;
        RECT 299.990 1304.140 300.310 1304.200 ;
        RECT 17.090 1304.000 300.310 1304.140 ;
        RECT 17.090 1303.940 17.410 1304.000 ;
        RECT 299.990 1303.940 300.310 1304.000 ;
      LAYER via ;
        RECT 17.120 1303.940 17.380 1304.200 ;
        RECT 300.020 1303.940 300.280 1304.200 ;
      LAYER met2 ;
        RECT 300.010 1366.275 300.290 1366.645 ;
        RECT 300.080 1304.230 300.220 1366.275 ;
        RECT 17.120 1303.910 17.380 1304.230 ;
        RECT 300.020 1303.910 300.280 1304.230 ;
        RECT 17.180 1298.645 17.320 1303.910 ;
        RECT 17.110 1298.275 17.390 1298.645 ;
      LAYER via2 ;
        RECT 300.010 1366.320 300.290 1366.600 ;
        RECT 17.110 1298.320 17.390 1298.600 ;
      LAYER met3 ;
        RECT 299.985 1366.610 300.315 1366.625 ;
        RECT 310.000 1366.610 314.000 1367.000 ;
        RECT 299.985 1366.400 314.000 1366.610 ;
        RECT 299.985 1366.310 310.500 1366.400 ;
        RECT 299.985 1366.295 300.315 1366.310 ;
        RECT -4.800 1298.610 2.400 1299.060 ;
        RECT 17.085 1298.610 17.415 1298.625 ;
        RECT -4.800 1298.310 17.415 1298.610 ;
        RECT -4.800 1297.860 2.400 1298.310 ;
        RECT 17.085 1298.295 17.415 1298.310 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1048.800 17.410 1048.860 ;
        RECT 299.990 1048.800 300.310 1048.860 ;
        RECT 17.090 1048.660 300.310 1048.800 ;
        RECT 17.090 1048.600 17.410 1048.660 ;
        RECT 299.990 1048.600 300.310 1048.660 ;
      LAYER via ;
        RECT 17.120 1048.600 17.380 1048.860 ;
        RECT 300.020 1048.600 300.280 1048.860 ;
      LAYER met2 ;
        RECT 300.010 1152.075 300.290 1152.445 ;
        RECT 300.080 1048.890 300.220 1152.075 ;
        RECT 17.120 1048.570 17.380 1048.890 ;
        RECT 300.020 1048.570 300.280 1048.890 ;
        RECT 17.180 1047.045 17.320 1048.570 ;
        RECT 17.110 1046.675 17.390 1047.045 ;
      LAYER via2 ;
        RECT 300.010 1152.120 300.290 1152.400 ;
        RECT 17.110 1046.720 17.390 1047.000 ;
      LAYER met3 ;
        RECT 299.985 1152.410 300.315 1152.425 ;
        RECT 310.000 1152.410 314.000 1152.800 ;
        RECT 299.985 1152.200 314.000 1152.410 ;
        RECT 299.985 1152.110 310.500 1152.200 ;
        RECT 299.985 1152.095 300.315 1152.110 ;
        RECT -4.800 1047.010 2.400 1047.460 ;
        RECT 17.085 1047.010 17.415 1047.025 ;
        RECT -4.800 1046.710 17.415 1047.010 ;
        RECT -4.800 1046.260 2.400 1046.710 ;
        RECT 17.085 1046.695 17.415 1046.710 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 800.260 16.030 800.320 ;
        RECT 300.910 800.260 301.230 800.320 ;
        RECT 15.710 800.120 301.230 800.260 ;
        RECT 15.710 800.060 16.030 800.120 ;
        RECT 300.910 800.060 301.230 800.120 ;
      LAYER via ;
        RECT 15.740 800.060 16.000 800.320 ;
        RECT 300.940 800.060 301.200 800.320 ;
      LAYER met2 ;
        RECT 300.930 937.875 301.210 938.245 ;
        RECT 301.000 800.350 301.140 937.875 ;
        RECT 15.740 800.030 16.000 800.350 ;
        RECT 300.940 800.030 301.200 800.350 ;
        RECT 15.800 796.125 15.940 800.030 ;
        RECT 15.730 795.755 16.010 796.125 ;
      LAYER via2 ;
        RECT 300.930 937.920 301.210 938.200 ;
        RECT 15.730 795.800 16.010 796.080 ;
      LAYER met3 ;
        RECT 300.905 938.210 301.235 938.225 ;
        RECT 310.000 938.210 314.000 938.600 ;
        RECT 300.905 938.000 314.000 938.210 ;
        RECT 300.905 937.910 310.500 938.000 ;
        RECT 300.905 937.895 301.235 937.910 ;
        RECT -4.800 796.090 2.400 796.540 ;
        RECT 15.705 796.090 16.035 796.105 ;
        RECT -4.800 795.790 16.035 796.090 ;
        RECT -4.800 795.340 2.400 795.790 ;
        RECT 15.705 795.775 16.035 795.790 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 544.920 17.410 544.980 ;
        RECT 300.910 544.920 301.230 544.980 ;
        RECT 17.090 544.780 301.230 544.920 ;
        RECT 17.090 544.720 17.410 544.780 ;
        RECT 300.910 544.720 301.230 544.780 ;
      LAYER via ;
        RECT 17.120 544.720 17.380 544.980 ;
        RECT 300.940 544.720 301.200 544.980 ;
      LAYER met2 ;
        RECT 300.930 723.675 301.210 724.045 ;
        RECT 301.000 545.010 301.140 723.675 ;
        RECT 17.120 544.690 17.380 545.010 ;
        RECT 300.940 544.690 301.200 545.010 ;
        RECT 17.180 544.525 17.320 544.690 ;
        RECT 17.110 544.155 17.390 544.525 ;
      LAYER via2 ;
        RECT 300.930 723.720 301.210 724.000 ;
        RECT 17.110 544.200 17.390 544.480 ;
      LAYER met3 ;
        RECT 300.905 724.010 301.235 724.025 ;
        RECT 310.000 724.010 314.000 724.400 ;
        RECT 300.905 723.800 314.000 724.010 ;
        RECT 300.905 723.710 310.500 723.800 ;
        RECT 300.905 723.695 301.235 723.710 ;
        RECT -4.800 544.490 2.400 544.940 ;
        RECT 17.085 544.490 17.415 544.505 ;
        RECT -4.800 544.190 17.415 544.490 ;
        RECT -4.800 543.740 2.400 544.190 ;
        RECT 17.085 544.175 17.415 544.190 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 296.720 15.570 296.780 ;
        RECT 301.370 296.720 301.690 296.780 ;
        RECT 15.250 296.580 301.690 296.720 ;
        RECT 15.250 296.520 15.570 296.580 ;
        RECT 301.370 296.520 301.690 296.580 ;
      LAYER via ;
        RECT 15.280 296.520 15.540 296.780 ;
        RECT 301.400 296.520 301.660 296.780 ;
      LAYER met2 ;
        RECT 301.390 509.475 301.670 509.845 ;
        RECT 301.460 296.810 301.600 509.475 ;
        RECT 15.280 296.490 15.540 296.810 ;
        RECT 301.400 296.490 301.660 296.810 ;
        RECT 15.340 292.925 15.480 296.490 ;
        RECT 15.270 292.555 15.550 292.925 ;
      LAYER via2 ;
        RECT 301.390 509.520 301.670 509.800 ;
        RECT 15.270 292.600 15.550 292.880 ;
      LAYER met3 ;
        RECT 301.365 509.810 301.695 509.825 ;
        RECT 310.000 509.810 314.000 510.200 ;
        RECT 301.365 509.600 314.000 509.810 ;
        RECT 301.365 509.510 310.500 509.600 ;
        RECT 301.365 509.495 301.695 509.510 ;
        RECT -4.800 292.890 2.400 293.340 ;
        RECT 15.245 292.890 15.575 292.905 ;
        RECT -4.800 292.590 15.575 292.890 ;
        RECT -4.800 292.140 2.400 292.590 ;
        RECT 15.245 292.575 15.575 292.590 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 48.180 17.410 48.240 ;
        RECT 299.990 48.180 300.310 48.240 ;
        RECT 17.090 48.040 300.310 48.180 ;
        RECT 17.090 47.980 17.410 48.040 ;
        RECT 299.990 47.980 300.310 48.040 ;
      LAYER via ;
        RECT 17.120 47.980 17.380 48.240 ;
        RECT 300.020 47.980 300.280 48.240 ;
      LAYER met2 ;
        RECT 300.010 295.275 300.290 295.645 ;
        RECT 300.080 48.270 300.220 295.275 ;
        RECT 17.120 47.950 17.380 48.270 ;
        RECT 300.020 47.950 300.280 48.270 ;
        RECT 17.180 42.005 17.320 47.950 ;
        RECT 17.110 41.635 17.390 42.005 ;
      LAYER via2 ;
        RECT 300.010 295.320 300.290 295.600 ;
        RECT 17.110 41.680 17.390 41.960 ;
      LAYER met3 ;
        RECT 299.985 295.610 300.315 295.625 ;
        RECT 310.000 295.610 314.000 296.000 ;
        RECT 299.985 295.400 314.000 295.610 ;
        RECT 299.985 295.310 310.500 295.400 ;
        RECT 299.985 295.295 300.315 295.310 ;
        RECT -4.800 41.970 2.400 42.420 ;
        RECT 17.085 41.970 17.415 41.985 ;
        RECT -4.800 41.670 17.415 41.970 ;
        RECT -4.800 41.220 2.400 41.670 ;
        RECT 17.085 41.655 17.415 41.670 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 903.960 2619.170 904.020 ;
        RECT 2900.830 903.960 2901.150 904.020 ;
        RECT 2618.850 903.820 2901.150 903.960 ;
        RECT 2618.850 903.760 2619.170 903.820 ;
        RECT 2900.830 903.760 2901.150 903.820 ;
      LAYER via ;
        RECT 2618.880 903.760 2619.140 904.020 ;
        RECT 2900.860 903.760 2901.120 904.020 ;
      LAYER met2 ;
        RECT 2618.870 1026.275 2619.150 1026.645 ;
        RECT 2618.940 904.050 2619.080 1026.275 ;
        RECT 2618.880 903.730 2619.140 904.050 ;
        RECT 2900.860 903.730 2901.120 904.050 ;
        RECT 2900.920 899.485 2901.060 903.730 ;
        RECT 2900.850 899.115 2901.130 899.485 ;
      LAYER via2 ;
        RECT 2618.870 1026.320 2619.150 1026.600 ;
        RECT 2900.850 899.160 2901.130 899.440 ;
      LAYER met3 ;
        RECT 2606.000 1026.610 2610.000 1027.000 ;
        RECT 2618.845 1026.610 2619.175 1026.625 ;
        RECT 2606.000 1026.400 2619.175 1026.610 ;
        RECT 2609.580 1026.310 2619.175 1026.400 ;
        RECT 2618.845 1026.295 2619.175 1026.310 ;
        RECT 2900.825 899.450 2901.155 899.465 ;
        RECT 2917.600 899.450 2924.800 899.900 ;
        RECT 2900.825 899.150 2924.800 899.450 ;
        RECT 2900.825 899.135 2901.155 899.150 ;
        RECT 2917.600 898.700 2924.800 899.150 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1138.560 2618.710 1138.620 ;
        RECT 2900.830 1138.560 2901.150 1138.620 ;
        RECT 2618.390 1138.420 2901.150 1138.560 ;
        RECT 2618.390 1138.360 2618.710 1138.420 ;
        RECT 2900.830 1138.360 2901.150 1138.420 ;
      LAYER via ;
        RECT 2618.420 1138.360 2618.680 1138.620 ;
        RECT 2900.860 1138.360 2901.120 1138.620 ;
      LAYER met2 ;
        RECT 2618.410 1226.195 2618.690 1226.565 ;
        RECT 2618.480 1138.650 2618.620 1226.195 ;
        RECT 2618.420 1138.330 2618.680 1138.650 ;
        RECT 2900.860 1138.330 2901.120 1138.650 ;
        RECT 2900.920 1134.085 2901.060 1138.330 ;
        RECT 2900.850 1133.715 2901.130 1134.085 ;
      LAYER via2 ;
        RECT 2618.410 1226.240 2618.690 1226.520 ;
        RECT 2900.850 1133.760 2901.130 1134.040 ;
      LAYER met3 ;
        RECT 2606.000 1226.530 2610.000 1226.920 ;
        RECT 2618.385 1226.530 2618.715 1226.545 ;
        RECT 2606.000 1226.320 2618.715 1226.530 ;
        RECT 2609.580 1226.230 2618.715 1226.320 ;
        RECT 2618.385 1226.215 2618.715 1226.230 ;
        RECT 2900.825 1134.050 2901.155 1134.065 ;
        RECT 2917.600 1134.050 2924.800 1134.500 ;
        RECT 2900.825 1133.750 2924.800 1134.050 ;
        RECT 2900.825 1133.735 2901.155 1133.750 ;
        RECT 2917.600 1133.300 2924.800 1133.750 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1373.160 2618.710 1373.220 ;
        RECT 2900.830 1373.160 2901.150 1373.220 ;
        RECT 2618.390 1373.020 2901.150 1373.160 ;
        RECT 2618.390 1372.960 2618.710 1373.020 ;
        RECT 2900.830 1372.960 2901.150 1373.020 ;
      LAYER via ;
        RECT 2618.420 1372.960 2618.680 1373.220 ;
        RECT 2900.860 1372.960 2901.120 1373.220 ;
      LAYER met2 ;
        RECT 2618.410 1426.115 2618.690 1426.485 ;
        RECT 2618.480 1373.250 2618.620 1426.115 ;
        RECT 2618.420 1372.930 2618.680 1373.250 ;
        RECT 2900.860 1372.930 2901.120 1373.250 ;
        RECT 2900.920 1368.685 2901.060 1372.930 ;
        RECT 2900.850 1368.315 2901.130 1368.685 ;
      LAYER via2 ;
        RECT 2618.410 1426.160 2618.690 1426.440 ;
        RECT 2900.850 1368.360 2901.130 1368.640 ;
      LAYER met3 ;
        RECT 2606.000 1426.450 2610.000 1426.840 ;
        RECT 2618.385 1426.450 2618.715 1426.465 ;
        RECT 2606.000 1426.240 2618.715 1426.450 ;
        RECT 2609.580 1426.150 2618.715 1426.240 ;
        RECT 2618.385 1426.135 2618.715 1426.150 ;
        RECT 2900.825 1368.650 2901.155 1368.665 ;
        RECT 2917.600 1368.650 2924.800 1369.100 ;
        RECT 2900.825 1368.350 2924.800 1368.650 ;
        RECT 2900.825 1368.335 2901.155 1368.350 ;
        RECT 2917.600 1367.900 2924.800 1368.350 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.630 1607.760 2615.950 1607.820 ;
        RECT 2900.830 1607.760 2901.150 1607.820 ;
        RECT 2615.630 1607.620 2901.150 1607.760 ;
        RECT 2615.630 1607.560 2615.950 1607.620 ;
        RECT 2900.830 1607.560 2901.150 1607.620 ;
      LAYER via ;
        RECT 2615.660 1607.560 2615.920 1607.820 ;
        RECT 2900.860 1607.560 2901.120 1607.820 ;
      LAYER met2 ;
        RECT 2615.650 1626.035 2615.930 1626.405 ;
        RECT 2615.720 1607.850 2615.860 1626.035 ;
        RECT 2615.660 1607.530 2615.920 1607.850 ;
        RECT 2900.860 1607.530 2901.120 1607.850 ;
        RECT 2900.920 1603.285 2901.060 1607.530 ;
        RECT 2900.850 1602.915 2901.130 1603.285 ;
      LAYER via2 ;
        RECT 2615.650 1626.080 2615.930 1626.360 ;
        RECT 2900.850 1602.960 2901.130 1603.240 ;
      LAYER met3 ;
        RECT 2606.000 1626.370 2610.000 1626.760 ;
        RECT 2615.625 1626.370 2615.955 1626.385 ;
        RECT 2606.000 1626.160 2615.955 1626.370 ;
        RECT 2609.580 1626.070 2615.955 1626.160 ;
        RECT 2615.625 1626.055 2615.955 1626.070 ;
        RECT 2900.825 1603.250 2901.155 1603.265 ;
        RECT 2917.600 1603.250 2924.800 1603.700 ;
        RECT 2900.825 1602.950 2924.800 1603.250 ;
        RECT 2900.825 1602.935 2901.155 1602.950 ;
        RECT 2917.600 1602.500 2924.800 1602.950 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2616.550 1835.560 2616.870 1835.620 ;
        RECT 2900.830 1835.560 2901.150 1835.620 ;
        RECT 2616.550 1835.420 2901.150 1835.560 ;
        RECT 2616.550 1835.360 2616.870 1835.420 ;
        RECT 2900.830 1835.360 2901.150 1835.420 ;
      LAYER via ;
        RECT 2616.580 1835.360 2616.840 1835.620 ;
        RECT 2900.860 1835.360 2901.120 1835.620 ;
      LAYER met2 ;
        RECT 2900.850 1837.515 2901.130 1837.885 ;
        RECT 2900.920 1835.650 2901.060 1837.515 ;
        RECT 2616.580 1835.330 2616.840 1835.650 ;
        RECT 2900.860 1835.330 2901.120 1835.650 ;
        RECT 2616.640 1827.005 2616.780 1835.330 ;
        RECT 2616.570 1826.635 2616.850 1827.005 ;
      LAYER via2 ;
        RECT 2900.850 1837.560 2901.130 1837.840 ;
        RECT 2616.570 1826.680 2616.850 1826.960 ;
      LAYER met3 ;
        RECT 2900.825 1837.850 2901.155 1837.865 ;
        RECT 2917.600 1837.850 2924.800 1838.300 ;
        RECT 2900.825 1837.550 2924.800 1837.850 ;
        RECT 2900.825 1837.535 2901.155 1837.550 ;
        RECT 2917.600 1837.100 2924.800 1837.550 ;
        RECT 2606.000 1826.970 2610.000 1827.360 ;
        RECT 2616.545 1826.970 2616.875 1826.985 ;
        RECT 2606.000 1826.760 2616.875 1826.970 ;
        RECT 2609.580 1826.670 2616.875 1826.760 ;
        RECT 2616.545 1826.655 2616.875 1826.670 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2070.160 2618.710 2070.220 ;
        RECT 2900.830 2070.160 2901.150 2070.220 ;
        RECT 2618.390 2070.020 2901.150 2070.160 ;
        RECT 2618.390 2069.960 2618.710 2070.020 ;
        RECT 2900.830 2069.960 2901.150 2070.020 ;
      LAYER via ;
        RECT 2618.420 2069.960 2618.680 2070.220 ;
        RECT 2900.860 2069.960 2901.120 2070.220 ;
      LAYER met2 ;
        RECT 2900.850 2072.115 2901.130 2072.485 ;
        RECT 2900.920 2070.250 2901.060 2072.115 ;
        RECT 2618.420 2069.930 2618.680 2070.250 ;
        RECT 2900.860 2069.930 2901.120 2070.250 ;
        RECT 2618.480 2026.925 2618.620 2069.930 ;
        RECT 2618.410 2026.555 2618.690 2026.925 ;
      LAYER via2 ;
        RECT 2900.850 2072.160 2901.130 2072.440 ;
        RECT 2618.410 2026.600 2618.690 2026.880 ;
      LAYER met3 ;
        RECT 2900.825 2072.450 2901.155 2072.465 ;
        RECT 2917.600 2072.450 2924.800 2072.900 ;
        RECT 2900.825 2072.150 2924.800 2072.450 ;
        RECT 2900.825 2072.135 2901.155 2072.150 ;
        RECT 2917.600 2071.700 2924.800 2072.150 ;
        RECT 2606.000 2026.890 2610.000 2027.280 ;
        RECT 2618.385 2026.890 2618.715 2026.905 ;
        RECT 2606.000 2026.680 2618.715 2026.890 ;
        RECT 2609.580 2026.590 2618.715 2026.680 ;
        RECT 2618.385 2026.575 2618.715 2026.590 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2304.760 2619.170 2304.820 ;
        RECT 2900.830 2304.760 2901.150 2304.820 ;
        RECT 2618.850 2304.620 2901.150 2304.760 ;
        RECT 2618.850 2304.560 2619.170 2304.620 ;
        RECT 2900.830 2304.560 2901.150 2304.620 ;
      LAYER via ;
        RECT 2618.880 2304.560 2619.140 2304.820 ;
        RECT 2900.860 2304.560 2901.120 2304.820 ;
      LAYER met2 ;
        RECT 2900.850 2306.715 2901.130 2307.085 ;
        RECT 2900.920 2304.850 2901.060 2306.715 ;
        RECT 2618.880 2304.530 2619.140 2304.850 ;
        RECT 2900.860 2304.530 2901.120 2304.850 ;
        RECT 2618.940 2226.845 2619.080 2304.530 ;
        RECT 2618.870 2226.475 2619.150 2226.845 ;
      LAYER via2 ;
        RECT 2900.850 2306.760 2901.130 2307.040 ;
        RECT 2618.870 2226.520 2619.150 2226.800 ;
      LAYER met3 ;
        RECT 2900.825 2307.050 2901.155 2307.065 ;
        RECT 2917.600 2307.050 2924.800 2307.500 ;
        RECT 2900.825 2306.750 2924.800 2307.050 ;
        RECT 2900.825 2306.735 2901.155 2306.750 ;
        RECT 2917.600 2306.300 2924.800 2306.750 ;
        RECT 2606.000 2226.810 2610.000 2227.200 ;
        RECT 2618.845 2226.810 2619.175 2226.825 ;
        RECT 2606.000 2226.600 2619.175 2226.810 ;
        RECT 2609.580 2226.510 2619.175 2226.600 ;
        RECT 2618.845 2226.495 2619.175 2226.510 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 124.000 2619.170 124.060 ;
        RECT 2900.830 124.000 2901.150 124.060 ;
        RECT 2618.850 123.860 2901.150 124.000 ;
        RECT 2618.850 123.800 2619.170 123.860 ;
        RECT 2900.830 123.800 2901.150 123.860 ;
      LAYER via ;
        RECT 2618.880 123.800 2619.140 124.060 ;
        RECT 2900.860 123.800 2901.120 124.060 ;
      LAYER met2 ;
        RECT 2618.870 359.875 2619.150 360.245 ;
        RECT 2618.940 124.090 2619.080 359.875 ;
        RECT 2618.880 123.770 2619.140 124.090 ;
        RECT 2900.860 123.770 2901.120 124.090 ;
        RECT 2900.920 117.485 2901.060 123.770 ;
        RECT 2900.850 117.115 2901.130 117.485 ;
      LAYER via2 ;
        RECT 2618.870 359.920 2619.150 360.200 ;
        RECT 2900.850 117.160 2901.130 117.440 ;
      LAYER met3 ;
        RECT 2606.000 360.210 2610.000 360.600 ;
        RECT 2618.845 360.210 2619.175 360.225 ;
        RECT 2606.000 360.000 2619.175 360.210 ;
        RECT 2609.580 359.910 2619.175 360.000 ;
        RECT 2618.845 359.895 2619.175 359.910 ;
        RECT 2900.825 117.450 2901.155 117.465 ;
        RECT 2917.600 117.450 2924.800 117.900 ;
        RECT 2900.825 117.150 2924.800 117.450 ;
        RECT 2900.825 117.135 2901.155 117.150 ;
        RECT 2917.600 116.700 2924.800 117.150 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2463.540 2619.170 2463.600 ;
        RECT 2900.830 2463.540 2901.150 2463.600 ;
        RECT 2618.850 2463.400 2901.150 2463.540 ;
        RECT 2618.850 2463.340 2619.170 2463.400 ;
        RECT 2900.830 2463.340 2901.150 2463.400 ;
      LAYER via ;
        RECT 2618.880 2463.340 2619.140 2463.600 ;
        RECT 2900.860 2463.340 2901.120 2463.600 ;
      LAYER met2 ;
        RECT 2618.880 2463.310 2619.140 2463.630 ;
        RECT 2900.860 2463.485 2901.120 2463.630 ;
        RECT 2618.940 2360.125 2619.080 2463.310 ;
        RECT 2900.850 2463.115 2901.130 2463.485 ;
        RECT 2618.870 2359.755 2619.150 2360.125 ;
      LAYER via2 ;
        RECT 2900.850 2463.160 2901.130 2463.440 ;
        RECT 2618.870 2359.800 2619.150 2360.080 ;
      LAYER met3 ;
        RECT 2900.825 2463.450 2901.155 2463.465 ;
        RECT 2917.600 2463.450 2924.800 2463.900 ;
        RECT 2900.825 2463.150 2924.800 2463.450 ;
        RECT 2900.825 2463.135 2901.155 2463.150 ;
        RECT 2917.600 2462.700 2924.800 2463.150 ;
        RECT 2606.000 2360.090 2610.000 2360.480 ;
        RECT 2618.845 2360.090 2619.175 2360.105 ;
        RECT 2606.000 2359.880 2619.175 2360.090 ;
        RECT 2609.580 2359.790 2619.175 2359.880 ;
        RECT 2618.845 2359.775 2619.175 2359.790 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2617.470 2698.140 2617.790 2698.200 ;
        RECT 2900.830 2698.140 2901.150 2698.200 ;
        RECT 2617.470 2698.000 2901.150 2698.140 ;
        RECT 2617.470 2697.940 2617.790 2698.000 ;
        RECT 2900.830 2697.940 2901.150 2698.000 ;
      LAYER via ;
        RECT 2617.500 2697.940 2617.760 2698.200 ;
        RECT 2900.860 2697.940 2901.120 2698.200 ;
      LAYER met2 ;
        RECT 2617.500 2697.910 2617.760 2698.230 ;
        RECT 2900.860 2698.085 2901.120 2698.230 ;
        RECT 2617.560 2691.170 2617.700 2697.910 ;
        RECT 2900.850 2697.715 2901.130 2698.085 ;
        RECT 2617.560 2691.030 2618.620 2691.170 ;
        RECT 2618.480 2560.045 2618.620 2691.030 ;
        RECT 2618.410 2559.675 2618.690 2560.045 ;
      LAYER via2 ;
        RECT 2900.850 2697.760 2901.130 2698.040 ;
        RECT 2618.410 2559.720 2618.690 2560.000 ;
      LAYER met3 ;
        RECT 2900.825 2698.050 2901.155 2698.065 ;
        RECT 2917.600 2698.050 2924.800 2698.500 ;
        RECT 2900.825 2697.750 2924.800 2698.050 ;
        RECT 2900.825 2697.735 2901.155 2697.750 ;
        RECT 2917.600 2697.300 2924.800 2697.750 ;
        RECT 2606.000 2560.010 2610.000 2560.400 ;
        RECT 2618.385 2560.010 2618.715 2560.025 ;
        RECT 2606.000 2559.800 2618.715 2560.010 ;
        RECT 2609.580 2559.710 2618.715 2559.800 ;
        RECT 2618.385 2559.695 2618.715 2559.710 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2932.740 2618.710 2932.800 ;
        RECT 2900.830 2932.740 2901.150 2932.800 ;
        RECT 2618.390 2932.600 2901.150 2932.740 ;
        RECT 2618.390 2932.540 2618.710 2932.600 ;
        RECT 2900.830 2932.540 2901.150 2932.600 ;
      LAYER via ;
        RECT 2618.420 2932.540 2618.680 2932.800 ;
        RECT 2900.860 2932.540 2901.120 2932.800 ;
      LAYER met2 ;
        RECT 2618.420 2932.510 2618.680 2932.830 ;
        RECT 2900.860 2932.685 2901.120 2932.830 ;
        RECT 2618.480 2759.965 2618.620 2932.510 ;
        RECT 2900.850 2932.315 2901.130 2932.685 ;
        RECT 2618.410 2759.595 2618.690 2759.965 ;
      LAYER via2 ;
        RECT 2900.850 2932.360 2901.130 2932.640 ;
        RECT 2618.410 2759.640 2618.690 2759.920 ;
      LAYER met3 ;
        RECT 2900.825 2932.650 2901.155 2932.665 ;
        RECT 2917.600 2932.650 2924.800 2933.100 ;
        RECT 2900.825 2932.350 2924.800 2932.650 ;
        RECT 2900.825 2932.335 2901.155 2932.350 ;
        RECT 2917.600 2931.900 2924.800 2932.350 ;
        RECT 2606.000 2759.930 2610.000 2760.320 ;
        RECT 2618.385 2759.930 2618.715 2759.945 ;
        RECT 2606.000 2759.720 2618.715 2759.930 ;
        RECT 2609.580 2759.630 2618.715 2759.720 ;
        RECT 2618.385 2759.615 2618.715 2759.630 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 3167.340 2618.710 3167.400 ;
        RECT 2900.830 3167.340 2901.150 3167.400 ;
        RECT 2618.390 3167.200 2901.150 3167.340 ;
        RECT 2618.390 3167.140 2618.710 3167.200 ;
        RECT 2900.830 3167.140 2901.150 3167.200 ;
      LAYER via ;
        RECT 2618.420 3167.140 2618.680 3167.400 ;
        RECT 2900.860 3167.140 2901.120 3167.400 ;
      LAYER met2 ;
        RECT 2618.420 3167.110 2618.680 3167.430 ;
        RECT 2900.860 3167.285 2901.120 3167.430 ;
        RECT 2618.480 2959.885 2618.620 3167.110 ;
        RECT 2900.850 3166.915 2901.130 3167.285 ;
        RECT 2618.410 2959.515 2618.690 2959.885 ;
      LAYER via2 ;
        RECT 2900.850 3166.960 2901.130 3167.240 ;
        RECT 2618.410 2959.560 2618.690 2959.840 ;
      LAYER met3 ;
        RECT 2900.825 3167.250 2901.155 3167.265 ;
        RECT 2917.600 3167.250 2924.800 3167.700 ;
        RECT 2900.825 3166.950 2924.800 3167.250 ;
        RECT 2900.825 3166.935 2901.155 3166.950 ;
        RECT 2917.600 3166.500 2924.800 3166.950 ;
        RECT 2606.000 2959.850 2610.000 2960.240 ;
        RECT 2618.385 2959.850 2618.715 2959.865 ;
        RECT 2606.000 2959.640 2618.715 2959.850 ;
        RECT 2609.580 2959.550 2618.715 2959.640 ;
        RECT 2618.385 2959.535 2618.715 2959.550 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3401.940 2619.170 3402.000 ;
        RECT 2900.830 3401.940 2901.150 3402.000 ;
        RECT 2618.850 3401.800 2901.150 3401.940 ;
        RECT 2618.850 3401.740 2619.170 3401.800 ;
        RECT 2900.830 3401.740 2901.150 3401.800 ;
      LAYER via ;
        RECT 2618.880 3401.740 2619.140 3402.000 ;
        RECT 2900.860 3401.740 2901.120 3402.000 ;
      LAYER met2 ;
        RECT 2618.880 3401.710 2619.140 3402.030 ;
        RECT 2900.860 3401.885 2901.120 3402.030 ;
        RECT 2618.940 3159.805 2619.080 3401.710 ;
        RECT 2900.850 3401.515 2901.130 3401.885 ;
        RECT 2618.870 3159.435 2619.150 3159.805 ;
      LAYER via2 ;
        RECT 2900.850 3401.560 2901.130 3401.840 ;
        RECT 2618.870 3159.480 2619.150 3159.760 ;
      LAYER met3 ;
        RECT 2900.825 3401.850 2901.155 3401.865 ;
        RECT 2917.600 3401.850 2924.800 3402.300 ;
        RECT 2900.825 3401.550 2924.800 3401.850 ;
        RECT 2900.825 3401.535 2901.155 3401.550 ;
        RECT 2917.600 3401.100 2924.800 3401.550 ;
        RECT 2606.000 3159.770 2610.000 3160.160 ;
        RECT 2618.845 3159.770 2619.175 3159.785 ;
        RECT 2606.000 3159.560 2619.175 3159.770 ;
        RECT 2609.580 3159.470 2619.175 3159.560 ;
        RECT 2618.845 3159.455 2619.175 3159.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2483.610 3501.900 2483.930 3501.960 ;
        RECT 2757.310 3501.900 2757.630 3501.960 ;
        RECT 2483.610 3501.760 2757.630 3501.900 ;
        RECT 2483.610 3501.700 2483.930 3501.760 ;
        RECT 2757.310 3501.700 2757.630 3501.760 ;
      LAYER via ;
        RECT 2483.640 3501.700 2483.900 3501.960 ;
        RECT 2757.340 3501.700 2757.600 3501.960 ;
      LAYER met2 ;
        RECT 2757.190 3517.600 2757.750 3524.800 ;
        RECT 2757.400 3501.990 2757.540 3517.600 ;
        RECT 2483.640 3501.670 2483.900 3501.990 ;
        RECT 2757.340 3501.670 2757.600 3501.990 ;
        RECT 2481.750 3259.650 2482.030 3260.000 ;
        RECT 2483.700 3259.650 2483.840 3501.670 ;
        RECT 2481.750 3259.510 2483.840 3259.650 ;
        RECT 2481.750 3256.000 2482.030 3259.510 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2228.310 3501.900 2228.630 3501.960 ;
        RECT 2433.010 3501.900 2433.330 3501.960 ;
        RECT 2228.310 3501.760 2433.330 3501.900 ;
        RECT 2228.310 3501.700 2228.630 3501.760 ;
        RECT 2433.010 3501.700 2433.330 3501.760 ;
      LAYER via ;
        RECT 2228.340 3501.700 2228.600 3501.960 ;
        RECT 2433.040 3501.700 2433.300 3501.960 ;
      LAYER met2 ;
        RECT 2432.890 3517.600 2433.450 3524.800 ;
        RECT 2433.100 3501.990 2433.240 3517.600 ;
        RECT 2228.340 3501.670 2228.600 3501.990 ;
        RECT 2433.040 3501.670 2433.300 3501.990 ;
        RECT 2226.450 3259.650 2226.730 3260.000 ;
        RECT 2228.400 3259.650 2228.540 3501.670 ;
        RECT 2226.450 3259.510 2228.540 3259.650 ;
        RECT 2226.450 3256.000 2226.730 3259.510 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 3501.900 1973.330 3501.960 ;
        RECT 2108.710 3501.900 2109.030 3501.960 ;
        RECT 1973.010 3501.760 2109.030 3501.900 ;
        RECT 1973.010 3501.700 1973.330 3501.760 ;
        RECT 2108.710 3501.700 2109.030 3501.760 ;
      LAYER via ;
        RECT 1973.040 3501.700 1973.300 3501.960 ;
        RECT 2108.740 3501.700 2109.000 3501.960 ;
      LAYER met2 ;
        RECT 2108.590 3517.600 2109.150 3524.800 ;
        RECT 2108.800 3501.990 2108.940 3517.600 ;
        RECT 1973.040 3501.670 1973.300 3501.990 ;
        RECT 2108.740 3501.670 2109.000 3501.990 ;
        RECT 1970.690 3258.970 1970.970 3260.000 ;
        RECT 1973.100 3258.970 1973.240 3501.670 ;
        RECT 1970.690 3258.830 1973.240 3258.970 ;
        RECT 1970.690 3256.000 1970.970 3258.830 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1717.710 3501.560 1718.030 3501.620 ;
        RECT 1783.950 3501.560 1784.270 3501.620 ;
        RECT 1717.710 3501.420 1784.270 3501.560 ;
        RECT 1717.710 3501.360 1718.030 3501.420 ;
        RECT 1783.950 3501.360 1784.270 3501.420 ;
      LAYER via ;
        RECT 1717.740 3501.360 1718.000 3501.620 ;
        RECT 1783.980 3501.360 1784.240 3501.620 ;
      LAYER met2 ;
        RECT 1783.830 3517.600 1784.390 3524.800 ;
        RECT 1784.040 3501.650 1784.180 3517.600 ;
        RECT 1717.740 3501.330 1718.000 3501.650 ;
        RECT 1783.980 3501.330 1784.240 3501.650 ;
        RECT 1714.930 3258.970 1715.210 3260.000 ;
        RECT 1717.800 3258.970 1717.940 3501.330 ;
        RECT 1714.930 3258.830 1717.940 3258.970 ;
        RECT 1714.930 3256.000 1715.210 3258.830 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1455.970 3498.500 1456.290 3498.560 ;
        RECT 1459.650 3498.500 1459.970 3498.560 ;
        RECT 1455.970 3498.360 1459.970 3498.500 ;
        RECT 1455.970 3498.300 1456.290 3498.360 ;
        RECT 1459.650 3498.300 1459.970 3498.360 ;
      LAYER via ;
        RECT 1456.000 3498.300 1456.260 3498.560 ;
        RECT 1459.680 3498.300 1459.940 3498.560 ;
      LAYER met2 ;
        RECT 1459.530 3517.600 1460.090 3524.800 ;
        RECT 1459.740 3498.590 1459.880 3517.600 ;
        RECT 1456.000 3498.270 1456.260 3498.590 ;
        RECT 1459.680 3498.270 1459.940 3498.590 ;
        RECT 1456.060 3258.970 1456.200 3498.270 ;
        RECT 1459.630 3258.970 1459.910 3260.000 ;
        RECT 1456.060 3258.830 1459.910 3258.970 ;
        RECT 1459.630 3256.000 1459.910 3258.830 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 358.600 2618.710 358.660 ;
        RECT 2900.830 358.600 2901.150 358.660 ;
        RECT 2618.390 358.460 2901.150 358.600 ;
        RECT 2618.390 358.400 2618.710 358.460 ;
        RECT 2900.830 358.400 2901.150 358.460 ;
      LAYER via ;
        RECT 2618.420 358.400 2618.680 358.660 ;
        RECT 2900.860 358.400 2901.120 358.660 ;
      LAYER met2 ;
        RECT 2618.410 559.795 2618.690 560.165 ;
        RECT 2618.480 358.690 2618.620 559.795 ;
        RECT 2618.420 358.370 2618.680 358.690 ;
        RECT 2900.860 358.370 2901.120 358.690 ;
        RECT 2900.920 352.085 2901.060 358.370 ;
        RECT 2900.850 351.715 2901.130 352.085 ;
      LAYER via2 ;
        RECT 2618.410 559.840 2618.690 560.120 ;
        RECT 2900.850 351.760 2901.130 352.040 ;
      LAYER met3 ;
        RECT 2606.000 560.130 2610.000 560.520 ;
        RECT 2618.385 560.130 2618.715 560.145 ;
        RECT 2606.000 559.920 2618.715 560.130 ;
        RECT 2609.580 559.830 2618.715 559.920 ;
        RECT 2618.385 559.815 2618.715 559.830 ;
        RECT 2900.825 352.050 2901.155 352.065 ;
        RECT 2917.600 352.050 2924.800 352.500 ;
        RECT 2900.825 351.750 2924.800 352.050 ;
        RECT 2900.825 351.735 2901.155 351.750 ;
        RECT 2917.600 351.300 2924.800 351.750 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1135.350 3498.500 1135.670 3498.560 ;
        RECT 1138.110 3498.500 1138.430 3498.560 ;
        RECT 1135.350 3498.360 1138.430 3498.500 ;
        RECT 1135.350 3498.300 1135.670 3498.360 ;
        RECT 1138.110 3498.300 1138.430 3498.360 ;
        RECT 1138.110 3274.100 1138.430 3274.160 ;
        RECT 1203.890 3274.100 1204.210 3274.160 ;
        RECT 1138.110 3273.960 1204.210 3274.100 ;
        RECT 1138.110 3273.900 1138.430 3273.960 ;
        RECT 1203.890 3273.900 1204.210 3273.960 ;
      LAYER via ;
        RECT 1135.380 3498.300 1135.640 3498.560 ;
        RECT 1138.140 3498.300 1138.400 3498.560 ;
        RECT 1138.140 3273.900 1138.400 3274.160 ;
        RECT 1203.920 3273.900 1204.180 3274.160 ;
      LAYER met2 ;
        RECT 1135.230 3517.600 1135.790 3524.800 ;
        RECT 1135.440 3498.590 1135.580 3517.600 ;
        RECT 1135.380 3498.270 1135.640 3498.590 ;
        RECT 1138.140 3498.270 1138.400 3498.590 ;
        RECT 1138.200 3274.190 1138.340 3498.270 ;
        RECT 1138.140 3273.870 1138.400 3274.190 ;
        RECT 1203.920 3273.870 1204.180 3274.190 ;
        RECT 1203.980 3260.000 1204.120 3273.870 ;
        RECT 1203.870 3256.000 1204.150 3260.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 810.590 3498.500 810.910 3498.560 ;
        RECT 813.810 3498.500 814.130 3498.560 ;
        RECT 810.590 3498.360 814.130 3498.500 ;
        RECT 810.590 3498.300 810.910 3498.360 ;
        RECT 813.810 3498.300 814.130 3498.360 ;
        RECT 813.810 3274.440 814.130 3274.500 ;
        RECT 948.590 3274.440 948.910 3274.500 ;
        RECT 813.810 3274.300 948.910 3274.440 ;
        RECT 813.810 3274.240 814.130 3274.300 ;
        RECT 948.590 3274.240 948.910 3274.300 ;
      LAYER via ;
        RECT 810.620 3498.300 810.880 3498.560 ;
        RECT 813.840 3498.300 814.100 3498.560 ;
        RECT 813.840 3274.240 814.100 3274.500 ;
        RECT 948.620 3274.240 948.880 3274.500 ;
      LAYER met2 ;
        RECT 810.470 3517.600 811.030 3524.800 ;
        RECT 810.680 3498.590 810.820 3517.600 ;
        RECT 810.620 3498.270 810.880 3498.590 ;
        RECT 813.840 3498.270 814.100 3498.590 ;
        RECT 813.900 3274.530 814.040 3498.270 ;
        RECT 813.840 3274.210 814.100 3274.530 ;
        RECT 948.620 3274.210 948.880 3274.530 ;
        RECT 948.680 3260.000 948.820 3274.210 ;
        RECT 948.570 3256.000 948.850 3260.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 486.290 3498.500 486.610 3498.560 ;
        RECT 489.510 3498.500 489.830 3498.560 ;
        RECT 486.290 3498.360 489.830 3498.500 ;
        RECT 486.290 3498.300 486.610 3498.360 ;
        RECT 489.510 3498.300 489.830 3498.360 ;
        RECT 489.510 3274.440 489.830 3274.500 ;
        RECT 692.830 3274.440 693.150 3274.500 ;
        RECT 489.510 3274.300 693.150 3274.440 ;
        RECT 489.510 3274.240 489.830 3274.300 ;
        RECT 692.830 3274.240 693.150 3274.300 ;
      LAYER via ;
        RECT 486.320 3498.300 486.580 3498.560 ;
        RECT 489.540 3498.300 489.800 3498.560 ;
        RECT 489.540 3274.240 489.800 3274.500 ;
        RECT 692.860 3274.240 693.120 3274.500 ;
      LAYER met2 ;
        RECT 486.170 3517.600 486.730 3524.800 ;
        RECT 486.380 3498.590 486.520 3517.600 ;
        RECT 486.320 3498.270 486.580 3498.590 ;
        RECT 489.540 3498.270 489.800 3498.590 ;
        RECT 489.600 3274.530 489.740 3498.270 ;
        RECT 489.540 3274.210 489.800 3274.530 ;
        RECT 692.860 3274.210 693.120 3274.530 ;
        RECT 692.920 3260.000 693.060 3274.210 ;
        RECT 692.810 3256.000 693.090 3260.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 161.990 3498.500 162.310 3498.560 ;
        RECT 165.210 3498.500 165.530 3498.560 ;
        RECT 161.990 3498.360 165.530 3498.500 ;
        RECT 161.990 3498.300 162.310 3498.360 ;
        RECT 165.210 3498.300 165.530 3498.360 ;
        RECT 165.210 3274.440 165.530 3274.500 ;
        RECT 437.530 3274.440 437.850 3274.500 ;
        RECT 165.210 3274.300 437.850 3274.440 ;
        RECT 165.210 3274.240 165.530 3274.300 ;
        RECT 437.530 3274.240 437.850 3274.300 ;
      LAYER via ;
        RECT 162.020 3498.300 162.280 3498.560 ;
        RECT 165.240 3498.300 165.500 3498.560 ;
        RECT 165.240 3274.240 165.500 3274.500 ;
        RECT 437.560 3274.240 437.820 3274.500 ;
      LAYER met2 ;
        RECT 161.870 3517.600 162.430 3524.800 ;
        RECT 162.080 3498.590 162.220 3517.600 ;
        RECT 162.020 3498.270 162.280 3498.590 ;
        RECT 165.240 3498.270 165.500 3498.590 ;
        RECT 165.300 3274.530 165.440 3498.270 ;
        RECT 165.240 3274.210 165.500 3274.530 ;
        RECT 437.560 3274.210 437.820 3274.530 ;
        RECT 437.620 3260.000 437.760 3274.210 ;
        RECT 437.510 3256.000 437.790 3260.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 3153.060 17.870 3153.120 ;
        RECT 296.770 3153.060 297.090 3153.120 ;
        RECT 17.550 3152.920 297.090 3153.060 ;
        RECT 17.550 3152.860 17.870 3152.920 ;
        RECT 296.770 3152.860 297.090 3152.920 ;
      LAYER via ;
        RECT 17.580 3152.860 17.840 3153.120 ;
        RECT 296.800 3152.860 297.060 3153.120 ;
      LAYER met2 ;
        RECT 17.570 3393.355 17.850 3393.725 ;
        RECT 17.640 3153.150 17.780 3393.355 ;
        RECT 17.580 3152.830 17.840 3153.150 ;
        RECT 296.800 3152.830 297.060 3153.150 ;
        RECT 296.860 3152.325 297.000 3152.830 ;
        RECT 296.790 3151.955 297.070 3152.325 ;
      LAYER via2 ;
        RECT 17.570 3393.400 17.850 3393.680 ;
        RECT 296.790 3152.000 297.070 3152.280 ;
      LAYER met3 ;
        RECT -4.800 3393.690 2.400 3394.140 ;
        RECT 17.545 3393.690 17.875 3393.705 ;
        RECT -4.800 3393.390 17.875 3393.690 ;
        RECT -4.800 3392.940 2.400 3393.390 ;
        RECT 17.545 3393.375 17.875 3393.390 ;
        RECT 296.765 3152.290 297.095 3152.305 ;
        RECT 310.000 3152.290 314.000 3152.680 ;
        RECT 296.765 3152.080 314.000 3152.290 ;
        RECT 296.765 3151.990 310.500 3152.080 ;
        RECT 296.765 3151.975 297.095 3151.990 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2939.200 17.410 2939.260 ;
        RECT 296.770 2939.200 297.090 2939.260 ;
        RECT 17.090 2939.060 297.090 2939.200 ;
        RECT 17.090 2939.000 17.410 2939.060 ;
        RECT 296.770 2939.000 297.090 2939.060 ;
      LAYER via ;
        RECT 17.120 2939.000 17.380 2939.260 ;
        RECT 296.800 2939.000 297.060 2939.260 ;
      LAYER met2 ;
        RECT 17.110 3141.755 17.390 3142.125 ;
        RECT 17.180 2939.290 17.320 3141.755 ;
        RECT 17.120 2938.970 17.380 2939.290 ;
        RECT 296.800 2938.970 297.060 2939.290 ;
        RECT 296.860 2938.125 297.000 2938.970 ;
        RECT 296.790 2937.755 297.070 2938.125 ;
      LAYER via2 ;
        RECT 17.110 3141.800 17.390 3142.080 ;
        RECT 296.790 2937.800 297.070 2938.080 ;
      LAYER met3 ;
        RECT -4.800 3142.090 2.400 3142.540 ;
        RECT 17.085 3142.090 17.415 3142.105 ;
        RECT -4.800 3141.790 17.415 3142.090 ;
        RECT -4.800 3141.340 2.400 3141.790 ;
        RECT 17.085 3141.775 17.415 3141.790 ;
        RECT 296.765 2938.090 297.095 2938.105 ;
        RECT 310.000 2938.090 314.000 2938.480 ;
        RECT 296.765 2937.880 314.000 2938.090 ;
        RECT 296.765 2937.790 310.500 2937.880 ;
        RECT 296.765 2937.775 297.095 2937.790 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2725.340 17.410 2725.400 ;
        RECT 296.770 2725.340 297.090 2725.400 ;
        RECT 17.090 2725.200 297.090 2725.340 ;
        RECT 17.090 2725.140 17.410 2725.200 ;
        RECT 296.770 2725.140 297.090 2725.200 ;
      LAYER via ;
        RECT 17.120 2725.140 17.380 2725.400 ;
        RECT 296.800 2725.140 297.060 2725.400 ;
      LAYER met2 ;
        RECT 17.110 2890.835 17.390 2891.205 ;
        RECT 17.180 2725.430 17.320 2890.835 ;
        RECT 17.120 2725.110 17.380 2725.430 ;
        RECT 296.800 2725.110 297.060 2725.430 ;
        RECT 296.860 2723.925 297.000 2725.110 ;
        RECT 296.790 2723.555 297.070 2723.925 ;
      LAYER via2 ;
        RECT 17.110 2890.880 17.390 2891.160 ;
        RECT 296.790 2723.600 297.070 2723.880 ;
      LAYER met3 ;
        RECT -4.800 2891.170 2.400 2891.620 ;
        RECT 17.085 2891.170 17.415 2891.185 ;
        RECT -4.800 2890.870 17.415 2891.170 ;
        RECT -4.800 2890.420 2.400 2890.870 ;
        RECT 17.085 2890.855 17.415 2890.870 ;
        RECT 296.765 2723.890 297.095 2723.905 ;
        RECT 310.000 2723.890 314.000 2724.280 ;
        RECT 296.765 2723.680 314.000 2723.890 ;
        RECT 296.765 2723.590 310.500 2723.680 ;
        RECT 296.765 2723.575 297.095 2723.590 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2511.480 17.410 2511.540 ;
        RECT 296.770 2511.480 297.090 2511.540 ;
        RECT 17.090 2511.340 297.090 2511.480 ;
        RECT 17.090 2511.280 17.410 2511.340 ;
        RECT 296.770 2511.280 297.090 2511.340 ;
      LAYER via ;
        RECT 17.120 2511.280 17.380 2511.540 ;
        RECT 296.800 2511.280 297.060 2511.540 ;
      LAYER met2 ;
        RECT 17.110 2639.235 17.390 2639.605 ;
        RECT 17.180 2511.570 17.320 2639.235 ;
        RECT 17.120 2511.250 17.380 2511.570 ;
        RECT 296.800 2511.250 297.060 2511.570 ;
        RECT 296.860 2509.725 297.000 2511.250 ;
        RECT 296.790 2509.355 297.070 2509.725 ;
      LAYER via2 ;
        RECT 17.110 2639.280 17.390 2639.560 ;
        RECT 296.790 2509.400 297.070 2509.680 ;
      LAYER met3 ;
        RECT -4.800 2639.570 2.400 2640.020 ;
        RECT 17.085 2639.570 17.415 2639.585 ;
        RECT -4.800 2639.270 17.415 2639.570 ;
        RECT -4.800 2638.820 2.400 2639.270 ;
        RECT 17.085 2639.255 17.415 2639.270 ;
        RECT 296.765 2509.690 297.095 2509.705 ;
        RECT 310.000 2509.690 314.000 2510.080 ;
        RECT 296.765 2509.480 314.000 2509.690 ;
        RECT 296.765 2509.390 310.500 2509.480 ;
        RECT 296.765 2509.375 297.095 2509.390 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2297.620 17.870 2297.680 ;
        RECT 296.770 2297.620 297.090 2297.680 ;
        RECT 17.550 2297.480 297.090 2297.620 ;
        RECT 17.550 2297.420 17.870 2297.480 ;
        RECT 296.770 2297.420 297.090 2297.480 ;
      LAYER via ;
        RECT 17.580 2297.420 17.840 2297.680 ;
        RECT 296.800 2297.420 297.060 2297.680 ;
      LAYER met2 ;
        RECT 17.570 2387.635 17.850 2388.005 ;
        RECT 17.640 2297.710 17.780 2387.635 ;
        RECT 17.580 2297.390 17.840 2297.710 ;
        RECT 296.800 2297.390 297.060 2297.710 ;
        RECT 296.860 2295.525 297.000 2297.390 ;
        RECT 296.790 2295.155 297.070 2295.525 ;
      LAYER via2 ;
        RECT 17.570 2387.680 17.850 2387.960 ;
        RECT 296.790 2295.200 297.070 2295.480 ;
      LAYER met3 ;
        RECT -4.800 2387.970 2.400 2388.420 ;
        RECT 17.545 2387.970 17.875 2387.985 ;
        RECT -4.800 2387.670 17.875 2387.970 ;
        RECT -4.800 2387.220 2.400 2387.670 ;
        RECT 17.545 2387.655 17.875 2387.670 ;
        RECT 296.765 2295.490 297.095 2295.505 ;
        RECT 310.000 2295.490 314.000 2295.880 ;
        RECT 296.765 2295.280 314.000 2295.490 ;
        RECT 296.765 2295.190 310.500 2295.280 ;
        RECT 296.765 2295.175 297.095 2295.190 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2083.760 17.410 2083.820 ;
        RECT 296.770 2083.760 297.090 2083.820 ;
        RECT 17.090 2083.620 297.090 2083.760 ;
        RECT 17.090 2083.560 17.410 2083.620 ;
        RECT 296.770 2083.560 297.090 2083.620 ;
      LAYER via ;
        RECT 17.120 2083.560 17.380 2083.820 ;
        RECT 296.800 2083.560 297.060 2083.820 ;
      LAYER met2 ;
        RECT 17.110 2136.035 17.390 2136.405 ;
        RECT 17.180 2083.850 17.320 2136.035 ;
        RECT 17.120 2083.530 17.380 2083.850 ;
        RECT 296.800 2083.530 297.060 2083.850 ;
        RECT 296.860 2081.325 297.000 2083.530 ;
        RECT 296.790 2080.955 297.070 2081.325 ;
      LAYER via2 ;
        RECT 17.110 2136.080 17.390 2136.360 ;
        RECT 296.790 2081.000 297.070 2081.280 ;
      LAYER met3 ;
        RECT -4.800 2136.370 2.400 2136.820 ;
        RECT 17.085 2136.370 17.415 2136.385 ;
        RECT -4.800 2136.070 17.415 2136.370 ;
        RECT -4.800 2135.620 2.400 2136.070 ;
        RECT 17.085 2136.055 17.415 2136.070 ;
        RECT 296.765 2081.290 297.095 2081.305 ;
        RECT 310.000 2081.290 314.000 2081.680 ;
        RECT 296.765 2081.080 314.000 2081.290 ;
        RECT 296.765 2080.990 310.500 2081.080 ;
        RECT 296.765 2080.975 297.095 2080.990 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 593.200 2618.710 593.260 ;
        RECT 2900.830 593.200 2901.150 593.260 ;
        RECT 2618.390 593.060 2901.150 593.200 ;
        RECT 2618.390 593.000 2618.710 593.060 ;
        RECT 2900.830 593.000 2901.150 593.060 ;
      LAYER via ;
        RECT 2618.420 593.000 2618.680 593.260 ;
        RECT 2900.860 593.000 2901.120 593.260 ;
      LAYER met2 ;
        RECT 2618.410 759.715 2618.690 760.085 ;
        RECT 2618.480 593.290 2618.620 759.715 ;
        RECT 2618.420 592.970 2618.680 593.290 ;
        RECT 2900.860 592.970 2901.120 593.290 ;
        RECT 2900.920 586.685 2901.060 592.970 ;
        RECT 2900.850 586.315 2901.130 586.685 ;
      LAYER via2 ;
        RECT 2618.410 759.760 2618.690 760.040 ;
        RECT 2900.850 586.360 2901.130 586.640 ;
      LAYER met3 ;
        RECT 2606.000 760.050 2610.000 760.440 ;
        RECT 2618.385 760.050 2618.715 760.065 ;
        RECT 2606.000 759.840 2618.715 760.050 ;
        RECT 2609.580 759.750 2618.715 759.840 ;
        RECT 2618.385 759.735 2618.715 759.750 ;
        RECT 2900.825 586.650 2901.155 586.665 ;
        RECT 2917.600 586.650 2924.800 587.100 ;
        RECT 2900.825 586.350 2924.800 586.650 ;
        RECT 2900.825 586.335 2901.155 586.350 ;
        RECT 2917.600 585.900 2924.800 586.350 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1869.900 17.410 1869.960 ;
        RECT 296.770 1869.900 297.090 1869.960 ;
        RECT 17.090 1869.760 297.090 1869.900 ;
        RECT 17.090 1869.700 17.410 1869.760 ;
        RECT 296.770 1869.700 297.090 1869.760 ;
      LAYER via ;
        RECT 17.120 1869.700 17.380 1869.960 ;
        RECT 296.800 1869.700 297.060 1869.960 ;
      LAYER met2 ;
        RECT 17.110 1885.115 17.390 1885.485 ;
        RECT 17.180 1869.990 17.320 1885.115 ;
        RECT 17.120 1869.670 17.380 1869.990 ;
        RECT 296.800 1869.670 297.060 1869.990 ;
        RECT 296.860 1867.125 297.000 1869.670 ;
        RECT 296.790 1866.755 297.070 1867.125 ;
      LAYER via2 ;
        RECT 17.110 1885.160 17.390 1885.440 ;
        RECT 296.790 1866.800 297.070 1867.080 ;
      LAYER met3 ;
        RECT -4.800 1885.450 2.400 1885.900 ;
        RECT 17.085 1885.450 17.415 1885.465 ;
        RECT -4.800 1885.150 17.415 1885.450 ;
        RECT -4.800 1884.700 2.400 1885.150 ;
        RECT 17.085 1885.135 17.415 1885.150 ;
        RECT 296.765 1867.090 297.095 1867.105 ;
        RECT 310.000 1867.090 314.000 1867.480 ;
        RECT 296.765 1866.880 314.000 1867.090 ;
        RECT 296.765 1866.790 310.500 1866.880 ;
        RECT 296.765 1866.775 297.095 1866.790 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1635.300 16.950 1635.360 ;
        RECT 296.770 1635.300 297.090 1635.360 ;
        RECT 16.630 1635.160 297.090 1635.300 ;
        RECT 16.630 1635.100 16.950 1635.160 ;
        RECT 296.770 1635.100 297.090 1635.160 ;
      LAYER via ;
        RECT 16.660 1635.100 16.920 1635.360 ;
        RECT 296.800 1635.100 297.060 1635.360 ;
      LAYER met2 ;
        RECT 296.790 1651.875 297.070 1652.245 ;
        RECT 296.860 1635.390 297.000 1651.875 ;
        RECT 16.660 1635.070 16.920 1635.390 ;
        RECT 296.800 1635.070 297.060 1635.390 ;
        RECT 16.720 1633.885 16.860 1635.070 ;
        RECT 16.650 1633.515 16.930 1633.885 ;
      LAYER via2 ;
        RECT 296.790 1651.920 297.070 1652.200 ;
        RECT 16.650 1633.560 16.930 1633.840 ;
      LAYER met3 ;
        RECT 296.765 1652.210 297.095 1652.225 ;
        RECT 310.000 1652.210 314.000 1652.600 ;
        RECT 296.765 1652.000 314.000 1652.210 ;
        RECT 296.765 1651.910 310.500 1652.000 ;
        RECT 296.765 1651.895 297.095 1651.910 ;
        RECT -4.800 1633.850 2.400 1634.300 ;
        RECT 16.625 1633.850 16.955 1633.865 ;
        RECT -4.800 1633.550 16.955 1633.850 ;
        RECT -4.800 1633.100 2.400 1633.550 ;
        RECT 16.625 1633.535 16.955 1633.550 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1386.760 17.410 1386.820 ;
        RECT 299.990 1386.760 300.310 1386.820 ;
        RECT 17.090 1386.620 300.310 1386.760 ;
        RECT 17.090 1386.560 17.410 1386.620 ;
        RECT 299.990 1386.560 300.310 1386.620 ;
      LAYER via ;
        RECT 17.120 1386.560 17.380 1386.820 ;
        RECT 300.020 1386.560 300.280 1386.820 ;
      LAYER met2 ;
        RECT 300.010 1437.675 300.290 1438.045 ;
        RECT 300.080 1386.850 300.220 1437.675 ;
        RECT 17.120 1386.530 17.380 1386.850 ;
        RECT 300.020 1386.530 300.280 1386.850 ;
        RECT 17.180 1382.285 17.320 1386.530 ;
        RECT 17.110 1381.915 17.390 1382.285 ;
      LAYER via2 ;
        RECT 300.010 1437.720 300.290 1438.000 ;
        RECT 17.110 1381.960 17.390 1382.240 ;
      LAYER met3 ;
        RECT 299.985 1438.010 300.315 1438.025 ;
        RECT 310.000 1438.010 314.000 1438.400 ;
        RECT 299.985 1437.800 314.000 1438.010 ;
        RECT 299.985 1437.710 310.500 1437.800 ;
        RECT 299.985 1437.695 300.315 1437.710 ;
        RECT -4.800 1382.250 2.400 1382.700 ;
        RECT 17.085 1382.250 17.415 1382.265 ;
        RECT -4.800 1381.950 17.415 1382.250 ;
        RECT -4.800 1381.500 2.400 1381.950 ;
        RECT 17.085 1381.935 17.415 1381.950 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1131.420 17.410 1131.480 ;
        RECT 300.450 1131.420 300.770 1131.480 ;
        RECT 17.090 1131.280 300.770 1131.420 ;
        RECT 17.090 1131.220 17.410 1131.280 ;
        RECT 300.450 1131.220 300.770 1131.280 ;
      LAYER via ;
        RECT 17.120 1131.220 17.380 1131.480 ;
        RECT 300.480 1131.220 300.740 1131.480 ;
      LAYER met2 ;
        RECT 300.470 1223.475 300.750 1223.845 ;
        RECT 300.540 1131.510 300.680 1223.475 ;
        RECT 17.120 1131.365 17.380 1131.510 ;
        RECT 17.110 1130.995 17.390 1131.365 ;
        RECT 300.480 1131.190 300.740 1131.510 ;
      LAYER via2 ;
        RECT 300.470 1223.520 300.750 1223.800 ;
        RECT 17.110 1131.040 17.390 1131.320 ;
      LAYER met3 ;
        RECT 300.445 1223.810 300.775 1223.825 ;
        RECT 310.000 1223.810 314.000 1224.200 ;
        RECT 300.445 1223.600 314.000 1223.810 ;
        RECT 300.445 1223.510 310.500 1223.600 ;
        RECT 300.445 1223.495 300.775 1223.510 ;
        RECT -4.800 1131.330 2.400 1131.780 ;
        RECT 17.085 1131.330 17.415 1131.345 ;
        RECT -4.800 1131.030 17.415 1131.330 ;
        RECT -4.800 1130.580 2.400 1131.030 ;
        RECT 17.085 1131.015 17.415 1131.030 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 883.220 17.410 883.280 ;
        RECT 299.990 883.220 300.310 883.280 ;
        RECT 17.090 883.080 300.310 883.220 ;
        RECT 17.090 883.020 17.410 883.080 ;
        RECT 299.990 883.020 300.310 883.080 ;
      LAYER via ;
        RECT 17.120 883.020 17.380 883.280 ;
        RECT 300.020 883.020 300.280 883.280 ;
      LAYER met2 ;
        RECT 300.010 1009.275 300.290 1009.645 ;
        RECT 300.080 883.310 300.220 1009.275 ;
        RECT 17.120 882.990 17.380 883.310 ;
        RECT 300.020 882.990 300.280 883.310 ;
        RECT 17.180 879.765 17.320 882.990 ;
        RECT 17.110 879.395 17.390 879.765 ;
      LAYER via2 ;
        RECT 300.010 1009.320 300.290 1009.600 ;
        RECT 17.110 879.440 17.390 879.720 ;
      LAYER met3 ;
        RECT 299.985 1009.610 300.315 1009.625 ;
        RECT 310.000 1009.610 314.000 1010.000 ;
        RECT 299.985 1009.400 314.000 1009.610 ;
        RECT 299.985 1009.310 310.500 1009.400 ;
        RECT 299.985 1009.295 300.315 1009.310 ;
        RECT -4.800 879.730 2.400 880.180 ;
        RECT 17.085 879.730 17.415 879.745 ;
        RECT -4.800 879.430 17.415 879.730 ;
        RECT -4.800 878.980 2.400 879.430 ;
        RECT 17.085 879.415 17.415 879.430 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 634.680 16.490 634.740 ;
        RECT 299.990 634.680 300.310 634.740 ;
        RECT 16.170 634.540 300.310 634.680 ;
        RECT 16.170 634.480 16.490 634.540 ;
        RECT 299.990 634.480 300.310 634.540 ;
      LAYER via ;
        RECT 16.200 634.480 16.460 634.740 ;
        RECT 300.020 634.480 300.280 634.740 ;
      LAYER met2 ;
        RECT 300.010 795.075 300.290 795.445 ;
        RECT 300.080 634.770 300.220 795.075 ;
        RECT 16.200 634.450 16.460 634.770 ;
        RECT 300.020 634.450 300.280 634.770 ;
        RECT 16.260 628.165 16.400 634.450 ;
        RECT 16.190 627.795 16.470 628.165 ;
      LAYER via2 ;
        RECT 300.010 795.120 300.290 795.400 ;
        RECT 16.190 627.840 16.470 628.120 ;
      LAYER met3 ;
        RECT 299.985 795.410 300.315 795.425 ;
        RECT 310.000 795.410 314.000 795.800 ;
        RECT 299.985 795.200 314.000 795.410 ;
        RECT 299.985 795.110 310.500 795.200 ;
        RECT 299.985 795.095 300.315 795.110 ;
        RECT -4.800 628.130 2.400 628.580 ;
        RECT 16.165 628.130 16.495 628.145 ;
        RECT -4.800 627.830 16.495 628.130 ;
        RECT -4.800 627.380 2.400 627.830 ;
        RECT 16.165 627.815 16.495 627.830 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 379.340 17.410 379.400 ;
        RECT 299.990 379.340 300.310 379.400 ;
        RECT 17.090 379.200 300.310 379.340 ;
        RECT 17.090 379.140 17.410 379.200 ;
        RECT 299.990 379.140 300.310 379.200 ;
      LAYER via ;
        RECT 17.120 379.140 17.380 379.400 ;
        RECT 300.020 379.140 300.280 379.400 ;
      LAYER met2 ;
        RECT 300.010 580.875 300.290 581.245 ;
        RECT 300.080 379.430 300.220 580.875 ;
        RECT 17.120 379.110 17.380 379.430 ;
        RECT 300.020 379.110 300.280 379.430 ;
        RECT 17.180 376.565 17.320 379.110 ;
        RECT 17.110 376.195 17.390 376.565 ;
      LAYER via2 ;
        RECT 300.010 580.920 300.290 581.200 ;
        RECT 17.110 376.240 17.390 376.520 ;
      LAYER met3 ;
        RECT 299.985 581.210 300.315 581.225 ;
        RECT 310.000 581.210 314.000 581.600 ;
        RECT 299.985 581.000 314.000 581.210 ;
        RECT 299.985 580.910 310.500 581.000 ;
        RECT 299.985 580.895 300.315 580.910 ;
        RECT -4.800 376.530 2.400 376.980 ;
        RECT 17.085 376.530 17.415 376.545 ;
        RECT -4.800 376.230 17.415 376.530 ;
        RECT -4.800 375.780 2.400 376.230 ;
        RECT 17.085 376.215 17.415 376.230 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 131.140 17.410 131.200 ;
        RECT 300.450 131.140 300.770 131.200 ;
        RECT 17.090 131.000 300.770 131.140 ;
        RECT 17.090 130.940 17.410 131.000 ;
        RECT 300.450 130.940 300.770 131.000 ;
      LAYER via ;
        RECT 17.120 130.940 17.380 131.200 ;
        RECT 300.480 130.940 300.740 131.200 ;
      LAYER met2 ;
        RECT 300.470 366.675 300.750 367.045 ;
        RECT 300.540 131.230 300.680 366.675 ;
        RECT 17.120 130.910 17.380 131.230 ;
        RECT 300.480 130.910 300.740 131.230 ;
        RECT 17.180 125.645 17.320 130.910 ;
        RECT 17.110 125.275 17.390 125.645 ;
      LAYER via2 ;
        RECT 300.470 366.720 300.750 367.000 ;
        RECT 17.110 125.320 17.390 125.600 ;
      LAYER met3 ;
        RECT 300.445 367.010 300.775 367.025 ;
        RECT 310.000 367.010 314.000 367.400 ;
        RECT 300.445 366.800 314.000 367.010 ;
        RECT 300.445 366.710 310.500 366.800 ;
        RECT 300.445 366.695 300.775 366.710 ;
        RECT -4.800 125.610 2.400 126.060 ;
        RECT 17.085 125.610 17.415 125.625 ;
        RECT -4.800 125.310 17.415 125.610 ;
        RECT -4.800 124.860 2.400 125.310 ;
        RECT 17.085 125.295 17.415 125.310 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 827.800 2618.710 827.860 ;
        RECT 2900.830 827.800 2901.150 827.860 ;
        RECT 2618.390 827.660 2901.150 827.800 ;
        RECT 2618.390 827.600 2618.710 827.660 ;
        RECT 2900.830 827.600 2901.150 827.660 ;
      LAYER via ;
        RECT 2618.420 827.600 2618.680 827.860 ;
        RECT 2900.860 827.600 2901.120 827.860 ;
      LAYER met2 ;
        RECT 2618.410 959.635 2618.690 960.005 ;
        RECT 2618.480 827.890 2618.620 959.635 ;
        RECT 2618.420 827.570 2618.680 827.890 ;
        RECT 2900.860 827.570 2901.120 827.890 ;
        RECT 2900.920 821.285 2901.060 827.570 ;
        RECT 2900.850 820.915 2901.130 821.285 ;
      LAYER via2 ;
        RECT 2618.410 959.680 2618.690 959.960 ;
        RECT 2900.850 820.960 2901.130 821.240 ;
      LAYER met3 ;
        RECT 2606.000 959.970 2610.000 960.360 ;
        RECT 2618.385 959.970 2618.715 959.985 ;
        RECT 2606.000 959.760 2618.715 959.970 ;
        RECT 2609.580 959.670 2618.715 959.760 ;
        RECT 2618.385 959.655 2618.715 959.670 ;
        RECT 2900.825 821.250 2901.155 821.265 ;
        RECT 2917.600 821.250 2924.800 821.700 ;
        RECT 2900.825 820.950 2924.800 821.250 ;
        RECT 2900.825 820.935 2901.155 820.950 ;
        RECT 2917.600 820.500 2924.800 820.950 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1062.400 2619.170 1062.460 ;
        RECT 2900.830 1062.400 2901.150 1062.460 ;
        RECT 2618.850 1062.260 2901.150 1062.400 ;
        RECT 2618.850 1062.200 2619.170 1062.260 ;
        RECT 2900.830 1062.200 2901.150 1062.260 ;
      LAYER via ;
        RECT 2618.880 1062.200 2619.140 1062.460 ;
        RECT 2900.860 1062.200 2901.120 1062.460 ;
      LAYER met2 ;
        RECT 2618.870 1159.555 2619.150 1159.925 ;
        RECT 2618.940 1062.490 2619.080 1159.555 ;
        RECT 2618.880 1062.170 2619.140 1062.490 ;
        RECT 2900.860 1062.170 2901.120 1062.490 ;
        RECT 2900.920 1055.885 2901.060 1062.170 ;
        RECT 2900.850 1055.515 2901.130 1055.885 ;
      LAYER via2 ;
        RECT 2618.870 1159.600 2619.150 1159.880 ;
        RECT 2900.850 1055.560 2901.130 1055.840 ;
      LAYER met3 ;
        RECT 2606.000 1159.890 2610.000 1160.280 ;
        RECT 2618.845 1159.890 2619.175 1159.905 ;
        RECT 2606.000 1159.680 2619.175 1159.890 ;
        RECT 2609.580 1159.590 2619.175 1159.680 ;
        RECT 2618.845 1159.575 2619.175 1159.590 ;
        RECT 2900.825 1055.850 2901.155 1055.865 ;
        RECT 2917.600 1055.850 2924.800 1056.300 ;
        RECT 2900.825 1055.550 2924.800 1055.850 ;
        RECT 2900.825 1055.535 2901.155 1055.550 ;
        RECT 2917.600 1055.100 2924.800 1055.550 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1297.000 2618.710 1297.060 ;
        RECT 2900.830 1297.000 2901.150 1297.060 ;
        RECT 2618.390 1296.860 2901.150 1297.000 ;
        RECT 2618.390 1296.800 2618.710 1296.860 ;
        RECT 2900.830 1296.800 2901.150 1296.860 ;
      LAYER via ;
        RECT 2618.420 1296.800 2618.680 1297.060 ;
        RECT 2900.860 1296.800 2901.120 1297.060 ;
      LAYER met2 ;
        RECT 2618.410 1359.475 2618.690 1359.845 ;
        RECT 2618.480 1297.090 2618.620 1359.475 ;
        RECT 2618.420 1296.770 2618.680 1297.090 ;
        RECT 2900.860 1296.770 2901.120 1297.090 ;
        RECT 2900.920 1290.485 2901.060 1296.770 ;
        RECT 2900.850 1290.115 2901.130 1290.485 ;
      LAYER via2 ;
        RECT 2618.410 1359.520 2618.690 1359.800 ;
        RECT 2900.850 1290.160 2901.130 1290.440 ;
      LAYER met3 ;
        RECT 2606.000 1359.810 2610.000 1360.200 ;
        RECT 2618.385 1359.810 2618.715 1359.825 ;
        RECT 2606.000 1359.600 2618.715 1359.810 ;
        RECT 2609.580 1359.510 2618.715 1359.600 ;
        RECT 2618.385 1359.495 2618.715 1359.510 ;
        RECT 2900.825 1290.450 2901.155 1290.465 ;
        RECT 2917.600 1290.450 2924.800 1290.900 ;
        RECT 2900.825 1290.150 2924.800 1290.450 ;
        RECT 2900.825 1290.135 2901.155 1290.150 ;
        RECT 2917.600 1289.700 2924.800 1290.150 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1531.600 2618.710 1531.660 ;
        RECT 2900.830 1531.600 2901.150 1531.660 ;
        RECT 2618.390 1531.460 2901.150 1531.600 ;
        RECT 2618.390 1531.400 2618.710 1531.460 ;
        RECT 2900.830 1531.400 2901.150 1531.460 ;
      LAYER via ;
        RECT 2618.420 1531.400 2618.680 1531.660 ;
        RECT 2900.860 1531.400 2901.120 1531.660 ;
      LAYER met2 ;
        RECT 2618.410 1559.395 2618.690 1559.765 ;
        RECT 2618.480 1531.690 2618.620 1559.395 ;
        RECT 2618.420 1531.370 2618.680 1531.690 ;
        RECT 2900.860 1531.370 2901.120 1531.690 ;
        RECT 2900.920 1525.085 2901.060 1531.370 ;
        RECT 2900.850 1524.715 2901.130 1525.085 ;
      LAYER via2 ;
        RECT 2618.410 1559.440 2618.690 1559.720 ;
        RECT 2900.850 1524.760 2901.130 1525.040 ;
      LAYER met3 ;
        RECT 2606.000 1559.730 2610.000 1560.120 ;
        RECT 2618.385 1559.730 2618.715 1559.745 ;
        RECT 2606.000 1559.520 2618.715 1559.730 ;
        RECT 2609.580 1559.430 2618.715 1559.520 ;
        RECT 2618.385 1559.415 2618.715 1559.430 ;
        RECT 2900.825 1525.050 2901.155 1525.065 ;
        RECT 2917.600 1525.050 2924.800 1525.500 ;
        RECT 2900.825 1524.750 2924.800 1525.050 ;
        RECT 2900.825 1524.735 2901.155 1524.750 ;
        RECT 2917.600 1524.300 2924.800 1524.750 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1762.800 2621.930 1762.860 ;
        RECT 2900.830 1762.800 2901.150 1762.860 ;
        RECT 2621.610 1762.660 2901.150 1762.800 ;
        RECT 2621.610 1762.600 2621.930 1762.660 ;
        RECT 2900.830 1762.600 2901.150 1762.660 ;
      LAYER via ;
        RECT 2621.640 1762.600 2621.900 1762.860 ;
        RECT 2900.860 1762.600 2901.120 1762.860 ;
      LAYER met2 ;
        RECT 2621.640 1762.570 2621.900 1762.890 ;
        RECT 2900.860 1762.570 2901.120 1762.890 ;
        RECT 2621.700 1759.685 2621.840 1762.570 ;
        RECT 2900.920 1759.685 2901.060 1762.570 ;
        RECT 2621.630 1759.315 2621.910 1759.685 ;
        RECT 2900.850 1759.315 2901.130 1759.685 ;
      LAYER via2 ;
        RECT 2621.630 1759.360 2621.910 1759.640 ;
        RECT 2900.850 1759.360 2901.130 1759.640 ;
      LAYER met3 ;
        RECT 2606.000 1759.650 2610.000 1760.040 ;
        RECT 2621.605 1759.650 2621.935 1759.665 ;
        RECT 2606.000 1759.440 2621.935 1759.650 ;
        RECT 2609.580 1759.350 2621.935 1759.440 ;
        RECT 2621.605 1759.335 2621.935 1759.350 ;
        RECT 2900.825 1759.650 2901.155 1759.665 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2900.825 1759.350 2924.800 1759.650 ;
        RECT 2900.825 1759.335 2901.155 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1994.340 2618.710 1994.400 ;
        RECT 2900.830 1994.340 2901.150 1994.400 ;
        RECT 2618.390 1994.200 2901.150 1994.340 ;
        RECT 2618.390 1994.140 2618.710 1994.200 ;
        RECT 2900.830 1994.140 2901.150 1994.200 ;
      LAYER via ;
        RECT 2618.420 1994.140 2618.680 1994.400 ;
        RECT 2900.860 1994.140 2901.120 1994.400 ;
      LAYER met2 ;
        RECT 2618.420 1994.110 2618.680 1994.430 ;
        RECT 2900.860 1994.285 2901.120 1994.430 ;
        RECT 2618.480 1960.285 2618.620 1994.110 ;
        RECT 2900.850 1993.915 2901.130 1994.285 ;
        RECT 2618.410 1959.915 2618.690 1960.285 ;
      LAYER via2 ;
        RECT 2900.850 1993.960 2901.130 1994.240 ;
        RECT 2618.410 1959.960 2618.690 1960.240 ;
      LAYER met3 ;
        RECT 2900.825 1994.250 2901.155 1994.265 ;
        RECT 2917.600 1994.250 2924.800 1994.700 ;
        RECT 2900.825 1993.950 2924.800 1994.250 ;
        RECT 2900.825 1993.935 2901.155 1993.950 ;
        RECT 2917.600 1993.500 2924.800 1993.950 ;
        RECT 2606.000 1960.250 2610.000 1960.640 ;
        RECT 2618.385 1960.250 2618.715 1960.265 ;
        RECT 2606.000 1960.040 2618.715 1960.250 ;
        RECT 2609.580 1959.950 2618.715 1960.040 ;
        RECT 2618.385 1959.935 2618.715 1959.950 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2228.940 2618.710 2229.000 ;
        RECT 2900.830 2228.940 2901.150 2229.000 ;
        RECT 2618.390 2228.800 2901.150 2228.940 ;
        RECT 2618.390 2228.740 2618.710 2228.800 ;
        RECT 2900.830 2228.740 2901.150 2228.800 ;
      LAYER via ;
        RECT 2618.420 2228.740 2618.680 2229.000 ;
        RECT 2900.860 2228.740 2901.120 2229.000 ;
      LAYER met2 ;
        RECT 2618.420 2228.710 2618.680 2229.030 ;
        RECT 2900.860 2228.885 2901.120 2229.030 ;
        RECT 2618.480 2160.205 2618.620 2228.710 ;
        RECT 2900.850 2228.515 2901.130 2228.885 ;
        RECT 2618.410 2159.835 2618.690 2160.205 ;
      LAYER via2 ;
        RECT 2900.850 2228.560 2901.130 2228.840 ;
        RECT 2618.410 2159.880 2618.690 2160.160 ;
      LAYER met3 ;
        RECT 2900.825 2228.850 2901.155 2228.865 ;
        RECT 2917.600 2228.850 2924.800 2229.300 ;
        RECT 2900.825 2228.550 2924.800 2228.850 ;
        RECT 2900.825 2228.535 2901.155 2228.550 ;
        RECT 2917.600 2228.100 2924.800 2228.550 ;
        RECT 2606.000 2160.170 2610.000 2160.560 ;
        RECT 2618.385 2160.170 2618.715 2160.185 ;
        RECT 2606.000 2159.960 2618.715 2160.170 ;
        RECT 2609.580 2159.870 2618.715 2159.960 ;
        RECT 2618.385 2159.855 2618.715 2159.870 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 24.040 633.350 24.100 ;
        RECT 807.370 24.040 807.690 24.100 ;
        RECT 633.030 23.900 807.690 24.040 ;
        RECT 633.030 23.840 633.350 23.900 ;
        RECT 807.370 23.840 807.690 23.900 ;
      LAYER via ;
        RECT 633.060 23.840 633.320 24.100 ;
        RECT 807.400 23.840 807.660 24.100 ;
      LAYER met2 ;
        RECT 809.650 260.170 809.930 264.000 ;
        RECT 807.460 260.030 809.930 260.170 ;
        RECT 807.460 24.130 807.600 260.030 ;
        RECT 809.650 260.000 809.930 260.030 ;
        RECT 633.060 23.810 633.320 24.130 ;
        RECT 807.400 23.810 807.660 24.130 ;
        RECT 633.120 2.400 633.260 23.810 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2217.730 243.680 2218.050 243.740 ;
        RECT 2231.990 243.680 2232.310 243.740 ;
        RECT 2217.730 243.540 2232.310 243.680 ;
        RECT 2217.730 243.480 2218.050 243.540 ;
        RECT 2231.990 243.480 2232.310 243.540 ;
        RECT 2231.990 31.180 2232.310 31.240 ;
        RECT 2417.370 31.180 2417.690 31.240 ;
        RECT 2231.990 31.040 2417.690 31.180 ;
        RECT 2231.990 30.980 2232.310 31.040 ;
        RECT 2417.370 30.980 2417.690 31.040 ;
      LAYER via ;
        RECT 2217.760 243.480 2218.020 243.740 ;
        RECT 2232.020 243.480 2232.280 243.740 ;
        RECT 2232.020 30.980 2232.280 31.240 ;
        RECT 2417.400 30.980 2417.660 31.240 ;
      LAYER met2 ;
        RECT 2217.710 260.000 2217.990 264.000 ;
        RECT 2217.820 243.770 2217.960 260.000 ;
        RECT 2217.760 243.450 2218.020 243.770 ;
        RECT 2232.020 243.450 2232.280 243.770 ;
        RECT 2232.080 31.270 2232.220 243.450 ;
        RECT 2232.020 30.950 2232.280 31.270 ;
        RECT 2417.400 30.950 2417.660 31.270 ;
        RECT 2417.460 2.400 2417.600 30.950 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2235.210 38.320 2235.530 38.380 ;
        RECT 2434.850 38.320 2435.170 38.380 ;
        RECT 2235.210 38.180 2435.170 38.320 ;
        RECT 2235.210 38.120 2235.530 38.180 ;
        RECT 2434.850 38.120 2435.170 38.180 ;
      LAYER via ;
        RECT 2235.240 38.120 2235.500 38.380 ;
        RECT 2434.880 38.120 2435.140 38.380 ;
      LAYER met2 ;
        RECT 2231.970 260.170 2232.250 264.000 ;
        RECT 2231.970 260.030 2235.440 260.170 ;
        RECT 2231.970 260.000 2232.250 260.030 ;
        RECT 2235.300 38.410 2235.440 260.030 ;
        RECT 2235.240 38.090 2235.500 38.410 ;
        RECT 2434.880 38.090 2435.140 38.410 ;
        RECT 2434.940 2.400 2435.080 38.090 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2249.010 45.120 2249.330 45.180 ;
        RECT 2452.790 45.120 2453.110 45.180 ;
        RECT 2249.010 44.980 2453.110 45.120 ;
        RECT 2249.010 44.920 2249.330 44.980 ;
        RECT 2452.790 44.920 2453.110 44.980 ;
      LAYER via ;
        RECT 2249.040 44.920 2249.300 45.180 ;
        RECT 2452.820 44.920 2453.080 45.180 ;
      LAYER met2 ;
        RECT 2246.230 260.170 2246.510 264.000 ;
        RECT 2246.230 260.030 2249.240 260.170 ;
        RECT 2246.230 260.000 2246.510 260.030 ;
        RECT 2249.100 45.210 2249.240 260.030 ;
        RECT 2249.040 44.890 2249.300 45.210 ;
        RECT 2452.820 44.890 2453.080 45.210 ;
        RECT 2452.880 2.400 2453.020 44.890 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2262.810 51.580 2263.130 51.640 ;
        RECT 2470.730 51.580 2471.050 51.640 ;
        RECT 2262.810 51.440 2471.050 51.580 ;
        RECT 2262.810 51.380 2263.130 51.440 ;
        RECT 2470.730 51.380 2471.050 51.440 ;
      LAYER via ;
        RECT 2262.840 51.380 2263.100 51.640 ;
        RECT 2470.760 51.380 2471.020 51.640 ;
      LAYER met2 ;
        RECT 2260.030 260.170 2260.310 264.000 ;
        RECT 2260.030 260.030 2263.040 260.170 ;
        RECT 2260.030 260.000 2260.310 260.030 ;
        RECT 2262.900 51.670 2263.040 260.030 ;
        RECT 2262.840 51.350 2263.100 51.670 ;
        RECT 2470.760 51.350 2471.020 51.670 ;
        RECT 2470.820 2.400 2470.960 51.350 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2274.310 245.040 2274.630 245.100 ;
        RECT 2411.390 245.040 2411.710 245.100 ;
        RECT 2274.310 244.900 2411.710 245.040 ;
        RECT 2274.310 244.840 2274.630 244.900 ;
        RECT 2411.390 244.840 2411.710 244.900 ;
        RECT 2411.390 30.840 2411.710 30.900 ;
        RECT 2488.670 30.840 2488.990 30.900 ;
        RECT 2411.390 30.700 2488.990 30.840 ;
        RECT 2411.390 30.640 2411.710 30.700 ;
        RECT 2488.670 30.640 2488.990 30.700 ;
      LAYER via ;
        RECT 2274.340 244.840 2274.600 245.100 ;
        RECT 2411.420 244.840 2411.680 245.100 ;
        RECT 2411.420 30.640 2411.680 30.900 ;
        RECT 2488.700 30.640 2488.960 30.900 ;
      LAYER met2 ;
        RECT 2274.290 260.000 2274.570 264.000 ;
        RECT 2274.400 245.130 2274.540 260.000 ;
        RECT 2274.340 244.810 2274.600 245.130 ;
        RECT 2411.420 244.810 2411.680 245.130 ;
        RECT 2411.480 30.930 2411.620 244.810 ;
        RECT 2411.420 30.610 2411.680 30.930 ;
        RECT 2488.700 30.610 2488.960 30.930 ;
        RECT 2488.760 2.400 2488.900 30.610 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2290.410 58.720 2290.730 58.780 ;
        RECT 2504.770 58.720 2505.090 58.780 ;
        RECT 2290.410 58.580 2505.090 58.720 ;
        RECT 2290.410 58.520 2290.730 58.580 ;
        RECT 2504.770 58.520 2505.090 58.580 ;
      LAYER via ;
        RECT 2290.440 58.520 2290.700 58.780 ;
        RECT 2504.800 58.520 2505.060 58.780 ;
      LAYER met2 ;
        RECT 2288.090 260.170 2288.370 264.000 ;
        RECT 2288.090 260.030 2290.640 260.170 ;
        RECT 2288.090 260.000 2288.370 260.030 ;
        RECT 2290.500 58.810 2290.640 260.030 ;
        RECT 2290.440 58.490 2290.700 58.810 ;
        RECT 2504.800 58.490 2505.060 58.810 ;
        RECT 2504.860 16.730 2505.000 58.490 ;
        RECT 2504.860 16.590 2506.380 16.730 ;
        RECT 2506.240 2.400 2506.380 16.590 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2303.750 65.860 2304.070 65.920 ;
        RECT 2518.570 65.860 2518.890 65.920 ;
        RECT 2303.750 65.720 2518.890 65.860 ;
        RECT 2303.750 65.660 2304.070 65.720 ;
        RECT 2518.570 65.660 2518.890 65.720 ;
      LAYER via ;
        RECT 2303.780 65.660 2304.040 65.920 ;
        RECT 2518.600 65.660 2518.860 65.920 ;
      LAYER met2 ;
        RECT 2302.350 260.170 2302.630 264.000 ;
        RECT 2302.350 260.030 2303.980 260.170 ;
        RECT 2302.350 260.000 2302.630 260.030 ;
        RECT 2303.840 65.950 2303.980 260.030 ;
        RECT 2303.780 65.630 2304.040 65.950 ;
        RECT 2518.600 65.630 2518.860 65.950 ;
        RECT 2518.660 16.730 2518.800 65.630 ;
        RECT 2518.660 16.590 2524.320 16.730 ;
        RECT 2524.180 2.400 2524.320 16.590 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2317.550 72.320 2317.870 72.380 ;
        RECT 2539.270 72.320 2539.590 72.380 ;
        RECT 2317.550 72.180 2539.590 72.320 ;
        RECT 2317.550 72.120 2317.870 72.180 ;
        RECT 2539.270 72.120 2539.590 72.180 ;
      LAYER via ;
        RECT 2317.580 72.120 2317.840 72.380 ;
        RECT 2539.300 72.120 2539.560 72.380 ;
      LAYER met2 ;
        RECT 2316.610 260.170 2316.890 264.000 ;
        RECT 2316.610 260.030 2317.780 260.170 ;
        RECT 2316.610 260.000 2316.890 260.030 ;
        RECT 2317.640 72.410 2317.780 260.030 ;
        RECT 2317.580 72.090 2317.840 72.410 ;
        RECT 2539.300 72.090 2539.560 72.410 ;
        RECT 2539.360 16.730 2539.500 72.090 ;
        RECT 2539.360 16.590 2542.260 16.730 ;
        RECT 2542.120 2.400 2542.260 16.590 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2331.810 37.980 2332.130 38.040 ;
        RECT 2559.970 37.980 2560.290 38.040 ;
        RECT 2331.810 37.840 2560.290 37.980 ;
        RECT 2331.810 37.780 2332.130 37.840 ;
        RECT 2559.970 37.780 2560.290 37.840 ;
      LAYER via ;
        RECT 2331.840 37.780 2332.100 38.040 ;
        RECT 2560.000 37.780 2560.260 38.040 ;
      LAYER met2 ;
        RECT 2330.410 260.170 2330.690 264.000 ;
        RECT 2330.410 260.030 2332.040 260.170 ;
        RECT 2330.410 260.000 2330.690 260.030 ;
        RECT 2331.900 38.070 2332.040 260.030 ;
        RECT 2331.840 37.750 2332.100 38.070 ;
        RECT 2560.000 37.750 2560.260 38.070 ;
        RECT 2560.060 2.400 2560.200 37.750 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2344.690 243.680 2345.010 243.740 ;
        RECT 2349.290 243.680 2349.610 243.740 ;
        RECT 2344.690 243.540 2349.610 243.680 ;
        RECT 2344.690 243.480 2345.010 243.540 ;
        RECT 2349.290 243.480 2349.610 243.540 ;
        RECT 2349.290 79.460 2349.610 79.520 ;
        RECT 2573.770 79.460 2574.090 79.520 ;
        RECT 2349.290 79.320 2574.090 79.460 ;
        RECT 2349.290 79.260 2349.610 79.320 ;
        RECT 2573.770 79.260 2574.090 79.320 ;
      LAYER via ;
        RECT 2344.720 243.480 2344.980 243.740 ;
        RECT 2349.320 243.480 2349.580 243.740 ;
        RECT 2349.320 79.260 2349.580 79.520 ;
        RECT 2573.800 79.260 2574.060 79.520 ;
      LAYER met2 ;
        RECT 2344.670 260.000 2344.950 264.000 ;
        RECT 2344.780 243.770 2344.920 260.000 ;
        RECT 2344.720 243.450 2344.980 243.770 ;
        RECT 2349.320 243.450 2349.580 243.770 ;
        RECT 2349.380 79.550 2349.520 243.450 ;
        RECT 2349.320 79.230 2349.580 79.550 ;
        RECT 2573.800 79.230 2574.060 79.550 ;
        RECT 2573.860 16.730 2574.000 79.230 ;
        RECT 2573.860 16.590 2578.140 16.730 ;
        RECT 2578.000 2.400 2578.140 16.590 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 811.510 24.040 811.830 24.100 ;
        RECT 945.830 24.040 946.150 24.100 ;
        RECT 811.510 23.900 946.150 24.040 ;
        RECT 811.510 23.840 811.830 23.900 ;
        RECT 945.830 23.840 946.150 23.900 ;
      LAYER via ;
        RECT 811.540 23.840 811.800 24.100 ;
        RECT 945.860 23.840 946.120 24.100 ;
      LAYER met2 ;
        RECT 950.410 260.850 950.690 264.000 ;
        RECT 946.840 260.710 950.690 260.850 ;
        RECT 946.840 62.290 946.980 260.710 ;
        RECT 950.410 260.000 950.690 260.710 ;
        RECT 945.920 62.150 946.980 62.290 ;
        RECT 945.920 24.130 946.060 62.150 ;
        RECT 811.540 23.810 811.800 24.130 ;
        RECT 945.860 23.810 946.120 24.130 ;
        RECT 811.600 2.400 811.740 23.810 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2358.950 26.760 2359.270 26.820 ;
        RECT 2595.390 26.760 2595.710 26.820 ;
        RECT 2358.950 26.620 2595.710 26.760 ;
        RECT 2358.950 26.560 2359.270 26.620 ;
        RECT 2595.390 26.560 2595.710 26.620 ;
      LAYER via ;
        RECT 2358.980 26.560 2359.240 26.820 ;
        RECT 2595.420 26.560 2595.680 26.820 ;
      LAYER met2 ;
        RECT 2358.470 260.170 2358.750 264.000 ;
        RECT 2358.470 260.030 2359.180 260.170 ;
        RECT 2358.470 260.000 2358.750 260.030 ;
        RECT 2359.040 26.850 2359.180 260.030 ;
        RECT 2358.980 26.530 2359.240 26.850 ;
        RECT 2595.420 26.530 2595.680 26.850 ;
        RECT 2595.480 2.400 2595.620 26.530 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2372.750 26.420 2373.070 26.480 ;
        RECT 2613.330 26.420 2613.650 26.480 ;
        RECT 2372.750 26.280 2613.650 26.420 ;
        RECT 2372.750 26.220 2373.070 26.280 ;
        RECT 2613.330 26.220 2613.650 26.280 ;
      LAYER via ;
        RECT 2372.780 26.220 2373.040 26.480 ;
        RECT 2613.360 26.220 2613.620 26.480 ;
      LAYER met2 ;
        RECT 2372.730 260.000 2373.010 264.000 ;
        RECT 2372.840 26.510 2372.980 260.000 ;
        RECT 2372.780 26.190 2373.040 26.510 ;
        RECT 2613.360 26.190 2613.620 26.510 ;
        RECT 2613.420 2.400 2613.560 26.190 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2387.010 25.740 2387.330 25.800 ;
        RECT 2631.270 25.740 2631.590 25.800 ;
        RECT 2387.010 25.600 2631.590 25.740 ;
        RECT 2387.010 25.540 2387.330 25.600 ;
        RECT 2631.270 25.540 2631.590 25.600 ;
      LAYER via ;
        RECT 2387.040 25.540 2387.300 25.800 ;
        RECT 2631.300 25.540 2631.560 25.800 ;
      LAYER met2 ;
        RECT 2386.990 260.000 2387.270 264.000 ;
        RECT 2387.100 25.830 2387.240 260.000 ;
        RECT 2387.040 25.510 2387.300 25.830 ;
        RECT 2631.300 25.510 2631.560 25.830 ;
        RECT 2631.360 2.400 2631.500 25.510 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.350 25.400 2400.670 25.460 ;
        RECT 2649.210 25.400 2649.530 25.460 ;
        RECT 2400.350 25.260 2649.530 25.400 ;
        RECT 2400.350 25.200 2400.670 25.260 ;
        RECT 2649.210 25.200 2649.530 25.260 ;
      LAYER via ;
        RECT 2400.380 25.200 2400.640 25.460 ;
        RECT 2649.240 25.200 2649.500 25.460 ;
      LAYER met2 ;
        RECT 2400.790 260.170 2401.070 264.000 ;
        RECT 2400.440 260.030 2401.070 260.170 ;
        RECT 2400.440 25.490 2400.580 260.030 ;
        RECT 2400.790 260.000 2401.070 260.030 ;
        RECT 2400.380 25.170 2400.640 25.490 ;
        RECT 2649.240 25.170 2649.500 25.490 ;
        RECT 2649.300 2.400 2649.440 25.170 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2415.070 244.020 2415.390 244.080 ;
        RECT 2421.510 244.020 2421.830 244.080 ;
        RECT 2415.070 243.880 2421.830 244.020 ;
        RECT 2415.070 243.820 2415.390 243.880 ;
        RECT 2421.510 243.820 2421.830 243.880 ;
        RECT 2421.510 26.080 2421.830 26.140 ;
        RECT 2667.150 26.080 2667.470 26.140 ;
        RECT 2421.510 25.940 2667.470 26.080 ;
        RECT 2421.510 25.880 2421.830 25.940 ;
        RECT 2667.150 25.880 2667.470 25.940 ;
      LAYER via ;
        RECT 2415.100 243.820 2415.360 244.080 ;
        RECT 2421.540 243.820 2421.800 244.080 ;
        RECT 2421.540 25.880 2421.800 26.140 ;
        RECT 2667.180 25.880 2667.440 26.140 ;
      LAYER met2 ;
        RECT 2415.050 260.000 2415.330 264.000 ;
        RECT 2415.160 244.110 2415.300 260.000 ;
        RECT 2415.100 243.790 2415.360 244.110 ;
        RECT 2421.540 243.790 2421.800 244.110 ;
        RECT 2421.600 26.170 2421.740 243.790 ;
        RECT 2421.540 25.850 2421.800 26.170 ;
        RECT 2667.180 25.850 2667.440 26.170 ;
        RECT 2667.240 2.400 2667.380 25.850 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2429.330 242.660 2429.650 242.720 ;
        RECT 2435.310 242.660 2435.630 242.720 ;
        RECT 2429.330 242.520 2435.630 242.660 ;
        RECT 2429.330 242.460 2429.650 242.520 ;
        RECT 2435.310 242.460 2435.630 242.520 ;
        RECT 2435.310 24.720 2435.630 24.780 ;
        RECT 2684.630 24.720 2684.950 24.780 ;
        RECT 2435.310 24.580 2684.950 24.720 ;
        RECT 2435.310 24.520 2435.630 24.580 ;
        RECT 2684.630 24.520 2684.950 24.580 ;
      LAYER via ;
        RECT 2429.360 242.460 2429.620 242.720 ;
        RECT 2435.340 242.460 2435.600 242.720 ;
        RECT 2435.340 24.520 2435.600 24.780 ;
        RECT 2684.660 24.520 2684.920 24.780 ;
      LAYER met2 ;
        RECT 2429.310 260.000 2429.590 264.000 ;
        RECT 2429.420 242.750 2429.560 260.000 ;
        RECT 2429.360 242.430 2429.620 242.750 ;
        RECT 2435.340 242.430 2435.600 242.750 ;
        RECT 2435.400 24.810 2435.540 242.430 ;
        RECT 2435.340 24.490 2435.600 24.810 ;
        RECT 2684.660 24.490 2684.920 24.810 ;
        RECT 2684.720 2.400 2684.860 24.490 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2448.265 193.205 2448.435 240.975 ;
        RECT 2497.945 23.545 2498.115 25.075 ;
        RECT 2545.785 23.545 2545.955 25.075 ;
        RECT 2594.545 23.545 2594.715 25.075 ;
        RECT 2642.385 23.545 2642.555 25.075 ;
      LAYER mcon ;
        RECT 2448.265 240.805 2448.435 240.975 ;
        RECT 2497.945 24.905 2498.115 25.075 ;
        RECT 2545.785 24.905 2545.955 25.075 ;
        RECT 2594.545 24.905 2594.715 25.075 ;
        RECT 2642.385 24.905 2642.555 25.075 ;
      LAYER met1 ;
        RECT 2444.970 241.640 2445.290 241.700 ;
        RECT 2448.190 241.640 2448.510 241.700 ;
        RECT 2444.970 241.500 2448.510 241.640 ;
        RECT 2444.970 241.440 2445.290 241.500 ;
        RECT 2448.190 241.440 2448.510 241.500 ;
        RECT 2448.190 240.960 2448.510 241.020 ;
        RECT 2447.995 240.820 2448.510 240.960 ;
        RECT 2448.190 240.760 2448.510 240.820 ;
        RECT 2448.205 193.360 2448.495 193.405 ;
        RECT 2449.110 193.360 2449.430 193.420 ;
        RECT 2448.205 193.220 2449.430 193.360 ;
        RECT 2448.205 193.175 2448.495 193.220 ;
        RECT 2449.110 193.160 2449.430 193.220 ;
        RECT 2448.190 158.680 2448.510 158.740 ;
        RECT 2449.110 158.680 2449.430 158.740 ;
        RECT 2448.190 158.540 2449.430 158.680 ;
        RECT 2448.190 158.480 2448.510 158.540 ;
        RECT 2449.110 158.480 2449.430 158.540 ;
        RECT 2702.570 25.740 2702.890 25.800 ;
        RECT 2666.780 25.600 2702.890 25.740 ;
        RECT 2448.190 25.060 2448.510 25.120 ;
        RECT 2497.885 25.060 2498.175 25.105 ;
        RECT 2448.190 24.920 2498.175 25.060 ;
        RECT 2448.190 24.860 2448.510 24.920 ;
        RECT 2497.885 24.875 2498.175 24.920 ;
        RECT 2545.725 25.060 2546.015 25.105 ;
        RECT 2594.485 25.060 2594.775 25.105 ;
        RECT 2545.725 24.920 2594.775 25.060 ;
        RECT 2545.725 24.875 2546.015 24.920 ;
        RECT 2594.485 24.875 2594.775 24.920 ;
        RECT 2642.325 25.060 2642.615 25.105 ;
        RECT 2666.780 25.060 2666.920 25.600 ;
        RECT 2702.570 25.540 2702.890 25.600 ;
        RECT 2642.325 24.920 2666.920 25.060 ;
        RECT 2642.325 24.875 2642.615 24.920 ;
        RECT 2497.885 23.700 2498.175 23.745 ;
        RECT 2545.725 23.700 2546.015 23.745 ;
        RECT 2497.885 23.560 2546.015 23.700 ;
        RECT 2497.885 23.515 2498.175 23.560 ;
        RECT 2545.725 23.515 2546.015 23.560 ;
        RECT 2594.485 23.700 2594.775 23.745 ;
        RECT 2642.325 23.700 2642.615 23.745 ;
        RECT 2594.485 23.560 2642.615 23.700 ;
        RECT 2594.485 23.515 2594.775 23.560 ;
        RECT 2642.325 23.515 2642.615 23.560 ;
      LAYER via ;
        RECT 2445.000 241.440 2445.260 241.700 ;
        RECT 2448.220 241.440 2448.480 241.700 ;
        RECT 2448.220 240.760 2448.480 241.020 ;
        RECT 2449.140 193.160 2449.400 193.420 ;
        RECT 2448.220 158.480 2448.480 158.740 ;
        RECT 2449.140 158.480 2449.400 158.740 ;
        RECT 2448.220 24.860 2448.480 25.120 ;
        RECT 2702.600 25.540 2702.860 25.800 ;
      LAYER met2 ;
        RECT 2443.110 260.170 2443.390 264.000 ;
        RECT 2443.110 260.030 2445.200 260.170 ;
        RECT 2443.110 260.000 2443.390 260.030 ;
        RECT 2445.060 241.730 2445.200 260.030 ;
        RECT 2445.000 241.410 2445.260 241.730 ;
        RECT 2448.220 241.410 2448.480 241.730 ;
        RECT 2448.280 241.050 2448.420 241.410 ;
        RECT 2448.220 240.730 2448.480 241.050 ;
        RECT 2449.140 193.130 2449.400 193.450 ;
        RECT 2449.200 158.770 2449.340 193.130 ;
        RECT 2448.220 158.450 2448.480 158.770 ;
        RECT 2449.140 158.450 2449.400 158.770 ;
        RECT 2448.280 134.370 2448.420 158.450 ;
        RECT 2448.280 134.230 2448.880 134.370 ;
        RECT 2448.740 62.290 2448.880 134.230 ;
        RECT 2448.280 62.150 2448.880 62.290 ;
        RECT 2448.280 25.150 2448.420 62.150 ;
        RECT 2702.600 25.510 2702.860 25.830 ;
        RECT 2448.220 24.830 2448.480 25.150 ;
        RECT 2702.660 2.400 2702.800 25.510 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2457.390 242.660 2457.710 242.720 ;
        RECT 2462.910 242.660 2463.230 242.720 ;
        RECT 2457.390 242.520 2463.230 242.660 ;
        RECT 2457.390 242.460 2457.710 242.520 ;
        RECT 2462.910 242.460 2463.230 242.520 ;
        RECT 2462.910 24.380 2463.230 24.440 ;
        RECT 2720.510 24.380 2720.830 24.440 ;
        RECT 2462.910 24.240 2720.830 24.380 ;
        RECT 2462.910 24.180 2463.230 24.240 ;
        RECT 2720.510 24.180 2720.830 24.240 ;
      LAYER via ;
        RECT 2457.420 242.460 2457.680 242.720 ;
        RECT 2462.940 242.460 2463.200 242.720 ;
        RECT 2462.940 24.180 2463.200 24.440 ;
        RECT 2720.540 24.180 2720.800 24.440 ;
      LAYER met2 ;
        RECT 2457.370 260.000 2457.650 264.000 ;
        RECT 2457.480 242.750 2457.620 260.000 ;
        RECT 2457.420 242.430 2457.680 242.750 ;
        RECT 2462.940 242.430 2463.200 242.750 ;
        RECT 2463.000 24.470 2463.140 242.430 ;
        RECT 2462.940 24.150 2463.200 24.470 ;
        RECT 2720.540 24.150 2720.800 24.470 ;
        RECT 2720.600 2.400 2720.740 24.150 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2471.190 241.640 2471.510 241.700 ;
        RECT 2475.330 241.640 2475.650 241.700 ;
        RECT 2471.190 241.500 2475.650 241.640 ;
        RECT 2471.190 241.440 2471.510 241.500 ;
        RECT 2475.330 241.440 2475.650 241.500 ;
        RECT 2475.330 158.680 2475.650 158.740 ;
        RECT 2476.250 158.680 2476.570 158.740 ;
        RECT 2475.330 158.540 2476.570 158.680 ;
        RECT 2475.330 158.480 2475.650 158.540 ;
        RECT 2476.250 158.480 2476.570 158.540 ;
        RECT 2476.250 110.540 2476.570 110.800 ;
        RECT 2476.340 110.120 2476.480 110.540 ;
        RECT 2476.250 109.860 2476.570 110.120 ;
        RECT 2475.790 24.040 2476.110 24.100 ;
        RECT 2738.450 24.040 2738.770 24.100 ;
        RECT 2475.790 23.900 2738.770 24.040 ;
        RECT 2475.790 23.840 2476.110 23.900 ;
        RECT 2738.450 23.840 2738.770 23.900 ;
      LAYER via ;
        RECT 2471.220 241.440 2471.480 241.700 ;
        RECT 2475.360 241.440 2475.620 241.700 ;
        RECT 2475.360 158.480 2475.620 158.740 ;
        RECT 2476.280 158.480 2476.540 158.740 ;
        RECT 2476.280 110.540 2476.540 110.800 ;
        RECT 2476.280 109.860 2476.540 110.120 ;
        RECT 2475.820 23.840 2476.080 24.100 ;
        RECT 2738.480 23.840 2738.740 24.100 ;
      LAYER met2 ;
        RECT 2471.170 260.000 2471.450 264.000 ;
        RECT 2471.280 241.730 2471.420 260.000 ;
        RECT 2471.220 241.410 2471.480 241.730 ;
        RECT 2475.360 241.410 2475.620 241.730 ;
        RECT 2475.420 241.130 2475.560 241.410 ;
        RECT 2474.960 240.990 2475.560 241.130 ;
        RECT 2474.960 206.450 2475.100 240.990 ;
        RECT 2474.960 206.310 2475.560 206.450 ;
        RECT 2475.420 158.770 2475.560 206.310 ;
        RECT 2475.360 158.450 2475.620 158.770 ;
        RECT 2476.280 158.450 2476.540 158.770 ;
        RECT 2476.340 110.830 2476.480 158.450 ;
        RECT 2476.280 110.510 2476.540 110.830 ;
        RECT 2476.280 109.830 2476.540 110.150 ;
        RECT 2476.340 62.290 2476.480 109.830 ;
        RECT 2475.880 62.150 2476.480 62.290 ;
        RECT 2475.880 24.130 2476.020 62.150 ;
        RECT 2475.820 23.810 2476.080 24.130 ;
        RECT 2738.480 23.810 2738.740 24.130 ;
        RECT 2738.540 2.400 2738.680 23.810 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2485.450 237.900 2485.770 237.960 ;
        RECT 2753.170 237.900 2753.490 237.960 ;
        RECT 2485.450 237.760 2753.490 237.900 ;
        RECT 2485.450 237.700 2485.770 237.760 ;
        RECT 2753.170 237.700 2753.490 237.760 ;
      LAYER via ;
        RECT 2485.480 237.700 2485.740 237.960 ;
        RECT 2753.200 237.700 2753.460 237.960 ;
      LAYER met2 ;
        RECT 2485.430 260.000 2485.710 264.000 ;
        RECT 2485.540 237.990 2485.680 260.000 ;
        RECT 2485.480 237.670 2485.740 237.990 ;
        RECT 2753.200 237.670 2753.460 237.990 ;
        RECT 2753.260 17.410 2753.400 237.670 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 829.450 30.840 829.770 30.900 ;
        RECT 959.630 30.840 959.950 30.900 ;
        RECT 829.450 30.700 959.950 30.840 ;
        RECT 829.450 30.640 829.770 30.700 ;
        RECT 959.630 30.640 959.950 30.700 ;
      LAYER via ;
        RECT 829.480 30.640 829.740 30.900 ;
        RECT 959.660 30.640 959.920 30.900 ;
      LAYER met2 ;
        RECT 964.670 260.170 964.950 264.000 ;
        RECT 963.400 260.030 964.950 260.170 ;
        RECT 963.400 230.250 963.540 260.030 ;
        RECT 964.670 260.000 964.950 260.030 ;
        RECT 960.180 230.110 963.540 230.250 ;
        RECT 960.180 110.570 960.320 230.110 ;
        RECT 959.720 110.430 960.320 110.570 ;
        RECT 959.720 30.930 959.860 110.430 ;
        RECT 829.480 30.610 829.740 30.930 ;
        RECT 959.660 30.610 959.920 30.930 ;
        RECT 829.540 2.400 829.680 30.610 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2499.710 231.100 2500.030 231.160 ;
        RECT 2773.870 231.100 2774.190 231.160 ;
        RECT 2499.710 230.960 2774.190 231.100 ;
        RECT 2499.710 230.900 2500.030 230.960 ;
        RECT 2773.870 230.900 2774.190 230.960 ;
      LAYER via ;
        RECT 2499.740 230.900 2500.000 231.160 ;
        RECT 2773.900 230.900 2774.160 231.160 ;
      LAYER met2 ;
        RECT 2499.690 260.000 2499.970 264.000 ;
        RECT 2499.800 231.190 2499.940 260.000 ;
        RECT 2499.740 230.870 2500.000 231.190 ;
        RECT 2773.900 230.870 2774.160 231.190 ;
        RECT 2773.960 2.400 2774.100 230.870 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2513.510 224.300 2513.830 224.360 ;
        RECT 2787.670 224.300 2787.990 224.360 ;
        RECT 2513.510 224.160 2787.990 224.300 ;
        RECT 2513.510 224.100 2513.830 224.160 ;
        RECT 2787.670 224.100 2787.990 224.160 ;
      LAYER via ;
        RECT 2513.540 224.100 2513.800 224.360 ;
        RECT 2787.700 224.100 2787.960 224.360 ;
      LAYER met2 ;
        RECT 2513.490 260.000 2513.770 264.000 ;
        RECT 2513.600 224.390 2513.740 260.000 ;
        RECT 2513.540 224.070 2513.800 224.390 ;
        RECT 2787.700 224.070 2787.960 224.390 ;
        RECT 2787.760 17.410 2787.900 224.070 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2527.770 241.640 2528.090 241.700 ;
        RECT 2531.910 241.640 2532.230 241.700 ;
        RECT 2527.770 241.500 2532.230 241.640 ;
        RECT 2527.770 241.440 2528.090 241.500 ;
        RECT 2531.910 241.440 2532.230 241.500 ;
        RECT 2531.910 30.840 2532.230 30.900 ;
        RECT 2809.750 30.840 2810.070 30.900 ;
        RECT 2531.910 30.700 2810.070 30.840 ;
        RECT 2531.910 30.640 2532.230 30.700 ;
        RECT 2809.750 30.640 2810.070 30.700 ;
      LAYER via ;
        RECT 2527.800 241.440 2528.060 241.700 ;
        RECT 2531.940 241.440 2532.200 241.700 ;
        RECT 2531.940 30.640 2532.200 30.900 ;
        RECT 2809.780 30.640 2810.040 30.900 ;
      LAYER met2 ;
        RECT 2527.750 260.000 2528.030 264.000 ;
        RECT 2527.860 241.730 2528.000 260.000 ;
        RECT 2527.800 241.410 2528.060 241.730 ;
        RECT 2531.940 241.410 2532.200 241.730 ;
        RECT 2532.000 30.930 2532.140 241.410 ;
        RECT 2531.940 30.610 2532.200 30.930 ;
        RECT 2809.780 30.610 2810.040 30.930 ;
        RECT 2809.840 2.400 2809.980 30.610 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2541.570 241.640 2541.890 241.700 ;
        RECT 2545.710 241.640 2546.030 241.700 ;
        RECT 2541.570 241.500 2546.030 241.640 ;
        RECT 2541.570 241.440 2541.890 241.500 ;
        RECT 2545.710 241.440 2546.030 241.500 ;
        RECT 2545.710 217.160 2546.030 217.220 ;
        RECT 2822.170 217.160 2822.490 217.220 ;
        RECT 2545.710 217.020 2822.490 217.160 ;
        RECT 2545.710 216.960 2546.030 217.020 ;
        RECT 2822.170 216.960 2822.490 217.020 ;
      LAYER via ;
        RECT 2541.600 241.440 2541.860 241.700 ;
        RECT 2545.740 241.440 2546.000 241.700 ;
        RECT 2545.740 216.960 2546.000 217.220 ;
        RECT 2822.200 216.960 2822.460 217.220 ;
      LAYER met2 ;
        RECT 2541.550 260.000 2541.830 264.000 ;
        RECT 2541.660 241.730 2541.800 260.000 ;
        RECT 2541.600 241.410 2541.860 241.730 ;
        RECT 2545.740 241.410 2546.000 241.730 ;
        RECT 2545.800 217.250 2545.940 241.410 ;
        RECT 2545.740 216.930 2546.000 217.250 ;
        RECT 2822.200 216.930 2822.460 217.250 ;
        RECT 2822.260 17.410 2822.400 216.930 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2555.830 244.020 2556.150 244.080 ;
        RECT 2559.510 244.020 2559.830 244.080 ;
        RECT 2555.830 243.880 2559.830 244.020 ;
        RECT 2555.830 243.820 2556.150 243.880 ;
        RECT 2559.510 243.820 2559.830 243.880 ;
        RECT 2559.510 210.360 2559.830 210.420 ;
        RECT 2842.870 210.360 2843.190 210.420 ;
        RECT 2559.510 210.220 2843.190 210.360 ;
        RECT 2559.510 210.160 2559.830 210.220 ;
        RECT 2842.870 210.160 2843.190 210.220 ;
      LAYER via ;
        RECT 2555.860 243.820 2556.120 244.080 ;
        RECT 2559.540 243.820 2559.800 244.080 ;
        RECT 2559.540 210.160 2559.800 210.420 ;
        RECT 2842.900 210.160 2843.160 210.420 ;
      LAYER met2 ;
        RECT 2555.810 260.000 2556.090 264.000 ;
        RECT 2555.920 244.110 2556.060 260.000 ;
        RECT 2555.860 243.790 2556.120 244.110 ;
        RECT 2559.540 243.790 2559.800 244.110 ;
        RECT 2559.600 210.450 2559.740 243.790 ;
        RECT 2559.540 210.130 2559.800 210.450 ;
        RECT 2842.900 210.130 2843.160 210.450 ;
        RECT 2842.960 17.410 2843.100 210.130 ;
        RECT 2842.960 17.270 2845.400 17.410 ;
        RECT 2845.260 2.400 2845.400 17.270 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 44.780 2573.630 44.840 ;
        RECT 2863.110 44.780 2863.430 44.840 ;
        RECT 2573.310 44.640 2863.430 44.780 ;
        RECT 2573.310 44.580 2573.630 44.640 ;
        RECT 2863.110 44.580 2863.430 44.640 ;
      LAYER via ;
        RECT 2573.340 44.580 2573.600 44.840 ;
        RECT 2863.140 44.580 2863.400 44.840 ;
      LAYER met2 ;
        RECT 2570.070 260.170 2570.350 264.000 ;
        RECT 2570.070 260.030 2573.540 260.170 ;
        RECT 2570.070 260.000 2570.350 260.030 ;
        RECT 2573.400 44.870 2573.540 260.030 ;
        RECT 2573.340 44.550 2573.600 44.870 ;
        RECT 2863.140 44.550 2863.400 44.870 ;
        RECT 2863.200 2.400 2863.340 44.550 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2587.110 58.720 2587.430 58.780 ;
        RECT 2873.690 58.720 2874.010 58.780 ;
        RECT 2587.110 58.580 2874.010 58.720 ;
        RECT 2587.110 58.520 2587.430 58.580 ;
        RECT 2873.690 58.520 2874.010 58.580 ;
        RECT 2873.690 17.580 2874.010 17.640 ;
        RECT 2881.050 17.580 2881.370 17.640 ;
        RECT 2873.690 17.440 2881.370 17.580 ;
        RECT 2873.690 17.380 2874.010 17.440 ;
        RECT 2881.050 17.380 2881.370 17.440 ;
      LAYER via ;
        RECT 2587.140 58.520 2587.400 58.780 ;
        RECT 2873.720 58.520 2873.980 58.780 ;
        RECT 2873.720 17.380 2873.980 17.640 ;
        RECT 2881.080 17.380 2881.340 17.640 ;
      LAYER met2 ;
        RECT 2583.870 260.170 2584.150 264.000 ;
        RECT 2583.870 260.030 2587.340 260.170 ;
        RECT 2583.870 260.000 2584.150 260.030 ;
        RECT 2587.200 58.810 2587.340 260.030 ;
        RECT 2587.140 58.490 2587.400 58.810 ;
        RECT 2873.720 58.490 2873.980 58.810 ;
        RECT 2873.780 17.670 2873.920 58.490 ;
        RECT 2873.720 17.350 2873.980 17.670 ;
        RECT 2881.080 17.350 2881.340 17.670 ;
        RECT 2881.140 2.400 2881.280 17.350 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2600.910 51.580 2601.230 51.640 ;
        RECT 2898.070 51.580 2898.390 51.640 ;
        RECT 2600.910 51.440 2898.390 51.580 ;
        RECT 2600.910 51.380 2601.230 51.440 ;
        RECT 2898.070 51.380 2898.390 51.440 ;
        RECT 2898.070 2.960 2898.390 3.020 ;
        RECT 2898.990 2.960 2899.310 3.020 ;
        RECT 2898.070 2.820 2899.310 2.960 ;
        RECT 2898.070 2.760 2898.390 2.820 ;
        RECT 2898.990 2.760 2899.310 2.820 ;
      LAYER via ;
        RECT 2600.940 51.380 2601.200 51.640 ;
        RECT 2898.100 51.380 2898.360 51.640 ;
        RECT 2898.100 2.760 2898.360 3.020 ;
        RECT 2899.020 2.760 2899.280 3.020 ;
      LAYER met2 ;
        RECT 2598.130 260.170 2598.410 264.000 ;
        RECT 2598.130 260.030 2601.140 260.170 ;
        RECT 2598.130 260.000 2598.410 260.030 ;
        RECT 2601.000 51.670 2601.140 260.030 ;
        RECT 2600.940 51.350 2601.200 51.670 ;
        RECT 2898.100 51.350 2898.360 51.670 ;
        RECT 2898.160 3.050 2898.300 51.350 ;
        RECT 2898.100 2.730 2898.360 3.050 ;
        RECT 2899.020 2.730 2899.280 3.050 ;
        RECT 2899.080 2.400 2899.220 2.730 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 973.890 207.300 974.210 207.360 ;
        RECT 977.110 207.300 977.430 207.360 ;
        RECT 973.890 207.160 977.430 207.300 ;
        RECT 973.890 207.100 974.210 207.160 ;
        RECT 977.110 207.100 977.430 207.160 ;
        RECT 846.930 37.980 847.250 38.040 ;
        RECT 973.430 37.980 973.750 38.040 ;
        RECT 846.930 37.840 973.750 37.980 ;
        RECT 846.930 37.780 847.250 37.840 ;
        RECT 973.430 37.780 973.750 37.840 ;
      LAYER via ;
        RECT 973.920 207.100 974.180 207.360 ;
        RECT 977.140 207.100 977.400 207.360 ;
        RECT 846.960 37.780 847.220 38.040 ;
        RECT 973.460 37.780 973.720 38.040 ;
      LAYER met2 ;
        RECT 978.470 260.170 978.750 264.000 ;
        RECT 977.200 260.030 978.750 260.170 ;
        RECT 977.200 207.390 977.340 260.030 ;
        RECT 978.470 260.000 978.750 260.030 ;
        RECT 973.920 207.070 974.180 207.390 ;
        RECT 977.140 207.070 977.400 207.390 ;
        RECT 973.980 110.570 974.120 207.070 ;
        RECT 973.520 110.430 974.120 110.570 ;
        RECT 973.520 38.070 973.660 110.430 ;
        RECT 846.960 37.750 847.220 38.070 ;
        RECT 973.460 37.750 973.720 38.070 ;
        RECT 847.020 2.400 847.160 37.750 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 987.305 157.845 987.475 193.035 ;
      LAYER mcon ;
        RECT 987.305 192.865 987.475 193.035 ;
      LAYER met1 ;
        RECT 987.230 193.020 987.550 193.080 ;
        RECT 987.035 192.880 987.550 193.020 ;
        RECT 987.230 192.820 987.550 192.880 ;
        RECT 987.230 158.000 987.550 158.060 ;
        RECT 987.035 157.860 987.550 158.000 ;
        RECT 987.230 157.800 987.550 157.860 ;
        RECT 864.870 44.780 865.190 44.840 ;
        RECT 987.230 44.780 987.550 44.840 ;
        RECT 864.870 44.640 987.550 44.780 ;
        RECT 864.870 44.580 865.190 44.640 ;
        RECT 987.230 44.580 987.550 44.640 ;
      LAYER via ;
        RECT 987.260 192.820 987.520 193.080 ;
        RECT 987.260 157.800 987.520 158.060 ;
        RECT 864.900 44.580 865.160 44.840 ;
        RECT 987.260 44.580 987.520 44.840 ;
      LAYER met2 ;
        RECT 992.730 260.850 993.010 264.000 ;
        RECT 989.620 260.710 993.010 260.850 ;
        RECT 989.620 256.090 989.760 260.710 ;
        RECT 992.730 260.000 993.010 260.710 ;
        RECT 989.160 255.950 989.760 256.090 ;
        RECT 989.160 207.810 989.300 255.950 ;
        RECT 987.780 207.670 989.300 207.810 ;
        RECT 987.780 207.130 987.920 207.670 ;
        RECT 987.320 206.990 987.920 207.130 ;
        RECT 987.320 193.110 987.460 206.990 ;
        RECT 987.260 192.790 987.520 193.110 ;
        RECT 987.260 157.770 987.520 158.090 ;
        RECT 987.320 44.870 987.460 157.770 ;
        RECT 864.900 44.550 865.160 44.870 ;
        RECT 987.260 44.550 987.520 44.870 ;
        RECT 864.960 2.400 865.100 44.550 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1002.485 157.845 1002.655 210.375 ;
      LAYER mcon ;
        RECT 1002.485 210.205 1002.655 210.375 ;
      LAYER met1 ;
        RECT 1002.425 210.360 1002.715 210.405 ;
        RECT 1005.630 210.360 1005.950 210.420 ;
        RECT 1002.425 210.220 1005.950 210.360 ;
        RECT 1002.425 210.175 1002.715 210.220 ;
        RECT 1005.630 210.160 1005.950 210.220 ;
        RECT 1002.410 158.000 1002.730 158.060 ;
        RECT 1002.215 157.860 1002.730 158.000 ;
        RECT 1002.410 157.800 1002.730 157.860 ;
        RECT 1001.490 120.940 1001.810 121.000 ;
        RECT 1002.410 120.940 1002.730 121.000 ;
        RECT 1001.490 120.800 1002.730 120.940 ;
        RECT 1001.490 120.740 1001.810 120.800 ;
        RECT 1002.410 120.740 1002.730 120.800 ;
        RECT 882.810 51.580 883.130 51.640 ;
        RECT 1001.950 51.580 1002.270 51.640 ;
        RECT 882.810 51.440 1002.270 51.580 ;
        RECT 882.810 51.380 883.130 51.440 ;
        RECT 1001.950 51.380 1002.270 51.440 ;
      LAYER via ;
        RECT 1005.660 210.160 1005.920 210.420 ;
        RECT 1002.440 157.800 1002.700 158.060 ;
        RECT 1001.520 120.740 1001.780 121.000 ;
        RECT 1002.440 120.740 1002.700 121.000 ;
        RECT 882.840 51.380 883.100 51.640 ;
        RECT 1001.980 51.380 1002.240 51.640 ;
      LAYER met2 ;
        RECT 1006.990 260.170 1007.270 264.000 ;
        RECT 1005.720 260.030 1007.270 260.170 ;
        RECT 1005.720 210.450 1005.860 260.030 ;
        RECT 1006.990 260.000 1007.270 260.030 ;
        RECT 1005.660 210.130 1005.920 210.450 ;
        RECT 1002.440 157.770 1002.700 158.090 ;
        RECT 1002.500 121.030 1002.640 157.770 ;
        RECT 1001.520 120.710 1001.780 121.030 ;
        RECT 1002.440 120.710 1002.700 121.030 ;
        RECT 1001.580 62.290 1001.720 120.710 ;
        RECT 1001.580 62.150 1002.180 62.290 ;
        RECT 1002.040 51.670 1002.180 62.150 ;
        RECT 882.840 51.350 883.100 51.670 ;
        RECT 1001.980 51.350 1002.240 51.670 ;
        RECT 882.900 2.400 883.040 51.350 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1015.825 144.925 1015.995 193.035 ;
        RECT 1015.825 58.565 1015.995 96.475 ;
      LAYER mcon ;
        RECT 1015.825 192.865 1015.995 193.035 ;
        RECT 1015.825 96.305 1015.995 96.475 ;
      LAYER met1 ;
        RECT 1015.765 193.020 1016.055 193.065 ;
        RECT 1016.210 193.020 1016.530 193.080 ;
        RECT 1015.765 192.880 1016.530 193.020 ;
        RECT 1015.765 192.835 1016.055 192.880 ;
        RECT 1016.210 192.820 1016.530 192.880 ;
        RECT 1015.750 145.080 1016.070 145.140 ;
        RECT 1015.555 144.940 1016.070 145.080 ;
        RECT 1015.750 144.880 1016.070 144.940 ;
        RECT 1014.830 110.400 1015.150 110.460 ;
        RECT 1015.750 110.400 1016.070 110.460 ;
        RECT 1014.830 110.260 1016.070 110.400 ;
        RECT 1014.830 110.200 1015.150 110.260 ;
        RECT 1015.750 110.200 1016.070 110.260 ;
        RECT 1015.750 96.460 1016.070 96.520 ;
        RECT 1015.555 96.320 1016.070 96.460 ;
        RECT 1015.750 96.260 1016.070 96.320 ;
        RECT 903.510 58.720 903.830 58.780 ;
        RECT 1015.765 58.720 1016.055 58.765 ;
        RECT 903.510 58.580 1016.055 58.720 ;
        RECT 903.510 58.520 903.830 58.580 ;
        RECT 1015.765 58.535 1016.055 58.580 ;
        RECT 900.750 18.260 901.070 18.320 ;
        RECT 903.510 18.260 903.830 18.320 ;
        RECT 900.750 18.120 903.830 18.260 ;
        RECT 900.750 18.060 901.070 18.120 ;
        RECT 903.510 18.060 903.830 18.120 ;
      LAYER via ;
        RECT 1016.240 192.820 1016.500 193.080 ;
        RECT 1015.780 144.880 1016.040 145.140 ;
        RECT 1014.860 110.200 1015.120 110.460 ;
        RECT 1015.780 110.200 1016.040 110.460 ;
        RECT 1015.780 96.260 1016.040 96.520 ;
        RECT 903.540 58.520 903.800 58.780 ;
        RECT 900.780 18.060 901.040 18.320 ;
        RECT 903.540 18.060 903.800 18.320 ;
      LAYER met2 ;
        RECT 1020.790 260.170 1021.070 264.000 ;
        RECT 1019.520 260.030 1021.070 260.170 ;
        RECT 1019.520 194.325 1019.660 260.030 ;
        RECT 1020.790 260.000 1021.070 260.030 ;
        RECT 1019.450 193.955 1019.730 194.325 ;
        RECT 1015.770 193.530 1016.050 193.645 ;
        RECT 1015.770 193.390 1016.440 193.530 ;
        RECT 1015.770 193.275 1016.050 193.390 ;
        RECT 1016.300 193.110 1016.440 193.390 ;
        RECT 1016.240 192.790 1016.500 193.110 ;
        RECT 1015.780 144.850 1016.040 145.170 ;
        RECT 1015.840 110.570 1015.980 144.850 ;
        RECT 1014.920 110.490 1015.980 110.570 ;
        RECT 1014.860 110.430 1016.040 110.490 ;
        RECT 1014.860 110.170 1015.120 110.430 ;
        RECT 1015.780 110.170 1016.040 110.430 ;
        RECT 1015.840 96.550 1015.980 110.170 ;
        RECT 1015.780 96.230 1016.040 96.550 ;
        RECT 903.540 58.490 903.800 58.810 ;
        RECT 903.600 18.350 903.740 58.490 ;
        RECT 900.780 18.030 901.040 18.350 ;
        RECT 903.540 18.030 903.800 18.350 ;
        RECT 900.840 2.400 900.980 18.030 ;
        RECT 900.630 -4.800 901.190 2.400 ;
      LAYER via2 ;
        RECT 1019.450 194.000 1019.730 194.280 ;
        RECT 1015.770 193.320 1016.050 193.600 ;
      LAYER met3 ;
        RECT 1019.425 194.290 1019.755 194.305 ;
        RECT 1015.070 193.990 1019.755 194.290 ;
        RECT 1015.070 193.610 1015.370 193.990 ;
        RECT 1019.425 193.975 1019.755 193.990 ;
        RECT 1015.745 193.610 1016.075 193.625 ;
        RECT 1015.070 193.310 1016.075 193.610 ;
        RECT 1015.745 193.295 1016.075 193.310 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1024.490 243.680 1024.810 243.740 ;
        RECT 1035.070 243.680 1035.390 243.740 ;
        RECT 1024.490 243.540 1035.390 243.680 ;
        RECT 1024.490 243.480 1024.810 243.540 ;
        RECT 1035.070 243.480 1035.390 243.540 ;
        RECT 918.690 24.380 919.010 24.440 ;
        RECT 1024.490 24.380 1024.810 24.440 ;
        RECT 918.690 24.240 1024.810 24.380 ;
        RECT 918.690 24.180 919.010 24.240 ;
        RECT 1024.490 24.180 1024.810 24.240 ;
      LAYER via ;
        RECT 1024.520 243.480 1024.780 243.740 ;
        RECT 1035.100 243.480 1035.360 243.740 ;
        RECT 918.720 24.180 918.980 24.440 ;
        RECT 1024.520 24.180 1024.780 24.440 ;
      LAYER met2 ;
        RECT 1035.050 260.000 1035.330 264.000 ;
        RECT 1035.160 243.770 1035.300 260.000 ;
        RECT 1024.520 243.450 1024.780 243.770 ;
        RECT 1035.100 243.450 1035.360 243.770 ;
        RECT 1024.580 24.470 1024.720 243.450 ;
        RECT 918.720 24.150 918.980 24.470 ;
        RECT 1024.520 24.150 1024.780 24.470 ;
        RECT 918.780 2.400 918.920 24.150 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1045.190 248.440 1045.510 248.500 ;
        RECT 1049.330 248.440 1049.650 248.500 ;
        RECT 1045.190 248.300 1049.650 248.440 ;
        RECT 1045.190 248.240 1045.510 248.300 ;
        RECT 1049.330 248.240 1049.650 248.300 ;
        RECT 938.010 65.520 938.330 65.580 ;
        RECT 1045.190 65.520 1045.510 65.580 ;
        RECT 938.010 65.380 1045.510 65.520 ;
        RECT 938.010 65.320 938.330 65.380 ;
        RECT 1045.190 65.320 1045.510 65.380 ;
        RECT 936.170 2.960 936.490 3.020 ;
        RECT 938.010 2.960 938.330 3.020 ;
        RECT 936.170 2.820 938.330 2.960 ;
        RECT 936.170 2.760 936.490 2.820 ;
        RECT 938.010 2.760 938.330 2.820 ;
      LAYER via ;
        RECT 1045.220 248.240 1045.480 248.500 ;
        RECT 1049.360 248.240 1049.620 248.500 ;
        RECT 938.040 65.320 938.300 65.580 ;
        RECT 1045.220 65.320 1045.480 65.580 ;
        RECT 936.200 2.760 936.460 3.020 ;
        RECT 938.040 2.760 938.300 3.020 ;
      LAYER met2 ;
        RECT 1049.310 260.000 1049.590 264.000 ;
        RECT 1049.420 248.530 1049.560 260.000 ;
        RECT 1045.220 248.210 1045.480 248.530 ;
        RECT 1049.360 248.210 1049.620 248.530 ;
        RECT 1045.280 65.610 1045.420 248.210 ;
        RECT 938.040 65.290 938.300 65.610 ;
        RECT 1045.220 65.290 1045.480 65.610 ;
        RECT 938.100 3.050 938.240 65.290 ;
        RECT 936.200 2.730 936.460 3.050 ;
        RECT 938.040 2.730 938.300 3.050 ;
        RECT 936.260 2.400 936.400 2.730 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.110 260.000 1063.390 264.000 ;
        RECT 1063.220 16.845 1063.360 260.000 ;
        RECT 954.130 16.475 954.410 16.845 ;
        RECT 1063.150 16.475 1063.430 16.845 ;
        RECT 954.200 2.400 954.340 16.475 ;
        RECT 953.990 -4.800 954.550 2.400 ;
      LAYER via2 ;
        RECT 954.130 16.520 954.410 16.800 ;
        RECT 1063.150 16.520 1063.430 16.800 ;
      LAYER met3 ;
        RECT 954.105 16.810 954.435 16.825 ;
        RECT 1063.125 16.810 1063.455 16.825 ;
        RECT 954.105 16.510 1063.455 16.810 ;
        RECT 954.105 16.495 954.435 16.510 ;
        RECT 1063.125 16.495 1063.455 16.510 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.370 260.170 1077.650 264.000 ;
        RECT 1077.020 260.030 1077.650 260.170 ;
        RECT 1077.020 17.525 1077.160 260.030 ;
        RECT 1077.370 260.000 1077.650 260.030 ;
        RECT 972.070 17.155 972.350 17.525 ;
        RECT 1076.950 17.155 1077.230 17.525 ;
        RECT 972.140 2.400 972.280 17.155 ;
        RECT 971.930 -4.800 972.490 2.400 ;
      LAYER via2 ;
        RECT 972.070 17.200 972.350 17.480 ;
        RECT 1076.950 17.200 1077.230 17.480 ;
      LAYER met3 ;
        RECT 972.045 17.490 972.375 17.505 ;
        RECT 1076.925 17.490 1077.255 17.505 ;
        RECT 972.045 17.190 1077.255 17.490 ;
        RECT 972.045 17.175 972.375 17.190 ;
        RECT 1076.925 17.175 1077.255 17.190 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 31.180 651.290 31.240 ;
        RECT 821.170 31.180 821.490 31.240 ;
        RECT 650.970 31.040 821.490 31.180 ;
        RECT 650.970 30.980 651.290 31.040 ;
        RECT 821.170 30.980 821.490 31.040 ;
      LAYER via ;
        RECT 651.000 30.980 651.260 31.240 ;
        RECT 821.200 30.980 821.460 31.240 ;
      LAYER met2 ;
        RECT 823.910 260.170 824.190 264.000 ;
        RECT 821.260 260.030 824.190 260.170 ;
        RECT 821.260 31.270 821.400 260.030 ;
        RECT 823.910 260.000 824.190 260.030 ;
        RECT 651.000 30.950 651.260 31.270 ;
        RECT 821.200 30.950 821.460 31.270 ;
        RECT 651.060 2.400 651.200 30.950 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1069.645 17.425 1069.815 19.635 ;
      LAYER mcon ;
        RECT 1069.645 19.465 1069.815 19.635 ;
      LAYER met1 ;
        RECT 1069.585 19.620 1069.875 19.665 ;
        RECT 1090.730 19.620 1091.050 19.680 ;
        RECT 1069.585 19.480 1091.050 19.620 ;
        RECT 1069.585 19.435 1069.875 19.480 ;
        RECT 1090.730 19.420 1091.050 19.480 ;
        RECT 989.990 17.580 990.310 17.640 ;
        RECT 1069.585 17.580 1069.875 17.625 ;
        RECT 989.990 17.440 1069.875 17.580 ;
        RECT 989.990 17.380 990.310 17.440 ;
        RECT 1069.585 17.395 1069.875 17.440 ;
      LAYER via ;
        RECT 1090.760 19.420 1091.020 19.680 ;
        RECT 990.020 17.380 990.280 17.640 ;
      LAYER met2 ;
        RECT 1091.170 260.170 1091.450 264.000 ;
        RECT 1090.820 260.030 1091.450 260.170 ;
        RECT 1090.820 19.710 1090.960 260.030 ;
        RECT 1091.170 260.000 1091.450 260.030 ;
        RECT 1090.760 19.390 1091.020 19.710 ;
        RECT 990.020 17.350 990.280 17.670 ;
        RECT 990.080 2.400 990.220 17.350 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1036.065 15.725 1036.235 20.655 ;
        RECT 1048.945 18.785 1049.115 20.655 ;
        RECT 1077.005 19.125 1077.175 19.975 ;
      LAYER mcon ;
        RECT 1036.065 20.485 1036.235 20.655 ;
        RECT 1048.945 20.485 1049.115 20.655 ;
        RECT 1077.005 19.805 1077.175 19.975 ;
      LAYER met1 ;
        RECT 1036.005 20.640 1036.295 20.685 ;
        RECT 1048.885 20.640 1049.175 20.685 ;
        RECT 1036.005 20.500 1049.175 20.640 ;
        RECT 1036.005 20.455 1036.295 20.500 ;
        RECT 1048.885 20.455 1049.175 20.500 ;
        RECT 1076.945 19.960 1077.235 20.005 ;
        RECT 1076.945 19.820 1091.420 19.960 ;
        RECT 1076.945 19.775 1077.235 19.820 ;
        RECT 1091.280 19.620 1091.420 19.820 ;
        RECT 1104.530 19.620 1104.850 19.680 ;
        RECT 1091.280 19.480 1104.850 19.620 ;
        RECT 1104.530 19.420 1104.850 19.480 ;
        RECT 1076.945 19.280 1077.235 19.325 ;
        RECT 1050.340 19.140 1077.235 19.280 ;
        RECT 1048.885 18.940 1049.175 18.985 ;
        RECT 1050.340 18.940 1050.480 19.140 ;
        RECT 1076.945 19.095 1077.235 19.140 ;
        RECT 1048.885 18.800 1050.480 18.940 ;
        RECT 1048.885 18.755 1049.175 18.800 ;
        RECT 1007.470 15.880 1007.790 15.940 ;
        RECT 1036.005 15.880 1036.295 15.925 ;
        RECT 1007.470 15.740 1036.295 15.880 ;
        RECT 1007.470 15.680 1007.790 15.740 ;
        RECT 1036.005 15.695 1036.295 15.740 ;
      LAYER via ;
        RECT 1104.560 19.420 1104.820 19.680 ;
        RECT 1007.500 15.680 1007.760 15.940 ;
      LAYER met2 ;
        RECT 1105.430 260.170 1105.710 264.000 ;
        RECT 1104.620 260.030 1105.710 260.170 ;
        RECT 1104.620 19.710 1104.760 260.030 ;
        RECT 1105.430 260.000 1105.710 260.030 ;
        RECT 1104.560 19.390 1104.820 19.710 ;
        RECT 1007.500 15.650 1007.760 15.970 ;
        RECT 1007.560 2.400 1007.700 15.650 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1042.505 15.385 1042.675 18.275 ;
      LAYER mcon ;
        RECT 1042.505 18.105 1042.675 18.275 ;
      LAYER met1 ;
        RECT 1118.790 18.600 1119.110 18.660 ;
        RECT 1106.000 18.460 1119.110 18.600 ;
        RECT 1042.445 18.260 1042.735 18.305 ;
        RECT 1106.000 18.260 1106.140 18.460 ;
        RECT 1118.790 18.400 1119.110 18.460 ;
        RECT 1042.445 18.120 1106.140 18.260 ;
        RECT 1042.445 18.075 1042.735 18.120 ;
        RECT 1025.410 15.540 1025.730 15.600 ;
        RECT 1042.445 15.540 1042.735 15.585 ;
        RECT 1025.410 15.400 1042.735 15.540 ;
        RECT 1025.410 15.340 1025.730 15.400 ;
        RECT 1042.445 15.355 1042.735 15.400 ;
      LAYER via ;
        RECT 1118.820 18.400 1119.080 18.660 ;
        RECT 1025.440 15.340 1025.700 15.600 ;
      LAYER met2 ;
        RECT 1119.690 260.170 1119.970 264.000 ;
        RECT 1118.880 260.030 1119.970 260.170 ;
        RECT 1118.880 18.690 1119.020 260.030 ;
        RECT 1119.690 260.000 1119.970 260.030 ;
        RECT 1118.820 18.370 1119.080 18.690 ;
        RECT 1025.440 15.310 1025.700 15.630 ;
        RECT 1025.500 2.400 1025.640 15.310 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1132.130 18.940 1132.450 19.000 ;
        RECT 1105.540 18.800 1132.450 18.940 ;
        RECT 1043.350 18.600 1043.670 18.660 ;
        RECT 1105.540 18.600 1105.680 18.800 ;
        RECT 1132.130 18.740 1132.450 18.800 ;
        RECT 1043.350 18.460 1105.680 18.600 ;
        RECT 1043.350 18.400 1043.670 18.460 ;
      LAYER via ;
        RECT 1043.380 18.400 1043.640 18.660 ;
        RECT 1132.160 18.740 1132.420 19.000 ;
      LAYER met2 ;
        RECT 1133.490 260.170 1133.770 264.000 ;
        RECT 1132.220 260.030 1133.770 260.170 ;
        RECT 1132.220 19.030 1132.360 260.030 ;
        RECT 1133.490 260.000 1133.770 260.030 ;
        RECT 1132.160 18.710 1132.420 19.030 ;
        RECT 1043.380 18.370 1043.640 18.690 ;
        RECT 1043.440 2.400 1043.580 18.370 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1061.290 17.240 1061.610 17.300 ;
        RECT 1145.470 17.240 1145.790 17.300 ;
        RECT 1061.290 17.100 1145.790 17.240 ;
        RECT 1061.290 17.040 1061.610 17.100 ;
        RECT 1145.470 17.040 1145.790 17.100 ;
      LAYER via ;
        RECT 1061.320 17.040 1061.580 17.300 ;
        RECT 1145.500 17.040 1145.760 17.300 ;
      LAYER met2 ;
        RECT 1147.750 260.170 1148.030 264.000 ;
        RECT 1145.560 260.030 1148.030 260.170 ;
        RECT 1145.560 17.330 1145.700 260.030 ;
        RECT 1147.750 260.000 1148.030 260.030 ;
        RECT 1061.320 17.010 1061.580 17.330 ;
        RECT 1145.500 17.010 1145.760 17.330 ;
        RECT 1061.380 2.400 1061.520 17.010 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.230 19.280 1079.550 19.340 ;
        RECT 1159.270 19.280 1159.590 19.340 ;
        RECT 1079.230 19.140 1159.590 19.280 ;
        RECT 1079.230 19.080 1079.550 19.140 ;
        RECT 1159.270 19.080 1159.590 19.140 ;
      LAYER via ;
        RECT 1079.260 19.080 1079.520 19.340 ;
        RECT 1159.300 19.080 1159.560 19.340 ;
      LAYER met2 ;
        RECT 1161.550 260.170 1161.830 264.000 ;
        RECT 1159.360 260.030 1161.830 260.170 ;
        RECT 1159.360 19.370 1159.500 260.030 ;
        RECT 1161.550 260.000 1161.830 260.030 ;
        RECT 1079.260 19.050 1079.520 19.370 ;
        RECT 1159.300 19.050 1159.560 19.370 ;
        RECT 1079.320 2.400 1079.460 19.050 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.070 17.920 1173.390 17.980 ;
        RECT 1156.140 17.780 1173.390 17.920 ;
        RECT 1096.710 17.580 1097.030 17.640 ;
        RECT 1156.140 17.580 1156.280 17.780 ;
        RECT 1173.070 17.720 1173.390 17.780 ;
        RECT 1096.710 17.440 1156.280 17.580 ;
        RECT 1096.710 17.380 1097.030 17.440 ;
      LAYER via ;
        RECT 1096.740 17.380 1097.000 17.640 ;
        RECT 1173.100 17.720 1173.360 17.980 ;
      LAYER met2 ;
        RECT 1175.810 260.170 1176.090 264.000 ;
        RECT 1173.160 260.030 1176.090 260.170 ;
        RECT 1173.160 18.010 1173.300 260.030 ;
        RECT 1175.810 260.000 1176.090 260.030 ;
        RECT 1173.100 17.690 1173.360 18.010 ;
        RECT 1096.740 17.350 1097.000 17.670 ;
        RECT 1096.800 2.400 1096.940 17.350 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1155.665 17.765 1155.835 18.615 ;
      LAYER mcon ;
        RECT 1155.665 18.445 1155.835 18.615 ;
      LAYER met1 ;
        RECT 1155.605 18.600 1155.895 18.645 ;
        RECT 1186.870 18.600 1187.190 18.660 ;
        RECT 1155.605 18.460 1187.190 18.600 ;
        RECT 1155.605 18.415 1155.895 18.460 ;
        RECT 1186.870 18.400 1187.190 18.460 ;
        RECT 1114.650 18.260 1114.970 18.320 ;
        RECT 1114.650 18.120 1131.900 18.260 ;
        RECT 1114.650 18.060 1114.970 18.120 ;
        RECT 1131.760 17.920 1131.900 18.120 ;
        RECT 1155.605 17.920 1155.895 17.965 ;
        RECT 1131.760 17.780 1155.895 17.920 ;
        RECT 1155.605 17.735 1155.895 17.780 ;
      LAYER via ;
        RECT 1186.900 18.400 1187.160 18.660 ;
        RECT 1114.680 18.060 1114.940 18.320 ;
      LAYER met2 ;
        RECT 1190.070 260.170 1190.350 264.000 ;
        RECT 1186.960 260.030 1190.350 260.170 ;
        RECT 1186.960 18.690 1187.100 260.030 ;
        RECT 1190.070 260.000 1190.350 260.030 ;
        RECT 1186.900 18.370 1187.160 18.690 ;
        RECT 1114.680 18.030 1114.940 18.350 ;
        RECT 1114.740 2.400 1114.880 18.030 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1145.545 18.445 1145.715 19.975 ;
      LAYER mcon ;
        RECT 1145.545 19.805 1145.715 19.975 ;
      LAYER met1 ;
        RECT 1145.485 19.960 1145.775 20.005 ;
        RECT 1200.670 19.960 1200.990 20.020 ;
        RECT 1145.485 19.820 1200.990 19.960 ;
        RECT 1145.485 19.775 1145.775 19.820 ;
        RECT 1200.670 19.760 1200.990 19.820 ;
        RECT 1132.590 18.600 1132.910 18.660 ;
        RECT 1145.485 18.600 1145.775 18.645 ;
        RECT 1132.590 18.460 1145.775 18.600 ;
        RECT 1132.590 18.400 1132.910 18.460 ;
        RECT 1145.485 18.415 1145.775 18.460 ;
      LAYER via ;
        RECT 1200.700 19.760 1200.960 20.020 ;
        RECT 1132.620 18.400 1132.880 18.660 ;
      LAYER met2 ;
        RECT 1203.870 260.170 1204.150 264.000 ;
        RECT 1200.760 260.030 1204.150 260.170 ;
        RECT 1200.760 20.050 1200.900 260.030 ;
        RECT 1203.870 260.000 1204.150 260.030 ;
        RECT 1200.700 19.730 1200.960 20.050 ;
        RECT 1132.620 18.370 1132.880 18.690 ;
        RECT 1132.680 2.400 1132.820 18.370 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1150.530 17.240 1150.850 17.300 ;
        RECT 1214.930 17.240 1215.250 17.300 ;
        RECT 1150.530 17.100 1215.250 17.240 ;
        RECT 1150.530 17.040 1150.850 17.100 ;
        RECT 1214.930 17.040 1215.250 17.100 ;
      LAYER via ;
        RECT 1150.560 17.040 1150.820 17.300 ;
        RECT 1214.960 17.040 1215.220 17.300 ;
      LAYER met2 ;
        RECT 1218.130 260.170 1218.410 264.000 ;
        RECT 1215.020 260.030 1218.410 260.170 ;
        RECT 1215.020 17.330 1215.160 260.030 ;
        RECT 1218.130 260.000 1218.410 260.030 ;
        RECT 1150.560 17.010 1150.820 17.330 ;
        RECT 1214.960 17.010 1215.220 17.330 ;
        RECT 1150.620 2.400 1150.760 17.010 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.450 38.320 668.770 38.380 ;
        RECT 834.970 38.320 835.290 38.380 ;
        RECT 668.450 38.180 835.290 38.320 ;
        RECT 668.450 38.120 668.770 38.180 ;
        RECT 834.970 38.120 835.290 38.180 ;
      LAYER via ;
        RECT 668.480 38.120 668.740 38.380 ;
        RECT 835.000 38.120 835.260 38.380 ;
      LAYER met2 ;
        RECT 837.710 260.170 837.990 264.000 ;
        RECT 835.060 260.030 837.990 260.170 ;
        RECT 835.060 38.410 835.200 260.030 ;
        RECT 837.710 260.000 837.990 260.030 ;
        RECT 668.480 38.090 668.740 38.410 ;
        RECT 835.000 38.090 835.260 38.410 ;
        RECT 668.540 7.890 668.680 38.090 ;
        RECT 668.540 7.750 669.140 7.890 ;
        RECT 669.000 2.400 669.140 7.750 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 246.740 1172.930 246.800 ;
        RECT 1232.410 246.740 1232.730 246.800 ;
        RECT 1172.610 246.600 1232.730 246.740 ;
        RECT 1172.610 246.540 1172.930 246.600 ;
        RECT 1232.410 246.540 1232.730 246.600 ;
        RECT 1168.470 17.580 1168.790 17.640 ;
        RECT 1172.610 17.580 1172.930 17.640 ;
        RECT 1168.470 17.440 1172.930 17.580 ;
        RECT 1168.470 17.380 1168.790 17.440 ;
        RECT 1172.610 17.380 1172.930 17.440 ;
      LAYER via ;
        RECT 1172.640 246.540 1172.900 246.800 ;
        RECT 1232.440 246.540 1232.700 246.800 ;
        RECT 1168.500 17.380 1168.760 17.640 ;
        RECT 1172.640 17.380 1172.900 17.640 ;
      LAYER met2 ;
        RECT 1232.390 260.000 1232.670 264.000 ;
        RECT 1232.500 246.830 1232.640 260.000 ;
        RECT 1172.640 246.510 1172.900 246.830 ;
        RECT 1232.440 246.510 1232.700 246.830 ;
        RECT 1172.700 17.670 1172.840 246.510 ;
        RECT 1168.500 17.350 1168.760 17.670 ;
        RECT 1172.640 17.350 1172.900 17.670 ;
        RECT 1168.560 2.400 1168.700 17.350 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 247.080 1186.730 247.140 ;
        RECT 1246.210 247.080 1246.530 247.140 ;
        RECT 1186.410 246.940 1246.530 247.080 ;
        RECT 1186.410 246.880 1186.730 246.940 ;
        RECT 1246.210 246.880 1246.530 246.940 ;
      LAYER via ;
        RECT 1186.440 246.880 1186.700 247.140 ;
        RECT 1246.240 246.880 1246.500 247.140 ;
      LAYER met2 ;
        RECT 1246.190 260.000 1246.470 264.000 ;
        RECT 1246.300 247.170 1246.440 260.000 ;
        RECT 1186.440 246.850 1186.700 247.170 ;
        RECT 1246.240 246.850 1246.500 247.170 ;
        RECT 1186.500 17.410 1186.640 246.850 ;
        RECT 1186.040 17.270 1186.640 17.410 ;
        RECT 1186.040 2.400 1186.180 17.270 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 248.100 1207.430 248.160 ;
        RECT 1260.470 248.100 1260.790 248.160 ;
        RECT 1207.110 247.960 1260.790 248.100 ;
        RECT 1207.110 247.900 1207.430 247.960 ;
        RECT 1260.470 247.900 1260.790 247.960 ;
        RECT 1203.890 17.580 1204.210 17.640 ;
        RECT 1207.110 17.580 1207.430 17.640 ;
        RECT 1203.890 17.440 1207.430 17.580 ;
        RECT 1203.890 17.380 1204.210 17.440 ;
        RECT 1207.110 17.380 1207.430 17.440 ;
      LAYER via ;
        RECT 1207.140 247.900 1207.400 248.160 ;
        RECT 1260.500 247.900 1260.760 248.160 ;
        RECT 1203.920 17.380 1204.180 17.640 ;
        RECT 1207.140 17.380 1207.400 17.640 ;
      LAYER met2 ;
        RECT 1260.450 260.000 1260.730 264.000 ;
        RECT 1260.560 248.190 1260.700 260.000 ;
        RECT 1207.140 247.870 1207.400 248.190 ;
        RECT 1260.500 247.870 1260.760 248.190 ;
        RECT 1207.200 17.670 1207.340 247.870 ;
        RECT 1203.920 17.350 1204.180 17.670 ;
        RECT 1207.140 17.350 1207.400 17.670 ;
        RECT 1203.980 2.400 1204.120 17.350 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.810 248.440 1228.130 248.500 ;
        RECT 1274.270 248.440 1274.590 248.500 ;
        RECT 1227.810 248.300 1274.590 248.440 ;
        RECT 1227.810 248.240 1228.130 248.300 ;
        RECT 1274.270 248.240 1274.590 248.300 ;
        RECT 1221.830 17.580 1222.150 17.640 ;
        RECT 1227.350 17.580 1227.670 17.640 ;
        RECT 1221.830 17.440 1227.670 17.580 ;
        RECT 1221.830 17.380 1222.150 17.440 ;
        RECT 1227.350 17.380 1227.670 17.440 ;
      LAYER via ;
        RECT 1227.840 248.240 1228.100 248.500 ;
        RECT 1274.300 248.240 1274.560 248.500 ;
        RECT 1221.860 17.380 1222.120 17.640 ;
        RECT 1227.380 17.380 1227.640 17.640 ;
      LAYER met2 ;
        RECT 1274.250 260.000 1274.530 264.000 ;
        RECT 1274.360 248.530 1274.500 260.000 ;
        RECT 1227.840 248.210 1228.100 248.530 ;
        RECT 1274.300 248.210 1274.560 248.530 ;
        RECT 1227.900 245.890 1228.040 248.210 ;
        RECT 1227.440 245.750 1228.040 245.890 ;
        RECT 1227.440 17.670 1227.580 245.750 ;
        RECT 1221.860 17.350 1222.120 17.670 ;
        RECT 1227.380 17.350 1227.640 17.670 ;
        RECT 1221.920 2.400 1222.060 17.350 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 247.760 1241.930 247.820 ;
        RECT 1288.530 247.760 1288.850 247.820 ;
        RECT 1241.610 247.620 1288.850 247.760 ;
        RECT 1241.610 247.560 1241.930 247.620 ;
        RECT 1288.530 247.560 1288.850 247.620 ;
      LAYER via ;
        RECT 1241.640 247.560 1241.900 247.820 ;
        RECT 1288.560 247.560 1288.820 247.820 ;
      LAYER met2 ;
        RECT 1288.510 260.000 1288.790 264.000 ;
        RECT 1288.620 247.850 1288.760 260.000 ;
        RECT 1241.640 247.530 1241.900 247.850 ;
        RECT 1288.560 247.530 1288.820 247.850 ;
        RECT 1241.700 16.730 1241.840 247.530 ;
        RECT 1239.860 16.590 1241.840 16.730 ;
        RECT 1239.860 2.400 1240.000 16.590 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 245.040 1262.630 245.100 ;
        RECT 1302.790 245.040 1303.110 245.100 ;
        RECT 1262.310 244.900 1303.110 245.040 ;
        RECT 1262.310 244.840 1262.630 244.900 ;
        RECT 1302.790 244.840 1303.110 244.900 ;
        RECT 1257.250 17.580 1257.570 17.640 ;
        RECT 1262.310 17.580 1262.630 17.640 ;
        RECT 1257.250 17.440 1262.630 17.580 ;
        RECT 1257.250 17.380 1257.570 17.440 ;
        RECT 1262.310 17.380 1262.630 17.440 ;
      LAYER via ;
        RECT 1262.340 244.840 1262.600 245.100 ;
        RECT 1302.820 244.840 1303.080 245.100 ;
        RECT 1257.280 17.380 1257.540 17.640 ;
        RECT 1262.340 17.380 1262.600 17.640 ;
      LAYER met2 ;
        RECT 1302.770 260.000 1303.050 264.000 ;
        RECT 1302.880 245.130 1303.020 260.000 ;
        RECT 1262.340 244.810 1262.600 245.130 ;
        RECT 1302.820 244.810 1303.080 245.130 ;
        RECT 1262.400 17.670 1262.540 244.810 ;
        RECT 1257.280 17.350 1257.540 17.670 ;
        RECT 1262.340 17.350 1262.600 17.670 ;
        RECT 1257.340 2.400 1257.480 17.350 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 247.420 1276.430 247.480 ;
        RECT 1316.590 247.420 1316.910 247.480 ;
        RECT 1276.110 247.280 1316.910 247.420 ;
        RECT 1276.110 247.220 1276.430 247.280 ;
        RECT 1316.590 247.220 1316.910 247.280 ;
      LAYER via ;
        RECT 1276.140 247.220 1276.400 247.480 ;
        RECT 1316.620 247.220 1316.880 247.480 ;
      LAYER met2 ;
        RECT 1316.570 260.000 1316.850 264.000 ;
        RECT 1316.680 247.510 1316.820 260.000 ;
        RECT 1276.140 247.190 1276.400 247.510 ;
        RECT 1316.620 247.190 1316.880 247.510 ;
        RECT 1276.200 17.410 1276.340 247.190 ;
        RECT 1275.280 17.270 1276.340 17.410 ;
        RECT 1275.280 2.400 1275.420 17.270 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 244.020 1297.130 244.080 ;
        RECT 1330.850 244.020 1331.170 244.080 ;
        RECT 1296.810 243.880 1331.170 244.020 ;
        RECT 1296.810 243.820 1297.130 243.880 ;
        RECT 1330.850 243.820 1331.170 243.880 ;
        RECT 1293.130 15.540 1293.450 15.600 ;
        RECT 1296.810 15.540 1297.130 15.600 ;
        RECT 1293.130 15.400 1297.130 15.540 ;
        RECT 1293.130 15.340 1293.450 15.400 ;
        RECT 1296.810 15.340 1297.130 15.400 ;
      LAYER via ;
        RECT 1296.840 243.820 1297.100 244.080 ;
        RECT 1330.880 243.820 1331.140 244.080 ;
        RECT 1293.160 15.340 1293.420 15.600 ;
        RECT 1296.840 15.340 1297.100 15.600 ;
      LAYER met2 ;
        RECT 1330.830 260.000 1331.110 264.000 ;
        RECT 1330.940 244.110 1331.080 260.000 ;
        RECT 1296.840 243.790 1297.100 244.110 ;
        RECT 1330.880 243.790 1331.140 244.110 ;
        RECT 1296.900 15.630 1297.040 243.790 ;
        RECT 1293.160 15.310 1293.420 15.630 ;
        RECT 1296.840 15.310 1297.100 15.630 ;
        RECT 1293.220 2.400 1293.360 15.310 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1317.510 242.660 1317.830 242.720 ;
        RECT 1344.650 242.660 1344.970 242.720 ;
        RECT 1317.510 242.520 1344.970 242.660 ;
        RECT 1317.510 242.460 1317.830 242.520 ;
        RECT 1344.650 242.460 1344.970 242.520 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 1317.510 17.580 1317.830 17.640 ;
        RECT 1311.070 17.440 1317.830 17.580 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
        RECT 1317.510 17.380 1317.830 17.440 ;
      LAYER via ;
        RECT 1317.540 242.460 1317.800 242.720 ;
        RECT 1344.680 242.460 1344.940 242.720 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
        RECT 1317.540 17.380 1317.800 17.640 ;
      LAYER met2 ;
        RECT 1344.630 260.000 1344.910 264.000 ;
        RECT 1344.740 242.750 1344.880 260.000 ;
        RECT 1317.540 242.430 1317.800 242.750 ;
        RECT 1344.680 242.430 1344.940 242.750 ;
        RECT 1317.600 17.670 1317.740 242.430 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 1317.540 17.350 1317.800 17.670 ;
        RECT 1311.160 2.400 1311.300 17.350 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 246.400 1331.630 246.460 ;
        RECT 1358.910 246.400 1359.230 246.460 ;
        RECT 1331.310 246.260 1359.230 246.400 ;
        RECT 1331.310 246.200 1331.630 246.260 ;
        RECT 1358.910 246.200 1359.230 246.260 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1329.010 17.440 1331.630 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
      LAYER via ;
        RECT 1331.340 246.200 1331.600 246.460 ;
        RECT 1358.940 246.200 1359.200 246.460 ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1331.340 17.380 1331.600 17.640 ;
      LAYER met2 ;
        RECT 1358.890 260.000 1359.170 264.000 ;
        RECT 1359.000 246.490 1359.140 260.000 ;
        RECT 1331.340 246.170 1331.600 246.490 ;
        RECT 1358.940 246.170 1359.200 246.490 ;
        RECT 1331.400 17.670 1331.540 246.170 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 838.190 241.640 838.510 241.700 ;
        RECT 851.990 241.640 852.310 241.700 ;
        RECT 838.190 241.500 852.310 241.640 ;
        RECT 838.190 241.440 838.510 241.500 ;
        RECT 851.990 241.440 852.310 241.500 ;
        RECT 686.390 44.780 686.710 44.840 ;
        RECT 838.190 44.780 838.510 44.840 ;
        RECT 686.390 44.640 838.510 44.780 ;
        RECT 686.390 44.580 686.710 44.640 ;
        RECT 838.190 44.580 838.510 44.640 ;
      LAYER via ;
        RECT 838.220 241.440 838.480 241.700 ;
        RECT 852.020 241.440 852.280 241.700 ;
        RECT 686.420 44.580 686.680 44.840 ;
        RECT 838.220 44.580 838.480 44.840 ;
      LAYER met2 ;
        RECT 851.970 260.000 852.250 264.000 ;
        RECT 852.080 241.730 852.220 260.000 ;
        RECT 838.220 241.410 838.480 241.730 ;
        RECT 852.020 241.410 852.280 241.730 ;
        RECT 838.280 44.870 838.420 241.410 ;
        RECT 686.420 44.550 686.680 44.870 ;
        RECT 838.220 44.550 838.480 44.870 ;
        RECT 686.480 2.400 686.620 44.550 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.010 243.000 1352.330 243.060 ;
        RECT 1373.170 243.000 1373.490 243.060 ;
        RECT 1352.010 242.860 1373.490 243.000 ;
        RECT 1352.010 242.800 1352.330 242.860 ;
        RECT 1373.170 242.800 1373.490 242.860 ;
        RECT 1346.490 15.200 1346.810 15.260 ;
        RECT 1352.010 15.200 1352.330 15.260 ;
        RECT 1346.490 15.060 1352.330 15.200 ;
        RECT 1346.490 15.000 1346.810 15.060 ;
        RECT 1352.010 15.000 1352.330 15.060 ;
      LAYER via ;
        RECT 1352.040 242.800 1352.300 243.060 ;
        RECT 1373.200 242.800 1373.460 243.060 ;
        RECT 1346.520 15.000 1346.780 15.260 ;
        RECT 1352.040 15.000 1352.300 15.260 ;
      LAYER met2 ;
        RECT 1373.150 260.000 1373.430 264.000 ;
        RECT 1373.260 243.090 1373.400 260.000 ;
        RECT 1352.040 242.770 1352.300 243.090 ;
        RECT 1373.200 242.770 1373.460 243.090 ;
        RECT 1352.100 15.290 1352.240 242.770 ;
        RECT 1346.520 14.970 1346.780 15.290 ;
        RECT 1352.040 14.970 1352.300 15.290 ;
        RECT 1346.580 2.400 1346.720 14.970 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 245.380 1366.130 245.440 ;
        RECT 1386.970 245.380 1387.290 245.440 ;
        RECT 1365.810 245.240 1387.290 245.380 ;
        RECT 1365.810 245.180 1366.130 245.240 ;
        RECT 1386.970 245.180 1387.290 245.240 ;
      LAYER via ;
        RECT 1365.840 245.180 1366.100 245.440 ;
        RECT 1387.000 245.180 1387.260 245.440 ;
      LAYER met2 ;
        RECT 1386.950 260.000 1387.230 264.000 ;
        RECT 1387.060 245.470 1387.200 260.000 ;
        RECT 1365.840 245.150 1366.100 245.470 ;
        RECT 1387.000 245.150 1387.260 245.470 ;
        RECT 1365.900 17.410 1366.040 245.150 ;
        RECT 1364.520 17.270 1366.040 17.410 ;
        RECT 1364.520 2.400 1364.660 17.270 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.510 245.720 1386.830 245.780 ;
        RECT 1401.230 245.720 1401.550 245.780 ;
        RECT 1386.510 245.580 1401.550 245.720 ;
        RECT 1386.510 245.520 1386.830 245.580 ;
        RECT 1401.230 245.520 1401.550 245.580 ;
        RECT 1382.370 17.580 1382.690 17.640 ;
        RECT 1386.510 17.580 1386.830 17.640 ;
        RECT 1382.370 17.440 1386.830 17.580 ;
        RECT 1382.370 17.380 1382.690 17.440 ;
        RECT 1386.510 17.380 1386.830 17.440 ;
      LAYER via ;
        RECT 1386.540 245.520 1386.800 245.780 ;
        RECT 1401.260 245.520 1401.520 245.780 ;
        RECT 1382.400 17.380 1382.660 17.640 ;
        RECT 1386.540 17.380 1386.800 17.640 ;
      LAYER met2 ;
        RECT 1401.210 260.000 1401.490 264.000 ;
        RECT 1401.320 245.810 1401.460 260.000 ;
        RECT 1386.540 245.490 1386.800 245.810 ;
        RECT 1401.260 245.490 1401.520 245.810 ;
        RECT 1386.600 17.670 1386.740 245.490 ;
        RECT 1382.400 17.350 1382.660 17.670 ;
        RECT 1386.540 17.350 1386.800 17.670 ;
        RECT 1382.460 2.400 1382.600 17.350 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1399.850 243.000 1400.170 243.060 ;
        RECT 1415.030 243.000 1415.350 243.060 ;
        RECT 1399.850 242.860 1415.350 243.000 ;
        RECT 1399.850 242.800 1400.170 242.860 ;
        RECT 1415.030 242.800 1415.350 242.860 ;
      LAYER via ;
        RECT 1399.880 242.800 1400.140 243.060 ;
        RECT 1415.060 242.800 1415.320 243.060 ;
      LAYER met2 ;
        RECT 1415.010 260.000 1415.290 264.000 ;
        RECT 1415.120 243.090 1415.260 260.000 ;
        RECT 1399.880 242.770 1400.140 243.090 ;
        RECT 1415.060 242.770 1415.320 243.090 ;
        RECT 1399.940 24.210 1400.080 242.770 ;
        RECT 1399.940 24.070 1400.540 24.210 ;
        RECT 1400.400 2.400 1400.540 24.070 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 241.640 1421.330 241.700 ;
        RECT 1429.290 241.640 1429.610 241.700 ;
        RECT 1421.010 241.500 1429.610 241.640 ;
        RECT 1421.010 241.440 1421.330 241.500 ;
        RECT 1429.290 241.440 1429.610 241.500 ;
        RECT 1418.250 15.540 1418.570 15.600 ;
        RECT 1421.010 15.540 1421.330 15.600 ;
        RECT 1418.250 15.400 1421.330 15.540 ;
        RECT 1418.250 15.340 1418.570 15.400 ;
        RECT 1421.010 15.340 1421.330 15.400 ;
      LAYER via ;
        RECT 1421.040 241.440 1421.300 241.700 ;
        RECT 1429.320 241.440 1429.580 241.700 ;
        RECT 1418.280 15.340 1418.540 15.600 ;
        RECT 1421.040 15.340 1421.300 15.600 ;
      LAYER met2 ;
        RECT 1429.270 260.000 1429.550 264.000 ;
        RECT 1429.380 241.730 1429.520 260.000 ;
        RECT 1421.040 241.410 1421.300 241.730 ;
        RECT 1429.320 241.410 1429.580 241.730 ;
        RECT 1421.100 15.630 1421.240 241.410 ;
        RECT 1418.280 15.310 1418.540 15.630 ;
        RECT 1421.040 15.310 1421.300 15.630 ;
        RECT 1418.340 2.400 1418.480 15.310 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1440.790 182.820 1441.110 182.880 ;
        RECT 1441.710 182.820 1442.030 182.880 ;
        RECT 1440.790 182.680 1442.030 182.820 ;
        RECT 1440.790 182.620 1441.110 182.680 ;
        RECT 1441.710 182.620 1442.030 182.680 ;
        RECT 1435.730 20.640 1436.050 20.700 ;
        RECT 1441.710 20.640 1442.030 20.700 ;
        RECT 1435.730 20.500 1442.030 20.640 ;
        RECT 1435.730 20.440 1436.050 20.500 ;
        RECT 1441.710 20.440 1442.030 20.500 ;
      LAYER via ;
        RECT 1440.820 182.620 1441.080 182.880 ;
        RECT 1441.740 182.620 1442.000 182.880 ;
        RECT 1435.760 20.440 1436.020 20.700 ;
        RECT 1441.740 20.440 1442.000 20.700 ;
      LAYER met2 ;
        RECT 1443.530 260.170 1443.810 264.000 ;
        RECT 1442.260 260.030 1443.810 260.170 ;
        RECT 1442.260 241.810 1442.400 260.030 ;
        RECT 1443.530 260.000 1443.810 260.030 ;
        RECT 1440.880 241.670 1442.400 241.810 ;
        RECT 1440.880 182.910 1441.020 241.670 ;
        RECT 1440.820 182.590 1441.080 182.910 ;
        RECT 1441.740 182.590 1442.000 182.910 ;
        RECT 1441.800 20.730 1441.940 182.590 ;
        RECT 1435.760 20.410 1436.020 20.730 ;
        RECT 1441.740 20.410 1442.000 20.730 ;
        RECT 1435.820 2.400 1435.960 20.410 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1455.125 138.125 1455.295 185.895 ;
      LAYER mcon ;
        RECT 1455.125 185.725 1455.295 185.895 ;
      LAYER met1 ;
        RECT 1454.590 241.640 1454.910 241.700 ;
        RECT 1457.350 241.640 1457.670 241.700 ;
        RECT 1454.590 241.500 1457.670 241.640 ;
        RECT 1454.590 241.440 1454.910 241.500 ;
        RECT 1457.350 241.440 1457.670 241.500 ;
        RECT 1454.130 185.880 1454.450 185.940 ;
        RECT 1455.065 185.880 1455.355 185.925 ;
        RECT 1454.130 185.740 1455.355 185.880 ;
        RECT 1454.130 185.680 1454.450 185.740 ;
        RECT 1455.065 185.695 1455.355 185.740 ;
        RECT 1455.050 138.280 1455.370 138.340 ;
        RECT 1454.855 138.140 1455.370 138.280 ;
        RECT 1455.050 138.080 1455.370 138.140 ;
        RECT 1453.210 93.060 1453.530 93.120 ;
        RECT 1455.510 93.060 1455.830 93.120 ;
        RECT 1453.210 92.920 1455.830 93.060 ;
        RECT 1453.210 92.860 1453.530 92.920 ;
        RECT 1455.510 92.860 1455.830 92.920 ;
      LAYER via ;
        RECT 1454.620 241.440 1454.880 241.700 ;
        RECT 1457.380 241.440 1457.640 241.700 ;
        RECT 1454.160 185.680 1454.420 185.940 ;
        RECT 1455.080 138.080 1455.340 138.340 ;
        RECT 1453.240 92.860 1453.500 93.120 ;
        RECT 1455.540 92.860 1455.800 93.120 ;
      LAYER met2 ;
        RECT 1457.330 260.000 1457.610 264.000 ;
        RECT 1457.440 241.730 1457.580 260.000 ;
        RECT 1454.620 241.410 1454.880 241.730 ;
        RECT 1457.380 241.410 1457.640 241.730 ;
        RECT 1454.680 210.530 1454.820 241.410 ;
        RECT 1454.220 210.390 1454.820 210.530 ;
        RECT 1454.220 185.970 1454.360 210.390 ;
        RECT 1454.160 185.650 1454.420 185.970 ;
        RECT 1455.080 138.050 1455.340 138.370 ;
        RECT 1455.140 137.770 1455.280 138.050 ;
        RECT 1455.140 137.630 1455.740 137.770 ;
        RECT 1455.600 93.150 1455.740 137.630 ;
        RECT 1453.240 92.830 1453.500 93.150 ;
        RECT 1455.540 92.830 1455.800 93.150 ;
        RECT 1453.300 13.330 1453.440 92.830 ;
        RECT 1453.300 13.190 1453.900 13.330 ;
        RECT 1453.760 2.400 1453.900 13.190 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1469.845 186.405 1470.015 234.515 ;
        RECT 1469.845 89.845 1470.015 137.955 ;
      LAYER mcon ;
        RECT 1469.845 234.345 1470.015 234.515 ;
        RECT 1469.845 137.785 1470.015 137.955 ;
      LAYER met1 ;
        RECT 1469.770 234.500 1470.090 234.560 ;
        RECT 1469.575 234.360 1470.090 234.500 ;
        RECT 1469.770 234.300 1470.090 234.360 ;
        RECT 1469.770 186.560 1470.090 186.620 ;
        RECT 1469.575 186.420 1470.090 186.560 ;
        RECT 1469.770 186.360 1470.090 186.420 ;
        RECT 1469.770 137.940 1470.090 138.000 ;
        RECT 1469.575 137.800 1470.090 137.940 ;
        RECT 1469.770 137.740 1470.090 137.800 ;
        RECT 1469.770 90.000 1470.090 90.060 ;
        RECT 1469.575 89.860 1470.090 90.000 ;
        RECT 1469.770 89.800 1470.090 89.860 ;
      LAYER via ;
        RECT 1469.800 234.300 1470.060 234.560 ;
        RECT 1469.800 186.360 1470.060 186.620 ;
        RECT 1469.800 137.740 1470.060 138.000 ;
        RECT 1469.800 89.800 1470.060 90.060 ;
      LAYER met2 ;
        RECT 1471.590 260.170 1471.870 264.000 ;
        RECT 1469.860 260.030 1471.870 260.170 ;
        RECT 1469.860 234.590 1470.000 260.030 ;
        RECT 1471.590 260.000 1471.870 260.030 ;
        RECT 1469.800 234.270 1470.060 234.590 ;
        RECT 1469.800 186.330 1470.060 186.650 ;
        RECT 1469.860 138.030 1470.000 186.330 ;
        RECT 1469.800 137.710 1470.060 138.030 ;
        RECT 1469.800 89.770 1470.060 90.090 ;
        RECT 1469.860 73.170 1470.000 89.770 ;
        RECT 1469.860 73.030 1471.840 73.170 ;
        RECT 1471.700 2.400 1471.840 73.030 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1484.030 20.640 1484.350 20.700 ;
        RECT 1489.550 20.640 1489.870 20.700 ;
        RECT 1484.030 20.500 1489.870 20.640 ;
        RECT 1484.030 20.440 1484.350 20.500 ;
        RECT 1489.550 20.440 1489.870 20.500 ;
      LAYER via ;
        RECT 1484.060 20.440 1484.320 20.700 ;
        RECT 1489.580 20.440 1489.840 20.700 ;
      LAYER met2 ;
        RECT 1485.850 260.170 1486.130 264.000 ;
        RECT 1484.120 260.030 1486.130 260.170 ;
        RECT 1484.120 20.730 1484.260 260.030 ;
        RECT 1485.850 260.000 1486.130 260.030 ;
        RECT 1484.060 20.410 1484.320 20.730 ;
        RECT 1489.580 20.410 1489.840 20.730 ;
        RECT 1489.640 2.400 1489.780 20.410 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1499.670 244.020 1499.990 244.080 ;
        RECT 1505.190 244.020 1505.510 244.080 ;
        RECT 1499.670 243.880 1505.510 244.020 ;
        RECT 1499.670 243.820 1499.990 243.880 ;
        RECT 1505.190 243.820 1505.510 243.880 ;
        RECT 1504.730 61.440 1505.050 61.500 ;
        RECT 1507.030 61.440 1507.350 61.500 ;
        RECT 1504.730 61.300 1507.350 61.440 ;
        RECT 1504.730 61.240 1505.050 61.300 ;
        RECT 1507.030 61.240 1507.350 61.300 ;
      LAYER via ;
        RECT 1499.700 243.820 1499.960 244.080 ;
        RECT 1505.220 243.820 1505.480 244.080 ;
        RECT 1504.760 61.240 1505.020 61.500 ;
        RECT 1507.060 61.240 1507.320 61.500 ;
      LAYER met2 ;
        RECT 1499.650 260.000 1499.930 264.000 ;
        RECT 1499.760 244.110 1499.900 260.000 ;
        RECT 1499.700 243.790 1499.960 244.110 ;
        RECT 1505.220 243.790 1505.480 244.110 ;
        RECT 1505.280 72.490 1505.420 243.790 ;
        RECT 1504.820 72.350 1505.420 72.490 ;
        RECT 1504.820 61.530 1504.960 72.350 ;
        RECT 1504.760 61.210 1505.020 61.530 ;
        RECT 1507.060 61.210 1507.320 61.530 ;
        RECT 1507.120 2.400 1507.260 61.210 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 709.850 51.580 710.170 51.640 ;
        RECT 862.570 51.580 862.890 51.640 ;
        RECT 709.850 51.440 862.890 51.580 ;
        RECT 709.850 51.380 710.170 51.440 ;
        RECT 862.570 51.380 862.890 51.440 ;
        RECT 704.330 17.920 704.650 17.980 ;
        RECT 709.850 17.920 710.170 17.980 ;
        RECT 704.330 17.780 710.170 17.920 ;
        RECT 704.330 17.720 704.650 17.780 ;
        RECT 709.850 17.720 710.170 17.780 ;
      LAYER via ;
        RECT 709.880 51.380 710.140 51.640 ;
        RECT 862.600 51.380 862.860 51.640 ;
        RECT 704.360 17.720 704.620 17.980 ;
        RECT 709.880 17.720 710.140 17.980 ;
      LAYER met2 ;
        RECT 866.230 260.170 866.510 264.000 ;
        RECT 862.660 260.030 866.510 260.170 ;
        RECT 862.660 51.670 862.800 260.030 ;
        RECT 866.230 260.000 866.510 260.030 ;
        RECT 709.880 51.350 710.140 51.670 ;
        RECT 862.600 51.350 862.860 51.670 ;
        RECT 709.940 18.010 710.080 51.350 ;
        RECT 704.360 17.690 704.620 18.010 ;
        RECT 709.880 17.690 710.140 18.010 ;
        RECT 704.420 2.400 704.560 17.690 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.610 17.240 1517.930 17.300 ;
        RECT 1524.970 17.240 1525.290 17.300 ;
        RECT 1517.610 17.100 1525.290 17.240 ;
        RECT 1517.610 17.040 1517.930 17.100 ;
        RECT 1524.970 17.040 1525.290 17.100 ;
      LAYER via ;
        RECT 1517.640 17.040 1517.900 17.300 ;
        RECT 1525.000 17.040 1525.260 17.300 ;
      LAYER met2 ;
        RECT 1513.910 260.170 1514.190 264.000 ;
        RECT 1513.910 260.030 1517.840 260.170 ;
        RECT 1513.910 260.000 1514.190 260.030 ;
        RECT 1517.700 17.330 1517.840 260.030 ;
        RECT 1517.640 17.010 1517.900 17.330 ;
        RECT 1525.000 17.010 1525.260 17.330 ;
        RECT 1525.060 2.400 1525.200 17.010 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.410 20.640 1531.730 20.700 ;
        RECT 1542.910 20.640 1543.230 20.700 ;
        RECT 1531.410 20.500 1543.230 20.640 ;
        RECT 1531.410 20.440 1531.730 20.500 ;
        RECT 1542.910 20.440 1543.230 20.500 ;
      LAYER via ;
        RECT 1531.440 20.440 1531.700 20.700 ;
        RECT 1542.940 20.440 1543.200 20.700 ;
      LAYER met2 ;
        RECT 1527.710 260.170 1527.990 264.000 ;
        RECT 1527.710 260.030 1531.640 260.170 ;
        RECT 1527.710 260.000 1527.990 260.030 ;
        RECT 1531.500 20.730 1531.640 260.030 ;
        RECT 1531.440 20.410 1531.700 20.730 ;
        RECT 1542.940 20.410 1543.200 20.730 ;
        RECT 1543.000 2.400 1543.140 20.410 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 17.920 1545.530 17.980 ;
        RECT 1560.850 17.920 1561.170 17.980 ;
        RECT 1545.210 17.780 1561.170 17.920 ;
        RECT 1545.210 17.720 1545.530 17.780 ;
        RECT 1560.850 17.720 1561.170 17.780 ;
      LAYER via ;
        RECT 1545.240 17.720 1545.500 17.980 ;
        RECT 1560.880 17.720 1561.140 17.980 ;
      LAYER met2 ;
        RECT 1541.970 260.170 1542.250 264.000 ;
        RECT 1541.970 260.030 1545.440 260.170 ;
        RECT 1541.970 260.000 1542.250 260.030 ;
        RECT 1545.300 18.010 1545.440 260.030 ;
        RECT 1545.240 17.690 1545.500 18.010 ;
        RECT 1560.880 17.690 1561.140 18.010 ;
        RECT 1560.940 2.400 1561.080 17.690 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1556.250 244.020 1556.570 244.080 ;
        RECT 1562.690 244.020 1563.010 244.080 ;
        RECT 1556.250 243.880 1563.010 244.020 ;
        RECT 1556.250 243.820 1556.570 243.880 ;
        RECT 1562.690 243.820 1563.010 243.880 ;
        RECT 1562.690 16.220 1563.010 16.280 ;
        RECT 1578.790 16.220 1579.110 16.280 ;
        RECT 1562.690 16.080 1579.110 16.220 ;
        RECT 1562.690 16.020 1563.010 16.080 ;
        RECT 1578.790 16.020 1579.110 16.080 ;
      LAYER via ;
        RECT 1556.280 243.820 1556.540 244.080 ;
        RECT 1562.720 243.820 1562.980 244.080 ;
        RECT 1562.720 16.020 1562.980 16.280 ;
        RECT 1578.820 16.020 1579.080 16.280 ;
      LAYER met2 ;
        RECT 1556.230 260.000 1556.510 264.000 ;
        RECT 1556.340 244.110 1556.480 260.000 ;
        RECT 1556.280 243.790 1556.540 244.110 ;
        RECT 1562.720 243.790 1562.980 244.110 ;
        RECT 1562.780 16.310 1562.920 243.790 ;
        RECT 1562.720 15.990 1562.980 16.310 ;
        RECT 1578.820 15.990 1579.080 16.310 ;
        RECT 1578.880 2.400 1579.020 15.990 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1570.050 244.020 1570.370 244.080 ;
        RECT 1576.490 244.020 1576.810 244.080 ;
        RECT 1570.050 243.880 1576.810 244.020 ;
        RECT 1570.050 243.820 1570.370 243.880 ;
        RECT 1576.490 243.820 1576.810 243.880 ;
        RECT 1576.490 18.940 1576.810 19.000 ;
        RECT 1596.270 18.940 1596.590 19.000 ;
        RECT 1576.490 18.800 1596.590 18.940 ;
        RECT 1576.490 18.740 1576.810 18.800 ;
        RECT 1596.270 18.740 1596.590 18.800 ;
      LAYER via ;
        RECT 1570.080 243.820 1570.340 244.080 ;
        RECT 1576.520 243.820 1576.780 244.080 ;
        RECT 1576.520 18.740 1576.780 19.000 ;
        RECT 1596.300 18.740 1596.560 19.000 ;
      LAYER met2 ;
        RECT 1570.030 260.000 1570.310 264.000 ;
        RECT 1570.140 244.110 1570.280 260.000 ;
        RECT 1570.080 243.790 1570.340 244.110 ;
        RECT 1576.520 243.790 1576.780 244.110 ;
        RECT 1576.580 19.030 1576.720 243.790 ;
        RECT 1576.520 18.710 1576.780 19.030 ;
        RECT 1596.300 18.710 1596.560 19.030 ;
        RECT 1596.360 2.400 1596.500 18.710 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1586.610 16.220 1586.930 16.280 ;
        RECT 1614.210 16.220 1614.530 16.280 ;
        RECT 1586.610 16.080 1614.530 16.220 ;
        RECT 1586.610 16.020 1586.930 16.080 ;
        RECT 1614.210 16.020 1614.530 16.080 ;
      LAYER via ;
        RECT 1586.640 16.020 1586.900 16.280 ;
        RECT 1614.240 16.020 1614.500 16.280 ;
      LAYER met2 ;
        RECT 1584.290 260.170 1584.570 264.000 ;
        RECT 1584.290 260.030 1586.840 260.170 ;
        RECT 1584.290 260.000 1584.570 260.030 ;
        RECT 1586.700 16.310 1586.840 260.030 ;
        RECT 1586.640 15.990 1586.900 16.310 ;
        RECT 1614.240 15.990 1614.500 16.310 ;
        RECT 1614.300 2.400 1614.440 15.990 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 19.960 1600.730 20.020 ;
        RECT 1632.150 19.960 1632.470 20.020 ;
        RECT 1600.410 19.820 1632.470 19.960 ;
        RECT 1600.410 19.760 1600.730 19.820 ;
        RECT 1632.150 19.760 1632.470 19.820 ;
      LAYER via ;
        RECT 1600.440 19.760 1600.700 20.020 ;
        RECT 1632.180 19.760 1632.440 20.020 ;
      LAYER met2 ;
        RECT 1598.090 260.170 1598.370 264.000 ;
        RECT 1598.090 260.030 1600.640 260.170 ;
        RECT 1598.090 260.000 1598.370 260.030 ;
        RECT 1600.500 20.050 1600.640 260.030 ;
        RECT 1600.440 19.730 1600.700 20.050 ;
        RECT 1632.180 19.730 1632.440 20.050 ;
        RECT 1632.240 2.400 1632.380 19.730 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 17.240 1614.530 17.300 ;
        RECT 1650.090 17.240 1650.410 17.300 ;
        RECT 1614.210 17.100 1650.410 17.240 ;
        RECT 1614.210 17.040 1614.530 17.100 ;
        RECT 1650.090 17.040 1650.410 17.100 ;
      LAYER via ;
        RECT 1614.240 17.040 1614.500 17.300 ;
        RECT 1650.120 17.040 1650.380 17.300 ;
      LAYER met2 ;
        RECT 1612.350 260.170 1612.630 264.000 ;
        RECT 1612.350 260.030 1614.440 260.170 ;
        RECT 1612.350 260.000 1612.630 260.030 ;
        RECT 1614.300 17.330 1614.440 260.030 ;
        RECT 1614.240 17.010 1614.500 17.330 ;
        RECT 1650.120 17.010 1650.380 17.330 ;
        RECT 1650.180 2.400 1650.320 17.010 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1628.010 18.600 1628.330 18.660 ;
        RECT 1668.030 18.600 1668.350 18.660 ;
        RECT 1628.010 18.460 1668.350 18.600 ;
        RECT 1628.010 18.400 1628.330 18.460 ;
        RECT 1668.030 18.400 1668.350 18.460 ;
      LAYER via ;
        RECT 1628.040 18.400 1628.300 18.660 ;
        RECT 1668.060 18.400 1668.320 18.660 ;
      LAYER met2 ;
        RECT 1626.610 260.170 1626.890 264.000 ;
        RECT 1626.610 260.030 1628.240 260.170 ;
        RECT 1626.610 260.000 1626.890 260.030 ;
        RECT 1628.100 18.690 1628.240 260.030 ;
        RECT 1628.040 18.370 1628.300 18.690 ;
        RECT 1668.060 18.370 1668.320 18.690 ;
        RECT 1668.120 2.400 1668.260 18.370 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.510 17.580 1685.830 17.640 ;
        RECT 1662.600 17.440 1685.830 17.580 ;
        RECT 1641.350 16.900 1641.670 16.960 ;
        RECT 1662.600 16.900 1662.740 17.440 ;
        RECT 1685.510 17.380 1685.830 17.440 ;
        RECT 1641.350 16.760 1662.740 16.900 ;
        RECT 1641.350 16.700 1641.670 16.760 ;
      LAYER via ;
        RECT 1641.380 16.700 1641.640 16.960 ;
        RECT 1685.540 17.380 1685.800 17.640 ;
      LAYER met2 ;
        RECT 1640.410 260.170 1640.690 264.000 ;
        RECT 1640.410 260.030 1641.580 260.170 ;
        RECT 1640.410 260.000 1640.690 260.030 ;
        RECT 1641.440 16.990 1641.580 260.030 ;
        RECT 1685.540 17.350 1685.800 17.670 ;
        RECT 1641.380 16.670 1641.640 16.990 ;
        RECT 1685.600 2.400 1685.740 17.350 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 58.720 724.430 58.780 ;
        RECT 876.370 58.720 876.690 58.780 ;
        RECT 724.110 58.580 876.690 58.720 ;
        RECT 724.110 58.520 724.430 58.580 ;
        RECT 876.370 58.520 876.690 58.580 ;
      LAYER via ;
        RECT 724.140 58.520 724.400 58.780 ;
        RECT 876.400 58.520 876.660 58.780 ;
      LAYER met2 ;
        RECT 880.030 260.170 880.310 264.000 ;
        RECT 876.460 260.030 880.310 260.170 ;
        RECT 876.460 58.810 876.600 260.030 ;
        RECT 880.030 260.000 880.310 260.030 ;
        RECT 724.140 58.490 724.400 58.810 ;
        RECT 876.400 58.490 876.660 58.810 ;
        RECT 724.200 3.130 724.340 58.490 ;
        RECT 722.360 2.990 724.340 3.130 ;
        RECT 722.360 2.400 722.500 2.990 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.450 17.240 1703.770 17.300 ;
        RECT 1663.060 17.100 1703.770 17.240 ;
        RECT 1655.150 16.560 1655.470 16.620 ;
        RECT 1663.060 16.560 1663.200 17.100 ;
        RECT 1703.450 17.040 1703.770 17.100 ;
        RECT 1655.150 16.420 1663.200 16.560 ;
        RECT 1655.150 16.360 1655.470 16.420 ;
      LAYER via ;
        RECT 1655.180 16.360 1655.440 16.620 ;
        RECT 1703.480 17.040 1703.740 17.300 ;
      LAYER met2 ;
        RECT 1654.670 260.170 1654.950 264.000 ;
        RECT 1654.670 260.030 1655.380 260.170 ;
        RECT 1654.670 260.000 1654.950 260.030 ;
        RECT 1655.240 16.650 1655.380 260.030 ;
        RECT 1703.480 17.010 1703.740 17.330 ;
        RECT 1655.180 16.330 1655.440 16.650 ;
        RECT 1703.540 2.400 1703.680 17.010 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.950 18.600 1669.270 18.660 ;
        RECT 1721.390 18.600 1721.710 18.660 ;
        RECT 1668.950 18.460 1721.710 18.600 ;
        RECT 1668.950 18.400 1669.270 18.460 ;
        RECT 1721.390 18.400 1721.710 18.460 ;
      LAYER via ;
        RECT 1668.980 18.400 1669.240 18.660 ;
        RECT 1721.420 18.400 1721.680 18.660 ;
      LAYER met2 ;
        RECT 1668.470 260.170 1668.750 264.000 ;
        RECT 1668.470 260.030 1669.180 260.170 ;
        RECT 1668.470 260.000 1668.750 260.030 ;
        RECT 1669.040 18.690 1669.180 260.030 ;
        RECT 1668.980 18.370 1669.240 18.690 ;
        RECT 1721.420 18.370 1721.680 18.690 ;
        RECT 1721.480 2.400 1721.620 18.370 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1682.750 18.260 1683.070 18.320 ;
        RECT 1739.330 18.260 1739.650 18.320 ;
        RECT 1682.750 18.120 1739.650 18.260 ;
        RECT 1682.750 18.060 1683.070 18.120 ;
        RECT 1739.330 18.060 1739.650 18.120 ;
      LAYER via ;
        RECT 1682.780 18.060 1683.040 18.320 ;
        RECT 1739.360 18.060 1739.620 18.320 ;
      LAYER met2 ;
        RECT 1682.730 260.000 1683.010 264.000 ;
        RECT 1682.840 18.350 1682.980 260.000 ;
        RECT 1682.780 18.030 1683.040 18.350 ;
        RECT 1739.360 18.030 1739.620 18.350 ;
        RECT 1739.420 2.400 1739.560 18.030 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1696.550 17.920 1696.870 17.980 ;
        RECT 1756.810 17.920 1757.130 17.980 ;
        RECT 1696.550 17.780 1757.130 17.920 ;
        RECT 1696.550 17.720 1696.870 17.780 ;
        RECT 1756.810 17.720 1757.130 17.780 ;
      LAYER via ;
        RECT 1696.580 17.720 1696.840 17.980 ;
        RECT 1756.840 17.720 1757.100 17.980 ;
      LAYER met2 ;
        RECT 1696.990 260.170 1697.270 264.000 ;
        RECT 1696.640 260.030 1697.270 260.170 ;
        RECT 1696.640 18.010 1696.780 260.030 ;
        RECT 1696.990 260.000 1697.270 260.030 ;
        RECT 1696.580 17.690 1696.840 18.010 ;
        RECT 1756.840 17.690 1757.100 18.010 ;
        RECT 1756.900 2.400 1757.040 17.690 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.350 17.240 1710.670 17.300 ;
        RECT 1774.750 17.240 1775.070 17.300 ;
        RECT 1710.350 17.100 1775.070 17.240 ;
        RECT 1710.350 17.040 1710.670 17.100 ;
        RECT 1774.750 17.040 1775.070 17.100 ;
      LAYER via ;
        RECT 1710.380 17.040 1710.640 17.300 ;
        RECT 1774.780 17.040 1775.040 17.300 ;
      LAYER met2 ;
        RECT 1710.790 260.170 1711.070 264.000 ;
        RECT 1710.440 260.030 1711.070 260.170 ;
        RECT 1710.440 17.330 1710.580 260.030 ;
        RECT 1710.790 260.000 1711.070 260.030 ;
        RECT 1710.380 17.010 1710.640 17.330 ;
        RECT 1774.780 17.010 1775.040 17.330 ;
        RECT 1774.840 2.400 1774.980 17.010 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1725.070 244.020 1725.390 244.080 ;
        RECT 1731.050 244.020 1731.370 244.080 ;
        RECT 1725.070 243.880 1731.370 244.020 ;
        RECT 1725.070 243.820 1725.390 243.880 ;
        RECT 1731.050 243.820 1731.370 243.880 ;
        RECT 1731.050 16.900 1731.370 16.960 ;
        RECT 1792.690 16.900 1793.010 16.960 ;
        RECT 1731.050 16.760 1793.010 16.900 ;
        RECT 1731.050 16.700 1731.370 16.760 ;
        RECT 1792.690 16.700 1793.010 16.760 ;
      LAYER via ;
        RECT 1725.100 243.820 1725.360 244.080 ;
        RECT 1731.080 243.820 1731.340 244.080 ;
        RECT 1731.080 16.700 1731.340 16.960 ;
        RECT 1792.720 16.700 1792.980 16.960 ;
      LAYER met2 ;
        RECT 1725.050 260.000 1725.330 264.000 ;
        RECT 1725.160 244.110 1725.300 260.000 ;
        RECT 1725.100 243.790 1725.360 244.110 ;
        RECT 1731.080 243.790 1731.340 244.110 ;
        RECT 1731.140 16.990 1731.280 243.790 ;
        RECT 1731.080 16.670 1731.340 16.990 ;
        RECT 1792.720 16.670 1792.980 16.990 ;
        RECT 1792.780 2.400 1792.920 16.670 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.330 244.020 1739.650 244.080 ;
        RECT 1744.850 244.020 1745.170 244.080 ;
        RECT 1739.330 243.880 1745.170 244.020 ;
        RECT 1739.330 243.820 1739.650 243.880 ;
        RECT 1744.850 243.820 1745.170 243.880 ;
        RECT 1744.850 18.600 1745.170 18.660 ;
        RECT 1810.630 18.600 1810.950 18.660 ;
        RECT 1744.850 18.460 1810.950 18.600 ;
        RECT 1744.850 18.400 1745.170 18.460 ;
        RECT 1810.630 18.400 1810.950 18.460 ;
      LAYER via ;
        RECT 1739.360 243.820 1739.620 244.080 ;
        RECT 1744.880 243.820 1745.140 244.080 ;
        RECT 1744.880 18.400 1745.140 18.660 ;
        RECT 1810.660 18.400 1810.920 18.660 ;
      LAYER met2 ;
        RECT 1739.310 260.000 1739.590 264.000 ;
        RECT 1739.420 244.110 1739.560 260.000 ;
        RECT 1739.360 243.790 1739.620 244.110 ;
        RECT 1744.880 243.790 1745.140 244.110 ;
        RECT 1744.940 18.690 1745.080 243.790 ;
        RECT 1744.880 18.370 1745.140 18.690 ;
        RECT 1810.660 18.370 1810.920 18.690 ;
        RECT 1810.720 2.400 1810.860 18.370 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1753.130 245.040 1753.450 245.100 ;
        RECT 1829.030 245.040 1829.350 245.100 ;
        RECT 1753.130 244.900 1829.350 245.040 ;
        RECT 1753.130 244.840 1753.450 244.900 ;
        RECT 1829.030 244.840 1829.350 244.900 ;
      LAYER via ;
        RECT 1753.160 244.840 1753.420 245.100 ;
        RECT 1829.060 244.840 1829.320 245.100 ;
      LAYER met2 ;
        RECT 1753.110 260.000 1753.390 264.000 ;
        RECT 1753.220 245.130 1753.360 260.000 ;
        RECT 1753.160 244.810 1753.420 245.130 ;
        RECT 1829.060 244.810 1829.320 245.130 ;
        RECT 1829.120 3.130 1829.260 244.810 ;
        RECT 1828.660 2.990 1829.260 3.130 ;
        RECT 1828.660 2.400 1828.800 2.990 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1767.390 244.020 1767.710 244.080 ;
        RECT 1772.450 244.020 1772.770 244.080 ;
        RECT 1767.390 243.880 1772.770 244.020 ;
        RECT 1767.390 243.820 1767.710 243.880 ;
        RECT 1772.450 243.820 1772.770 243.880 ;
        RECT 1772.450 17.920 1772.770 17.980 ;
        RECT 1846.050 17.920 1846.370 17.980 ;
        RECT 1772.450 17.780 1846.370 17.920 ;
        RECT 1772.450 17.720 1772.770 17.780 ;
        RECT 1846.050 17.720 1846.370 17.780 ;
      LAYER via ;
        RECT 1767.420 243.820 1767.680 244.080 ;
        RECT 1772.480 243.820 1772.740 244.080 ;
        RECT 1772.480 17.720 1772.740 17.980 ;
        RECT 1846.080 17.720 1846.340 17.980 ;
      LAYER met2 ;
        RECT 1767.370 260.000 1767.650 264.000 ;
        RECT 1767.480 244.110 1767.620 260.000 ;
        RECT 1767.420 243.790 1767.680 244.110 ;
        RECT 1772.480 243.790 1772.740 244.110 ;
        RECT 1772.540 18.010 1772.680 243.790 ;
        RECT 1772.480 17.690 1772.740 18.010 ;
        RECT 1846.080 17.690 1846.340 18.010 ;
        RECT 1846.140 2.400 1846.280 17.690 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1781.190 244.020 1781.510 244.080 ;
        RECT 1786.250 244.020 1786.570 244.080 ;
        RECT 1781.190 243.880 1786.570 244.020 ;
        RECT 1781.190 243.820 1781.510 243.880 ;
        RECT 1786.250 243.820 1786.570 243.880 ;
        RECT 1786.250 24.040 1786.570 24.100 ;
        RECT 1863.990 24.040 1864.310 24.100 ;
        RECT 1786.250 23.900 1864.310 24.040 ;
        RECT 1786.250 23.840 1786.570 23.900 ;
        RECT 1863.990 23.840 1864.310 23.900 ;
      LAYER via ;
        RECT 1781.220 243.820 1781.480 244.080 ;
        RECT 1786.280 243.820 1786.540 244.080 ;
        RECT 1786.280 23.840 1786.540 24.100 ;
        RECT 1864.020 23.840 1864.280 24.100 ;
      LAYER met2 ;
        RECT 1781.170 260.000 1781.450 264.000 ;
        RECT 1781.280 244.110 1781.420 260.000 ;
        RECT 1781.220 243.790 1781.480 244.110 ;
        RECT 1786.280 243.790 1786.540 244.110 ;
        RECT 1786.340 24.130 1786.480 243.790 ;
        RECT 1786.280 23.810 1786.540 24.130 ;
        RECT 1864.020 23.810 1864.280 24.130 ;
        RECT 1864.080 2.400 1864.220 23.810 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 744.810 65.520 745.130 65.580 ;
        RECT 890.170 65.520 890.490 65.580 ;
        RECT 744.810 65.380 890.490 65.520 ;
        RECT 744.810 65.320 745.130 65.380 ;
        RECT 890.170 65.320 890.490 65.380 ;
        RECT 740.210 17.580 740.530 17.640 ;
        RECT 744.810 17.580 745.130 17.640 ;
        RECT 740.210 17.440 745.130 17.580 ;
        RECT 740.210 17.380 740.530 17.440 ;
        RECT 744.810 17.380 745.130 17.440 ;
      LAYER via ;
        RECT 744.840 65.320 745.100 65.580 ;
        RECT 890.200 65.320 890.460 65.580 ;
        RECT 740.240 17.380 740.500 17.640 ;
        RECT 744.840 17.380 745.100 17.640 ;
      LAYER met2 ;
        RECT 894.290 260.170 894.570 264.000 ;
        RECT 890.260 260.030 894.570 260.170 ;
        RECT 890.260 65.610 890.400 260.030 ;
        RECT 894.290 260.000 894.570 260.030 ;
        RECT 744.840 65.290 745.100 65.610 ;
        RECT 890.200 65.290 890.460 65.610 ;
        RECT 744.900 17.670 745.040 65.290 ;
        RECT 740.240 17.350 740.500 17.670 ;
        RECT 744.840 17.350 745.100 17.670 ;
        RECT 740.300 2.400 740.440 17.350 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1795.450 244.020 1795.770 244.080 ;
        RECT 1800.050 244.020 1800.370 244.080 ;
        RECT 1795.450 243.880 1800.370 244.020 ;
        RECT 1795.450 243.820 1795.770 243.880 ;
        RECT 1800.050 243.820 1800.370 243.880 ;
        RECT 1800.050 30.840 1800.370 30.900 ;
        RECT 1881.930 30.840 1882.250 30.900 ;
        RECT 1800.050 30.700 1882.250 30.840 ;
        RECT 1800.050 30.640 1800.370 30.700 ;
        RECT 1881.930 30.640 1882.250 30.700 ;
      LAYER via ;
        RECT 1795.480 243.820 1795.740 244.080 ;
        RECT 1800.080 243.820 1800.340 244.080 ;
        RECT 1800.080 30.640 1800.340 30.900 ;
        RECT 1881.960 30.640 1882.220 30.900 ;
      LAYER met2 ;
        RECT 1795.430 260.000 1795.710 264.000 ;
        RECT 1795.540 244.110 1795.680 260.000 ;
        RECT 1795.480 243.790 1795.740 244.110 ;
        RECT 1800.080 243.790 1800.340 244.110 ;
        RECT 1800.140 30.930 1800.280 243.790 ;
        RECT 1800.080 30.610 1800.340 30.930 ;
        RECT 1881.960 30.610 1882.220 30.930 ;
        RECT 1882.020 2.400 1882.160 30.610 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1809.710 244.020 1810.030 244.080 ;
        RECT 1813.850 244.020 1814.170 244.080 ;
        RECT 1809.710 243.880 1814.170 244.020 ;
        RECT 1809.710 243.820 1810.030 243.880 ;
        RECT 1813.850 243.820 1814.170 243.880 ;
        RECT 1813.850 37.980 1814.170 38.040 ;
        RECT 1899.870 37.980 1900.190 38.040 ;
        RECT 1813.850 37.840 1900.190 37.980 ;
        RECT 1813.850 37.780 1814.170 37.840 ;
        RECT 1899.870 37.780 1900.190 37.840 ;
      LAYER via ;
        RECT 1809.740 243.820 1810.000 244.080 ;
        RECT 1813.880 243.820 1814.140 244.080 ;
        RECT 1813.880 37.780 1814.140 38.040 ;
        RECT 1899.900 37.780 1900.160 38.040 ;
      LAYER met2 ;
        RECT 1809.690 260.000 1809.970 264.000 ;
        RECT 1809.800 244.110 1809.940 260.000 ;
        RECT 1809.740 243.790 1810.000 244.110 ;
        RECT 1813.880 243.790 1814.140 244.110 ;
        RECT 1813.940 38.070 1814.080 243.790 ;
        RECT 1813.880 37.750 1814.140 38.070 ;
        RECT 1899.900 37.750 1900.160 38.070 ;
        RECT 1899.960 2.400 1900.100 37.750 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1823.510 242.660 1823.830 242.720 ;
        RECT 1866.290 242.660 1866.610 242.720 ;
        RECT 1823.510 242.520 1866.610 242.660 ;
        RECT 1823.510 242.460 1823.830 242.520 ;
        RECT 1866.290 242.460 1866.610 242.520 ;
        RECT 1866.290 24.380 1866.610 24.440 ;
        RECT 1916.890 24.380 1917.210 24.440 ;
        RECT 1866.290 24.240 1917.210 24.380 ;
        RECT 1866.290 24.180 1866.610 24.240 ;
        RECT 1916.890 24.180 1917.210 24.240 ;
      LAYER via ;
        RECT 1823.540 242.460 1823.800 242.720 ;
        RECT 1866.320 242.460 1866.580 242.720 ;
        RECT 1866.320 24.180 1866.580 24.440 ;
        RECT 1916.920 24.180 1917.180 24.440 ;
      LAYER met2 ;
        RECT 1823.490 260.000 1823.770 264.000 ;
        RECT 1823.600 242.750 1823.740 260.000 ;
        RECT 1823.540 242.430 1823.800 242.750 ;
        RECT 1866.320 242.430 1866.580 242.750 ;
        RECT 1866.380 24.470 1866.520 242.430 ;
        RECT 1866.320 24.150 1866.580 24.470 ;
        RECT 1916.920 24.150 1917.180 24.470 ;
        RECT 1916.980 18.090 1917.120 24.150 ;
        RECT 1916.980 17.950 1918.040 18.090 ;
        RECT 1917.900 2.400 1918.040 17.950 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1837.770 244.020 1838.090 244.080 ;
        RECT 1841.910 244.020 1842.230 244.080 ;
        RECT 1837.770 243.880 1842.230 244.020 ;
        RECT 1837.770 243.820 1838.090 243.880 ;
        RECT 1841.910 243.820 1842.230 243.880 ;
        RECT 1841.910 113.800 1842.230 113.860 ;
        RECT 1932.070 113.800 1932.390 113.860 ;
        RECT 1841.910 113.660 1932.390 113.800 ;
        RECT 1841.910 113.600 1842.230 113.660 ;
        RECT 1932.070 113.600 1932.390 113.660 ;
        RECT 1932.070 2.960 1932.390 3.020 ;
        RECT 1935.290 2.960 1935.610 3.020 ;
        RECT 1932.070 2.820 1935.610 2.960 ;
        RECT 1932.070 2.760 1932.390 2.820 ;
        RECT 1935.290 2.760 1935.610 2.820 ;
      LAYER via ;
        RECT 1837.800 243.820 1838.060 244.080 ;
        RECT 1841.940 243.820 1842.200 244.080 ;
        RECT 1841.940 113.600 1842.200 113.860 ;
        RECT 1932.100 113.600 1932.360 113.860 ;
        RECT 1932.100 2.760 1932.360 3.020 ;
        RECT 1935.320 2.760 1935.580 3.020 ;
      LAYER met2 ;
        RECT 1837.750 260.000 1838.030 264.000 ;
        RECT 1837.860 244.110 1838.000 260.000 ;
        RECT 1837.800 243.790 1838.060 244.110 ;
        RECT 1841.940 243.790 1842.200 244.110 ;
        RECT 1842.000 113.890 1842.140 243.790 ;
        RECT 1841.940 113.570 1842.200 113.890 ;
        RECT 1932.100 113.570 1932.360 113.890 ;
        RECT 1932.160 3.050 1932.300 113.570 ;
        RECT 1932.100 2.730 1932.360 3.050 ;
        RECT 1935.320 2.730 1935.580 3.050 ;
        RECT 1935.380 2.400 1935.520 2.730 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1851.570 244.020 1851.890 244.080 ;
        RECT 1855.710 244.020 1856.030 244.080 ;
        RECT 1851.570 243.880 1856.030 244.020 ;
        RECT 1851.570 243.820 1851.890 243.880 ;
        RECT 1855.710 243.820 1856.030 243.880 ;
        RECT 1855.710 44.780 1856.030 44.840 ;
        RECT 1953.230 44.780 1953.550 44.840 ;
        RECT 1855.710 44.640 1953.550 44.780 ;
        RECT 1855.710 44.580 1856.030 44.640 ;
        RECT 1953.230 44.580 1953.550 44.640 ;
      LAYER via ;
        RECT 1851.600 243.820 1851.860 244.080 ;
        RECT 1855.740 243.820 1856.000 244.080 ;
        RECT 1855.740 44.580 1856.000 44.840 ;
        RECT 1953.260 44.580 1953.520 44.840 ;
      LAYER met2 ;
        RECT 1851.550 260.000 1851.830 264.000 ;
        RECT 1851.660 244.110 1851.800 260.000 ;
        RECT 1851.600 243.790 1851.860 244.110 ;
        RECT 1855.740 243.790 1856.000 244.110 ;
        RECT 1855.800 44.870 1855.940 243.790 ;
        RECT 1855.740 44.550 1856.000 44.870 ;
        RECT 1953.260 44.550 1953.520 44.870 ;
        RECT 1953.320 2.400 1953.460 44.550 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1865.830 245.040 1866.150 245.100 ;
        RECT 1955.990 245.040 1956.310 245.100 ;
        RECT 1865.830 244.900 1956.310 245.040 ;
        RECT 1865.830 244.840 1866.150 244.900 ;
        RECT 1955.990 244.840 1956.310 244.900 ;
        RECT 1955.990 23.360 1956.310 23.420 ;
        RECT 1971.170 23.360 1971.490 23.420 ;
        RECT 1955.990 23.220 1971.490 23.360 ;
        RECT 1955.990 23.160 1956.310 23.220 ;
        RECT 1971.170 23.160 1971.490 23.220 ;
      LAYER via ;
        RECT 1865.860 244.840 1866.120 245.100 ;
        RECT 1956.020 244.840 1956.280 245.100 ;
        RECT 1956.020 23.160 1956.280 23.420 ;
        RECT 1971.200 23.160 1971.460 23.420 ;
      LAYER met2 ;
        RECT 1865.810 260.000 1866.090 264.000 ;
        RECT 1865.920 245.130 1866.060 260.000 ;
        RECT 1865.860 244.810 1866.120 245.130 ;
        RECT 1956.020 244.810 1956.280 245.130 ;
        RECT 1956.080 23.450 1956.220 244.810 ;
        RECT 1956.020 23.130 1956.280 23.450 ;
        RECT 1971.200 23.130 1971.460 23.450 ;
        RECT 1971.260 2.400 1971.400 23.130 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1883.310 30.840 1883.630 30.900 ;
        RECT 1989.110 30.840 1989.430 30.900 ;
        RECT 1883.310 30.700 1989.430 30.840 ;
        RECT 1883.310 30.640 1883.630 30.700 ;
        RECT 1989.110 30.640 1989.430 30.700 ;
      LAYER via ;
        RECT 1883.340 30.640 1883.600 30.900 ;
        RECT 1989.140 30.640 1989.400 30.900 ;
      LAYER met2 ;
        RECT 1880.070 260.170 1880.350 264.000 ;
        RECT 1880.070 260.030 1883.540 260.170 ;
        RECT 1880.070 260.000 1880.350 260.030 ;
        RECT 1883.400 30.930 1883.540 260.030 ;
        RECT 1883.340 30.610 1883.600 30.930 ;
        RECT 1989.140 30.610 1989.400 30.930 ;
        RECT 1989.200 2.400 1989.340 30.610 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1893.890 243.680 1894.210 243.740 ;
        RECT 1907.690 243.680 1908.010 243.740 ;
        RECT 1893.890 243.540 1908.010 243.680 ;
        RECT 1893.890 243.480 1894.210 243.540 ;
        RECT 1907.690 243.480 1908.010 243.540 ;
        RECT 1907.690 24.040 1908.010 24.100 ;
        RECT 2006.590 24.040 2006.910 24.100 ;
        RECT 1907.690 23.900 2006.910 24.040 ;
        RECT 1907.690 23.840 1908.010 23.900 ;
        RECT 2006.590 23.840 2006.910 23.900 ;
      LAYER via ;
        RECT 1893.920 243.480 1894.180 243.740 ;
        RECT 1907.720 243.480 1907.980 243.740 ;
        RECT 1907.720 23.840 1907.980 24.100 ;
        RECT 2006.620 23.840 2006.880 24.100 ;
      LAYER met2 ;
        RECT 1893.870 260.000 1894.150 264.000 ;
        RECT 1893.980 243.770 1894.120 260.000 ;
        RECT 1893.920 243.450 1894.180 243.770 ;
        RECT 1907.720 243.450 1907.980 243.770 ;
        RECT 1907.780 24.130 1907.920 243.450 ;
        RECT 1907.720 23.810 1907.980 24.130 ;
        RECT 2006.620 23.810 2006.880 24.130 ;
        RECT 2006.680 2.400 2006.820 23.810 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1910.910 38.320 1911.230 38.380 ;
        RECT 2024.530 38.320 2024.850 38.380 ;
        RECT 1910.910 38.180 2024.850 38.320 ;
        RECT 1910.910 38.120 1911.230 38.180 ;
        RECT 2024.530 38.120 2024.850 38.180 ;
      LAYER via ;
        RECT 1910.940 38.120 1911.200 38.380 ;
        RECT 2024.560 38.120 2024.820 38.380 ;
      LAYER met2 ;
        RECT 1908.130 260.170 1908.410 264.000 ;
        RECT 1908.130 260.030 1911.140 260.170 ;
        RECT 1908.130 260.000 1908.410 260.030 ;
        RECT 1911.000 38.410 1911.140 260.030 ;
        RECT 1910.940 38.090 1911.200 38.410 ;
        RECT 2024.560 38.090 2024.820 38.410 ;
        RECT 2024.620 2.400 2024.760 38.090 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.710 51.580 1925.030 51.640 ;
        RECT 2042.930 51.580 2043.250 51.640 ;
        RECT 1924.710 51.440 2043.250 51.580 ;
        RECT 1924.710 51.380 1925.030 51.440 ;
        RECT 2042.930 51.380 2043.250 51.440 ;
      LAYER via ;
        RECT 1924.740 51.380 1925.000 51.640 ;
        RECT 2042.960 51.380 2043.220 51.640 ;
      LAYER met2 ;
        RECT 1922.390 260.170 1922.670 264.000 ;
        RECT 1922.390 260.030 1924.940 260.170 ;
        RECT 1922.390 260.000 1922.670 260.030 ;
        RECT 1924.800 51.670 1924.940 260.030 ;
        RECT 1924.740 51.350 1925.000 51.670 ;
        RECT 2042.960 51.350 2043.220 51.670 ;
        RECT 2043.020 17.410 2043.160 51.350 ;
        RECT 2042.560 17.270 2043.160 17.410 ;
        RECT 2042.560 2.400 2042.700 17.270 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.610 72.320 758.930 72.380 ;
        RECT 903.970 72.320 904.290 72.380 ;
        RECT 758.610 72.180 904.290 72.320 ;
        RECT 758.610 72.120 758.930 72.180 ;
        RECT 903.970 72.120 904.290 72.180 ;
        RECT 757.690 2.960 758.010 3.020 ;
        RECT 758.610 2.960 758.930 3.020 ;
        RECT 757.690 2.820 758.930 2.960 ;
        RECT 757.690 2.760 758.010 2.820 ;
        RECT 758.610 2.760 758.930 2.820 ;
      LAYER via ;
        RECT 758.640 72.120 758.900 72.380 ;
        RECT 904.000 72.120 904.260 72.380 ;
        RECT 757.720 2.760 757.980 3.020 ;
        RECT 758.640 2.760 758.900 3.020 ;
      LAYER met2 ;
        RECT 908.090 260.170 908.370 264.000 ;
        RECT 904.060 260.030 908.370 260.170 ;
        RECT 904.060 72.410 904.200 260.030 ;
        RECT 908.090 260.000 908.370 260.030 ;
        RECT 758.640 72.090 758.900 72.410 ;
        RECT 904.000 72.090 904.260 72.410 ;
        RECT 758.700 3.050 758.840 72.090 ;
        RECT 757.720 2.730 757.980 3.050 ;
        RECT 758.640 2.730 758.900 3.050 ;
        RECT 757.780 2.400 757.920 2.730 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 58.720 1938.830 58.780 ;
        RECT 2056.270 58.720 2056.590 58.780 ;
        RECT 1938.510 58.580 2056.590 58.720 ;
        RECT 1938.510 58.520 1938.830 58.580 ;
        RECT 2056.270 58.520 2056.590 58.580 ;
      LAYER via ;
        RECT 1938.540 58.520 1938.800 58.780 ;
        RECT 2056.300 58.520 2056.560 58.780 ;
      LAYER met2 ;
        RECT 1936.190 260.170 1936.470 264.000 ;
        RECT 1936.190 260.030 1938.740 260.170 ;
        RECT 1936.190 260.000 1936.470 260.030 ;
        RECT 1938.600 58.810 1938.740 260.030 ;
        RECT 1938.540 58.490 1938.800 58.810 ;
        RECT 2056.300 58.490 2056.560 58.810 ;
        RECT 2056.360 16.730 2056.500 58.490 ;
        RECT 2056.360 16.590 2060.640 16.730 ;
        RECT 2060.500 2.400 2060.640 16.590 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1950.470 243.680 1950.790 243.740 ;
        RECT 1956.450 243.680 1956.770 243.740 ;
        RECT 1950.470 243.540 1956.770 243.680 ;
        RECT 1950.470 243.480 1950.790 243.540 ;
        RECT 1956.450 243.480 1956.770 243.540 ;
        RECT 1956.450 44.780 1956.770 44.840 ;
        RECT 2078.350 44.780 2078.670 44.840 ;
        RECT 1956.450 44.640 2078.670 44.780 ;
        RECT 1956.450 44.580 1956.770 44.640 ;
        RECT 2078.350 44.580 2078.670 44.640 ;
      LAYER via ;
        RECT 1950.500 243.480 1950.760 243.740 ;
        RECT 1956.480 243.480 1956.740 243.740 ;
        RECT 1956.480 44.580 1956.740 44.840 ;
        RECT 2078.380 44.580 2078.640 44.840 ;
      LAYER met2 ;
        RECT 1950.450 260.000 1950.730 264.000 ;
        RECT 1950.560 243.770 1950.700 260.000 ;
        RECT 1950.500 243.450 1950.760 243.770 ;
        RECT 1956.480 243.450 1956.740 243.770 ;
        RECT 1956.540 44.870 1956.680 243.450 ;
        RECT 1956.480 44.550 1956.740 44.870 ;
        RECT 2078.380 44.550 2078.640 44.870 ;
        RECT 2078.440 2.400 2078.580 44.550 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1964.270 248.100 1964.590 248.160 ;
        RECT 1969.790 248.100 1970.110 248.160 ;
        RECT 1964.270 247.960 1970.110 248.100 ;
        RECT 1964.270 247.900 1964.590 247.960 ;
        RECT 1969.790 247.900 1970.110 247.960 ;
        RECT 1969.790 24.380 1970.110 24.440 ;
        RECT 2095.830 24.380 2096.150 24.440 ;
        RECT 1969.790 24.240 2096.150 24.380 ;
        RECT 1969.790 24.180 1970.110 24.240 ;
        RECT 2095.830 24.180 2096.150 24.240 ;
      LAYER via ;
        RECT 1964.300 247.900 1964.560 248.160 ;
        RECT 1969.820 247.900 1970.080 248.160 ;
        RECT 1969.820 24.180 1970.080 24.440 ;
        RECT 2095.860 24.180 2096.120 24.440 ;
      LAYER met2 ;
        RECT 1964.250 260.000 1964.530 264.000 ;
        RECT 1964.360 248.190 1964.500 260.000 ;
        RECT 1964.300 247.870 1964.560 248.190 ;
        RECT 1969.820 247.870 1970.080 248.190 ;
        RECT 1969.880 24.470 1970.020 247.870 ;
        RECT 1969.820 24.150 1970.080 24.470 ;
        RECT 2095.860 24.150 2096.120 24.470 ;
        RECT 2095.920 2.400 2096.060 24.150 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.450 65.860 1979.770 65.920 ;
        RECT 2111.470 65.860 2111.790 65.920 ;
        RECT 1979.450 65.720 2111.790 65.860 ;
        RECT 1979.450 65.660 1979.770 65.720 ;
        RECT 2111.470 65.660 2111.790 65.720 ;
      LAYER via ;
        RECT 1979.480 65.660 1979.740 65.920 ;
        RECT 2111.500 65.660 2111.760 65.920 ;
      LAYER met2 ;
        RECT 1978.510 260.170 1978.790 264.000 ;
        RECT 1978.510 260.030 1979.680 260.170 ;
        RECT 1978.510 260.000 1978.790 260.030 ;
        RECT 1979.540 65.950 1979.680 260.030 ;
        RECT 1979.480 65.630 1979.740 65.950 ;
        RECT 2111.500 65.630 2111.760 65.950 ;
        RECT 2111.560 16.730 2111.700 65.630 ;
        RECT 2111.560 16.590 2114.000 16.730 ;
        RECT 2113.860 2.400 2114.000 16.590 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.250 30.840 1993.570 30.900 ;
        RECT 2131.250 30.840 2131.570 30.900 ;
        RECT 1993.250 30.700 2131.570 30.840 ;
        RECT 1993.250 30.640 1993.570 30.700 ;
        RECT 2131.250 30.640 2131.570 30.700 ;
      LAYER via ;
        RECT 1993.280 30.640 1993.540 30.900 ;
        RECT 2131.280 30.640 2131.540 30.900 ;
      LAYER met2 ;
        RECT 1992.770 260.170 1993.050 264.000 ;
        RECT 1992.770 260.030 1993.480 260.170 ;
        RECT 1992.770 260.000 1993.050 260.030 ;
        RECT 1993.340 30.930 1993.480 260.030 ;
        RECT 1993.280 30.610 1993.540 30.930 ;
        RECT 2131.280 30.610 2131.540 30.930 ;
        RECT 2131.340 17.410 2131.480 30.610 ;
        RECT 2131.340 17.270 2131.940 17.410 ;
        RECT 2131.800 2.400 2131.940 17.270 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2006.590 243.680 2006.910 243.740 ;
        RECT 2011.190 243.680 2011.510 243.740 ;
        RECT 2006.590 243.540 2011.510 243.680 ;
        RECT 2006.590 243.480 2006.910 243.540 ;
        RECT 2011.190 243.480 2011.510 243.540 ;
        RECT 2011.190 37.980 2011.510 38.040 ;
        RECT 2149.650 37.980 2149.970 38.040 ;
        RECT 2011.190 37.840 2149.970 37.980 ;
        RECT 2011.190 37.780 2011.510 37.840 ;
        RECT 2149.650 37.780 2149.970 37.840 ;
      LAYER via ;
        RECT 2006.620 243.480 2006.880 243.740 ;
        RECT 2011.220 243.480 2011.480 243.740 ;
        RECT 2011.220 37.780 2011.480 38.040 ;
        RECT 2149.680 37.780 2149.940 38.040 ;
      LAYER met2 ;
        RECT 2006.570 260.000 2006.850 264.000 ;
        RECT 2006.680 243.770 2006.820 260.000 ;
        RECT 2006.620 243.450 2006.880 243.770 ;
        RECT 2011.220 243.450 2011.480 243.770 ;
        RECT 2011.280 38.070 2011.420 243.450 ;
        RECT 2011.220 37.750 2011.480 38.070 ;
        RECT 2149.680 37.750 2149.940 38.070 ;
        RECT 2149.740 2.400 2149.880 37.750 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2020.850 72.660 2021.170 72.720 ;
        RECT 2167.130 72.660 2167.450 72.720 ;
        RECT 2020.850 72.520 2167.450 72.660 ;
        RECT 2020.850 72.460 2021.170 72.520 ;
        RECT 2167.130 72.460 2167.450 72.520 ;
      LAYER via ;
        RECT 2020.880 72.460 2021.140 72.720 ;
        RECT 2167.160 72.460 2167.420 72.720 ;
      LAYER met2 ;
        RECT 2020.830 260.000 2021.110 264.000 ;
        RECT 2020.940 72.750 2021.080 260.000 ;
        RECT 2020.880 72.430 2021.140 72.750 ;
        RECT 2167.160 72.430 2167.420 72.750 ;
        RECT 2167.220 2.960 2167.360 72.430 ;
        RECT 2167.220 2.820 2167.820 2.960 ;
        RECT 2167.680 2.400 2167.820 2.820 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2035.110 24.040 2035.430 24.100 ;
        RECT 2185.070 24.040 2185.390 24.100 ;
        RECT 2035.110 23.900 2185.390 24.040 ;
        RECT 2035.110 23.840 2035.430 23.900 ;
        RECT 2185.070 23.840 2185.390 23.900 ;
      LAYER via ;
        RECT 2035.140 23.840 2035.400 24.100 ;
        RECT 2185.100 23.840 2185.360 24.100 ;
      LAYER met2 ;
        RECT 2034.630 260.170 2034.910 264.000 ;
        RECT 2034.630 260.030 2035.340 260.170 ;
        RECT 2034.630 260.000 2034.910 260.030 ;
        RECT 2035.200 24.130 2035.340 260.030 ;
        RECT 2035.140 23.810 2035.400 24.130 ;
        RECT 2185.100 23.810 2185.360 24.130 ;
        RECT 2185.160 2.400 2185.300 23.810 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.450 51.580 2048.770 51.640 ;
        RECT 2201.170 51.580 2201.490 51.640 ;
        RECT 2048.450 51.440 2201.490 51.580 ;
        RECT 2048.450 51.380 2048.770 51.440 ;
        RECT 2201.170 51.380 2201.490 51.440 ;
      LAYER via ;
        RECT 2048.480 51.380 2048.740 51.640 ;
        RECT 2201.200 51.380 2201.460 51.640 ;
      LAYER met2 ;
        RECT 2048.890 260.170 2049.170 264.000 ;
        RECT 2048.540 260.030 2049.170 260.170 ;
        RECT 2048.540 51.670 2048.680 260.030 ;
        RECT 2048.890 260.000 2049.170 260.030 ;
        RECT 2048.480 51.350 2048.740 51.670 ;
        RECT 2201.200 51.350 2201.460 51.670 ;
        RECT 2201.260 3.130 2201.400 51.350 ;
        RECT 2201.260 2.990 2202.780 3.130 ;
        RECT 2202.640 2.960 2202.780 2.990 ;
        RECT 2202.640 2.820 2203.240 2.960 ;
        RECT 2203.100 2.400 2203.240 2.820 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2063.170 244.020 2063.490 244.080 ;
        RECT 2069.610 244.020 2069.930 244.080 ;
        RECT 2063.170 243.880 2069.930 244.020 ;
        RECT 2063.170 243.820 2063.490 243.880 ;
        RECT 2069.610 243.820 2069.930 243.880 ;
        RECT 2069.610 58.720 2069.930 58.780 ;
        RECT 2215.430 58.720 2215.750 58.780 ;
        RECT 2069.610 58.580 2215.750 58.720 ;
        RECT 2069.610 58.520 2069.930 58.580 ;
        RECT 2215.430 58.520 2215.750 58.580 ;
        RECT 2215.430 2.960 2215.750 3.020 ;
        RECT 2220.950 2.960 2221.270 3.020 ;
        RECT 2215.430 2.820 2221.270 2.960 ;
        RECT 2215.430 2.760 2215.750 2.820 ;
        RECT 2220.950 2.760 2221.270 2.820 ;
      LAYER via ;
        RECT 2063.200 243.820 2063.460 244.080 ;
        RECT 2069.640 243.820 2069.900 244.080 ;
        RECT 2069.640 58.520 2069.900 58.780 ;
        RECT 2215.460 58.520 2215.720 58.780 ;
        RECT 2215.460 2.760 2215.720 3.020 ;
        RECT 2220.980 2.760 2221.240 3.020 ;
      LAYER met2 ;
        RECT 2063.150 260.000 2063.430 264.000 ;
        RECT 2063.260 244.110 2063.400 260.000 ;
        RECT 2063.200 243.790 2063.460 244.110 ;
        RECT 2069.640 243.790 2069.900 244.110 ;
        RECT 2069.700 58.810 2069.840 243.790 ;
        RECT 2069.640 58.490 2069.900 58.810 ;
        RECT 2215.460 58.490 2215.720 58.810 ;
        RECT 2215.520 3.050 2215.660 58.490 ;
        RECT 2215.460 2.730 2215.720 3.050 ;
        RECT 2220.980 2.730 2221.240 3.050 ;
        RECT 2221.040 2.400 2221.180 2.730 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 237.900 779.630 237.960 ;
        RECT 922.370 237.900 922.690 237.960 ;
        RECT 779.310 237.760 922.690 237.900 ;
        RECT 779.310 237.700 779.630 237.760 ;
        RECT 922.370 237.700 922.690 237.760 ;
        RECT 775.630 20.640 775.950 20.700 ;
        RECT 779.310 20.640 779.630 20.700 ;
        RECT 775.630 20.500 779.630 20.640 ;
        RECT 775.630 20.440 775.950 20.500 ;
        RECT 779.310 20.440 779.630 20.500 ;
      LAYER via ;
        RECT 779.340 237.700 779.600 237.960 ;
        RECT 922.400 237.700 922.660 237.960 ;
        RECT 775.660 20.440 775.920 20.700 ;
        RECT 779.340 20.440 779.600 20.700 ;
      LAYER met2 ;
        RECT 922.350 260.000 922.630 264.000 ;
        RECT 922.460 237.990 922.600 260.000 ;
        RECT 779.340 237.670 779.600 237.990 ;
        RECT 922.400 237.670 922.660 237.990 ;
        RECT 779.400 20.730 779.540 237.670 ;
        RECT 775.660 20.410 775.920 20.730 ;
        RECT 779.340 20.410 779.600 20.730 ;
        RECT 775.720 2.400 775.860 20.410 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.970 244.020 2077.290 244.080 ;
        RECT 2083.410 244.020 2083.730 244.080 ;
        RECT 2076.970 243.880 2083.730 244.020 ;
        RECT 2076.970 243.820 2077.290 243.880 ;
        RECT 2083.410 243.820 2083.730 243.880 ;
        RECT 2083.410 44.780 2083.730 44.840 ;
        RECT 2238.890 44.780 2239.210 44.840 ;
        RECT 2083.410 44.640 2239.210 44.780 ;
        RECT 2083.410 44.580 2083.730 44.640 ;
        RECT 2238.890 44.580 2239.210 44.640 ;
      LAYER via ;
        RECT 2077.000 243.820 2077.260 244.080 ;
        RECT 2083.440 243.820 2083.700 244.080 ;
        RECT 2083.440 44.580 2083.700 44.840 ;
        RECT 2238.920 44.580 2239.180 44.840 ;
      LAYER met2 ;
        RECT 2076.950 260.000 2077.230 264.000 ;
        RECT 2077.060 244.110 2077.200 260.000 ;
        RECT 2077.000 243.790 2077.260 244.110 ;
        RECT 2083.440 243.790 2083.700 244.110 ;
        RECT 2083.500 44.870 2083.640 243.790 ;
        RECT 2083.440 44.550 2083.700 44.870 ;
        RECT 2238.920 44.550 2239.180 44.870 ;
        RECT 2238.980 2.400 2239.120 44.550 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2091.230 242.660 2091.550 242.720 ;
        RECT 2100.890 242.660 2101.210 242.720 ;
        RECT 2091.230 242.520 2101.210 242.660 ;
        RECT 2091.230 242.460 2091.550 242.520 ;
        RECT 2100.890 242.460 2101.210 242.520 ;
        RECT 2100.890 79.460 2101.210 79.520 ;
        RECT 2256.830 79.460 2257.150 79.520 ;
        RECT 2100.890 79.320 2257.150 79.460 ;
        RECT 2100.890 79.260 2101.210 79.320 ;
        RECT 2256.830 79.260 2257.150 79.320 ;
      LAYER via ;
        RECT 2091.260 242.460 2091.520 242.720 ;
        RECT 2100.920 242.460 2101.180 242.720 ;
        RECT 2100.920 79.260 2101.180 79.520 ;
        RECT 2256.860 79.260 2257.120 79.520 ;
      LAYER met2 ;
        RECT 2091.210 260.000 2091.490 264.000 ;
        RECT 2091.320 242.750 2091.460 260.000 ;
        RECT 2091.260 242.430 2091.520 242.750 ;
        RECT 2100.920 242.430 2101.180 242.750 ;
        RECT 2100.980 79.550 2101.120 242.430 ;
        RECT 2100.920 79.230 2101.180 79.550 ;
        RECT 2256.860 79.230 2257.120 79.550 ;
        RECT 2256.920 17.410 2257.060 79.230 ;
        RECT 2256.460 17.270 2257.060 17.410 ;
        RECT 2256.460 2.400 2256.600 17.270 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2105.030 244.020 2105.350 244.080 ;
        RECT 2111.010 244.020 2111.330 244.080 ;
        RECT 2105.030 243.880 2111.330 244.020 ;
        RECT 2105.030 243.820 2105.350 243.880 ;
        RECT 2111.010 243.820 2111.330 243.880 ;
        RECT 2111.010 65.520 2111.330 65.580 ;
        RECT 2270.170 65.520 2270.490 65.580 ;
        RECT 2111.010 65.380 2270.490 65.520 ;
        RECT 2111.010 65.320 2111.330 65.380 ;
        RECT 2270.170 65.320 2270.490 65.380 ;
      LAYER via ;
        RECT 2105.060 243.820 2105.320 244.080 ;
        RECT 2111.040 243.820 2111.300 244.080 ;
        RECT 2111.040 65.320 2111.300 65.580 ;
        RECT 2270.200 65.320 2270.460 65.580 ;
      LAYER met2 ;
        RECT 2105.010 260.000 2105.290 264.000 ;
        RECT 2105.120 244.110 2105.260 260.000 ;
        RECT 2105.060 243.790 2105.320 244.110 ;
        RECT 2111.040 243.790 2111.300 244.110 ;
        RECT 2111.100 65.610 2111.240 243.790 ;
        RECT 2111.040 65.290 2111.300 65.610 ;
        RECT 2270.200 65.290 2270.460 65.610 ;
        RECT 2270.260 16.730 2270.400 65.290 ;
        RECT 2270.260 16.590 2274.540 16.730 ;
        RECT 2274.400 2.400 2274.540 16.590 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2119.290 244.020 2119.610 244.080 ;
        RECT 2124.350 244.020 2124.670 244.080 ;
        RECT 2119.290 243.880 2124.670 244.020 ;
        RECT 2119.290 243.820 2119.610 243.880 ;
        RECT 2124.350 243.820 2124.670 243.880 ;
        RECT 2124.350 86.600 2124.670 86.660 ;
        RECT 2290.870 86.600 2291.190 86.660 ;
        RECT 2124.350 86.460 2291.190 86.600 ;
        RECT 2124.350 86.400 2124.670 86.460 ;
        RECT 2290.870 86.400 2291.190 86.460 ;
      LAYER via ;
        RECT 2119.320 243.820 2119.580 244.080 ;
        RECT 2124.380 243.820 2124.640 244.080 ;
        RECT 2124.380 86.400 2124.640 86.660 ;
        RECT 2290.900 86.400 2291.160 86.660 ;
      LAYER met2 ;
        RECT 2119.270 260.000 2119.550 264.000 ;
        RECT 2119.380 244.110 2119.520 260.000 ;
        RECT 2119.320 243.790 2119.580 244.110 ;
        RECT 2124.380 243.790 2124.640 244.110 ;
        RECT 2124.440 86.690 2124.580 243.790 ;
        RECT 2124.380 86.370 2124.640 86.690 ;
        RECT 2290.900 86.370 2291.160 86.690 ;
        RECT 2290.960 16.730 2291.100 86.370 ;
        RECT 2290.960 16.590 2292.480 16.730 ;
        RECT 2292.340 2.400 2292.480 16.590 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2190.665 96.645 2190.835 144.755 ;
      LAYER mcon ;
        RECT 2190.665 144.585 2190.835 144.755 ;
      LAYER met1 ;
        RECT 2133.550 245.720 2133.870 245.780 ;
        RECT 2190.590 245.720 2190.910 245.780 ;
        RECT 2133.550 245.580 2190.910 245.720 ;
        RECT 2133.550 245.520 2133.870 245.580 ;
        RECT 2190.590 245.520 2190.910 245.580 ;
        RECT 2190.590 144.740 2190.910 144.800 ;
        RECT 2190.395 144.600 2190.910 144.740 ;
        RECT 2190.590 144.540 2190.910 144.600 ;
        RECT 2190.605 96.800 2190.895 96.845 ;
        RECT 2191.510 96.800 2191.830 96.860 ;
        RECT 2190.605 96.660 2191.830 96.800 ;
        RECT 2190.605 96.615 2190.895 96.660 ;
        RECT 2191.510 96.600 2191.830 96.660 ;
        RECT 2191.510 24.040 2191.830 24.100 ;
        RECT 2310.190 24.040 2310.510 24.100 ;
        RECT 2191.510 23.900 2310.510 24.040 ;
        RECT 2191.510 23.840 2191.830 23.900 ;
        RECT 2310.190 23.840 2310.510 23.900 ;
      LAYER via ;
        RECT 2133.580 245.520 2133.840 245.780 ;
        RECT 2190.620 245.520 2190.880 245.780 ;
        RECT 2190.620 144.540 2190.880 144.800 ;
        RECT 2191.540 96.600 2191.800 96.860 ;
        RECT 2191.540 23.840 2191.800 24.100 ;
        RECT 2310.220 23.840 2310.480 24.100 ;
      LAYER met2 ;
        RECT 2133.530 260.000 2133.810 264.000 ;
        RECT 2133.640 245.810 2133.780 260.000 ;
        RECT 2133.580 245.490 2133.840 245.810 ;
        RECT 2190.620 245.490 2190.880 245.810 ;
        RECT 2190.680 144.830 2190.820 245.490 ;
        RECT 2190.620 144.510 2190.880 144.830 ;
        RECT 2191.540 96.570 2191.800 96.890 ;
        RECT 2191.600 24.130 2191.740 96.570 ;
        RECT 2191.540 23.810 2191.800 24.130 ;
        RECT 2310.220 23.810 2310.480 24.130 ;
        RECT 2310.280 2.400 2310.420 23.810 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2147.350 241.980 2147.670 242.040 ;
        RECT 2152.410 241.980 2152.730 242.040 ;
        RECT 2147.350 241.840 2152.730 241.980 ;
        RECT 2147.350 241.780 2147.670 241.840 ;
        RECT 2152.410 241.780 2152.730 241.840 ;
        RECT 2152.410 93.400 2152.730 93.460 ;
        RECT 2325.370 93.400 2325.690 93.460 ;
        RECT 2152.410 93.260 2325.690 93.400 ;
        RECT 2152.410 93.200 2152.730 93.260 ;
        RECT 2325.370 93.200 2325.690 93.260 ;
      LAYER via ;
        RECT 2147.380 241.780 2147.640 242.040 ;
        RECT 2152.440 241.780 2152.700 242.040 ;
        RECT 2152.440 93.200 2152.700 93.460 ;
        RECT 2325.400 93.200 2325.660 93.460 ;
      LAYER met2 ;
        RECT 2147.330 260.000 2147.610 264.000 ;
        RECT 2147.440 242.070 2147.580 260.000 ;
        RECT 2147.380 241.750 2147.640 242.070 ;
        RECT 2152.440 241.750 2152.700 242.070 ;
        RECT 2152.500 93.490 2152.640 241.750 ;
        RECT 2152.440 93.170 2152.700 93.490 ;
        RECT 2325.400 93.170 2325.660 93.490 ;
        RECT 2325.460 16.730 2325.600 93.170 ;
        RECT 2325.460 16.590 2328.360 16.730 ;
        RECT 2328.220 2.400 2328.360 16.590 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2161.610 244.020 2161.930 244.080 ;
        RECT 2169.890 244.020 2170.210 244.080 ;
        RECT 2161.610 243.880 2170.210 244.020 ;
        RECT 2161.610 243.820 2161.930 243.880 ;
        RECT 2169.890 243.820 2170.210 243.880 ;
        RECT 2169.890 99.860 2170.210 99.920 ;
        RECT 2339.630 99.860 2339.950 99.920 ;
        RECT 2169.890 99.720 2339.950 99.860 ;
        RECT 2169.890 99.660 2170.210 99.720 ;
        RECT 2339.630 99.660 2339.950 99.720 ;
        RECT 2339.630 17.580 2339.950 17.640 ;
        RECT 2345.610 17.580 2345.930 17.640 ;
        RECT 2339.630 17.440 2345.930 17.580 ;
        RECT 2339.630 17.380 2339.950 17.440 ;
        RECT 2345.610 17.380 2345.930 17.440 ;
      LAYER via ;
        RECT 2161.640 243.820 2161.900 244.080 ;
        RECT 2169.920 243.820 2170.180 244.080 ;
        RECT 2169.920 99.660 2170.180 99.920 ;
        RECT 2339.660 99.660 2339.920 99.920 ;
        RECT 2339.660 17.380 2339.920 17.640 ;
        RECT 2345.640 17.380 2345.900 17.640 ;
      LAYER met2 ;
        RECT 2161.590 260.000 2161.870 264.000 ;
        RECT 2161.700 244.110 2161.840 260.000 ;
        RECT 2161.640 243.790 2161.900 244.110 ;
        RECT 2169.920 243.790 2170.180 244.110 ;
        RECT 2169.980 99.950 2170.120 243.790 ;
        RECT 2169.920 99.630 2170.180 99.950 ;
        RECT 2339.660 99.630 2339.920 99.950 ;
        RECT 2339.720 17.670 2339.860 99.630 ;
        RECT 2339.660 17.350 2339.920 17.670 ;
        RECT 2345.640 17.350 2345.900 17.670 ;
        RECT 2345.700 2.400 2345.840 17.350 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2175.870 245.380 2176.190 245.440 ;
        RECT 2287.190 245.380 2287.510 245.440 ;
        RECT 2175.870 245.240 2287.510 245.380 ;
        RECT 2175.870 245.180 2176.190 245.240 ;
        RECT 2287.190 245.180 2287.510 245.240 ;
        RECT 2287.190 24.380 2287.510 24.440 ;
        RECT 2287.190 24.240 2311.340 24.380 ;
        RECT 2287.190 24.180 2287.510 24.240 ;
        RECT 2311.200 24.040 2311.340 24.240 ;
        RECT 2363.550 24.040 2363.870 24.100 ;
        RECT 2311.200 23.900 2363.870 24.040 ;
        RECT 2363.550 23.840 2363.870 23.900 ;
      LAYER via ;
        RECT 2175.900 245.180 2176.160 245.440 ;
        RECT 2287.220 245.180 2287.480 245.440 ;
        RECT 2287.220 24.180 2287.480 24.440 ;
        RECT 2363.580 23.840 2363.840 24.100 ;
      LAYER met2 ;
        RECT 2175.850 260.000 2176.130 264.000 ;
        RECT 2175.960 245.470 2176.100 260.000 ;
        RECT 2175.900 245.150 2176.160 245.470 ;
        RECT 2287.220 245.150 2287.480 245.470 ;
        RECT 2287.280 24.470 2287.420 245.150 ;
        RECT 2287.220 24.150 2287.480 24.470 ;
        RECT 2363.580 23.810 2363.840 24.130 ;
        RECT 2363.640 2.400 2363.780 23.810 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2189.670 244.020 2189.990 244.080 ;
        RECT 2193.810 244.020 2194.130 244.080 ;
        RECT 2189.670 243.880 2194.130 244.020 ;
        RECT 2189.670 243.820 2189.990 243.880 ;
        RECT 2193.810 243.820 2194.130 243.880 ;
        RECT 2193.810 107.340 2194.130 107.400 ;
        RECT 2380.570 107.340 2380.890 107.400 ;
        RECT 2193.810 107.200 2380.890 107.340 ;
        RECT 2193.810 107.140 2194.130 107.200 ;
        RECT 2380.570 107.140 2380.890 107.200 ;
      LAYER via ;
        RECT 2189.700 243.820 2189.960 244.080 ;
        RECT 2193.840 243.820 2194.100 244.080 ;
        RECT 2193.840 107.140 2194.100 107.400 ;
        RECT 2380.600 107.140 2380.860 107.400 ;
      LAYER met2 ;
        RECT 2189.650 260.000 2189.930 264.000 ;
        RECT 2189.760 244.110 2189.900 260.000 ;
        RECT 2189.700 243.790 2189.960 244.110 ;
        RECT 2193.840 243.790 2194.100 244.110 ;
        RECT 2193.900 107.430 2194.040 243.790 ;
        RECT 2193.840 107.110 2194.100 107.430 ;
        RECT 2380.600 107.110 2380.860 107.430 ;
        RECT 2380.660 3.130 2380.800 107.110 ;
        RECT 2380.660 2.990 2381.720 3.130 ;
        RECT 2381.580 2.400 2381.720 2.990 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2207.610 30.840 2207.930 30.900 ;
        RECT 2399.430 30.840 2399.750 30.900 ;
        RECT 2207.610 30.700 2399.750 30.840 ;
        RECT 2207.610 30.640 2207.930 30.700 ;
        RECT 2399.430 30.640 2399.750 30.700 ;
      LAYER via ;
        RECT 2207.640 30.640 2207.900 30.900 ;
        RECT 2399.460 30.640 2399.720 30.900 ;
      LAYER met2 ;
        RECT 2203.910 260.170 2204.190 264.000 ;
        RECT 2203.910 260.030 2207.840 260.170 ;
        RECT 2203.910 260.000 2204.190 260.030 ;
        RECT 2207.700 30.930 2207.840 260.030 ;
        RECT 2207.640 30.610 2207.900 30.930 ;
        RECT 2399.460 30.610 2399.720 30.930 ;
        RECT 2399.520 2.400 2399.660 30.610 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 799.550 79.460 799.870 79.520 ;
        RECT 932.030 79.460 932.350 79.520 ;
        RECT 799.550 79.320 932.350 79.460 ;
        RECT 799.550 79.260 799.870 79.320 ;
        RECT 932.030 79.260 932.350 79.320 ;
        RECT 793.570 20.640 793.890 20.700 ;
        RECT 799.550 20.640 799.870 20.700 ;
        RECT 793.570 20.500 799.870 20.640 ;
        RECT 793.570 20.440 793.890 20.500 ;
        RECT 799.550 20.440 799.870 20.500 ;
      LAYER via ;
        RECT 799.580 79.260 799.840 79.520 ;
        RECT 932.060 79.260 932.320 79.520 ;
        RECT 793.600 20.440 793.860 20.700 ;
        RECT 799.580 20.440 799.840 20.700 ;
      LAYER met2 ;
        RECT 936.610 260.170 936.890 264.000 ;
        RECT 932.120 260.030 936.890 260.170 ;
        RECT 932.120 79.550 932.260 260.030 ;
        RECT 936.610 260.000 936.890 260.030 ;
        RECT 799.580 79.230 799.840 79.550 ;
        RECT 932.060 79.230 932.320 79.550 ;
        RECT 799.640 20.730 799.780 79.230 ;
        RECT 793.600 20.410 793.860 20.730 ;
        RECT 799.580 20.410 799.840 20.730 ;
        RECT 793.660 2.400 793.800 20.410 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 810.590 244.020 810.910 244.080 ;
        RECT 814.270 244.020 814.590 244.080 ;
        RECT 810.590 243.880 814.590 244.020 ;
        RECT 810.590 243.820 810.910 243.880 ;
        RECT 814.270 243.820 814.590 243.880 ;
        RECT 641.310 86.260 641.630 86.320 ;
        RECT 810.590 86.260 810.910 86.320 ;
        RECT 641.310 86.120 810.910 86.260 ;
        RECT 641.310 86.060 641.630 86.120 ;
        RECT 810.590 86.060 810.910 86.120 ;
        RECT 639.010 17.580 639.330 17.640 ;
        RECT 641.310 17.580 641.630 17.640 ;
        RECT 639.010 17.440 641.630 17.580 ;
        RECT 639.010 17.380 639.330 17.440 ;
        RECT 641.310 17.380 641.630 17.440 ;
      LAYER via ;
        RECT 810.620 243.820 810.880 244.080 ;
        RECT 814.300 243.820 814.560 244.080 ;
        RECT 641.340 86.060 641.600 86.320 ;
        RECT 810.620 86.060 810.880 86.320 ;
        RECT 639.040 17.380 639.300 17.640 ;
        RECT 641.340 17.380 641.600 17.640 ;
      LAYER met2 ;
        RECT 814.250 260.000 814.530 264.000 ;
        RECT 814.360 244.110 814.500 260.000 ;
        RECT 810.620 243.790 810.880 244.110 ;
        RECT 814.300 243.790 814.560 244.110 ;
        RECT 810.680 86.350 810.820 243.790 ;
        RECT 641.340 86.030 641.600 86.350 ;
        RECT 810.620 86.030 810.880 86.350 ;
        RECT 641.400 17.670 641.540 86.030 ;
        RECT 639.040 17.350 639.300 17.670 ;
        RECT 641.340 17.350 641.600 17.670 ;
        RECT 639.100 2.400 639.240 17.350 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2222.790 244.020 2223.110 244.080 ;
        RECT 2227.850 244.020 2228.170 244.080 ;
        RECT 2222.790 243.880 2228.170 244.020 ;
        RECT 2222.790 243.820 2223.110 243.880 ;
        RECT 2227.850 243.820 2228.170 243.880 ;
        RECT 2227.850 114.140 2228.170 114.200 ;
        RECT 2421.970 114.140 2422.290 114.200 ;
        RECT 2227.850 114.000 2422.290 114.140 ;
        RECT 2227.850 113.940 2228.170 114.000 ;
        RECT 2421.970 113.940 2422.290 114.000 ;
      LAYER via ;
        RECT 2222.820 243.820 2223.080 244.080 ;
        RECT 2227.880 243.820 2228.140 244.080 ;
        RECT 2227.880 113.940 2228.140 114.200 ;
        RECT 2422.000 113.940 2422.260 114.200 ;
      LAYER met2 ;
        RECT 2222.770 260.000 2223.050 264.000 ;
        RECT 2222.880 244.110 2223.020 260.000 ;
        RECT 2222.820 243.790 2223.080 244.110 ;
        RECT 2227.880 243.790 2228.140 244.110 ;
        RECT 2227.940 114.230 2228.080 243.790 ;
        RECT 2227.880 113.910 2228.140 114.230 ;
        RECT 2422.000 113.910 2422.260 114.230 ;
        RECT 2422.060 16.730 2422.200 113.910 ;
        RECT 2422.060 16.590 2423.120 16.730 ;
        RECT 2422.980 2.400 2423.120 16.590 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2435.845 144.925 2436.015 193.035 ;
        RECT 2435.845 48.365 2436.015 96.475 ;
      LAYER mcon ;
        RECT 2435.845 192.865 2436.015 193.035 ;
        RECT 2435.845 96.305 2436.015 96.475 ;
      LAYER met1 ;
        RECT 2236.590 237.900 2236.910 237.960 ;
        RECT 2435.770 237.900 2436.090 237.960 ;
        RECT 2236.590 237.760 2436.090 237.900 ;
        RECT 2236.590 237.700 2236.910 237.760 ;
        RECT 2435.770 237.700 2436.090 237.760 ;
        RECT 2435.770 193.020 2436.090 193.080 ;
        RECT 2435.575 192.880 2436.090 193.020 ;
        RECT 2435.770 192.820 2436.090 192.880 ;
        RECT 2435.770 145.080 2436.090 145.140 ;
        RECT 2435.575 144.940 2436.090 145.080 ;
        RECT 2435.770 144.880 2436.090 144.940 ;
        RECT 2435.770 96.460 2436.090 96.520 ;
        RECT 2435.575 96.320 2436.090 96.460 ;
        RECT 2435.770 96.260 2436.090 96.320 ;
        RECT 2435.770 48.520 2436.090 48.580 ;
        RECT 2435.575 48.380 2436.090 48.520 ;
        RECT 2435.770 48.320 2436.090 48.380 ;
        RECT 2435.310 2.960 2435.630 3.020 ;
        RECT 2440.830 2.960 2441.150 3.020 ;
        RECT 2435.310 2.820 2441.150 2.960 ;
        RECT 2435.310 2.760 2435.630 2.820 ;
        RECT 2440.830 2.760 2441.150 2.820 ;
      LAYER via ;
        RECT 2236.620 237.700 2236.880 237.960 ;
        RECT 2435.800 237.700 2436.060 237.960 ;
        RECT 2435.800 192.820 2436.060 193.080 ;
        RECT 2435.800 144.880 2436.060 145.140 ;
        RECT 2435.800 96.260 2436.060 96.520 ;
        RECT 2435.800 48.320 2436.060 48.580 ;
        RECT 2435.340 2.760 2435.600 3.020 ;
        RECT 2440.860 2.760 2441.120 3.020 ;
      LAYER met2 ;
        RECT 2236.570 260.000 2236.850 264.000 ;
        RECT 2236.680 237.990 2236.820 260.000 ;
        RECT 2236.620 237.670 2236.880 237.990 ;
        RECT 2435.800 237.670 2436.060 237.990 ;
        RECT 2435.860 193.110 2436.000 237.670 ;
        RECT 2435.800 192.790 2436.060 193.110 ;
        RECT 2435.800 144.850 2436.060 145.170 ;
        RECT 2435.860 96.550 2436.000 144.850 ;
        RECT 2435.800 96.230 2436.060 96.550 ;
        RECT 2435.800 48.290 2436.060 48.610 ;
        RECT 2435.860 14.690 2436.000 48.290 ;
        RECT 2435.400 14.550 2436.000 14.690 ;
        RECT 2435.400 3.050 2435.540 14.550 ;
        RECT 2435.340 2.730 2435.600 3.050 ;
        RECT 2440.860 2.730 2441.120 3.050 ;
        RECT 2440.920 2.400 2441.060 2.730 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2250.850 248.440 2251.170 248.500 ;
        RECT 2259.590 248.440 2259.910 248.500 ;
        RECT 2250.850 248.300 2259.910 248.440 ;
        RECT 2250.850 248.240 2251.170 248.300 ;
        RECT 2259.590 248.240 2259.910 248.300 ;
        RECT 2259.590 120.600 2259.910 120.660 ;
        RECT 2456.470 120.600 2456.790 120.660 ;
        RECT 2259.590 120.460 2456.790 120.600 ;
        RECT 2259.590 120.400 2259.910 120.460 ;
        RECT 2456.470 120.400 2456.790 120.460 ;
        RECT 2456.010 2.960 2456.330 3.020 ;
        RECT 2458.770 2.960 2459.090 3.020 ;
        RECT 2456.010 2.820 2459.090 2.960 ;
        RECT 2456.010 2.760 2456.330 2.820 ;
        RECT 2458.770 2.760 2459.090 2.820 ;
      LAYER via ;
        RECT 2250.880 248.240 2251.140 248.500 ;
        RECT 2259.620 248.240 2259.880 248.500 ;
        RECT 2259.620 120.400 2259.880 120.660 ;
        RECT 2456.500 120.400 2456.760 120.660 ;
        RECT 2456.040 2.760 2456.300 3.020 ;
        RECT 2458.800 2.760 2459.060 3.020 ;
      LAYER met2 ;
        RECT 2250.830 260.000 2251.110 264.000 ;
        RECT 2250.940 248.530 2251.080 260.000 ;
        RECT 2250.880 248.210 2251.140 248.530 ;
        RECT 2259.620 248.210 2259.880 248.530 ;
        RECT 2259.680 120.690 2259.820 248.210 ;
        RECT 2259.620 120.370 2259.880 120.690 ;
        RECT 2456.500 120.370 2456.760 120.690 ;
        RECT 2456.560 14.690 2456.700 120.370 ;
        RECT 2456.100 14.550 2456.700 14.690 ;
        RECT 2456.100 3.050 2456.240 14.550 ;
        RECT 2456.040 2.730 2456.300 3.050 ;
        RECT 2458.800 2.730 2459.060 3.050 ;
        RECT 2458.860 2.400 2459.000 2.730 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2264.650 244.020 2264.970 244.080 ;
        RECT 2269.250 244.020 2269.570 244.080 ;
        RECT 2264.650 243.880 2269.570 244.020 ;
        RECT 2264.650 243.820 2264.970 243.880 ;
        RECT 2269.250 243.820 2269.570 243.880 ;
        RECT 2269.250 86.260 2269.570 86.320 ;
        RECT 2470.270 86.260 2470.590 86.320 ;
        RECT 2269.250 86.120 2470.590 86.260 ;
        RECT 2269.250 86.060 2269.570 86.120 ;
        RECT 2470.270 86.060 2470.590 86.120 ;
        RECT 2470.270 38.320 2470.590 38.380 ;
        RECT 2476.710 38.320 2477.030 38.380 ;
        RECT 2470.270 38.180 2477.030 38.320 ;
        RECT 2470.270 38.120 2470.590 38.180 ;
        RECT 2476.710 38.120 2477.030 38.180 ;
      LAYER via ;
        RECT 2264.680 243.820 2264.940 244.080 ;
        RECT 2269.280 243.820 2269.540 244.080 ;
        RECT 2269.280 86.060 2269.540 86.320 ;
        RECT 2470.300 86.060 2470.560 86.320 ;
        RECT 2470.300 38.120 2470.560 38.380 ;
        RECT 2476.740 38.120 2477.000 38.380 ;
      LAYER met2 ;
        RECT 2264.630 260.000 2264.910 264.000 ;
        RECT 2264.740 244.110 2264.880 260.000 ;
        RECT 2264.680 243.790 2264.940 244.110 ;
        RECT 2269.280 243.790 2269.540 244.110 ;
        RECT 2269.340 86.350 2269.480 243.790 ;
        RECT 2269.280 86.030 2269.540 86.350 ;
        RECT 2470.300 86.030 2470.560 86.350 ;
        RECT 2470.360 38.410 2470.500 86.030 ;
        RECT 2470.300 38.090 2470.560 38.410 ;
        RECT 2476.740 38.090 2477.000 38.410 ;
        RECT 2476.800 2.400 2476.940 38.090 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2278.910 231.100 2279.230 231.160 ;
        RECT 2490.970 231.100 2491.290 231.160 ;
        RECT 2278.910 230.960 2491.290 231.100 ;
        RECT 2278.910 230.900 2279.230 230.960 ;
        RECT 2490.970 230.900 2491.290 230.960 ;
      LAYER via ;
        RECT 2278.940 230.900 2279.200 231.160 ;
        RECT 2491.000 230.900 2491.260 231.160 ;
      LAYER met2 ;
        RECT 2278.890 260.000 2279.170 264.000 ;
        RECT 2279.000 231.190 2279.140 260.000 ;
        RECT 2278.940 230.870 2279.200 231.190 ;
        RECT 2491.000 230.870 2491.260 231.190 ;
        RECT 2491.060 16.730 2491.200 230.870 ;
        RECT 2491.060 16.590 2494.880 16.730 ;
        RECT 2494.740 2.400 2494.880 16.590 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2293.170 244.020 2293.490 244.080 ;
        RECT 2297.310 244.020 2297.630 244.080 ;
        RECT 2293.170 243.880 2297.630 244.020 ;
        RECT 2293.170 243.820 2293.490 243.880 ;
        RECT 2297.310 243.820 2297.630 243.880 ;
        RECT 2297.310 127.740 2297.630 127.800 ;
        RECT 2512.130 127.740 2512.450 127.800 ;
        RECT 2297.310 127.600 2512.450 127.740 ;
        RECT 2297.310 127.540 2297.630 127.600 ;
        RECT 2512.130 127.540 2512.450 127.600 ;
      LAYER via ;
        RECT 2293.200 243.820 2293.460 244.080 ;
        RECT 2297.340 243.820 2297.600 244.080 ;
        RECT 2297.340 127.540 2297.600 127.800 ;
        RECT 2512.160 127.540 2512.420 127.800 ;
      LAYER met2 ;
        RECT 2293.150 260.000 2293.430 264.000 ;
        RECT 2293.260 244.110 2293.400 260.000 ;
        RECT 2293.200 243.790 2293.460 244.110 ;
        RECT 2297.340 243.790 2297.600 244.110 ;
        RECT 2297.400 127.830 2297.540 243.790 ;
        RECT 2297.340 127.510 2297.600 127.830 ;
        RECT 2512.160 127.510 2512.420 127.830 ;
        RECT 2512.220 2.400 2512.360 127.510 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2306.970 243.680 2307.290 243.740 ;
        RECT 2321.690 243.680 2322.010 243.740 ;
        RECT 2306.970 243.540 2322.010 243.680 ;
        RECT 2306.970 243.480 2307.290 243.540 ;
        RECT 2321.690 243.480 2322.010 243.540 ;
        RECT 2321.690 134.540 2322.010 134.600 ;
        RECT 2525.470 134.540 2525.790 134.600 ;
        RECT 2321.690 134.400 2525.790 134.540 ;
        RECT 2321.690 134.340 2322.010 134.400 ;
        RECT 2525.470 134.340 2525.790 134.400 ;
      LAYER via ;
        RECT 2307.000 243.480 2307.260 243.740 ;
        RECT 2321.720 243.480 2321.980 243.740 ;
        RECT 2321.720 134.340 2321.980 134.600 ;
        RECT 2525.500 134.340 2525.760 134.600 ;
      LAYER met2 ;
        RECT 2306.950 260.000 2307.230 264.000 ;
        RECT 2307.060 243.770 2307.200 260.000 ;
        RECT 2307.000 243.450 2307.260 243.770 ;
        RECT 2321.720 243.450 2321.980 243.770 ;
        RECT 2321.780 134.630 2321.920 243.450 ;
        RECT 2321.720 134.310 2321.980 134.630 ;
        RECT 2525.500 134.310 2525.760 134.630 ;
        RECT 2525.560 16.730 2525.700 134.310 ;
        RECT 2525.560 16.590 2530.300 16.730 ;
        RECT 2530.160 2.400 2530.300 16.590 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2321.230 244.020 2321.550 244.080 ;
        RECT 2324.910 244.020 2325.230 244.080 ;
        RECT 2321.230 243.880 2325.230 244.020 ;
        RECT 2321.230 243.820 2321.550 243.880 ;
        RECT 2324.910 243.820 2325.230 243.880 ;
        RECT 2324.910 93.060 2325.230 93.120 ;
        RECT 2546.170 93.060 2546.490 93.120 ;
        RECT 2324.910 92.920 2546.490 93.060 ;
        RECT 2324.910 92.860 2325.230 92.920 ;
        RECT 2546.170 92.860 2546.490 92.920 ;
      LAYER via ;
        RECT 2321.260 243.820 2321.520 244.080 ;
        RECT 2324.940 243.820 2325.200 244.080 ;
        RECT 2324.940 92.860 2325.200 93.120 ;
        RECT 2546.200 92.860 2546.460 93.120 ;
      LAYER met2 ;
        RECT 2321.210 260.000 2321.490 264.000 ;
        RECT 2321.320 244.110 2321.460 260.000 ;
        RECT 2321.260 243.790 2321.520 244.110 ;
        RECT 2324.940 243.790 2325.200 244.110 ;
        RECT 2325.000 93.150 2325.140 243.790 ;
        RECT 2324.940 92.830 2325.200 93.150 ;
        RECT 2546.200 92.830 2546.460 93.150 ;
        RECT 2546.260 16.730 2546.400 92.830 ;
        RECT 2546.260 16.590 2548.240 16.730 ;
        RECT 2548.100 2.400 2548.240 16.590 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2335.030 244.020 2335.350 244.080 ;
        RECT 2338.710 244.020 2339.030 244.080 ;
        RECT 2335.030 243.880 2339.030 244.020 ;
        RECT 2335.030 243.820 2335.350 243.880 ;
        RECT 2338.710 243.820 2339.030 243.880 ;
        RECT 2338.710 44.780 2339.030 44.840 ;
        RECT 2565.950 44.780 2566.270 44.840 ;
        RECT 2338.710 44.640 2566.270 44.780 ;
        RECT 2338.710 44.580 2339.030 44.640 ;
        RECT 2565.950 44.580 2566.270 44.640 ;
      LAYER via ;
        RECT 2335.060 243.820 2335.320 244.080 ;
        RECT 2338.740 243.820 2339.000 244.080 ;
        RECT 2338.740 44.580 2339.000 44.840 ;
        RECT 2565.980 44.580 2566.240 44.840 ;
      LAYER met2 ;
        RECT 2335.010 260.000 2335.290 264.000 ;
        RECT 2335.120 244.110 2335.260 260.000 ;
        RECT 2335.060 243.790 2335.320 244.110 ;
        RECT 2338.740 243.790 2339.000 244.110 ;
        RECT 2338.800 44.870 2338.940 243.790 ;
        RECT 2338.740 44.550 2339.000 44.870 ;
        RECT 2565.980 44.550 2566.240 44.870 ;
        RECT 2566.040 2.400 2566.180 44.550 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2352.510 141.340 2352.830 141.400 ;
        RECT 2580.670 141.340 2580.990 141.400 ;
        RECT 2352.510 141.200 2580.990 141.340 ;
        RECT 2352.510 141.140 2352.830 141.200 ;
        RECT 2580.670 141.140 2580.990 141.200 ;
      LAYER via ;
        RECT 2352.540 141.140 2352.800 141.400 ;
        RECT 2580.700 141.140 2580.960 141.400 ;
      LAYER met2 ;
        RECT 2349.270 260.170 2349.550 264.000 ;
        RECT 2349.270 260.030 2352.740 260.170 ;
        RECT 2349.270 260.000 2349.550 260.030 ;
        RECT 2352.600 141.430 2352.740 260.030 ;
        RECT 2352.540 141.110 2352.800 141.430 ;
        RECT 2580.700 141.110 2580.960 141.430 ;
        RECT 2580.760 16.730 2580.900 141.110 ;
        RECT 2580.760 16.590 2584.120 16.730 ;
        RECT 2583.980 2.400 2584.120 16.590 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 820.710 86.260 821.030 86.320 ;
        RECT 952.270 86.260 952.590 86.320 ;
        RECT 820.710 86.120 952.590 86.260 ;
        RECT 820.710 86.060 821.030 86.120 ;
        RECT 952.270 86.060 952.590 86.120 ;
        RECT 817.490 20.640 817.810 20.700 ;
        RECT 820.710 20.640 821.030 20.700 ;
        RECT 817.490 20.500 821.030 20.640 ;
        RECT 817.490 20.440 817.810 20.500 ;
        RECT 820.710 20.440 821.030 20.500 ;
      LAYER via ;
        RECT 820.740 86.060 821.000 86.320 ;
        RECT 952.300 86.060 952.560 86.320 ;
        RECT 817.520 20.440 817.780 20.700 ;
        RECT 820.740 20.440 821.000 20.700 ;
      LAYER met2 ;
        RECT 955.010 260.170 955.290 264.000 ;
        RECT 952.360 260.030 955.290 260.170 ;
        RECT 952.360 86.350 952.500 260.030 ;
        RECT 955.010 260.000 955.290 260.030 ;
        RECT 820.740 86.030 821.000 86.350 ;
        RECT 952.300 86.030 952.560 86.350 ;
        RECT 820.800 20.730 820.940 86.030 ;
        RECT 817.520 20.410 817.780 20.730 ;
        RECT 820.740 20.410 821.000 20.730 ;
        RECT 817.580 2.400 817.720 20.410 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2363.550 243.680 2363.870 243.740 ;
        RECT 2376.890 243.680 2377.210 243.740 ;
        RECT 2363.550 243.540 2377.210 243.680 ;
        RECT 2363.550 243.480 2363.870 243.540 ;
        RECT 2376.890 243.480 2377.210 243.540 ;
        RECT 2376.890 99.860 2377.210 99.920 ;
        RECT 2601.830 99.860 2602.150 99.920 ;
        RECT 2376.890 99.720 2602.150 99.860 ;
        RECT 2376.890 99.660 2377.210 99.720 ;
        RECT 2601.830 99.660 2602.150 99.720 ;
      LAYER via ;
        RECT 2363.580 243.480 2363.840 243.740 ;
        RECT 2376.920 243.480 2377.180 243.740 ;
        RECT 2376.920 99.660 2377.180 99.920 ;
        RECT 2601.860 99.660 2602.120 99.920 ;
      LAYER met2 ;
        RECT 2363.530 260.000 2363.810 264.000 ;
        RECT 2363.640 243.770 2363.780 260.000 ;
        RECT 2363.580 243.450 2363.840 243.770 ;
        RECT 2376.920 243.450 2377.180 243.770 ;
        RECT 2376.980 99.950 2377.120 243.450 ;
        RECT 2376.920 99.630 2377.180 99.950 ;
        RECT 2601.860 99.630 2602.120 99.950 ;
        RECT 2601.920 17.410 2602.060 99.630 ;
        RECT 2601.460 17.270 2602.060 17.410 ;
        RECT 2601.460 2.400 2601.600 17.270 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2380.110 107.000 2380.430 107.060 ;
        RECT 2615.170 107.000 2615.490 107.060 ;
        RECT 2380.110 106.860 2615.490 107.000 ;
        RECT 2380.110 106.800 2380.430 106.860 ;
        RECT 2615.170 106.800 2615.490 106.860 ;
      LAYER via ;
        RECT 2380.140 106.800 2380.400 107.060 ;
        RECT 2615.200 106.800 2615.460 107.060 ;
      LAYER met2 ;
        RECT 2377.330 260.170 2377.610 264.000 ;
        RECT 2377.330 260.030 2380.340 260.170 ;
        RECT 2377.330 260.000 2377.610 260.030 ;
        RECT 2380.200 107.090 2380.340 260.030 ;
        RECT 2380.140 106.770 2380.400 107.090 ;
        RECT 2615.200 106.770 2615.460 107.090 ;
        RECT 2615.260 16.730 2615.400 106.770 ;
        RECT 2615.260 16.590 2619.540 16.730 ;
        RECT 2619.400 2.400 2619.540 16.590 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2393.910 155.280 2394.230 155.340 ;
        RECT 2635.870 155.280 2636.190 155.340 ;
        RECT 2393.910 155.140 2636.190 155.280 ;
        RECT 2393.910 155.080 2394.230 155.140 ;
        RECT 2635.870 155.080 2636.190 155.140 ;
      LAYER via ;
        RECT 2393.940 155.080 2394.200 155.340 ;
        RECT 2635.900 155.080 2636.160 155.340 ;
      LAYER met2 ;
        RECT 2391.590 260.170 2391.870 264.000 ;
        RECT 2391.590 260.030 2394.140 260.170 ;
        RECT 2391.590 260.000 2391.870 260.030 ;
        RECT 2394.000 155.370 2394.140 260.030 ;
        RECT 2393.940 155.050 2394.200 155.370 ;
        RECT 2635.900 155.050 2636.160 155.370 ;
        RECT 2635.960 16.730 2636.100 155.050 ;
        RECT 2635.960 16.590 2637.480 16.730 ;
        RECT 2637.340 2.400 2637.480 16.590 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2407.710 113.800 2408.030 113.860 ;
        RECT 2649.670 113.800 2649.990 113.860 ;
        RECT 2407.710 113.660 2649.990 113.800 ;
        RECT 2407.710 113.600 2408.030 113.660 ;
        RECT 2649.670 113.600 2649.990 113.660 ;
      LAYER via ;
        RECT 2407.740 113.600 2408.000 113.860 ;
        RECT 2649.700 113.600 2649.960 113.860 ;
      LAYER met2 ;
        RECT 2405.850 260.170 2406.130 264.000 ;
        RECT 2405.850 260.030 2407.940 260.170 ;
        RECT 2405.850 260.000 2406.130 260.030 ;
        RECT 2407.800 113.890 2407.940 260.030 ;
        RECT 2407.740 113.570 2408.000 113.890 ;
        RECT 2649.700 113.570 2649.960 113.890 ;
        RECT 2649.760 17.410 2649.900 113.570 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2421.050 203.560 2421.370 203.620 ;
        RECT 2670.370 203.560 2670.690 203.620 ;
        RECT 2421.050 203.420 2670.690 203.560 ;
        RECT 2421.050 203.360 2421.370 203.420 ;
        RECT 2670.370 203.360 2670.690 203.420 ;
      LAYER via ;
        RECT 2421.080 203.360 2421.340 203.620 ;
        RECT 2670.400 203.360 2670.660 203.620 ;
      LAYER met2 ;
        RECT 2419.650 260.170 2419.930 264.000 ;
        RECT 2419.650 260.030 2421.280 260.170 ;
        RECT 2419.650 260.000 2419.930 260.030 ;
        RECT 2421.140 203.650 2421.280 260.030 ;
        RECT 2421.080 203.330 2421.340 203.650 ;
        RECT 2670.400 203.330 2670.660 203.650 ;
        RECT 2670.460 17.410 2670.600 203.330 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2434.850 189.620 2435.170 189.680 ;
        RECT 2684.170 189.620 2684.490 189.680 ;
        RECT 2434.850 189.480 2684.490 189.620 ;
        RECT 2434.850 189.420 2435.170 189.480 ;
        RECT 2684.170 189.420 2684.490 189.480 ;
        RECT 2684.170 16.560 2684.490 16.620 ;
        RECT 2690.610 16.560 2690.930 16.620 ;
        RECT 2684.170 16.420 2690.930 16.560 ;
        RECT 2684.170 16.360 2684.490 16.420 ;
        RECT 2690.610 16.360 2690.930 16.420 ;
      LAYER via ;
        RECT 2434.880 189.420 2435.140 189.680 ;
        RECT 2684.200 189.420 2684.460 189.680 ;
        RECT 2684.200 16.360 2684.460 16.620 ;
        RECT 2690.640 16.360 2690.900 16.620 ;
      LAYER met2 ;
        RECT 2433.910 260.170 2434.190 264.000 ;
        RECT 2433.910 260.030 2435.080 260.170 ;
        RECT 2433.910 260.000 2434.190 260.030 ;
        RECT 2434.940 189.710 2435.080 260.030 ;
        RECT 2434.880 189.390 2435.140 189.710 ;
        RECT 2684.200 189.390 2684.460 189.710 ;
        RECT 2684.260 16.650 2684.400 189.390 ;
        RECT 2684.200 16.330 2684.460 16.650 ;
        RECT 2690.640 16.330 2690.900 16.650 ;
        RECT 2690.700 2.400 2690.840 16.330 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2448.650 207.100 2448.970 207.360 ;
        RECT 2448.740 206.680 2448.880 207.100 ;
        RECT 2448.650 206.420 2448.970 206.680 ;
        RECT 2448.650 148.140 2448.970 148.200 ;
        RECT 2704.870 148.140 2705.190 148.200 ;
        RECT 2448.650 148.000 2705.190 148.140 ;
        RECT 2448.650 147.940 2448.970 148.000 ;
        RECT 2704.870 147.940 2705.190 148.000 ;
      LAYER via ;
        RECT 2448.680 207.100 2448.940 207.360 ;
        RECT 2448.680 206.420 2448.940 206.680 ;
        RECT 2448.680 147.940 2448.940 148.200 ;
        RECT 2704.900 147.940 2705.160 148.200 ;
      LAYER met2 ;
        RECT 2447.710 260.170 2447.990 264.000 ;
        RECT 2447.710 260.030 2448.880 260.170 ;
        RECT 2447.710 260.000 2447.990 260.030 ;
        RECT 2448.740 207.390 2448.880 260.030 ;
        RECT 2448.680 207.070 2448.940 207.390 ;
        RECT 2448.680 206.390 2448.940 206.710 ;
        RECT 2448.740 148.230 2448.880 206.390 ;
        RECT 2448.680 147.910 2448.940 148.230 ;
        RECT 2704.900 147.910 2705.160 148.230 ;
        RECT 2704.960 17.410 2705.100 147.910 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2462.450 182.820 2462.770 182.880 ;
        RECT 2725.570 182.820 2725.890 182.880 ;
        RECT 2462.450 182.680 2725.890 182.820 ;
        RECT 2462.450 182.620 2462.770 182.680 ;
        RECT 2725.570 182.620 2725.890 182.680 ;
      LAYER via ;
        RECT 2462.480 182.620 2462.740 182.880 ;
        RECT 2725.600 182.620 2725.860 182.880 ;
      LAYER met2 ;
        RECT 2461.970 260.170 2462.250 264.000 ;
        RECT 2461.970 260.030 2462.680 260.170 ;
        RECT 2461.970 260.000 2462.250 260.030 ;
        RECT 2462.540 182.910 2462.680 260.030 ;
        RECT 2462.480 182.590 2462.740 182.910 ;
        RECT 2725.600 182.590 2725.860 182.910 ;
        RECT 2725.660 17.410 2725.800 182.590 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2475.790 241.640 2476.110 241.700 ;
        RECT 2480.390 241.640 2480.710 241.700 ;
        RECT 2475.790 241.500 2480.710 241.640 ;
        RECT 2475.790 241.440 2476.110 241.500 ;
        RECT 2480.390 241.440 2480.710 241.500 ;
        RECT 2480.390 86.260 2480.710 86.320 ;
        RECT 2739.370 86.260 2739.690 86.320 ;
        RECT 2480.390 86.120 2739.690 86.260 ;
        RECT 2480.390 86.060 2480.710 86.120 ;
        RECT 2739.370 86.060 2739.690 86.120 ;
      LAYER via ;
        RECT 2475.820 241.440 2476.080 241.700 ;
        RECT 2480.420 241.440 2480.680 241.700 ;
        RECT 2480.420 86.060 2480.680 86.320 ;
        RECT 2739.400 86.060 2739.660 86.320 ;
      LAYER met2 ;
        RECT 2476.230 260.000 2476.510 264.000 ;
        RECT 2476.340 248.610 2476.480 260.000 ;
        RECT 2475.880 248.470 2476.480 248.610 ;
        RECT 2475.880 241.730 2476.020 248.470 ;
        RECT 2475.820 241.410 2476.080 241.730 ;
        RECT 2480.420 241.410 2480.680 241.730 ;
        RECT 2480.480 86.350 2480.620 241.410 ;
        RECT 2480.420 86.030 2480.680 86.350 ;
        RECT 2739.400 86.030 2739.660 86.350 ;
        RECT 2739.460 17.410 2739.600 86.030 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2490.050 176.020 2490.370 176.080 ;
        RECT 2760.070 176.020 2760.390 176.080 ;
        RECT 2490.050 175.880 2760.390 176.020 ;
        RECT 2490.050 175.820 2490.370 175.880 ;
        RECT 2760.070 175.820 2760.390 175.880 ;
      LAYER via ;
        RECT 2490.080 175.820 2490.340 176.080 ;
        RECT 2760.100 175.820 2760.360 176.080 ;
      LAYER met2 ;
        RECT 2490.030 260.000 2490.310 264.000 ;
        RECT 2490.140 176.110 2490.280 260.000 ;
        RECT 2490.080 175.790 2490.340 176.110 ;
        RECT 2760.100 175.790 2760.360 176.110 ;
        RECT 2760.160 17.410 2760.300 175.790 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 835.430 20.300 835.750 20.360 ;
        RECT 966.070 20.300 966.390 20.360 ;
        RECT 835.430 20.160 966.390 20.300 ;
        RECT 835.430 20.100 835.750 20.160 ;
        RECT 966.070 20.100 966.390 20.160 ;
      LAYER via ;
        RECT 835.460 20.100 835.720 20.360 ;
        RECT 966.100 20.100 966.360 20.360 ;
      LAYER met2 ;
        RECT 969.270 260.170 969.550 264.000 ;
        RECT 966.160 260.030 969.550 260.170 ;
        RECT 966.160 20.390 966.300 260.030 ;
        RECT 969.270 260.000 969.550 260.030 ;
        RECT 835.460 20.070 835.720 20.390 ;
        RECT 966.100 20.070 966.360 20.390 ;
        RECT 835.520 2.400 835.660 20.070 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2504.310 65.520 2504.630 65.580 ;
        RECT 2774.330 65.520 2774.650 65.580 ;
        RECT 2504.310 65.380 2774.650 65.520 ;
        RECT 2504.310 65.320 2504.630 65.380 ;
        RECT 2774.330 65.320 2774.650 65.380 ;
      LAYER via ;
        RECT 2504.340 65.320 2504.600 65.580 ;
        RECT 2774.360 65.320 2774.620 65.580 ;
      LAYER met2 ;
        RECT 2504.290 260.000 2504.570 264.000 ;
        RECT 2504.400 65.610 2504.540 260.000 ;
        RECT 2504.340 65.290 2504.600 65.610 ;
        RECT 2774.360 65.290 2774.620 65.610 ;
        RECT 2774.420 17.410 2774.560 65.290 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2518.110 127.740 2518.430 127.800 ;
        RECT 2794.570 127.740 2794.890 127.800 ;
        RECT 2518.110 127.600 2794.890 127.740 ;
        RECT 2518.110 127.540 2518.430 127.600 ;
        RECT 2794.570 127.540 2794.890 127.600 ;
      LAYER via ;
        RECT 2518.140 127.540 2518.400 127.800 ;
        RECT 2794.600 127.540 2794.860 127.800 ;
      LAYER met2 ;
        RECT 2518.090 260.000 2518.370 264.000 ;
        RECT 2518.200 127.830 2518.340 260.000 ;
        RECT 2518.140 127.510 2518.400 127.830 ;
        RECT 2794.600 127.510 2794.860 127.830 ;
        RECT 2794.660 17.410 2794.800 127.510 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2532.370 244.020 2532.690 244.080 ;
        RECT 2538.350 244.020 2538.670 244.080 ;
        RECT 2532.370 243.880 2538.670 244.020 ;
        RECT 2532.370 243.820 2532.690 243.880 ;
        RECT 2538.350 243.820 2538.670 243.880 ;
        RECT 2538.350 168.880 2538.670 168.940 ;
        RECT 2815.730 168.880 2816.050 168.940 ;
        RECT 2538.350 168.740 2816.050 168.880 ;
        RECT 2538.350 168.680 2538.670 168.740 ;
        RECT 2815.730 168.680 2816.050 168.740 ;
      LAYER via ;
        RECT 2532.400 243.820 2532.660 244.080 ;
        RECT 2538.380 243.820 2538.640 244.080 ;
        RECT 2538.380 168.680 2538.640 168.940 ;
        RECT 2815.760 168.680 2816.020 168.940 ;
      LAYER met2 ;
        RECT 2532.350 260.000 2532.630 264.000 ;
        RECT 2532.460 244.110 2532.600 260.000 ;
        RECT 2532.400 243.790 2532.660 244.110 ;
        RECT 2538.380 243.790 2538.640 244.110 ;
        RECT 2538.440 168.970 2538.580 243.790 ;
        RECT 2538.380 168.650 2538.640 168.970 ;
        RECT 2815.760 168.650 2816.020 168.970 ;
        RECT 2815.820 2.400 2815.960 168.650 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2546.630 243.340 2546.950 243.400 ;
        RECT 2552.150 243.340 2552.470 243.400 ;
        RECT 2546.630 243.200 2552.470 243.340 ;
        RECT 2546.630 243.140 2546.950 243.200 ;
        RECT 2552.150 243.140 2552.470 243.200 ;
        RECT 2552.150 72.320 2552.470 72.380 ;
        RECT 2829.070 72.320 2829.390 72.380 ;
        RECT 2552.150 72.180 2829.390 72.320 ;
        RECT 2552.150 72.120 2552.470 72.180 ;
        RECT 2829.070 72.120 2829.390 72.180 ;
      LAYER via ;
        RECT 2546.660 243.140 2546.920 243.400 ;
        RECT 2552.180 243.140 2552.440 243.400 ;
        RECT 2552.180 72.120 2552.440 72.380 ;
        RECT 2829.100 72.120 2829.360 72.380 ;
      LAYER met2 ;
        RECT 2546.610 260.000 2546.890 264.000 ;
        RECT 2546.720 243.430 2546.860 260.000 ;
        RECT 2546.660 243.110 2546.920 243.430 ;
        RECT 2552.180 243.110 2552.440 243.430 ;
        RECT 2552.240 72.410 2552.380 243.110 ;
        RECT 2552.180 72.090 2552.440 72.410 ;
        RECT 2829.100 72.090 2829.360 72.410 ;
        RECT 2829.160 17.410 2829.300 72.090 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2560.430 243.340 2560.750 243.400 ;
        RECT 2565.950 243.340 2566.270 243.400 ;
        RECT 2560.430 243.200 2566.270 243.340 ;
        RECT 2560.430 243.140 2560.750 243.200 ;
        RECT 2565.950 243.140 2566.270 243.200 ;
        RECT 2565.950 59.880 2566.270 60.140 ;
        RECT 2566.040 59.060 2566.180 59.880 ;
        RECT 2566.410 59.060 2566.730 59.120 ;
        RECT 2566.040 58.920 2566.730 59.060 ;
        RECT 2566.410 58.860 2566.730 58.920 ;
        RECT 2566.410 18.600 2566.730 18.660 ;
        RECT 2851.150 18.600 2851.470 18.660 ;
        RECT 2566.410 18.460 2851.470 18.600 ;
        RECT 2566.410 18.400 2566.730 18.460 ;
        RECT 2851.150 18.400 2851.470 18.460 ;
      LAYER via ;
        RECT 2560.460 243.140 2560.720 243.400 ;
        RECT 2565.980 243.140 2566.240 243.400 ;
        RECT 2565.980 59.880 2566.240 60.140 ;
        RECT 2566.440 58.860 2566.700 59.120 ;
        RECT 2566.440 18.400 2566.700 18.660 ;
        RECT 2851.180 18.400 2851.440 18.660 ;
      LAYER met2 ;
        RECT 2560.410 260.000 2560.690 264.000 ;
        RECT 2560.520 243.430 2560.660 260.000 ;
        RECT 2560.460 243.110 2560.720 243.430 ;
        RECT 2565.980 243.110 2566.240 243.430 ;
        RECT 2566.040 60.170 2566.180 243.110 ;
        RECT 2565.980 59.850 2566.240 60.170 ;
        RECT 2566.440 58.830 2566.700 59.150 ;
        RECT 2566.500 18.690 2566.640 58.830 ;
        RECT 2566.440 18.370 2566.700 18.690 ;
        RECT 2851.180 18.370 2851.440 18.690 ;
        RECT 2851.240 2.400 2851.380 18.370 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2574.690 244.020 2575.010 244.080 ;
        RECT 2580.210 244.020 2580.530 244.080 ;
        RECT 2574.690 243.880 2580.530 244.020 ;
        RECT 2574.690 243.820 2575.010 243.880 ;
        RECT 2580.210 243.820 2580.530 243.880 ;
        RECT 2580.210 18.940 2580.530 19.000 ;
        RECT 2869.090 18.940 2869.410 19.000 ;
        RECT 2580.210 18.800 2869.410 18.940 ;
        RECT 2580.210 18.740 2580.530 18.800 ;
        RECT 2869.090 18.740 2869.410 18.800 ;
      LAYER via ;
        RECT 2574.720 243.820 2574.980 244.080 ;
        RECT 2580.240 243.820 2580.500 244.080 ;
        RECT 2580.240 18.740 2580.500 19.000 ;
        RECT 2869.120 18.740 2869.380 19.000 ;
      LAYER met2 ;
        RECT 2574.670 260.000 2574.950 264.000 ;
        RECT 2574.780 244.110 2574.920 260.000 ;
        RECT 2574.720 243.790 2574.980 244.110 ;
        RECT 2580.240 243.790 2580.500 244.110 ;
        RECT 2580.300 19.030 2580.440 243.790 ;
        RECT 2580.240 18.710 2580.500 19.030 ;
        RECT 2869.120 18.710 2869.380 19.030 ;
        RECT 2869.180 2.400 2869.320 18.710 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2588.490 244.020 2588.810 244.080 ;
        RECT 2594.010 244.020 2594.330 244.080 ;
        RECT 2588.490 243.880 2594.330 244.020 ;
        RECT 2588.490 243.820 2588.810 243.880 ;
        RECT 2594.010 243.820 2594.330 243.880 ;
        RECT 2594.010 18.260 2594.330 18.320 ;
        RECT 2887.030 18.260 2887.350 18.320 ;
        RECT 2594.010 18.120 2887.350 18.260 ;
        RECT 2594.010 18.060 2594.330 18.120 ;
        RECT 2887.030 18.060 2887.350 18.120 ;
      LAYER via ;
        RECT 2588.520 243.820 2588.780 244.080 ;
        RECT 2594.040 243.820 2594.300 244.080 ;
        RECT 2594.040 18.060 2594.300 18.320 ;
        RECT 2887.060 18.060 2887.320 18.320 ;
      LAYER met2 ;
        RECT 2588.470 260.000 2588.750 264.000 ;
        RECT 2588.580 244.110 2588.720 260.000 ;
        RECT 2588.520 243.790 2588.780 244.110 ;
        RECT 2594.040 243.790 2594.300 244.110 ;
        RECT 2594.100 18.350 2594.240 243.790 ;
        RECT 2594.040 18.030 2594.300 18.350 ;
        RECT 2887.060 18.030 2887.320 18.350 ;
        RECT 2887.120 2.400 2887.260 18.030 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2602.750 244.020 2603.070 244.080 ;
        RECT 2607.350 244.020 2607.670 244.080 ;
        RECT 2602.750 243.880 2607.670 244.020 ;
        RECT 2602.750 243.820 2603.070 243.880 ;
        RECT 2607.350 243.820 2607.670 243.880 ;
        RECT 2607.810 17.240 2608.130 17.300 ;
        RECT 2904.970 17.240 2905.290 17.300 ;
        RECT 2607.810 17.100 2905.290 17.240 ;
        RECT 2607.810 17.040 2608.130 17.100 ;
        RECT 2904.970 17.040 2905.290 17.100 ;
      LAYER via ;
        RECT 2602.780 243.820 2603.040 244.080 ;
        RECT 2607.380 243.820 2607.640 244.080 ;
        RECT 2607.840 17.040 2608.100 17.300 ;
        RECT 2905.000 17.040 2905.260 17.300 ;
      LAYER met2 ;
        RECT 2602.730 260.000 2603.010 264.000 ;
        RECT 2602.840 244.110 2602.980 260.000 ;
        RECT 2602.780 243.790 2603.040 244.110 ;
        RECT 2607.380 243.790 2607.640 244.110 ;
        RECT 2607.440 17.410 2607.580 243.790 ;
        RECT 2607.440 17.330 2608.040 17.410 ;
        RECT 2607.440 17.270 2608.100 17.330 ;
        RECT 2607.840 17.010 2608.100 17.270 ;
        RECT 2905.000 17.010 2905.260 17.330 ;
        RECT 2905.060 2.400 2905.200 17.010 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 852.910 20.640 853.230 20.700 ;
        RECT 979.870 20.640 980.190 20.700 ;
        RECT 852.910 20.500 980.190 20.640 ;
        RECT 852.910 20.440 853.230 20.500 ;
        RECT 979.870 20.440 980.190 20.500 ;
      LAYER via ;
        RECT 852.940 20.440 853.200 20.700 ;
        RECT 979.900 20.440 980.160 20.700 ;
      LAYER met2 ;
        RECT 983.530 260.170 983.810 264.000 ;
        RECT 979.960 260.030 983.810 260.170 ;
        RECT 979.960 20.730 980.100 260.030 ;
        RECT 983.530 260.000 983.810 260.030 ;
        RECT 852.940 20.410 853.200 20.730 ;
        RECT 979.900 20.410 980.160 20.730 ;
        RECT 853.000 2.400 853.140 20.410 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 16.560 871.170 16.620 ;
        RECT 993.670 16.560 993.990 16.620 ;
        RECT 870.850 16.420 993.990 16.560 ;
        RECT 870.850 16.360 871.170 16.420 ;
        RECT 993.670 16.360 993.990 16.420 ;
      LAYER via ;
        RECT 870.880 16.360 871.140 16.620 ;
        RECT 993.700 16.360 993.960 16.620 ;
      LAYER met2 ;
        RECT 997.330 260.170 997.610 264.000 ;
        RECT 993.760 260.030 997.610 260.170 ;
        RECT 993.760 16.650 993.900 260.030 ;
        RECT 997.330 260.000 997.610 260.030 ;
        RECT 870.880 16.330 871.140 16.650 ;
        RECT 993.700 16.330 993.960 16.650 ;
        RECT 870.940 2.400 871.080 16.330 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 888.790 17.920 889.110 17.980 ;
        RECT 1007.470 17.920 1007.790 17.980 ;
        RECT 888.790 17.780 1007.790 17.920 ;
        RECT 888.790 17.720 889.110 17.780 ;
        RECT 1007.470 17.720 1007.790 17.780 ;
      LAYER via ;
        RECT 888.820 17.720 889.080 17.980 ;
        RECT 1007.500 17.720 1007.760 17.980 ;
      LAYER met2 ;
        RECT 1011.590 260.170 1011.870 264.000 ;
        RECT 1007.560 260.030 1011.870 260.170 ;
        RECT 1007.560 18.010 1007.700 260.030 ;
        RECT 1011.590 260.000 1011.870 260.030 ;
        RECT 888.820 17.690 889.080 18.010 ;
        RECT 1007.500 17.690 1007.760 18.010 ;
        RECT 888.880 2.400 889.020 17.690 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 906.730 18.260 907.050 18.320 ;
        RECT 1021.270 18.260 1021.590 18.320 ;
        RECT 906.730 18.120 1021.590 18.260 ;
        RECT 906.730 18.060 907.050 18.120 ;
        RECT 1021.270 18.060 1021.590 18.120 ;
      LAYER via ;
        RECT 906.760 18.060 907.020 18.320 ;
        RECT 1021.300 18.060 1021.560 18.320 ;
      LAYER met2 ;
        RECT 1025.850 260.170 1026.130 264.000 ;
        RECT 1021.360 260.030 1026.130 260.170 ;
        RECT 1021.360 18.350 1021.500 260.030 ;
        RECT 1025.850 260.000 1026.130 260.030 ;
        RECT 906.760 18.030 907.020 18.350 ;
        RECT 1021.300 18.030 1021.560 18.350 ;
        RECT 906.820 2.400 906.960 18.030 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1003.865 18.445 1004.035 20.655 ;
      LAYER mcon ;
        RECT 1003.865 20.485 1004.035 20.655 ;
      LAYER met1 ;
        RECT 1003.805 20.640 1004.095 20.685 ;
        RECT 1035.530 20.640 1035.850 20.700 ;
        RECT 1003.805 20.500 1035.850 20.640 ;
        RECT 1003.805 20.455 1004.095 20.500 ;
        RECT 1035.530 20.440 1035.850 20.500 ;
        RECT 924.210 18.600 924.530 18.660 ;
        RECT 1003.805 18.600 1004.095 18.645 ;
        RECT 924.210 18.460 1004.095 18.600 ;
        RECT 924.210 18.400 924.530 18.460 ;
        RECT 1003.805 18.415 1004.095 18.460 ;
      LAYER via ;
        RECT 1035.560 20.440 1035.820 20.700 ;
        RECT 924.240 18.400 924.500 18.660 ;
      LAYER met2 ;
        RECT 1039.650 260.170 1039.930 264.000 ;
        RECT 1035.620 260.030 1039.930 260.170 ;
        RECT 1035.620 20.730 1035.760 260.030 ;
        RECT 1039.650 260.000 1039.930 260.030 ;
        RECT 1035.560 20.410 1035.820 20.730 ;
        RECT 924.240 18.370 924.500 18.690 ;
        RECT 924.300 2.400 924.440 18.370 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 942.150 19.280 942.470 19.340 ;
        RECT 1049.790 19.280 1050.110 19.340 ;
        RECT 942.150 19.140 1050.110 19.280 ;
        RECT 942.150 19.080 942.470 19.140 ;
        RECT 1049.790 19.080 1050.110 19.140 ;
      LAYER via ;
        RECT 942.180 19.080 942.440 19.340 ;
        RECT 1049.820 19.080 1050.080 19.340 ;
      LAYER met2 ;
        RECT 1053.910 260.170 1054.190 264.000 ;
        RECT 1049.880 260.030 1054.190 260.170 ;
        RECT 1049.880 19.370 1050.020 260.030 ;
        RECT 1053.910 260.000 1054.190 260.030 ;
        RECT 942.180 19.050 942.440 19.370 ;
        RECT 1049.820 19.050 1050.080 19.370 ;
        RECT 942.240 2.400 942.380 19.050 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1062.670 244.020 1062.990 244.080 ;
        RECT 1066.350 244.020 1066.670 244.080 ;
        RECT 1062.670 243.880 1066.670 244.020 ;
        RECT 1062.670 243.820 1062.990 243.880 ;
        RECT 1066.350 243.820 1066.670 243.880 ;
        RECT 960.090 19.620 960.410 19.680 ;
        RECT 1062.670 19.620 1062.990 19.680 ;
        RECT 960.090 19.480 1062.990 19.620 ;
        RECT 960.090 19.420 960.410 19.480 ;
        RECT 1062.670 19.420 1062.990 19.480 ;
      LAYER via ;
        RECT 1062.700 243.820 1062.960 244.080 ;
        RECT 1066.380 243.820 1066.640 244.080 ;
        RECT 960.120 19.420 960.380 19.680 ;
        RECT 1062.700 19.420 1062.960 19.680 ;
      LAYER met2 ;
        RECT 1067.710 260.170 1067.990 264.000 ;
        RECT 1066.440 260.030 1067.990 260.170 ;
        RECT 1066.440 244.110 1066.580 260.030 ;
        RECT 1067.710 260.000 1067.990 260.030 ;
        RECT 1062.700 243.790 1062.960 244.110 ;
        RECT 1066.380 243.790 1066.640 244.110 ;
        RECT 1062.760 19.710 1062.900 243.790 ;
        RECT 960.120 19.390 960.380 19.710 ;
        RECT 1062.700 19.390 1062.960 19.710 ;
        RECT 960.180 2.400 960.320 19.390 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1076.470 244.020 1076.790 244.080 ;
        RECT 1080.150 244.020 1080.470 244.080 ;
        RECT 1076.470 243.880 1080.470 244.020 ;
        RECT 1076.470 243.820 1076.790 243.880 ;
        RECT 1080.150 243.820 1080.470 243.880 ;
        RECT 978.030 19.960 978.350 20.020 ;
        RECT 1076.470 19.960 1076.790 20.020 ;
        RECT 978.030 19.820 1076.790 19.960 ;
        RECT 978.030 19.760 978.350 19.820 ;
        RECT 1076.470 19.760 1076.790 19.820 ;
      LAYER via ;
        RECT 1076.500 243.820 1076.760 244.080 ;
        RECT 1080.180 243.820 1080.440 244.080 ;
        RECT 978.060 19.760 978.320 20.020 ;
        RECT 1076.500 19.760 1076.760 20.020 ;
      LAYER met2 ;
        RECT 1081.970 260.170 1082.250 264.000 ;
        RECT 1080.240 260.030 1082.250 260.170 ;
        RECT 1080.240 244.110 1080.380 260.030 ;
        RECT 1081.970 260.000 1082.250 260.030 ;
        RECT 1076.500 243.790 1076.760 244.110 ;
        RECT 1080.180 243.790 1080.440 244.110 ;
        RECT 1076.560 20.050 1076.700 243.790 ;
        RECT 978.060 19.730 978.320 20.050 ;
        RECT 1076.500 19.730 1076.760 20.050 ;
        RECT 978.120 2.400 978.260 19.730 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 231.100 662.330 231.160 ;
        RECT 828.530 231.100 828.850 231.160 ;
        RECT 662.010 230.960 828.850 231.100 ;
        RECT 662.010 230.900 662.330 230.960 ;
        RECT 828.530 230.900 828.850 230.960 ;
        RECT 656.950 17.920 657.270 17.980 ;
        RECT 662.010 17.920 662.330 17.980 ;
        RECT 656.950 17.780 662.330 17.920 ;
        RECT 656.950 17.720 657.270 17.780 ;
        RECT 662.010 17.720 662.330 17.780 ;
      LAYER via ;
        RECT 662.040 230.900 662.300 231.160 ;
        RECT 828.560 230.900 828.820 231.160 ;
        RECT 656.980 17.720 657.240 17.980 ;
        RECT 662.040 17.720 662.300 17.980 ;
      LAYER met2 ;
        RECT 828.510 260.000 828.790 264.000 ;
        RECT 828.620 231.190 828.760 260.000 ;
        RECT 662.040 230.870 662.300 231.190 ;
        RECT 828.560 230.870 828.820 231.190 ;
        RECT 662.100 18.010 662.240 230.870 ;
        RECT 656.980 17.690 657.240 18.010 ;
        RECT 662.040 17.690 662.300 18.010 ;
        RECT 657.040 2.400 657.180 17.690 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 995.970 16.560 996.290 16.620 ;
        RECT 1091.650 16.560 1091.970 16.620 ;
        RECT 995.970 16.420 1091.970 16.560 ;
        RECT 995.970 16.360 996.290 16.420 ;
        RECT 1091.650 16.360 1091.970 16.420 ;
      LAYER via ;
        RECT 996.000 16.360 996.260 16.620 ;
        RECT 1091.680 16.360 1091.940 16.620 ;
      LAYER met2 ;
        RECT 1096.230 260.170 1096.510 264.000 ;
        RECT 1091.740 260.030 1096.510 260.170 ;
        RECT 1091.740 16.650 1091.880 260.030 ;
        RECT 1096.230 260.000 1096.510 260.030 ;
        RECT 996.000 16.330 996.260 16.650 ;
        RECT 1091.680 16.330 1091.940 16.650 ;
        RECT 996.060 2.400 996.200 16.330 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 245.040 1014.230 245.100 ;
        RECT 1110.050 245.040 1110.370 245.100 ;
        RECT 1013.910 244.900 1110.370 245.040 ;
        RECT 1013.910 244.840 1014.230 244.900 ;
        RECT 1110.050 244.840 1110.370 244.900 ;
      LAYER via ;
        RECT 1013.940 244.840 1014.200 245.100 ;
        RECT 1110.080 244.840 1110.340 245.100 ;
      LAYER met2 ;
        RECT 1110.030 260.000 1110.310 264.000 ;
        RECT 1110.140 245.130 1110.280 260.000 ;
        RECT 1013.940 244.810 1014.200 245.130 ;
        RECT 1110.080 244.810 1110.340 245.130 ;
        RECT 1014.000 3.130 1014.140 244.810 ;
        RECT 1013.540 2.990 1014.140 3.130 ;
        RECT 1013.540 2.400 1013.680 2.990 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.610 245.720 1034.930 245.780 ;
        RECT 1124.310 245.720 1124.630 245.780 ;
        RECT 1034.610 245.580 1124.630 245.720 ;
        RECT 1034.610 245.520 1034.930 245.580 ;
        RECT 1124.310 245.520 1124.630 245.580 ;
        RECT 1031.390 17.920 1031.710 17.980 ;
        RECT 1034.610 17.920 1034.930 17.980 ;
        RECT 1031.390 17.780 1034.930 17.920 ;
        RECT 1031.390 17.720 1031.710 17.780 ;
        RECT 1034.610 17.720 1034.930 17.780 ;
      LAYER via ;
        RECT 1034.640 245.520 1034.900 245.780 ;
        RECT 1124.340 245.520 1124.600 245.780 ;
        RECT 1031.420 17.720 1031.680 17.980 ;
        RECT 1034.640 17.720 1034.900 17.980 ;
      LAYER met2 ;
        RECT 1124.290 260.000 1124.570 264.000 ;
        RECT 1124.400 245.810 1124.540 260.000 ;
        RECT 1034.640 245.490 1034.900 245.810 ;
        RECT 1124.340 245.490 1124.600 245.810 ;
        RECT 1034.700 18.010 1034.840 245.490 ;
        RECT 1031.420 17.690 1031.680 18.010 ;
        RECT 1034.640 17.690 1034.900 18.010 ;
        RECT 1031.480 2.400 1031.620 17.690 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1131.670 244.020 1131.990 244.080 ;
        RECT 1136.270 244.020 1136.590 244.080 ;
        RECT 1131.670 243.880 1136.590 244.020 ;
        RECT 1131.670 243.820 1131.990 243.880 ;
        RECT 1136.270 243.820 1136.590 243.880 ;
        RECT 1049.330 15.880 1049.650 15.940 ;
        RECT 1131.670 15.880 1131.990 15.940 ;
        RECT 1049.330 15.740 1131.990 15.880 ;
        RECT 1049.330 15.680 1049.650 15.740 ;
        RECT 1131.670 15.680 1131.990 15.740 ;
      LAYER via ;
        RECT 1131.700 243.820 1131.960 244.080 ;
        RECT 1136.300 243.820 1136.560 244.080 ;
        RECT 1049.360 15.680 1049.620 15.940 ;
        RECT 1131.700 15.680 1131.960 15.940 ;
      LAYER met2 ;
        RECT 1138.090 260.170 1138.370 264.000 ;
        RECT 1136.360 260.030 1138.370 260.170 ;
        RECT 1136.360 244.110 1136.500 260.030 ;
        RECT 1138.090 260.000 1138.370 260.030 ;
        RECT 1131.700 243.790 1131.960 244.110 ;
        RECT 1136.300 243.790 1136.560 244.110 ;
        RECT 1131.760 15.970 1131.900 243.790 ;
        RECT 1049.360 15.650 1049.620 15.970 ;
        RECT 1131.700 15.650 1131.960 15.970 ;
        RECT 1049.420 2.400 1049.560 15.650 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 245.380 1069.430 245.440 ;
        RECT 1152.370 245.380 1152.690 245.440 ;
        RECT 1069.110 245.240 1152.690 245.380 ;
        RECT 1069.110 245.180 1069.430 245.240 ;
        RECT 1152.370 245.180 1152.690 245.240 ;
      LAYER via ;
        RECT 1069.140 245.180 1069.400 245.440 ;
        RECT 1152.400 245.180 1152.660 245.440 ;
      LAYER met2 ;
        RECT 1152.350 260.000 1152.630 264.000 ;
        RECT 1152.460 245.470 1152.600 260.000 ;
        RECT 1069.140 245.150 1069.400 245.470 ;
        RECT 1152.400 245.150 1152.660 245.470 ;
        RECT 1069.200 3.130 1069.340 245.150 ;
        RECT 1067.360 2.990 1069.340 3.130 ;
        RECT 1067.360 2.400 1067.500 2.990 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 246.740 1090.130 246.800 ;
        RECT 1166.630 246.740 1166.950 246.800 ;
        RECT 1089.810 246.600 1166.950 246.740 ;
        RECT 1089.810 246.540 1090.130 246.600 ;
        RECT 1166.630 246.540 1166.950 246.600 ;
        RECT 1085.210 17.580 1085.530 17.640 ;
        RECT 1089.810 17.580 1090.130 17.640 ;
        RECT 1085.210 17.440 1090.130 17.580 ;
        RECT 1085.210 17.380 1085.530 17.440 ;
        RECT 1089.810 17.380 1090.130 17.440 ;
      LAYER via ;
        RECT 1089.840 246.540 1090.100 246.800 ;
        RECT 1166.660 246.540 1166.920 246.800 ;
        RECT 1085.240 17.380 1085.500 17.640 ;
        RECT 1089.840 17.380 1090.100 17.640 ;
      LAYER met2 ;
        RECT 1166.610 260.000 1166.890 264.000 ;
        RECT 1166.720 246.830 1166.860 260.000 ;
        RECT 1089.840 246.510 1090.100 246.830 ;
        RECT 1166.660 246.510 1166.920 246.830 ;
        RECT 1089.900 17.670 1090.040 246.510 ;
        RECT 1085.240 17.350 1085.500 17.670 ;
        RECT 1089.840 17.350 1090.100 17.670 ;
        RECT 1085.300 2.400 1085.440 17.350 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.610 247.080 1103.930 247.140 ;
        RECT 1180.430 247.080 1180.750 247.140 ;
        RECT 1103.610 246.940 1180.750 247.080 ;
        RECT 1103.610 246.880 1103.930 246.940 ;
        RECT 1180.430 246.880 1180.750 246.940 ;
        RECT 1102.690 2.960 1103.010 3.020 ;
        RECT 1103.610 2.960 1103.930 3.020 ;
        RECT 1102.690 2.820 1103.930 2.960 ;
        RECT 1102.690 2.760 1103.010 2.820 ;
        RECT 1103.610 2.760 1103.930 2.820 ;
      LAYER via ;
        RECT 1103.640 246.880 1103.900 247.140 ;
        RECT 1180.460 246.880 1180.720 247.140 ;
        RECT 1102.720 2.760 1102.980 3.020 ;
        RECT 1103.640 2.760 1103.900 3.020 ;
      LAYER met2 ;
        RECT 1180.410 260.000 1180.690 264.000 ;
        RECT 1180.520 247.170 1180.660 260.000 ;
        RECT 1103.640 246.850 1103.900 247.170 ;
        RECT 1180.460 246.850 1180.720 247.170 ;
        RECT 1103.700 3.050 1103.840 246.850 ;
        RECT 1102.720 2.730 1102.980 3.050 ;
        RECT 1103.640 2.730 1103.900 3.050 ;
        RECT 1102.780 2.400 1102.920 2.730 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1120.630 19.620 1120.950 19.680 ;
        RECT 1194.230 19.620 1194.550 19.680 ;
        RECT 1120.630 19.480 1194.550 19.620 ;
        RECT 1120.630 19.420 1120.950 19.480 ;
        RECT 1194.230 19.420 1194.550 19.480 ;
      LAYER via ;
        RECT 1120.660 19.420 1120.920 19.680 ;
        RECT 1194.260 19.420 1194.520 19.680 ;
      LAYER met2 ;
        RECT 1194.670 260.170 1194.950 264.000 ;
        RECT 1194.320 260.030 1194.950 260.170 ;
        RECT 1194.320 19.710 1194.460 260.030 ;
        RECT 1194.670 260.000 1194.950 260.030 ;
        RECT 1120.660 19.390 1120.920 19.710 ;
        RECT 1194.260 19.390 1194.520 19.710 ;
        RECT 1120.720 2.400 1120.860 19.390 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 246.060 1145.330 246.120 ;
        RECT 1208.490 246.060 1208.810 246.120 ;
        RECT 1145.010 245.920 1208.810 246.060 ;
        RECT 1145.010 245.860 1145.330 245.920 ;
        RECT 1208.490 245.860 1208.810 245.920 ;
        RECT 1138.570 16.900 1138.890 16.960 ;
        RECT 1145.010 16.900 1145.330 16.960 ;
        RECT 1138.570 16.760 1145.330 16.900 ;
        RECT 1138.570 16.700 1138.890 16.760 ;
        RECT 1145.010 16.700 1145.330 16.760 ;
      LAYER via ;
        RECT 1145.040 245.860 1145.300 246.120 ;
        RECT 1208.520 245.860 1208.780 246.120 ;
        RECT 1138.600 16.700 1138.860 16.960 ;
        RECT 1145.040 16.700 1145.300 16.960 ;
      LAYER met2 ;
        RECT 1208.470 260.000 1208.750 264.000 ;
        RECT 1208.580 246.150 1208.720 260.000 ;
        RECT 1145.040 245.830 1145.300 246.150 ;
        RECT 1208.520 245.830 1208.780 246.150 ;
        RECT 1145.100 16.990 1145.240 245.830 ;
        RECT 1138.600 16.670 1138.860 16.990 ;
        RECT 1145.040 16.670 1145.300 16.990 ;
        RECT 1138.660 2.400 1138.800 16.670 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 245.380 1159.130 245.440 ;
        RECT 1222.750 245.380 1223.070 245.440 ;
        RECT 1158.810 245.240 1223.070 245.380 ;
        RECT 1158.810 245.180 1159.130 245.240 ;
        RECT 1222.750 245.180 1223.070 245.240 ;
        RECT 1156.510 17.580 1156.830 17.640 ;
        RECT 1158.810 17.580 1159.130 17.640 ;
        RECT 1156.510 17.440 1159.130 17.580 ;
        RECT 1156.510 17.380 1156.830 17.440 ;
        RECT 1158.810 17.380 1159.130 17.440 ;
      LAYER via ;
        RECT 1158.840 245.180 1159.100 245.440 ;
        RECT 1222.780 245.180 1223.040 245.440 ;
        RECT 1156.540 17.380 1156.800 17.640 ;
        RECT 1158.840 17.380 1159.100 17.640 ;
      LAYER met2 ;
        RECT 1222.730 260.000 1223.010 264.000 ;
        RECT 1222.840 245.470 1222.980 260.000 ;
        RECT 1158.840 245.150 1159.100 245.470 ;
        RECT 1222.780 245.150 1223.040 245.470 ;
        RECT 1158.900 17.670 1159.040 245.150 ;
        RECT 1156.540 17.350 1156.800 17.670 ;
        RECT 1158.840 17.350 1159.100 17.670 ;
        RECT 1156.600 2.400 1156.740 17.350 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 675.810 93.060 676.130 93.120 ;
        RECT 841.870 93.060 842.190 93.120 ;
        RECT 675.810 92.920 842.190 93.060 ;
        RECT 675.810 92.860 676.130 92.920 ;
        RECT 841.870 92.860 842.190 92.920 ;
      LAYER via ;
        RECT 675.840 92.860 676.100 93.120 ;
        RECT 841.900 92.860 842.160 93.120 ;
      LAYER met2 ;
        RECT 842.770 260.170 843.050 264.000 ;
        RECT 841.960 260.030 843.050 260.170 ;
        RECT 841.960 93.150 842.100 260.030 ;
        RECT 842.770 260.000 843.050 260.030 ;
        RECT 675.840 92.830 676.100 93.150 ;
        RECT 841.900 92.830 842.160 93.150 ;
        RECT 675.900 3.130 676.040 92.830 ;
        RECT 674.520 2.990 676.040 3.130 ;
        RECT 674.520 2.400 674.660 2.990 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1235.630 18.260 1235.950 18.320 ;
        RECT 1197.540 18.120 1235.950 18.260 ;
        RECT 1173.990 17.580 1174.310 17.640 ;
        RECT 1197.540 17.580 1197.680 18.120 ;
        RECT 1235.630 18.060 1235.950 18.120 ;
        RECT 1173.990 17.440 1197.680 17.580 ;
        RECT 1173.990 17.380 1174.310 17.440 ;
      LAYER via ;
        RECT 1174.020 17.380 1174.280 17.640 ;
        RECT 1235.660 18.060 1235.920 18.320 ;
      LAYER met2 ;
        RECT 1236.990 260.170 1237.270 264.000 ;
        RECT 1235.720 260.030 1237.270 260.170 ;
        RECT 1235.720 18.350 1235.860 260.030 ;
        RECT 1236.990 260.000 1237.270 260.030 ;
        RECT 1235.660 18.030 1235.920 18.350 ;
        RECT 1174.020 17.350 1174.280 17.670 ;
        RECT 1174.080 2.400 1174.220 17.350 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.310 247.420 1193.630 247.480 ;
        RECT 1250.810 247.420 1251.130 247.480 ;
        RECT 1193.310 247.280 1251.130 247.420 ;
        RECT 1193.310 247.220 1193.630 247.280 ;
        RECT 1250.810 247.220 1251.130 247.280 ;
        RECT 1191.930 2.960 1192.250 3.020 ;
        RECT 1193.310 2.960 1193.630 3.020 ;
        RECT 1191.930 2.820 1193.630 2.960 ;
        RECT 1191.930 2.760 1192.250 2.820 ;
        RECT 1193.310 2.760 1193.630 2.820 ;
      LAYER via ;
        RECT 1193.340 247.220 1193.600 247.480 ;
        RECT 1250.840 247.220 1251.100 247.480 ;
        RECT 1191.960 2.760 1192.220 3.020 ;
        RECT 1193.340 2.760 1193.600 3.020 ;
      LAYER met2 ;
        RECT 1250.790 260.000 1251.070 264.000 ;
        RECT 1250.900 247.510 1251.040 260.000 ;
        RECT 1193.340 247.190 1193.600 247.510 ;
        RECT 1250.840 247.190 1251.100 247.510 ;
        RECT 1193.400 3.050 1193.540 247.190 ;
        RECT 1191.960 2.730 1192.220 3.050 ;
        RECT 1193.340 2.730 1193.600 3.050 ;
        RECT 1192.020 2.400 1192.160 2.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1214.010 246.060 1214.330 246.120 ;
        RECT 1265.070 246.060 1265.390 246.120 ;
        RECT 1214.010 245.920 1265.390 246.060 ;
        RECT 1214.010 245.860 1214.330 245.920 ;
        RECT 1265.070 245.860 1265.390 245.920 ;
        RECT 1209.870 17.580 1210.190 17.640 ;
        RECT 1214.010 17.580 1214.330 17.640 ;
        RECT 1209.870 17.440 1214.330 17.580 ;
        RECT 1209.870 17.380 1210.190 17.440 ;
        RECT 1214.010 17.380 1214.330 17.440 ;
      LAYER via ;
        RECT 1214.040 245.860 1214.300 246.120 ;
        RECT 1265.100 245.860 1265.360 246.120 ;
        RECT 1209.900 17.380 1210.160 17.640 ;
        RECT 1214.040 17.380 1214.300 17.640 ;
      LAYER met2 ;
        RECT 1265.050 260.000 1265.330 264.000 ;
        RECT 1265.160 246.150 1265.300 260.000 ;
        RECT 1214.040 245.830 1214.300 246.150 ;
        RECT 1265.100 245.830 1265.360 246.150 ;
        RECT 1214.100 17.670 1214.240 245.830 ;
        RECT 1209.900 17.350 1210.160 17.670 ;
        RECT 1214.040 17.350 1214.300 17.670 ;
        RECT 1209.960 2.400 1210.100 17.350 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 245.380 1228.130 245.440 ;
        RECT 1279.330 245.380 1279.650 245.440 ;
        RECT 1227.810 245.240 1279.650 245.380 ;
        RECT 1227.810 245.180 1228.130 245.240 ;
        RECT 1279.330 245.180 1279.650 245.240 ;
      LAYER via ;
        RECT 1227.840 245.180 1228.100 245.440 ;
        RECT 1279.360 245.180 1279.620 245.440 ;
      LAYER met2 ;
        RECT 1279.310 260.000 1279.590 264.000 ;
        RECT 1279.420 245.470 1279.560 260.000 ;
        RECT 1227.840 245.150 1228.100 245.470 ;
        RECT 1279.360 245.150 1279.620 245.470 ;
        RECT 1227.900 2.400 1228.040 245.150 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 247.080 1248.830 247.140 ;
        RECT 1293.130 247.080 1293.450 247.140 ;
        RECT 1248.510 246.940 1293.450 247.080 ;
        RECT 1248.510 246.880 1248.830 246.940 ;
        RECT 1293.130 246.880 1293.450 246.940 ;
        RECT 1245.750 17.580 1246.070 17.640 ;
        RECT 1248.510 17.580 1248.830 17.640 ;
        RECT 1245.750 17.440 1248.830 17.580 ;
        RECT 1245.750 17.380 1246.070 17.440 ;
        RECT 1248.510 17.380 1248.830 17.440 ;
      LAYER via ;
        RECT 1248.540 246.880 1248.800 247.140 ;
        RECT 1293.160 246.880 1293.420 247.140 ;
        RECT 1245.780 17.380 1246.040 17.640 ;
        RECT 1248.540 17.380 1248.800 17.640 ;
      LAYER met2 ;
        RECT 1293.110 260.000 1293.390 264.000 ;
        RECT 1293.220 247.170 1293.360 260.000 ;
        RECT 1248.540 246.850 1248.800 247.170 ;
        RECT 1293.160 246.850 1293.420 247.170 ;
        RECT 1248.600 17.670 1248.740 246.850 ;
        RECT 1245.780 17.350 1246.040 17.670 ;
        RECT 1248.540 17.350 1248.800 17.670 ;
        RECT 1245.840 2.400 1245.980 17.350 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1269.210 246.060 1269.530 246.120 ;
        RECT 1307.390 246.060 1307.710 246.120 ;
        RECT 1269.210 245.920 1307.710 246.060 ;
        RECT 1269.210 245.860 1269.530 245.920 ;
        RECT 1307.390 245.860 1307.710 245.920 ;
        RECT 1263.230 17.580 1263.550 17.640 ;
        RECT 1269.210 17.580 1269.530 17.640 ;
        RECT 1263.230 17.440 1269.530 17.580 ;
        RECT 1263.230 17.380 1263.550 17.440 ;
        RECT 1269.210 17.380 1269.530 17.440 ;
      LAYER via ;
        RECT 1269.240 245.860 1269.500 246.120 ;
        RECT 1307.420 245.860 1307.680 246.120 ;
        RECT 1263.260 17.380 1263.520 17.640 ;
        RECT 1269.240 17.380 1269.500 17.640 ;
      LAYER met2 ;
        RECT 1307.370 260.000 1307.650 264.000 ;
        RECT 1307.480 246.150 1307.620 260.000 ;
        RECT 1269.240 245.830 1269.500 246.150 ;
        RECT 1307.420 245.830 1307.680 246.150 ;
        RECT 1269.300 17.670 1269.440 245.830 ;
        RECT 1263.260 17.350 1263.520 17.670 ;
        RECT 1269.240 17.350 1269.500 17.670 ;
        RECT 1263.320 2.400 1263.460 17.350 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 245.380 1283.330 245.440 ;
        RECT 1321.190 245.380 1321.510 245.440 ;
        RECT 1283.010 245.240 1321.510 245.380 ;
        RECT 1283.010 245.180 1283.330 245.240 ;
        RECT 1321.190 245.180 1321.510 245.240 ;
      LAYER via ;
        RECT 1283.040 245.180 1283.300 245.440 ;
        RECT 1321.220 245.180 1321.480 245.440 ;
      LAYER met2 ;
        RECT 1321.170 260.000 1321.450 264.000 ;
        RECT 1321.280 245.470 1321.420 260.000 ;
        RECT 1283.040 245.150 1283.300 245.470 ;
        RECT 1321.220 245.150 1321.480 245.470 ;
        RECT 1283.100 17.410 1283.240 245.150 ;
        RECT 1281.260 17.270 1283.240 17.410 ;
        RECT 1281.260 2.400 1281.400 17.270 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1307.390 241.980 1307.710 242.040 ;
        RECT 1335.450 241.980 1335.770 242.040 ;
        RECT 1307.390 241.840 1335.770 241.980 ;
        RECT 1307.390 241.780 1307.710 241.840 ;
        RECT 1335.450 241.780 1335.770 241.840 ;
        RECT 1299.110 17.580 1299.430 17.640 ;
        RECT 1307.390 17.580 1307.710 17.640 ;
        RECT 1299.110 17.440 1307.710 17.580 ;
        RECT 1299.110 17.380 1299.430 17.440 ;
        RECT 1307.390 17.380 1307.710 17.440 ;
      LAYER via ;
        RECT 1307.420 241.780 1307.680 242.040 ;
        RECT 1335.480 241.780 1335.740 242.040 ;
        RECT 1299.140 17.380 1299.400 17.640 ;
        RECT 1307.420 17.380 1307.680 17.640 ;
      LAYER met2 ;
        RECT 1335.430 260.000 1335.710 264.000 ;
        RECT 1335.540 242.070 1335.680 260.000 ;
        RECT 1307.420 241.750 1307.680 242.070 ;
        RECT 1335.480 241.750 1335.740 242.070 ;
        RECT 1307.480 17.670 1307.620 241.750 ;
        RECT 1299.140 17.350 1299.400 17.670 ;
        RECT 1307.420 17.350 1307.680 17.670 ;
        RECT 1299.200 2.400 1299.340 17.350 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 248.100 1317.370 248.160 ;
        RECT 1349.710 248.100 1350.030 248.160 ;
        RECT 1317.050 247.960 1350.030 248.100 ;
        RECT 1317.050 247.900 1317.370 247.960 ;
        RECT 1349.710 247.900 1350.030 247.960 ;
      LAYER via ;
        RECT 1317.080 247.900 1317.340 248.160 ;
        RECT 1349.740 247.900 1350.000 248.160 ;
      LAYER met2 ;
        RECT 1349.690 260.000 1349.970 264.000 ;
        RECT 1349.800 248.190 1349.940 260.000 ;
        RECT 1317.080 247.870 1317.340 248.190 ;
        RECT 1349.740 247.870 1350.000 248.190 ;
        RECT 1317.140 2.400 1317.280 247.870 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 245.720 1338.530 245.780 ;
        RECT 1363.510 245.720 1363.830 245.780 ;
        RECT 1338.210 245.580 1363.830 245.720 ;
        RECT 1338.210 245.520 1338.530 245.580 ;
        RECT 1363.510 245.520 1363.830 245.580 ;
        RECT 1334.990 17.240 1335.310 17.300 ;
        RECT 1338.210 17.240 1338.530 17.300 ;
        RECT 1334.990 17.100 1338.530 17.240 ;
        RECT 1334.990 17.040 1335.310 17.100 ;
        RECT 1338.210 17.040 1338.530 17.100 ;
      LAYER via ;
        RECT 1338.240 245.520 1338.500 245.780 ;
        RECT 1363.540 245.520 1363.800 245.780 ;
        RECT 1335.020 17.040 1335.280 17.300 ;
        RECT 1338.240 17.040 1338.500 17.300 ;
      LAYER met2 ;
        RECT 1363.490 260.000 1363.770 264.000 ;
        RECT 1363.600 245.810 1363.740 260.000 ;
        RECT 1338.240 245.490 1338.500 245.810 ;
        RECT 1363.540 245.490 1363.800 245.810 ;
        RECT 1338.300 17.330 1338.440 245.490 ;
        RECT 1335.020 17.010 1335.280 17.330 ;
        RECT 1338.240 17.010 1338.500 17.330 ;
        RECT 1335.080 2.400 1335.220 17.010 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 696.510 224.300 696.830 224.360 ;
        RECT 856.130 224.300 856.450 224.360 ;
        RECT 696.510 224.160 856.450 224.300 ;
        RECT 696.510 224.100 696.830 224.160 ;
        RECT 856.130 224.100 856.450 224.160 ;
        RECT 692.370 15.200 692.690 15.260 ;
        RECT 696.510 15.200 696.830 15.260 ;
        RECT 692.370 15.060 696.830 15.200 ;
        RECT 692.370 15.000 692.690 15.060 ;
        RECT 696.510 15.000 696.830 15.060 ;
      LAYER via ;
        RECT 696.540 224.100 696.800 224.360 ;
        RECT 856.160 224.100 856.420 224.360 ;
        RECT 692.400 15.000 692.660 15.260 ;
        RECT 696.540 15.000 696.800 15.260 ;
      LAYER met2 ;
        RECT 856.570 260.170 856.850 264.000 ;
        RECT 856.220 260.030 856.850 260.170 ;
        RECT 856.220 224.390 856.360 260.030 ;
        RECT 856.570 260.000 856.850 260.030 ;
        RECT 696.540 224.070 696.800 224.390 ;
        RECT 856.160 224.070 856.420 224.390 ;
        RECT 696.600 15.290 696.740 224.070 ;
        RECT 692.400 14.970 692.660 15.290 ;
        RECT 696.540 14.970 696.800 15.290 ;
        RECT 692.460 2.400 692.600 14.970 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1362.590 244.020 1362.910 244.080 ;
        RECT 1377.770 244.020 1378.090 244.080 ;
        RECT 1362.590 243.880 1378.090 244.020 ;
        RECT 1362.590 243.820 1362.910 243.880 ;
        RECT 1377.770 243.820 1378.090 243.880 ;
        RECT 1352.470 17.580 1352.790 17.640 ;
        RECT 1362.590 17.580 1362.910 17.640 ;
        RECT 1352.470 17.440 1362.910 17.580 ;
        RECT 1352.470 17.380 1352.790 17.440 ;
        RECT 1362.590 17.380 1362.910 17.440 ;
      LAYER via ;
        RECT 1362.620 243.820 1362.880 244.080 ;
        RECT 1377.800 243.820 1378.060 244.080 ;
        RECT 1352.500 17.380 1352.760 17.640 ;
        RECT 1362.620 17.380 1362.880 17.640 ;
      LAYER met2 ;
        RECT 1377.750 260.000 1378.030 264.000 ;
        RECT 1377.860 244.110 1378.000 260.000 ;
        RECT 1362.620 243.790 1362.880 244.110 ;
        RECT 1377.800 243.790 1378.060 244.110 ;
        RECT 1362.680 17.670 1362.820 243.790 ;
        RECT 1352.500 17.350 1352.760 17.670 ;
        RECT 1362.620 17.350 1362.880 17.670 ;
        RECT 1352.560 2.400 1352.700 17.350 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1372.710 248.100 1373.030 248.160 ;
        RECT 1391.570 248.100 1391.890 248.160 ;
        RECT 1372.710 247.960 1391.890 248.100 ;
        RECT 1372.710 247.900 1373.030 247.960 ;
        RECT 1391.570 247.900 1391.890 247.960 ;
        RECT 1370.410 17.580 1370.730 17.640 ;
        RECT 1372.710 17.580 1373.030 17.640 ;
        RECT 1370.410 17.440 1373.030 17.580 ;
        RECT 1370.410 17.380 1370.730 17.440 ;
        RECT 1372.710 17.380 1373.030 17.440 ;
      LAYER via ;
        RECT 1372.740 247.900 1373.000 248.160 ;
        RECT 1391.600 247.900 1391.860 248.160 ;
        RECT 1370.440 17.380 1370.700 17.640 ;
        RECT 1372.740 17.380 1373.000 17.640 ;
      LAYER met2 ;
        RECT 1391.550 260.000 1391.830 264.000 ;
        RECT 1391.660 248.190 1391.800 260.000 ;
        RECT 1372.740 247.870 1373.000 248.190 ;
        RECT 1391.600 247.870 1391.860 248.190 ;
        RECT 1372.800 17.670 1372.940 247.870 ;
        RECT 1370.440 17.350 1370.700 17.670 ;
        RECT 1372.740 17.350 1373.000 17.670 ;
        RECT 1370.500 2.400 1370.640 17.350 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1388.350 17.240 1388.670 17.300 ;
        RECT 1401.230 17.240 1401.550 17.300 ;
        RECT 1388.350 17.100 1401.550 17.240 ;
        RECT 1388.350 17.040 1388.670 17.100 ;
        RECT 1401.230 17.040 1401.550 17.100 ;
      LAYER via ;
        RECT 1388.380 17.040 1388.640 17.300 ;
        RECT 1401.260 17.040 1401.520 17.300 ;
      LAYER met2 ;
        RECT 1405.810 260.170 1406.090 264.000 ;
        RECT 1402.240 260.030 1406.090 260.170 ;
        RECT 1402.240 243.850 1402.380 260.030 ;
        RECT 1405.810 260.000 1406.090 260.030 ;
        RECT 1401.320 243.710 1402.380 243.850 ;
        RECT 1401.320 17.330 1401.460 243.710 ;
        RECT 1388.380 17.010 1388.640 17.330 ;
        RECT 1401.260 17.010 1401.520 17.330 ;
        RECT 1388.440 2.400 1388.580 17.010 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 244.020 1407.530 244.080 ;
        RECT 1420.090 244.020 1420.410 244.080 ;
        RECT 1407.210 243.880 1420.410 244.020 ;
        RECT 1407.210 243.820 1407.530 243.880 ;
        RECT 1420.090 243.820 1420.410 243.880 ;
      LAYER via ;
        RECT 1407.240 243.820 1407.500 244.080 ;
        RECT 1420.120 243.820 1420.380 244.080 ;
      LAYER met2 ;
        RECT 1420.070 260.000 1420.350 264.000 ;
        RECT 1420.180 244.110 1420.320 260.000 ;
        RECT 1407.240 243.790 1407.500 244.110 ;
        RECT 1420.120 243.790 1420.380 244.110 ;
        RECT 1407.300 24.210 1407.440 243.790 ;
        RECT 1406.380 24.070 1407.440 24.210 ;
        RECT 1406.380 2.400 1406.520 24.070 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1423.770 19.960 1424.090 20.020 ;
        RECT 1428.830 19.960 1429.150 20.020 ;
        RECT 1423.770 19.820 1429.150 19.960 ;
        RECT 1423.770 19.760 1424.090 19.820 ;
        RECT 1428.830 19.760 1429.150 19.820 ;
      LAYER via ;
        RECT 1423.800 19.760 1424.060 20.020 ;
        RECT 1428.860 19.760 1429.120 20.020 ;
      LAYER met2 ;
        RECT 1433.870 260.170 1434.150 264.000 ;
        RECT 1430.300 260.030 1434.150 260.170 ;
        RECT 1430.300 230.250 1430.440 260.030 ;
        RECT 1433.870 260.000 1434.150 260.030 ;
        RECT 1428.920 230.110 1430.440 230.250 ;
        RECT 1428.920 20.050 1429.060 230.110 ;
        RECT 1423.800 19.730 1424.060 20.050 ;
        RECT 1428.860 19.730 1429.120 20.050 ;
        RECT 1423.860 2.400 1424.000 19.730 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1448.150 241.640 1448.470 241.700 ;
        RECT 1441.340 241.500 1448.470 241.640 ;
        RECT 1441.340 241.360 1441.480 241.500 ;
        RECT 1448.150 241.440 1448.470 241.500 ;
        RECT 1441.250 241.100 1441.570 241.360 ;
      LAYER via ;
        RECT 1448.180 241.440 1448.440 241.700 ;
        RECT 1441.280 241.100 1441.540 241.360 ;
      LAYER met2 ;
        RECT 1448.130 260.000 1448.410 264.000 ;
        RECT 1448.240 241.730 1448.380 260.000 ;
        RECT 1448.180 241.410 1448.440 241.730 ;
        RECT 1441.280 241.070 1441.540 241.390 ;
        RECT 1441.340 20.130 1441.480 241.070 ;
        RECT 1441.340 19.990 1441.940 20.130 ;
        RECT 1441.800 2.400 1441.940 19.990 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1456.965 144.925 1457.135 193.035 ;
      LAYER mcon ;
        RECT 1456.965 192.865 1457.135 193.035 ;
      LAYER met1 ;
        RECT 1456.890 193.020 1457.210 193.080 ;
        RECT 1456.695 192.880 1457.210 193.020 ;
        RECT 1456.890 192.820 1457.210 192.880 ;
        RECT 1456.905 145.080 1457.195 145.125 ;
        RECT 1457.350 145.080 1457.670 145.140 ;
        RECT 1456.905 144.940 1457.670 145.080 ;
        RECT 1456.905 144.895 1457.195 144.940 ;
        RECT 1457.350 144.880 1457.670 144.940 ;
        RECT 1456.430 110.400 1456.750 110.460 ;
        RECT 1457.350 110.400 1457.670 110.460 ;
        RECT 1456.430 110.260 1457.670 110.400 ;
        RECT 1456.430 110.200 1456.750 110.260 ;
        RECT 1457.350 110.200 1457.670 110.260 ;
        RECT 1457.350 20.640 1457.670 20.700 ;
        RECT 1459.650 20.640 1459.970 20.700 ;
        RECT 1457.350 20.500 1459.970 20.640 ;
        RECT 1457.350 20.440 1457.670 20.500 ;
        RECT 1459.650 20.440 1459.970 20.500 ;
      LAYER via ;
        RECT 1456.920 192.820 1457.180 193.080 ;
        RECT 1457.380 144.880 1457.640 145.140 ;
        RECT 1456.460 110.200 1456.720 110.460 ;
        RECT 1457.380 110.200 1457.640 110.460 ;
        RECT 1457.380 20.440 1457.640 20.700 ;
        RECT 1459.680 20.440 1459.940 20.700 ;
      LAYER met2 ;
        RECT 1462.390 260.170 1462.670 264.000 ;
        RECT 1458.360 260.030 1462.670 260.170 ;
        RECT 1458.360 226.170 1458.500 260.030 ;
        RECT 1462.390 260.000 1462.670 260.030 ;
        RECT 1456.980 226.030 1458.500 226.170 ;
        RECT 1456.980 193.110 1457.120 226.030 ;
        RECT 1456.920 192.790 1457.180 193.110 ;
        RECT 1457.380 144.850 1457.640 145.170 ;
        RECT 1457.440 110.570 1457.580 144.850 ;
        RECT 1456.520 110.490 1457.580 110.570 ;
        RECT 1456.460 110.430 1457.640 110.490 ;
        RECT 1456.460 110.170 1456.720 110.430 ;
        RECT 1457.380 110.170 1457.640 110.430 ;
        RECT 1457.440 60.250 1457.580 110.170 ;
        RECT 1457.440 60.110 1458.040 60.250 ;
        RECT 1457.900 58.890 1458.040 60.110 ;
        RECT 1457.440 58.750 1458.040 58.890 ;
        RECT 1457.440 20.730 1457.580 58.750 ;
        RECT 1457.380 20.410 1457.640 20.730 ;
        RECT 1459.680 20.410 1459.940 20.730 ;
        RECT 1459.740 2.400 1459.880 20.410 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1476.190 260.000 1476.470 264.000 ;
        RECT 1476.300 20.130 1476.440 260.000 ;
        RECT 1476.300 19.990 1477.820 20.130 ;
        RECT 1477.680 2.400 1477.820 19.990 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1490.470 20.640 1490.790 20.700 ;
        RECT 1495.530 20.640 1495.850 20.700 ;
        RECT 1490.470 20.500 1495.850 20.640 ;
        RECT 1490.470 20.440 1490.790 20.500 ;
        RECT 1495.530 20.440 1495.850 20.500 ;
      LAYER via ;
        RECT 1490.500 20.440 1490.760 20.700 ;
        RECT 1495.560 20.440 1495.820 20.700 ;
      LAYER met2 ;
        RECT 1490.450 260.000 1490.730 264.000 ;
        RECT 1490.560 20.730 1490.700 260.000 ;
        RECT 1490.500 20.410 1490.760 20.730 ;
        RECT 1495.560 20.410 1495.820 20.730 ;
        RECT 1495.620 2.400 1495.760 20.410 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1504.270 241.640 1504.590 241.700 ;
        RECT 1510.710 241.640 1511.030 241.700 ;
        RECT 1504.270 241.500 1511.030 241.640 ;
        RECT 1504.270 241.440 1504.590 241.500 ;
        RECT 1510.710 241.440 1511.030 241.500 ;
        RECT 1510.710 17.580 1511.030 17.640 ;
        RECT 1513.010 17.580 1513.330 17.640 ;
        RECT 1510.710 17.440 1513.330 17.580 ;
        RECT 1510.710 17.380 1511.030 17.440 ;
        RECT 1513.010 17.380 1513.330 17.440 ;
      LAYER via ;
        RECT 1504.300 241.440 1504.560 241.700 ;
        RECT 1510.740 241.440 1511.000 241.700 ;
        RECT 1510.740 17.380 1511.000 17.640 ;
        RECT 1513.040 17.380 1513.300 17.640 ;
      LAYER met2 ;
        RECT 1504.250 260.000 1504.530 264.000 ;
        RECT 1504.360 241.730 1504.500 260.000 ;
        RECT 1504.300 241.410 1504.560 241.730 ;
        RECT 1510.740 241.410 1511.000 241.730 ;
        RECT 1510.800 17.670 1510.940 241.410 ;
        RECT 1510.740 17.350 1511.000 17.670 ;
        RECT 1513.040 17.350 1513.300 17.670 ;
        RECT 1513.100 2.400 1513.240 17.350 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 710.310 99.860 710.630 99.920 ;
        RECT 869.930 99.860 870.250 99.920 ;
        RECT 710.310 99.720 870.250 99.860 ;
        RECT 710.310 99.660 710.630 99.720 ;
        RECT 869.930 99.660 870.250 99.720 ;
      LAYER via ;
        RECT 710.340 99.660 710.600 99.920 ;
        RECT 869.960 99.660 870.220 99.920 ;
      LAYER met2 ;
        RECT 870.830 260.170 871.110 264.000 ;
        RECT 870.020 260.030 871.110 260.170 ;
        RECT 870.020 99.950 870.160 260.030 ;
        RECT 870.830 260.000 871.110 260.030 ;
        RECT 710.340 99.630 710.600 99.950 ;
        RECT 869.960 99.630 870.220 99.950 ;
        RECT 710.400 2.400 710.540 99.630 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1518.530 242.320 1518.850 242.380 ;
        RECT 1524.510 242.320 1524.830 242.380 ;
        RECT 1518.530 242.180 1524.830 242.320 ;
        RECT 1518.530 242.120 1518.850 242.180 ;
        RECT 1524.510 242.120 1524.830 242.180 ;
        RECT 1524.510 17.580 1524.830 17.640 ;
        RECT 1530.950 17.580 1531.270 17.640 ;
        RECT 1524.510 17.440 1531.270 17.580 ;
        RECT 1524.510 17.380 1524.830 17.440 ;
        RECT 1530.950 17.380 1531.270 17.440 ;
      LAYER via ;
        RECT 1518.560 242.120 1518.820 242.380 ;
        RECT 1524.540 242.120 1524.800 242.380 ;
        RECT 1524.540 17.380 1524.800 17.640 ;
        RECT 1530.980 17.380 1531.240 17.640 ;
      LAYER met2 ;
        RECT 1518.510 260.000 1518.790 264.000 ;
        RECT 1518.620 242.410 1518.760 260.000 ;
        RECT 1518.560 242.090 1518.820 242.410 ;
        RECT 1524.540 242.090 1524.800 242.410 ;
        RECT 1524.600 17.670 1524.740 242.090 ;
        RECT 1524.540 17.350 1524.800 17.670 ;
        RECT 1530.980 17.350 1531.240 17.670 ;
        RECT 1531.040 2.400 1531.180 17.350 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1532.790 243.340 1533.110 243.400 ;
        RECT 1546.590 243.340 1546.910 243.400 ;
        RECT 1532.790 243.200 1546.910 243.340 ;
        RECT 1532.790 243.140 1533.110 243.200 ;
        RECT 1546.590 243.140 1546.910 243.200 ;
      LAYER via ;
        RECT 1532.820 243.140 1533.080 243.400 ;
        RECT 1546.620 243.140 1546.880 243.400 ;
      LAYER met2 ;
        RECT 1532.770 260.000 1533.050 264.000 ;
        RECT 1532.880 243.430 1533.020 260.000 ;
        RECT 1532.820 243.110 1533.080 243.430 ;
        RECT 1546.620 243.110 1546.880 243.430 ;
        RECT 1546.680 7.210 1546.820 243.110 ;
        RECT 1546.680 7.070 1548.660 7.210 ;
        RECT 1548.520 3.130 1548.660 7.070 ;
        RECT 1548.520 2.990 1549.120 3.130 ;
        RECT 1548.980 2.400 1549.120 2.990 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1546.590 244.020 1546.910 244.080 ;
        RECT 1552.110 244.020 1552.430 244.080 ;
        RECT 1546.590 243.880 1552.430 244.020 ;
        RECT 1546.590 243.820 1546.910 243.880 ;
        RECT 1552.110 243.820 1552.430 243.880 ;
        RECT 1552.110 17.580 1552.430 17.640 ;
        RECT 1566.830 17.580 1567.150 17.640 ;
        RECT 1552.110 17.440 1567.150 17.580 ;
        RECT 1552.110 17.380 1552.430 17.440 ;
        RECT 1566.830 17.380 1567.150 17.440 ;
      LAYER via ;
        RECT 1546.620 243.820 1546.880 244.080 ;
        RECT 1552.140 243.820 1552.400 244.080 ;
        RECT 1552.140 17.380 1552.400 17.640 ;
        RECT 1566.860 17.380 1567.120 17.640 ;
      LAYER met2 ;
        RECT 1546.570 260.000 1546.850 264.000 ;
        RECT 1546.680 244.110 1546.820 260.000 ;
        RECT 1546.620 243.790 1546.880 244.110 ;
        RECT 1552.140 243.790 1552.400 244.110 ;
        RECT 1552.200 17.670 1552.340 243.790 ;
        RECT 1552.140 17.350 1552.400 17.670 ;
        RECT 1566.860 17.350 1567.120 17.670 ;
        RECT 1566.920 2.400 1567.060 17.350 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1560.850 243.680 1561.170 243.740 ;
        RECT 1565.910 243.680 1566.230 243.740 ;
        RECT 1560.850 243.540 1566.230 243.680 ;
        RECT 1560.850 243.480 1561.170 243.540 ;
        RECT 1565.910 243.480 1566.230 243.540 ;
        RECT 1584.770 17.580 1585.090 17.640 ;
        RECT 1567.380 17.440 1585.090 17.580 ;
        RECT 1565.910 17.240 1566.230 17.300 ;
        RECT 1567.380 17.240 1567.520 17.440 ;
        RECT 1584.770 17.380 1585.090 17.440 ;
        RECT 1565.910 17.100 1567.520 17.240 ;
        RECT 1565.910 17.040 1566.230 17.100 ;
      LAYER via ;
        RECT 1560.880 243.480 1561.140 243.740 ;
        RECT 1565.940 243.480 1566.200 243.740 ;
        RECT 1565.940 17.040 1566.200 17.300 ;
        RECT 1584.800 17.380 1585.060 17.640 ;
      LAYER met2 ;
        RECT 1560.830 260.000 1561.110 264.000 ;
        RECT 1560.940 243.770 1561.080 260.000 ;
        RECT 1560.880 243.450 1561.140 243.770 ;
        RECT 1565.940 243.450 1566.200 243.770 ;
        RECT 1566.000 17.330 1566.140 243.450 ;
        RECT 1584.800 17.350 1585.060 17.670 ;
        RECT 1565.940 17.010 1566.200 17.330 ;
        RECT 1584.860 2.400 1585.000 17.350 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1574.650 243.680 1574.970 243.740 ;
        RECT 1579.710 243.680 1580.030 243.740 ;
        RECT 1574.650 243.540 1580.030 243.680 ;
        RECT 1574.650 243.480 1574.970 243.540 ;
        RECT 1579.710 243.480 1580.030 243.540 ;
        RECT 1579.710 18.260 1580.030 18.320 ;
        RECT 1602.250 18.260 1602.570 18.320 ;
        RECT 1579.710 18.120 1602.570 18.260 ;
        RECT 1579.710 18.060 1580.030 18.120 ;
        RECT 1602.250 18.060 1602.570 18.120 ;
      LAYER via ;
        RECT 1574.680 243.480 1574.940 243.740 ;
        RECT 1579.740 243.480 1580.000 243.740 ;
        RECT 1579.740 18.060 1580.000 18.320 ;
        RECT 1602.280 18.060 1602.540 18.320 ;
      LAYER met2 ;
        RECT 1574.630 260.000 1574.910 264.000 ;
        RECT 1574.740 243.770 1574.880 260.000 ;
        RECT 1574.680 243.450 1574.940 243.770 ;
        RECT 1579.740 243.450 1580.000 243.770 ;
        RECT 1579.800 18.350 1579.940 243.450 ;
        RECT 1579.740 18.030 1580.000 18.350 ;
        RECT 1602.280 18.030 1602.540 18.350 ;
        RECT 1602.340 2.400 1602.480 18.030 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1588.910 244.020 1589.230 244.080 ;
        RECT 1604.090 244.020 1604.410 244.080 ;
        RECT 1588.910 243.880 1604.410 244.020 ;
        RECT 1588.910 243.820 1589.230 243.880 ;
        RECT 1604.090 243.820 1604.410 243.880 ;
        RECT 1604.090 16.560 1604.410 16.620 ;
        RECT 1620.190 16.560 1620.510 16.620 ;
        RECT 1604.090 16.420 1620.510 16.560 ;
        RECT 1604.090 16.360 1604.410 16.420 ;
        RECT 1620.190 16.360 1620.510 16.420 ;
      LAYER via ;
        RECT 1588.940 243.820 1589.200 244.080 ;
        RECT 1604.120 243.820 1604.380 244.080 ;
        RECT 1604.120 16.360 1604.380 16.620 ;
        RECT 1620.220 16.360 1620.480 16.620 ;
      LAYER met2 ;
        RECT 1588.890 260.000 1589.170 264.000 ;
        RECT 1589.000 244.110 1589.140 260.000 ;
        RECT 1588.940 243.790 1589.200 244.110 ;
        RECT 1604.120 243.790 1604.380 244.110 ;
        RECT 1604.180 16.650 1604.320 243.790 ;
        RECT 1604.120 16.330 1604.380 16.650 ;
        RECT 1620.220 16.330 1620.480 16.650 ;
        RECT 1620.280 2.400 1620.420 16.330 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1603.170 243.000 1603.490 243.060 ;
        RECT 1607.310 243.000 1607.630 243.060 ;
        RECT 1603.170 242.860 1607.630 243.000 ;
        RECT 1603.170 242.800 1603.490 242.860 ;
        RECT 1607.310 242.800 1607.630 242.860 ;
        RECT 1607.310 15.200 1607.630 15.260 ;
        RECT 1638.130 15.200 1638.450 15.260 ;
        RECT 1607.310 15.060 1638.450 15.200 ;
        RECT 1607.310 15.000 1607.630 15.060 ;
        RECT 1638.130 15.000 1638.450 15.060 ;
      LAYER via ;
        RECT 1603.200 242.800 1603.460 243.060 ;
        RECT 1607.340 242.800 1607.600 243.060 ;
        RECT 1607.340 15.000 1607.600 15.260 ;
        RECT 1638.160 15.000 1638.420 15.260 ;
      LAYER met2 ;
        RECT 1603.150 260.000 1603.430 264.000 ;
        RECT 1603.260 243.090 1603.400 260.000 ;
        RECT 1603.200 242.770 1603.460 243.090 ;
        RECT 1607.340 242.770 1607.600 243.090 ;
        RECT 1607.400 15.290 1607.540 242.770 ;
        RECT 1607.340 14.970 1607.600 15.290 ;
        RECT 1638.160 14.970 1638.420 15.290 ;
        RECT 1638.220 2.400 1638.360 14.970 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1616.970 243.000 1617.290 243.060 ;
        RECT 1621.110 243.000 1621.430 243.060 ;
        RECT 1616.970 242.860 1621.430 243.000 ;
        RECT 1616.970 242.800 1617.290 242.860 ;
        RECT 1621.110 242.800 1621.430 242.860 ;
        RECT 1621.110 18.260 1621.430 18.320 ;
        RECT 1656.070 18.260 1656.390 18.320 ;
        RECT 1621.110 18.120 1656.390 18.260 ;
        RECT 1621.110 18.060 1621.430 18.120 ;
        RECT 1656.070 18.060 1656.390 18.120 ;
      LAYER via ;
        RECT 1617.000 242.800 1617.260 243.060 ;
        RECT 1621.140 242.800 1621.400 243.060 ;
        RECT 1621.140 18.060 1621.400 18.320 ;
        RECT 1656.100 18.060 1656.360 18.320 ;
      LAYER met2 ;
        RECT 1616.950 260.000 1617.230 264.000 ;
        RECT 1617.060 243.090 1617.200 260.000 ;
        RECT 1617.000 242.770 1617.260 243.090 ;
        RECT 1621.140 242.770 1621.400 243.090 ;
        RECT 1621.200 18.350 1621.340 242.770 ;
        RECT 1621.140 18.030 1621.400 18.350 ;
        RECT 1656.100 18.030 1656.360 18.350 ;
        RECT 1656.160 2.400 1656.300 18.030 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1631.230 244.020 1631.550 244.080 ;
        RECT 1634.910 244.020 1635.230 244.080 ;
        RECT 1631.230 243.880 1635.230 244.020 ;
        RECT 1631.230 243.820 1631.550 243.880 ;
        RECT 1634.910 243.820 1635.230 243.880 ;
        RECT 1634.910 14.520 1635.230 14.580 ;
        RECT 1673.550 14.520 1673.870 14.580 ;
        RECT 1634.910 14.380 1673.870 14.520 ;
        RECT 1634.910 14.320 1635.230 14.380 ;
        RECT 1673.550 14.320 1673.870 14.380 ;
      LAYER via ;
        RECT 1631.260 243.820 1631.520 244.080 ;
        RECT 1634.940 243.820 1635.200 244.080 ;
        RECT 1634.940 14.320 1635.200 14.580 ;
        RECT 1673.580 14.320 1673.840 14.580 ;
      LAYER met2 ;
        RECT 1631.210 260.000 1631.490 264.000 ;
        RECT 1631.320 244.110 1631.460 260.000 ;
        RECT 1631.260 243.790 1631.520 244.110 ;
        RECT 1634.940 243.790 1635.200 244.110 ;
        RECT 1635.000 14.610 1635.140 243.790 ;
        RECT 1634.940 14.290 1635.200 14.610 ;
        RECT 1673.580 14.290 1673.840 14.610 ;
        RECT 1673.640 2.400 1673.780 14.290 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1645.030 244.020 1645.350 244.080 ;
        RECT 1648.710 244.020 1649.030 244.080 ;
        RECT 1645.030 243.880 1649.030 244.020 ;
        RECT 1645.030 243.820 1645.350 243.880 ;
        RECT 1648.710 243.820 1649.030 243.880 ;
        RECT 1648.710 17.920 1649.030 17.980 ;
        RECT 1691.490 17.920 1691.810 17.980 ;
        RECT 1648.710 17.780 1691.810 17.920 ;
        RECT 1648.710 17.720 1649.030 17.780 ;
        RECT 1691.490 17.720 1691.810 17.780 ;
      LAYER via ;
        RECT 1645.060 243.820 1645.320 244.080 ;
        RECT 1648.740 243.820 1649.000 244.080 ;
        RECT 1648.740 17.720 1649.000 17.980 ;
        RECT 1691.520 17.720 1691.780 17.980 ;
      LAYER met2 ;
        RECT 1645.010 260.000 1645.290 264.000 ;
        RECT 1645.120 244.110 1645.260 260.000 ;
        RECT 1645.060 243.790 1645.320 244.110 ;
        RECT 1648.740 243.790 1649.000 244.110 ;
        RECT 1648.800 18.010 1648.940 243.790 ;
        RECT 1648.740 17.690 1649.000 18.010 ;
        RECT 1691.520 17.690 1691.780 18.010 ;
        RECT 1691.580 2.400 1691.720 17.690 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 731.010 107.340 731.330 107.400 ;
        RECT 883.730 107.340 884.050 107.400 ;
        RECT 731.010 107.200 884.050 107.340 ;
        RECT 731.010 107.140 731.330 107.200 ;
        RECT 883.730 107.140 884.050 107.200 ;
        RECT 728.250 17.920 728.570 17.980 ;
        RECT 731.010 17.920 731.330 17.980 ;
        RECT 728.250 17.780 731.330 17.920 ;
        RECT 728.250 17.720 728.570 17.780 ;
        RECT 731.010 17.720 731.330 17.780 ;
      LAYER via ;
        RECT 731.040 107.140 731.300 107.400 ;
        RECT 883.760 107.140 884.020 107.400 ;
        RECT 728.280 17.720 728.540 17.980 ;
        RECT 731.040 17.720 731.300 17.980 ;
      LAYER met2 ;
        RECT 884.630 260.170 884.910 264.000 ;
        RECT 883.820 260.030 884.910 260.170 ;
        RECT 883.820 107.430 883.960 260.030 ;
        RECT 884.630 260.000 884.910 260.030 ;
        RECT 731.040 107.110 731.300 107.430 ;
        RECT 883.760 107.110 884.020 107.430 ;
        RECT 731.100 18.010 731.240 107.110 ;
        RECT 728.280 17.690 728.540 18.010 ;
        RECT 731.040 17.690 731.300 18.010 ;
        RECT 728.340 2.400 728.480 17.690 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 19.960 1662.830 20.020 ;
        RECT 1709.430 19.960 1709.750 20.020 ;
        RECT 1662.510 19.820 1709.750 19.960 ;
        RECT 1662.510 19.760 1662.830 19.820 ;
        RECT 1709.430 19.760 1709.750 19.820 ;
      LAYER via ;
        RECT 1662.540 19.760 1662.800 20.020 ;
        RECT 1709.460 19.760 1709.720 20.020 ;
      LAYER met2 ;
        RECT 1659.270 260.170 1659.550 264.000 ;
        RECT 1659.270 260.030 1662.740 260.170 ;
        RECT 1659.270 260.000 1659.550 260.030 ;
        RECT 1662.600 20.050 1662.740 260.030 ;
        RECT 1662.540 19.730 1662.800 20.050 ;
        RECT 1709.460 19.730 1709.720 20.050 ;
        RECT 1709.520 2.400 1709.660 19.730 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1676.310 19.620 1676.630 19.680 ;
        RECT 1727.370 19.620 1727.690 19.680 ;
        RECT 1676.310 19.480 1727.690 19.620 ;
        RECT 1676.310 19.420 1676.630 19.480 ;
        RECT 1727.370 19.420 1727.690 19.480 ;
      LAYER via ;
        RECT 1676.340 19.420 1676.600 19.680 ;
        RECT 1727.400 19.420 1727.660 19.680 ;
      LAYER met2 ;
        RECT 1673.530 260.170 1673.810 264.000 ;
        RECT 1673.530 260.030 1676.540 260.170 ;
        RECT 1673.530 260.000 1673.810 260.030 ;
        RECT 1676.400 19.710 1676.540 260.030 ;
        RECT 1676.340 19.390 1676.600 19.710 ;
        RECT 1727.400 19.390 1727.660 19.710 ;
        RECT 1727.460 2.400 1727.600 19.390 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1690.110 20.640 1690.430 20.700 ;
        RECT 1744.390 20.640 1744.710 20.700 ;
        RECT 1690.110 20.500 1744.710 20.640 ;
        RECT 1690.110 20.440 1690.430 20.500 ;
        RECT 1744.390 20.440 1744.710 20.500 ;
      LAYER via ;
        RECT 1690.140 20.440 1690.400 20.700 ;
        RECT 1744.420 20.440 1744.680 20.700 ;
      LAYER met2 ;
        RECT 1687.330 260.170 1687.610 264.000 ;
        RECT 1687.330 260.030 1690.340 260.170 ;
        RECT 1687.330 260.000 1687.610 260.030 ;
        RECT 1690.200 20.730 1690.340 260.030 ;
        RECT 1690.140 20.410 1690.400 20.730 ;
        RECT 1744.420 20.410 1744.680 20.730 ;
        RECT 1744.480 18.090 1744.620 20.410 ;
        RECT 1744.480 17.950 1745.540 18.090 ;
        RECT 1745.400 2.400 1745.540 17.950 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1703.910 16.560 1704.230 16.620 ;
        RECT 1762.790 16.560 1763.110 16.620 ;
        RECT 1703.910 16.420 1763.110 16.560 ;
        RECT 1703.910 16.360 1704.230 16.420 ;
        RECT 1762.790 16.360 1763.110 16.420 ;
      LAYER via ;
        RECT 1703.940 16.360 1704.200 16.620 ;
        RECT 1762.820 16.360 1763.080 16.620 ;
      LAYER met2 ;
        RECT 1701.590 260.170 1701.870 264.000 ;
        RECT 1701.590 260.030 1704.140 260.170 ;
        RECT 1701.590 260.000 1701.870 260.030 ;
        RECT 1704.000 16.650 1704.140 260.030 ;
        RECT 1703.940 16.330 1704.200 16.650 ;
        RECT 1762.820 16.330 1763.080 16.650 ;
        RECT 1762.880 2.400 1763.020 16.330 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1717.710 17.580 1718.030 17.640 ;
        RECT 1780.730 17.580 1781.050 17.640 ;
        RECT 1717.710 17.440 1781.050 17.580 ;
        RECT 1717.710 17.380 1718.030 17.440 ;
        RECT 1780.730 17.380 1781.050 17.440 ;
      LAYER via ;
        RECT 1717.740 17.380 1718.000 17.640 ;
        RECT 1780.760 17.380 1781.020 17.640 ;
      LAYER met2 ;
        RECT 1715.850 260.170 1716.130 264.000 ;
        RECT 1715.850 260.030 1717.940 260.170 ;
        RECT 1715.850 260.000 1716.130 260.030 ;
        RECT 1717.800 17.670 1717.940 260.030 ;
        RECT 1717.740 17.350 1718.000 17.670 ;
        RECT 1780.760 17.350 1781.020 17.670 ;
        RECT 1780.820 2.400 1780.960 17.350 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.510 19.960 1731.830 20.020 ;
        RECT 1798.670 19.960 1798.990 20.020 ;
        RECT 1731.510 19.820 1798.990 19.960 ;
        RECT 1731.510 19.760 1731.830 19.820 ;
        RECT 1798.670 19.760 1798.990 19.820 ;
      LAYER via ;
        RECT 1731.540 19.760 1731.800 20.020 ;
        RECT 1798.700 19.760 1798.960 20.020 ;
      LAYER met2 ;
        RECT 1729.650 260.170 1729.930 264.000 ;
        RECT 1729.650 260.030 1731.740 260.170 ;
        RECT 1729.650 260.000 1729.930 260.030 ;
        RECT 1731.600 20.050 1731.740 260.030 ;
        RECT 1731.540 19.730 1731.800 20.050 ;
        RECT 1798.700 19.730 1798.960 20.050 ;
        RECT 1798.760 2.400 1798.900 19.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1745.310 19.280 1745.630 19.340 ;
        RECT 1816.610 19.280 1816.930 19.340 ;
        RECT 1745.310 19.140 1816.930 19.280 ;
        RECT 1745.310 19.080 1745.630 19.140 ;
        RECT 1816.610 19.080 1816.930 19.140 ;
      LAYER via ;
        RECT 1745.340 19.080 1745.600 19.340 ;
        RECT 1816.640 19.080 1816.900 19.340 ;
      LAYER met2 ;
        RECT 1743.910 260.170 1744.190 264.000 ;
        RECT 1743.910 260.030 1745.540 260.170 ;
        RECT 1743.910 260.000 1744.190 260.030 ;
        RECT 1745.400 19.370 1745.540 260.030 ;
        RECT 1745.340 19.050 1745.600 19.370 ;
        RECT 1816.640 19.050 1816.900 19.370 ;
        RECT 1816.700 2.400 1816.840 19.050 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1759.110 18.940 1759.430 19.000 ;
        RECT 1834.550 18.940 1834.870 19.000 ;
        RECT 1759.110 18.800 1834.870 18.940 ;
        RECT 1759.110 18.740 1759.430 18.800 ;
        RECT 1834.550 18.740 1834.870 18.800 ;
      LAYER via ;
        RECT 1759.140 18.740 1759.400 19.000 ;
        RECT 1834.580 18.740 1834.840 19.000 ;
      LAYER met2 ;
        RECT 1757.710 260.170 1757.990 264.000 ;
        RECT 1757.710 260.030 1759.340 260.170 ;
        RECT 1757.710 260.000 1757.990 260.030 ;
        RECT 1759.200 19.030 1759.340 260.030 ;
        RECT 1759.140 18.710 1759.400 19.030 ;
        RECT 1834.580 18.710 1834.840 19.030 ;
        RECT 1834.640 2.400 1834.780 18.710 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 20.300 1773.230 20.360 ;
        RECT 1852.030 20.300 1852.350 20.360 ;
        RECT 1772.910 20.160 1852.350 20.300 ;
        RECT 1772.910 20.100 1773.230 20.160 ;
        RECT 1852.030 20.100 1852.350 20.160 ;
      LAYER via ;
        RECT 1772.940 20.100 1773.200 20.360 ;
        RECT 1852.060 20.100 1852.320 20.360 ;
      LAYER met2 ;
        RECT 1771.970 260.170 1772.250 264.000 ;
        RECT 1771.970 260.030 1773.140 260.170 ;
        RECT 1771.970 260.000 1772.250 260.030 ;
        RECT 1773.000 20.390 1773.140 260.030 ;
        RECT 1772.940 20.070 1773.200 20.390 ;
        RECT 1852.060 20.070 1852.320 20.390 ;
        RECT 1852.120 2.400 1852.260 20.070 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1786.710 17.580 1787.030 17.640 ;
        RECT 1869.970 17.580 1870.290 17.640 ;
        RECT 1786.710 17.440 1870.290 17.580 ;
        RECT 1786.710 17.380 1787.030 17.440 ;
        RECT 1869.970 17.380 1870.290 17.440 ;
      LAYER via ;
        RECT 1786.740 17.380 1787.000 17.640 ;
        RECT 1870.000 17.380 1870.260 17.640 ;
      LAYER met2 ;
        RECT 1786.230 260.170 1786.510 264.000 ;
        RECT 1786.230 260.030 1786.940 260.170 ;
        RECT 1786.230 260.000 1786.510 260.030 ;
        RECT 1786.800 17.670 1786.940 260.030 ;
        RECT 1786.740 17.350 1787.000 17.670 ;
        RECT 1870.000 17.350 1870.260 17.670 ;
        RECT 1870.060 2.400 1870.200 17.350 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 858.045 16.065 858.215 18.275 ;
      LAYER mcon ;
        RECT 858.045 18.105 858.215 18.275 ;
      LAYER met1 ;
        RECT 746.190 18.260 746.510 18.320 ;
        RECT 857.985 18.260 858.275 18.305 ;
        RECT 746.190 18.120 858.275 18.260 ;
        RECT 746.190 18.060 746.510 18.120 ;
        RECT 857.985 18.075 858.275 18.120 ;
        RECT 857.985 16.220 858.275 16.265 ;
        RECT 897.530 16.220 897.850 16.280 ;
        RECT 857.985 16.080 897.850 16.220 ;
        RECT 857.985 16.035 858.275 16.080 ;
        RECT 897.530 16.020 897.850 16.080 ;
      LAYER via ;
        RECT 746.220 18.060 746.480 18.320 ;
        RECT 897.560 16.020 897.820 16.280 ;
      LAYER met2 ;
        RECT 898.890 260.170 899.170 264.000 ;
        RECT 897.620 260.030 899.170 260.170 ;
        RECT 746.220 18.030 746.480 18.350 ;
        RECT 746.280 2.400 746.420 18.030 ;
        RECT 897.620 16.310 897.760 260.030 ;
        RECT 898.890 260.000 899.170 260.030 ;
        RECT 897.560 15.990 897.820 16.310 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.510 17.240 1800.830 17.300 ;
        RECT 1887.910 17.240 1888.230 17.300 ;
        RECT 1800.510 17.100 1888.230 17.240 ;
        RECT 1800.510 17.040 1800.830 17.100 ;
        RECT 1887.910 17.040 1888.230 17.100 ;
      LAYER via ;
        RECT 1800.540 17.040 1800.800 17.300 ;
        RECT 1887.940 17.040 1888.200 17.300 ;
      LAYER met2 ;
        RECT 1800.030 260.170 1800.310 264.000 ;
        RECT 1800.030 260.030 1800.740 260.170 ;
        RECT 1800.030 260.000 1800.310 260.030 ;
        RECT 1800.600 17.330 1800.740 260.030 ;
        RECT 1800.540 17.010 1800.800 17.330 ;
        RECT 1887.940 17.010 1888.200 17.330 ;
        RECT 1888.000 2.400 1888.140 17.010 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1814.310 18.600 1814.630 18.660 ;
        RECT 1905.850 18.600 1906.170 18.660 ;
        RECT 1814.310 18.460 1906.170 18.600 ;
        RECT 1814.310 18.400 1814.630 18.460 ;
        RECT 1905.850 18.400 1906.170 18.460 ;
      LAYER via ;
        RECT 1814.340 18.400 1814.600 18.660 ;
        RECT 1905.880 18.400 1906.140 18.660 ;
      LAYER met2 ;
        RECT 1814.290 260.000 1814.570 264.000 ;
        RECT 1814.400 18.690 1814.540 260.000 ;
        RECT 1814.340 18.370 1814.600 18.690 ;
        RECT 1905.880 18.370 1906.140 18.690 ;
        RECT 1905.940 2.400 1906.080 18.370 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1828.110 19.280 1828.430 19.340 ;
        RECT 1923.330 19.280 1923.650 19.340 ;
        RECT 1828.110 19.140 1923.650 19.280 ;
        RECT 1828.110 19.080 1828.430 19.140 ;
        RECT 1923.330 19.080 1923.650 19.140 ;
      LAYER via ;
        RECT 1828.140 19.080 1828.400 19.340 ;
        RECT 1923.360 19.080 1923.620 19.340 ;
      LAYER met2 ;
        RECT 1828.090 260.000 1828.370 264.000 ;
        RECT 1828.200 19.370 1828.340 260.000 ;
        RECT 1828.140 19.050 1828.400 19.370 ;
        RECT 1923.360 19.050 1923.620 19.370 ;
        RECT 1923.420 2.400 1923.560 19.050 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1842.370 244.020 1842.690 244.080 ;
        RECT 1848.350 244.020 1848.670 244.080 ;
        RECT 1842.370 243.880 1848.670 244.020 ;
        RECT 1842.370 243.820 1842.690 243.880 ;
        RECT 1848.350 243.820 1848.670 243.880 ;
        RECT 1848.350 18.940 1848.670 19.000 ;
        RECT 1941.270 18.940 1941.590 19.000 ;
        RECT 1848.350 18.800 1941.590 18.940 ;
        RECT 1848.350 18.740 1848.670 18.800 ;
        RECT 1941.270 18.740 1941.590 18.800 ;
      LAYER via ;
        RECT 1842.400 243.820 1842.660 244.080 ;
        RECT 1848.380 243.820 1848.640 244.080 ;
        RECT 1848.380 18.740 1848.640 19.000 ;
        RECT 1941.300 18.740 1941.560 19.000 ;
      LAYER met2 ;
        RECT 1842.350 260.000 1842.630 264.000 ;
        RECT 1842.460 244.110 1842.600 260.000 ;
        RECT 1842.400 243.790 1842.660 244.110 ;
        RECT 1848.380 243.790 1848.640 244.110 ;
        RECT 1848.440 19.030 1848.580 243.790 ;
        RECT 1848.380 18.710 1848.640 19.030 ;
        RECT 1941.300 18.710 1941.560 19.030 ;
        RECT 1941.360 2.400 1941.500 18.710 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1856.630 244.020 1856.950 244.080 ;
        RECT 1862.150 244.020 1862.470 244.080 ;
        RECT 1856.630 243.880 1862.470 244.020 ;
        RECT 1856.630 243.820 1856.950 243.880 ;
        RECT 1862.150 243.820 1862.470 243.880 ;
        RECT 1862.150 15.880 1862.470 15.940 ;
        RECT 1959.210 15.880 1959.530 15.940 ;
        RECT 1862.150 15.740 1959.530 15.880 ;
        RECT 1862.150 15.680 1862.470 15.740 ;
        RECT 1959.210 15.680 1959.530 15.740 ;
      LAYER via ;
        RECT 1856.660 243.820 1856.920 244.080 ;
        RECT 1862.180 243.820 1862.440 244.080 ;
        RECT 1862.180 15.680 1862.440 15.940 ;
        RECT 1959.240 15.680 1959.500 15.940 ;
      LAYER met2 ;
        RECT 1856.610 260.000 1856.890 264.000 ;
        RECT 1856.720 244.110 1856.860 260.000 ;
        RECT 1856.660 243.790 1856.920 244.110 ;
        RECT 1862.180 243.790 1862.440 244.110 ;
        RECT 1862.240 15.970 1862.380 243.790 ;
        RECT 1862.180 15.650 1862.440 15.970 ;
        RECT 1959.240 15.650 1959.500 15.970 ;
        RECT 1959.300 2.400 1959.440 15.650 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1870.430 244.020 1870.750 244.080 ;
        RECT 1876.410 244.020 1876.730 244.080 ;
        RECT 1870.430 243.880 1876.730 244.020 ;
        RECT 1870.430 243.820 1870.750 243.880 ;
        RECT 1876.410 243.820 1876.730 243.880 ;
        RECT 1876.410 16.220 1876.730 16.280 ;
        RECT 1977.150 16.220 1977.470 16.280 ;
        RECT 1876.410 16.080 1977.470 16.220 ;
        RECT 1876.410 16.020 1876.730 16.080 ;
        RECT 1977.150 16.020 1977.470 16.080 ;
      LAYER via ;
        RECT 1870.460 243.820 1870.720 244.080 ;
        RECT 1876.440 243.820 1876.700 244.080 ;
        RECT 1876.440 16.020 1876.700 16.280 ;
        RECT 1977.180 16.020 1977.440 16.280 ;
      LAYER met2 ;
        RECT 1870.410 260.000 1870.690 264.000 ;
        RECT 1870.520 244.110 1870.660 260.000 ;
        RECT 1870.460 243.790 1870.720 244.110 ;
        RECT 1876.440 243.790 1876.700 244.110 ;
        RECT 1876.500 16.310 1876.640 243.790 ;
        RECT 1876.440 15.990 1876.700 16.310 ;
        RECT 1977.180 15.990 1977.440 16.310 ;
        RECT 1977.240 2.400 1977.380 15.990 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1884.690 244.020 1885.010 244.080 ;
        RECT 1890.210 244.020 1890.530 244.080 ;
        RECT 1884.690 243.880 1890.530 244.020 ;
        RECT 1884.690 243.820 1885.010 243.880 ;
        RECT 1890.210 243.820 1890.530 243.880 ;
        RECT 1890.210 16.900 1890.530 16.960 ;
        RECT 1995.090 16.900 1995.410 16.960 ;
        RECT 1890.210 16.760 1995.410 16.900 ;
        RECT 1890.210 16.700 1890.530 16.760 ;
        RECT 1995.090 16.700 1995.410 16.760 ;
      LAYER via ;
        RECT 1884.720 243.820 1884.980 244.080 ;
        RECT 1890.240 243.820 1890.500 244.080 ;
        RECT 1890.240 16.700 1890.500 16.960 ;
        RECT 1995.120 16.700 1995.380 16.960 ;
      LAYER met2 ;
        RECT 1884.670 260.000 1884.950 264.000 ;
        RECT 1884.780 244.110 1884.920 260.000 ;
        RECT 1884.720 243.790 1884.980 244.110 ;
        RECT 1890.240 243.790 1890.500 244.110 ;
        RECT 1890.300 16.990 1890.440 243.790 ;
        RECT 1890.240 16.670 1890.500 16.990 ;
        RECT 1995.120 16.670 1995.380 16.990 ;
        RECT 1995.180 2.400 1995.320 16.670 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1898.490 244.020 1898.810 244.080 ;
        RECT 1904.010 244.020 1904.330 244.080 ;
        RECT 1898.490 243.880 1904.330 244.020 ;
        RECT 1898.490 243.820 1898.810 243.880 ;
        RECT 1904.010 243.820 1904.330 243.880 ;
        RECT 1904.010 16.560 1904.330 16.620 ;
        RECT 2012.570 16.560 2012.890 16.620 ;
        RECT 1904.010 16.420 2012.890 16.560 ;
        RECT 1904.010 16.360 1904.330 16.420 ;
        RECT 2012.570 16.360 2012.890 16.420 ;
      LAYER via ;
        RECT 1898.520 243.820 1898.780 244.080 ;
        RECT 1904.040 243.820 1904.300 244.080 ;
        RECT 1904.040 16.360 1904.300 16.620 ;
        RECT 2012.600 16.360 2012.860 16.620 ;
      LAYER met2 ;
        RECT 1898.470 260.000 1898.750 264.000 ;
        RECT 1898.580 244.110 1898.720 260.000 ;
        RECT 1898.520 243.790 1898.780 244.110 ;
        RECT 1904.040 243.790 1904.300 244.110 ;
        RECT 1904.100 16.650 1904.240 243.790 ;
        RECT 1904.040 16.330 1904.300 16.650 ;
        RECT 2012.600 16.330 2012.860 16.650 ;
        RECT 2012.660 2.400 2012.800 16.330 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1912.750 244.020 1913.070 244.080 ;
        RECT 1917.350 244.020 1917.670 244.080 ;
        RECT 1912.750 243.880 1917.670 244.020 ;
        RECT 1912.750 243.820 1913.070 243.880 ;
        RECT 1917.350 243.820 1917.670 243.880 ;
        RECT 1917.350 19.960 1917.670 20.020 ;
        RECT 2030.510 19.960 2030.830 20.020 ;
        RECT 1917.350 19.820 2030.830 19.960 ;
        RECT 1917.350 19.760 1917.670 19.820 ;
        RECT 2030.510 19.760 2030.830 19.820 ;
      LAYER via ;
        RECT 1912.780 243.820 1913.040 244.080 ;
        RECT 1917.380 243.820 1917.640 244.080 ;
        RECT 1917.380 19.760 1917.640 20.020 ;
        RECT 2030.540 19.760 2030.800 20.020 ;
      LAYER met2 ;
        RECT 1912.730 260.000 1913.010 264.000 ;
        RECT 1912.840 244.110 1912.980 260.000 ;
        RECT 1912.780 243.790 1913.040 244.110 ;
        RECT 1917.380 243.790 1917.640 244.110 ;
        RECT 1917.440 20.050 1917.580 243.790 ;
        RECT 1917.380 19.730 1917.640 20.050 ;
        RECT 2030.540 19.730 2030.800 20.050 ;
        RECT 2030.600 2.400 2030.740 19.730 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1927.010 244.020 1927.330 244.080 ;
        RECT 1931.150 244.020 1931.470 244.080 ;
        RECT 1927.010 243.880 1931.470 244.020 ;
        RECT 1927.010 243.820 1927.330 243.880 ;
        RECT 1931.150 243.820 1931.470 243.880 ;
        RECT 1931.150 20.640 1931.470 20.700 ;
        RECT 2048.450 20.640 2048.770 20.700 ;
        RECT 1931.150 20.500 2048.770 20.640 ;
        RECT 1931.150 20.440 1931.470 20.500 ;
        RECT 2048.450 20.440 2048.770 20.500 ;
      LAYER via ;
        RECT 1927.040 243.820 1927.300 244.080 ;
        RECT 1931.180 243.820 1931.440 244.080 ;
        RECT 1931.180 20.440 1931.440 20.700 ;
        RECT 2048.480 20.440 2048.740 20.700 ;
      LAYER met2 ;
        RECT 1926.990 260.000 1927.270 264.000 ;
        RECT 1927.100 244.110 1927.240 260.000 ;
        RECT 1927.040 243.790 1927.300 244.110 ;
        RECT 1931.180 243.790 1931.440 244.110 ;
        RECT 1931.240 20.730 1931.380 243.790 ;
        RECT 1931.180 20.410 1931.440 20.730 ;
        RECT 2048.480 20.410 2048.740 20.730 ;
        RECT 2048.540 2.400 2048.680 20.410 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 810.665 16.745 810.835 18.955 ;
      LAYER mcon ;
        RECT 810.665 18.785 810.835 18.955 ;
      LAYER met1 ;
        RECT 810.605 18.940 810.895 18.985 ;
        RECT 910.870 18.940 911.190 19.000 ;
        RECT 810.605 18.800 911.190 18.940 ;
        RECT 810.605 18.755 810.895 18.800 ;
        RECT 910.870 18.740 911.190 18.800 ;
        RECT 763.670 16.900 763.990 16.960 ;
        RECT 810.605 16.900 810.895 16.945 ;
        RECT 763.670 16.760 810.895 16.900 ;
        RECT 763.670 16.700 763.990 16.760 ;
        RECT 810.605 16.715 810.895 16.760 ;
      LAYER via ;
        RECT 910.900 18.740 911.160 19.000 ;
        RECT 763.700 16.700 763.960 16.960 ;
      LAYER met2 ;
        RECT 913.150 260.170 913.430 264.000 ;
        RECT 910.960 260.030 913.430 260.170 ;
        RECT 910.960 19.030 911.100 260.030 ;
        RECT 913.150 260.000 913.430 260.030 ;
        RECT 910.900 18.710 911.160 19.030 ;
        RECT 763.700 16.670 763.960 16.990 ;
        RECT 763.760 2.400 763.900 16.670 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1940.810 244.020 1941.130 244.080 ;
        RECT 1945.410 244.020 1945.730 244.080 ;
        RECT 1940.810 243.880 1945.730 244.020 ;
        RECT 1940.810 243.820 1941.130 243.880 ;
        RECT 1945.410 243.820 1945.730 243.880 ;
        RECT 1945.410 19.280 1945.730 19.340 ;
        RECT 2066.390 19.280 2066.710 19.340 ;
        RECT 1945.410 19.140 2066.710 19.280 ;
        RECT 1945.410 19.080 1945.730 19.140 ;
        RECT 2066.390 19.080 2066.710 19.140 ;
      LAYER via ;
        RECT 1940.840 243.820 1941.100 244.080 ;
        RECT 1945.440 243.820 1945.700 244.080 ;
        RECT 1945.440 19.080 1945.700 19.340 ;
        RECT 2066.420 19.080 2066.680 19.340 ;
      LAYER met2 ;
        RECT 1940.790 260.000 1941.070 264.000 ;
        RECT 1940.900 244.110 1941.040 260.000 ;
        RECT 1940.840 243.790 1941.100 244.110 ;
        RECT 1945.440 243.790 1945.700 244.110 ;
        RECT 1945.500 19.370 1945.640 243.790 ;
        RECT 1945.440 19.050 1945.700 19.370 ;
        RECT 2066.420 19.050 2066.680 19.370 ;
        RECT 2066.480 2.400 2066.620 19.050 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1955.070 245.380 1955.390 245.440 ;
        RECT 2084.330 245.380 2084.650 245.440 ;
        RECT 1955.070 245.240 2084.650 245.380 ;
        RECT 1955.070 245.180 1955.390 245.240 ;
        RECT 2084.330 245.180 2084.650 245.240 ;
      LAYER via ;
        RECT 1955.100 245.180 1955.360 245.440 ;
        RECT 2084.360 245.180 2084.620 245.440 ;
      LAYER met2 ;
        RECT 1955.050 260.000 1955.330 264.000 ;
        RECT 1955.160 245.470 1955.300 260.000 ;
        RECT 1955.100 245.150 1955.360 245.470 ;
        RECT 2084.360 245.150 2084.620 245.470 ;
        RECT 2084.420 2.400 2084.560 245.150 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 79.460 1973.330 79.520 ;
        RECT 2097.670 79.460 2097.990 79.520 ;
        RECT 1973.010 79.320 2097.990 79.460 ;
        RECT 1973.010 79.260 1973.330 79.320 ;
        RECT 2097.670 79.260 2097.990 79.320 ;
      LAYER via ;
        RECT 1973.040 79.260 1973.300 79.520 ;
        RECT 2097.700 79.260 2097.960 79.520 ;
      LAYER met2 ;
        RECT 1969.310 260.170 1969.590 264.000 ;
        RECT 1969.310 260.030 1973.240 260.170 ;
        RECT 1969.310 260.000 1969.590 260.030 ;
        RECT 1973.100 79.550 1973.240 260.030 ;
        RECT 1973.040 79.230 1973.300 79.550 ;
        RECT 2097.700 79.230 2097.960 79.550 ;
        RECT 2097.760 17.410 2097.900 79.230 ;
        RECT 2097.760 17.270 2102.040 17.410 ;
        RECT 2101.900 2.400 2102.040 17.270 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1983.130 243.340 1983.450 243.400 ;
        RECT 1997.390 243.340 1997.710 243.400 ;
        RECT 1983.130 243.200 1997.710 243.340 ;
        RECT 1983.130 243.140 1983.450 243.200 ;
        RECT 1997.390 243.140 1997.710 243.200 ;
        RECT 1997.390 86.260 1997.710 86.320 ;
        RECT 2118.370 86.260 2118.690 86.320 ;
        RECT 1997.390 86.120 2118.690 86.260 ;
        RECT 1997.390 86.060 1997.710 86.120 ;
        RECT 2118.370 86.060 2118.690 86.120 ;
      LAYER via ;
        RECT 1983.160 243.140 1983.420 243.400 ;
        RECT 1997.420 243.140 1997.680 243.400 ;
        RECT 1997.420 86.060 1997.680 86.320 ;
        RECT 2118.400 86.060 2118.660 86.320 ;
      LAYER met2 ;
        RECT 1983.110 260.000 1983.390 264.000 ;
        RECT 1983.220 243.430 1983.360 260.000 ;
        RECT 1983.160 243.110 1983.420 243.430 ;
        RECT 1997.420 243.110 1997.680 243.430 ;
        RECT 1997.480 86.350 1997.620 243.110 ;
        RECT 1997.420 86.030 1997.680 86.350 ;
        RECT 2118.400 86.030 2118.660 86.350 ;
        RECT 2118.460 16.730 2118.600 86.030 ;
        RECT 2118.460 16.590 2119.980 16.730 ;
        RECT 2119.840 2.400 2119.980 16.590 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2000.610 93.060 2000.930 93.120 ;
        RECT 2132.170 93.060 2132.490 93.120 ;
        RECT 2000.610 92.920 2132.490 93.060 ;
        RECT 2000.610 92.860 2000.930 92.920 ;
        RECT 2132.170 92.860 2132.490 92.920 ;
      LAYER via ;
        RECT 2000.640 92.860 2000.900 93.120 ;
        RECT 2132.200 92.860 2132.460 93.120 ;
      LAYER met2 ;
        RECT 1997.370 260.170 1997.650 264.000 ;
        RECT 1997.370 260.030 2000.840 260.170 ;
        RECT 1997.370 260.000 1997.650 260.030 ;
        RECT 2000.700 93.150 2000.840 260.030 ;
        RECT 2000.640 92.830 2000.900 93.150 ;
        RECT 2132.200 92.830 2132.460 93.150 ;
        RECT 2132.260 16.730 2132.400 92.830 ;
        RECT 2132.260 16.590 2137.920 16.730 ;
        RECT 2137.780 2.400 2137.920 16.590 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2014.410 113.800 2014.730 113.860 ;
        RECT 2152.870 113.800 2153.190 113.860 ;
        RECT 2014.410 113.660 2153.190 113.800 ;
        RECT 2014.410 113.600 2014.730 113.660 ;
        RECT 2152.870 113.600 2153.190 113.660 ;
      LAYER via ;
        RECT 2014.440 113.600 2014.700 113.860 ;
        RECT 2152.900 113.600 2153.160 113.860 ;
      LAYER met2 ;
        RECT 2011.170 260.170 2011.450 264.000 ;
        RECT 2011.170 260.030 2014.640 260.170 ;
        RECT 2011.170 260.000 2011.450 260.030 ;
        RECT 2014.500 113.890 2014.640 260.030 ;
        RECT 2014.440 113.570 2014.700 113.890 ;
        RECT 2152.900 113.570 2153.160 113.890 ;
        RECT 2152.960 16.730 2153.100 113.570 ;
        RECT 2152.960 16.590 2155.860 16.730 ;
        RECT 2155.720 2.400 2155.860 16.590 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2028.210 99.860 2028.530 99.920 ;
        RECT 2166.670 99.860 2166.990 99.920 ;
        RECT 2028.210 99.720 2166.990 99.860 ;
        RECT 2028.210 99.660 2028.530 99.720 ;
        RECT 2166.670 99.660 2166.990 99.720 ;
        RECT 2166.670 17.240 2166.990 17.300 ;
        RECT 2173.110 17.240 2173.430 17.300 ;
        RECT 2166.670 17.100 2173.430 17.240 ;
        RECT 2166.670 17.040 2166.990 17.100 ;
        RECT 2173.110 17.040 2173.430 17.100 ;
      LAYER via ;
        RECT 2028.240 99.660 2028.500 99.920 ;
        RECT 2166.700 99.660 2166.960 99.920 ;
        RECT 2166.700 17.040 2166.960 17.300 ;
        RECT 2173.140 17.040 2173.400 17.300 ;
      LAYER met2 ;
        RECT 2025.430 260.170 2025.710 264.000 ;
        RECT 2025.430 260.030 2028.440 260.170 ;
        RECT 2025.430 260.000 2025.710 260.030 ;
        RECT 2028.300 99.950 2028.440 260.030 ;
        RECT 2028.240 99.630 2028.500 99.950 ;
        RECT 2166.700 99.630 2166.960 99.950 ;
        RECT 2166.760 17.330 2166.900 99.630 ;
        RECT 2166.700 17.010 2166.960 17.330 ;
        RECT 2173.140 17.010 2173.400 17.330 ;
        RECT 2173.200 2.400 2173.340 17.010 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2039.710 243.680 2040.030 243.740 ;
        RECT 2052.590 243.680 2052.910 243.740 ;
        RECT 2039.710 243.540 2052.910 243.680 ;
        RECT 2039.710 243.480 2040.030 243.540 ;
        RECT 2052.590 243.480 2052.910 243.540 ;
        RECT 2052.590 107.000 2052.910 107.060 ;
        RECT 2187.370 107.000 2187.690 107.060 ;
        RECT 2052.590 106.860 2187.690 107.000 ;
        RECT 2052.590 106.800 2052.910 106.860 ;
        RECT 2187.370 106.800 2187.690 106.860 ;
        RECT 2187.370 2.960 2187.690 3.020 ;
        RECT 2191.050 2.960 2191.370 3.020 ;
        RECT 2187.370 2.820 2191.370 2.960 ;
        RECT 2187.370 2.760 2187.690 2.820 ;
        RECT 2191.050 2.760 2191.370 2.820 ;
      LAYER via ;
        RECT 2039.740 243.480 2040.000 243.740 ;
        RECT 2052.620 243.480 2052.880 243.740 ;
        RECT 2052.620 106.800 2052.880 107.060 ;
        RECT 2187.400 106.800 2187.660 107.060 ;
        RECT 2187.400 2.760 2187.660 3.020 ;
        RECT 2191.080 2.760 2191.340 3.020 ;
      LAYER met2 ;
        RECT 2039.690 260.000 2039.970 264.000 ;
        RECT 2039.800 243.770 2039.940 260.000 ;
        RECT 2039.740 243.450 2040.000 243.770 ;
        RECT 2052.620 243.450 2052.880 243.770 ;
        RECT 2052.680 107.090 2052.820 243.450 ;
        RECT 2052.620 106.770 2052.880 107.090 ;
        RECT 2187.400 106.770 2187.660 107.090 ;
        RECT 2187.460 3.050 2187.600 106.770 ;
        RECT 2187.400 2.730 2187.660 3.050 ;
        RECT 2191.080 2.730 2191.340 3.050 ;
        RECT 2191.140 2.400 2191.280 2.730 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2055.810 120.600 2056.130 120.660 ;
        RECT 2208.070 120.600 2208.390 120.660 ;
        RECT 2055.810 120.460 2208.390 120.600 ;
        RECT 2055.810 120.400 2056.130 120.460 ;
        RECT 2208.070 120.400 2208.390 120.460 ;
        RECT 2208.070 2.960 2208.390 3.020 ;
        RECT 2208.990 2.960 2209.310 3.020 ;
        RECT 2208.070 2.820 2209.310 2.960 ;
        RECT 2208.070 2.760 2208.390 2.820 ;
        RECT 2208.990 2.760 2209.310 2.820 ;
      LAYER via ;
        RECT 2055.840 120.400 2056.100 120.660 ;
        RECT 2208.100 120.400 2208.360 120.660 ;
        RECT 2208.100 2.760 2208.360 3.020 ;
        RECT 2209.020 2.760 2209.280 3.020 ;
      LAYER met2 ;
        RECT 2053.490 260.170 2053.770 264.000 ;
        RECT 2053.490 260.030 2056.040 260.170 ;
        RECT 2053.490 260.000 2053.770 260.030 ;
        RECT 2055.900 120.690 2056.040 260.030 ;
        RECT 2055.840 120.370 2056.100 120.690 ;
        RECT 2208.100 120.370 2208.360 120.690 ;
        RECT 2208.160 3.050 2208.300 120.370 ;
        RECT 2208.100 2.730 2208.360 3.050 ;
        RECT 2209.020 2.730 2209.280 3.050 ;
        RECT 2209.080 2.400 2209.220 2.730 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2069.150 127.740 2069.470 127.800 ;
        RECT 2221.870 127.740 2222.190 127.800 ;
        RECT 2069.150 127.600 2222.190 127.740 ;
        RECT 2069.150 127.540 2069.470 127.600 ;
        RECT 2221.870 127.540 2222.190 127.600 ;
        RECT 2221.870 2.960 2222.190 3.020 ;
        RECT 2226.930 2.960 2227.250 3.020 ;
        RECT 2221.870 2.820 2227.250 2.960 ;
        RECT 2221.870 2.760 2222.190 2.820 ;
        RECT 2226.930 2.760 2227.250 2.820 ;
      LAYER via ;
        RECT 2069.180 127.540 2069.440 127.800 ;
        RECT 2221.900 127.540 2222.160 127.800 ;
        RECT 2221.900 2.760 2222.160 3.020 ;
        RECT 2226.960 2.760 2227.220 3.020 ;
      LAYER met2 ;
        RECT 2067.750 260.170 2068.030 264.000 ;
        RECT 2067.750 260.030 2069.380 260.170 ;
        RECT 2067.750 260.000 2068.030 260.030 ;
        RECT 2069.240 127.830 2069.380 260.030 ;
        RECT 2069.180 127.510 2069.440 127.830 ;
        RECT 2221.900 127.510 2222.160 127.830 ;
        RECT 2221.960 3.050 2222.100 127.510 ;
        RECT 2221.900 2.730 2222.160 3.050 ;
        RECT 2226.960 2.730 2227.220 3.050 ;
        RECT 2227.020 2.400 2227.160 2.730 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 781.610 19.960 781.930 20.020 ;
        RECT 924.670 19.960 924.990 20.020 ;
        RECT 781.610 19.820 924.990 19.960 ;
        RECT 781.610 19.760 781.930 19.820 ;
        RECT 924.670 19.760 924.990 19.820 ;
      LAYER via ;
        RECT 781.640 19.760 781.900 20.020 ;
        RECT 924.700 19.760 924.960 20.020 ;
      LAYER met2 ;
        RECT 926.950 260.170 927.230 264.000 ;
        RECT 924.760 260.030 927.230 260.170 ;
        RECT 924.760 20.050 924.900 260.030 ;
        RECT 926.950 260.000 927.230 260.030 ;
        RECT 781.640 19.730 781.900 20.050 ;
        RECT 924.700 19.730 924.960 20.050 ;
        RECT 781.700 2.400 781.840 19.730 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2082.950 134.540 2083.270 134.600 ;
        RECT 2242.570 134.540 2242.890 134.600 ;
        RECT 2082.950 134.400 2242.890 134.540 ;
        RECT 2082.950 134.340 2083.270 134.400 ;
        RECT 2242.570 134.340 2242.890 134.400 ;
        RECT 2242.570 2.960 2242.890 3.020 ;
        RECT 2244.870 2.960 2245.190 3.020 ;
        RECT 2242.570 2.820 2245.190 2.960 ;
        RECT 2242.570 2.760 2242.890 2.820 ;
        RECT 2244.870 2.760 2245.190 2.820 ;
      LAYER via ;
        RECT 2082.980 134.340 2083.240 134.600 ;
        RECT 2242.600 134.340 2242.860 134.600 ;
        RECT 2242.600 2.760 2242.860 3.020 ;
        RECT 2244.900 2.760 2245.160 3.020 ;
      LAYER met2 ;
        RECT 2081.550 260.170 2081.830 264.000 ;
        RECT 2081.550 260.030 2083.180 260.170 ;
        RECT 2081.550 260.000 2081.830 260.030 ;
        RECT 2083.040 134.630 2083.180 260.030 ;
        RECT 2082.980 134.310 2083.240 134.630 ;
        RECT 2242.600 134.310 2242.860 134.630 ;
        RECT 2242.660 3.050 2242.800 134.310 ;
        RECT 2242.600 2.730 2242.860 3.050 ;
        RECT 2244.900 2.730 2245.160 3.050 ;
        RECT 2244.960 2.400 2245.100 2.730 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2095.830 246.740 2096.150 246.800 ;
        RECT 2114.690 246.740 2115.010 246.800 ;
        RECT 2095.830 246.600 2115.010 246.740 ;
        RECT 2095.830 246.540 2096.150 246.600 ;
        RECT 2114.690 246.540 2115.010 246.600 ;
        RECT 2114.690 141.340 2115.010 141.400 ;
        RECT 2256.370 141.340 2256.690 141.400 ;
        RECT 2114.690 141.200 2256.690 141.340 ;
        RECT 2114.690 141.140 2115.010 141.200 ;
        RECT 2256.370 141.140 2256.690 141.200 ;
        RECT 2256.370 18.600 2256.690 18.660 ;
        RECT 2262.350 18.600 2262.670 18.660 ;
        RECT 2256.370 18.460 2262.670 18.600 ;
        RECT 2256.370 18.400 2256.690 18.460 ;
        RECT 2262.350 18.400 2262.670 18.460 ;
      LAYER via ;
        RECT 2095.860 246.540 2096.120 246.800 ;
        RECT 2114.720 246.540 2114.980 246.800 ;
        RECT 2114.720 141.140 2114.980 141.400 ;
        RECT 2256.400 141.140 2256.660 141.400 ;
        RECT 2256.400 18.400 2256.660 18.660 ;
        RECT 2262.380 18.400 2262.640 18.660 ;
      LAYER met2 ;
        RECT 2095.810 260.000 2096.090 264.000 ;
        RECT 2095.920 246.830 2096.060 260.000 ;
        RECT 2095.860 246.510 2096.120 246.830 ;
        RECT 2114.720 246.510 2114.980 246.830 ;
        RECT 2114.780 141.430 2114.920 246.510 ;
        RECT 2114.720 141.110 2114.980 141.430 ;
        RECT 2256.400 141.110 2256.660 141.430 ;
        RECT 2256.460 18.690 2256.600 141.110 ;
        RECT 2256.400 18.370 2256.660 18.690 ;
        RECT 2262.380 18.370 2262.640 18.690 ;
        RECT 2262.440 2.400 2262.580 18.370 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2110.550 148.140 2110.870 148.200 ;
        RECT 2277.070 148.140 2277.390 148.200 ;
        RECT 2110.550 148.000 2277.390 148.140 ;
        RECT 2110.550 147.940 2110.870 148.000 ;
        RECT 2277.070 147.940 2277.390 148.000 ;
      LAYER via ;
        RECT 2110.580 147.940 2110.840 148.200 ;
        RECT 2277.100 147.940 2277.360 148.200 ;
      LAYER met2 ;
        RECT 2110.070 260.170 2110.350 264.000 ;
        RECT 2110.070 260.030 2110.780 260.170 ;
        RECT 2110.070 260.000 2110.350 260.030 ;
        RECT 2110.640 148.230 2110.780 260.030 ;
        RECT 2110.580 147.910 2110.840 148.230 ;
        RECT 2277.100 147.910 2277.360 148.230 ;
        RECT 2277.160 16.730 2277.300 147.910 ;
        RECT 2277.160 16.590 2280.520 16.730 ;
        RECT 2280.380 2.400 2280.520 16.590 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.810 72.320 2125.130 72.380 ;
        RECT 2298.230 72.320 2298.550 72.380 ;
        RECT 2124.810 72.180 2298.550 72.320 ;
        RECT 2124.810 72.120 2125.130 72.180 ;
        RECT 2298.230 72.120 2298.550 72.180 ;
      LAYER via ;
        RECT 2124.840 72.120 2125.100 72.380 ;
        RECT 2298.260 72.120 2298.520 72.380 ;
      LAYER met2 ;
        RECT 2123.870 260.170 2124.150 264.000 ;
        RECT 2123.870 260.030 2125.040 260.170 ;
        RECT 2123.870 260.000 2124.150 260.030 ;
        RECT 2124.900 72.410 2125.040 260.030 ;
        RECT 2124.840 72.090 2125.100 72.410 ;
        RECT 2298.260 72.090 2298.520 72.410 ;
        RECT 2298.320 2.400 2298.460 72.090 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.610 155.280 2138.930 155.340 ;
        RECT 2311.570 155.280 2311.890 155.340 ;
        RECT 2138.610 155.140 2311.890 155.280 ;
        RECT 2138.610 155.080 2138.930 155.140 ;
        RECT 2311.570 155.080 2311.890 155.140 ;
      LAYER via ;
        RECT 2138.640 155.080 2138.900 155.340 ;
        RECT 2311.600 155.080 2311.860 155.340 ;
      LAYER met2 ;
        RECT 2138.130 260.170 2138.410 264.000 ;
        RECT 2138.130 260.030 2138.840 260.170 ;
        RECT 2138.130 260.000 2138.410 260.030 ;
        RECT 2138.700 155.370 2138.840 260.030 ;
        RECT 2138.640 155.050 2138.900 155.370 ;
        RECT 2311.600 155.050 2311.860 155.370 ;
        RECT 2311.660 16.730 2311.800 155.050 ;
        RECT 2311.660 16.590 2316.400 16.730 ;
        RECT 2316.260 2.400 2316.400 16.590 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2151.950 162.080 2152.270 162.140 ;
        RECT 2332.270 162.080 2332.590 162.140 ;
        RECT 2151.950 161.940 2332.590 162.080 ;
        RECT 2151.950 161.880 2152.270 161.940 ;
        RECT 2332.270 161.880 2332.590 161.940 ;
      LAYER via ;
        RECT 2151.980 161.880 2152.240 162.140 ;
        RECT 2332.300 161.880 2332.560 162.140 ;
      LAYER met2 ;
        RECT 2152.390 260.170 2152.670 264.000 ;
        RECT 2152.040 260.030 2152.670 260.170 ;
        RECT 2152.040 162.170 2152.180 260.030 ;
        RECT 2152.390 260.000 2152.670 260.030 ;
        RECT 2151.980 161.850 2152.240 162.170 ;
        RECT 2332.300 161.850 2332.560 162.170 ;
        RECT 2332.360 16.730 2332.500 161.850 ;
        RECT 2332.360 16.590 2334.340 16.730 ;
        RECT 2334.200 2.400 2334.340 16.590 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2166.210 168.880 2166.530 168.940 ;
        RECT 2346.070 168.880 2346.390 168.940 ;
        RECT 2166.210 168.740 2346.390 168.880 ;
        RECT 2166.210 168.680 2166.530 168.740 ;
        RECT 2346.070 168.680 2346.390 168.740 ;
      LAYER via ;
        RECT 2166.240 168.680 2166.500 168.940 ;
        RECT 2346.100 168.680 2346.360 168.940 ;
      LAYER met2 ;
        RECT 2166.190 260.000 2166.470 264.000 ;
        RECT 2166.300 168.970 2166.440 260.000 ;
        RECT 2166.240 168.650 2166.500 168.970 ;
        RECT 2346.100 168.650 2346.360 168.970 ;
        RECT 2346.160 16.730 2346.300 168.650 ;
        RECT 2346.160 16.590 2351.820 16.730 ;
        RECT 2351.680 2.400 2351.820 16.590 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2180.470 244.020 2180.790 244.080 ;
        RECT 2186.450 244.020 2186.770 244.080 ;
        RECT 2180.470 243.880 2186.770 244.020 ;
        RECT 2180.470 243.820 2180.790 243.880 ;
        RECT 2186.450 243.820 2186.770 243.880 ;
        RECT 2186.450 17.240 2186.770 17.300 ;
        RECT 2369.530 17.240 2369.850 17.300 ;
        RECT 2186.450 17.100 2369.850 17.240 ;
        RECT 2186.450 17.040 2186.770 17.100 ;
        RECT 2369.530 17.040 2369.850 17.100 ;
      LAYER via ;
        RECT 2180.500 243.820 2180.760 244.080 ;
        RECT 2186.480 243.820 2186.740 244.080 ;
        RECT 2186.480 17.040 2186.740 17.300 ;
        RECT 2369.560 17.040 2369.820 17.300 ;
      LAYER met2 ;
        RECT 2180.450 260.000 2180.730 264.000 ;
        RECT 2180.560 244.110 2180.700 260.000 ;
        RECT 2180.500 243.790 2180.760 244.110 ;
        RECT 2186.480 243.790 2186.740 244.110 ;
        RECT 2186.540 17.330 2186.680 243.790 ;
        RECT 2186.480 17.010 2186.740 17.330 ;
        RECT 2369.560 17.010 2369.820 17.330 ;
        RECT 2369.620 2.400 2369.760 17.010 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2194.270 244.020 2194.590 244.080 ;
        RECT 2200.710 244.020 2201.030 244.080 ;
        RECT 2194.270 243.880 2201.030 244.020 ;
        RECT 2194.270 243.820 2194.590 243.880 ;
        RECT 2200.710 243.820 2201.030 243.880 ;
        RECT 2200.710 16.560 2201.030 16.620 ;
        RECT 2387.470 16.560 2387.790 16.620 ;
        RECT 2200.710 16.420 2387.790 16.560 ;
        RECT 2200.710 16.360 2201.030 16.420 ;
        RECT 2387.470 16.360 2387.790 16.420 ;
      LAYER via ;
        RECT 2194.300 243.820 2194.560 244.080 ;
        RECT 2200.740 243.820 2201.000 244.080 ;
        RECT 2200.740 16.360 2201.000 16.620 ;
        RECT 2387.500 16.360 2387.760 16.620 ;
      LAYER met2 ;
        RECT 2194.250 260.000 2194.530 264.000 ;
        RECT 2194.360 244.110 2194.500 260.000 ;
        RECT 2194.300 243.790 2194.560 244.110 ;
        RECT 2200.740 243.790 2201.000 244.110 ;
        RECT 2200.800 16.650 2200.940 243.790 ;
        RECT 2200.740 16.330 2201.000 16.650 ;
        RECT 2387.500 16.330 2387.760 16.650 ;
        RECT 2387.560 2.400 2387.700 16.330 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2208.530 244.020 2208.850 244.080 ;
        RECT 2214.050 244.020 2214.370 244.080 ;
        RECT 2208.530 243.880 2214.370 244.020 ;
        RECT 2208.530 243.820 2208.850 243.880 ;
        RECT 2214.050 243.820 2214.370 243.880 ;
        RECT 2214.050 20.640 2214.370 20.700 ;
        RECT 2405.410 20.640 2405.730 20.700 ;
        RECT 2214.050 20.500 2405.730 20.640 ;
        RECT 2214.050 20.440 2214.370 20.500 ;
        RECT 2405.410 20.440 2405.730 20.500 ;
      LAYER via ;
        RECT 2208.560 243.820 2208.820 244.080 ;
        RECT 2214.080 243.820 2214.340 244.080 ;
        RECT 2214.080 20.440 2214.340 20.700 ;
        RECT 2405.440 20.440 2405.700 20.700 ;
      LAYER met2 ;
        RECT 2208.510 260.000 2208.790 264.000 ;
        RECT 2208.620 244.110 2208.760 260.000 ;
        RECT 2208.560 243.790 2208.820 244.110 ;
        RECT 2214.080 243.790 2214.340 244.110 ;
        RECT 2214.140 20.730 2214.280 243.790 ;
        RECT 2214.080 20.410 2214.340 20.730 ;
        RECT 2405.440 20.410 2405.700 20.730 ;
        RECT 2405.500 2.400 2405.640 20.410 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 800.010 245.720 800.330 245.780 ;
        RECT 941.230 245.720 941.550 245.780 ;
        RECT 800.010 245.580 941.550 245.720 ;
        RECT 800.010 245.520 800.330 245.580 ;
        RECT 941.230 245.520 941.550 245.580 ;
      LAYER via ;
        RECT 800.040 245.520 800.300 245.780 ;
        RECT 941.260 245.520 941.520 245.780 ;
      LAYER met2 ;
        RECT 941.210 260.000 941.490 264.000 ;
        RECT 941.320 245.810 941.460 260.000 ;
        RECT 800.040 245.490 800.300 245.810 ;
        RECT 941.260 245.490 941.520 245.810 ;
        RECT 800.100 20.130 800.240 245.490 ;
        RECT 799.640 19.990 800.240 20.130 ;
        RECT 799.640 2.400 799.780 19.990 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 217.160 648.530 217.220 ;
        RECT 814.730 217.160 815.050 217.220 ;
        RECT 648.210 217.020 815.050 217.160 ;
        RECT 648.210 216.960 648.530 217.020 ;
        RECT 814.730 216.960 815.050 217.020 ;
        RECT 644.990 17.580 645.310 17.640 ;
        RECT 648.210 17.580 648.530 17.640 ;
        RECT 644.990 17.440 648.530 17.580 ;
        RECT 644.990 17.380 645.310 17.440 ;
        RECT 648.210 17.380 648.530 17.440 ;
      LAYER via ;
        RECT 648.240 216.960 648.500 217.220 ;
        RECT 814.760 216.960 815.020 217.220 ;
        RECT 645.020 17.380 645.280 17.640 ;
        RECT 648.240 17.380 648.500 17.640 ;
      LAYER met2 ;
        RECT 819.310 260.170 819.590 264.000 ;
        RECT 814.820 260.030 819.590 260.170 ;
        RECT 814.820 217.250 814.960 260.030 ;
        RECT 819.310 260.000 819.590 260.030 ;
        RECT 648.240 216.930 648.500 217.250 ;
        RECT 814.760 216.930 815.020 217.250 ;
        RECT 648.300 17.670 648.440 216.930 ;
        RECT 645.020 17.350 645.280 17.670 ;
        RECT 648.240 17.350 648.500 17.670 ;
        RECT 645.080 2.400 645.220 17.350 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2228.310 19.620 2228.630 19.680 ;
        RECT 2428.870 19.620 2429.190 19.680 ;
        RECT 2228.310 19.480 2429.190 19.620 ;
        RECT 2228.310 19.420 2228.630 19.480 ;
        RECT 2428.870 19.420 2429.190 19.480 ;
      LAYER via ;
        RECT 2228.340 19.420 2228.600 19.680 ;
        RECT 2428.900 19.420 2429.160 19.680 ;
      LAYER met2 ;
        RECT 2227.370 260.170 2227.650 264.000 ;
        RECT 2227.370 260.030 2228.540 260.170 ;
        RECT 2227.370 260.000 2227.650 260.030 ;
        RECT 2228.400 19.710 2228.540 260.030 ;
        RECT 2228.340 19.390 2228.600 19.710 ;
        RECT 2428.900 19.390 2429.160 19.710 ;
        RECT 2428.960 2.400 2429.100 19.390 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2241.650 19.960 2241.970 20.020 ;
        RECT 2446.810 19.960 2447.130 20.020 ;
        RECT 2241.650 19.820 2447.130 19.960 ;
        RECT 2241.650 19.760 2241.970 19.820 ;
        RECT 2446.810 19.760 2447.130 19.820 ;
      LAYER via ;
        RECT 2241.680 19.760 2241.940 20.020 ;
        RECT 2446.840 19.760 2447.100 20.020 ;
      LAYER met2 ;
        RECT 2241.170 260.170 2241.450 264.000 ;
        RECT 2241.170 260.030 2241.880 260.170 ;
        RECT 2241.170 260.000 2241.450 260.030 ;
        RECT 2241.740 20.050 2241.880 260.030 ;
        RECT 2241.680 19.730 2241.940 20.050 ;
        RECT 2446.840 19.730 2447.100 20.050 ;
        RECT 2446.900 2.400 2447.040 19.730 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2255.910 19.280 2256.230 19.340 ;
        RECT 2464.750 19.280 2465.070 19.340 ;
        RECT 2255.910 19.140 2465.070 19.280 ;
        RECT 2255.910 19.080 2256.230 19.140 ;
        RECT 2464.750 19.080 2465.070 19.140 ;
      LAYER via ;
        RECT 2255.940 19.080 2256.200 19.340 ;
        RECT 2464.780 19.080 2465.040 19.340 ;
      LAYER met2 ;
        RECT 2255.430 260.170 2255.710 264.000 ;
        RECT 2255.430 260.030 2256.140 260.170 ;
        RECT 2255.430 260.000 2255.710 260.030 ;
        RECT 2256.000 19.370 2256.140 260.030 ;
        RECT 2255.940 19.050 2256.200 19.370 ;
        RECT 2464.780 19.050 2465.040 19.370 ;
        RECT 2464.840 2.400 2464.980 19.050 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 18.600 2270.030 18.660 ;
        RECT 2482.690 18.600 2483.010 18.660 ;
        RECT 2269.710 18.460 2483.010 18.600 ;
        RECT 2269.710 18.400 2270.030 18.460 ;
        RECT 2482.690 18.400 2483.010 18.460 ;
      LAYER via ;
        RECT 2269.740 18.400 2270.000 18.660 ;
        RECT 2482.720 18.400 2482.980 18.660 ;
      LAYER met2 ;
        RECT 2269.690 260.000 2269.970 264.000 ;
        RECT 2269.800 18.690 2269.940 260.000 ;
        RECT 2269.740 18.370 2270.000 18.690 ;
        RECT 2482.720 18.370 2482.980 18.690 ;
        RECT 2482.780 2.400 2482.920 18.370 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2283.490 260.000 2283.770 264.000 ;
        RECT 2283.600 16.845 2283.740 260.000 ;
        RECT 2283.530 16.475 2283.810 16.845 ;
        RECT 2500.650 16.475 2500.930 16.845 ;
        RECT 2500.720 2.400 2500.860 16.475 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
      LAYER via2 ;
        RECT 2283.530 16.520 2283.810 16.800 ;
        RECT 2500.650 16.520 2500.930 16.800 ;
      LAYER met3 ;
        RECT 2283.505 16.810 2283.835 16.825 ;
        RECT 2500.625 16.810 2500.955 16.825 ;
        RECT 2283.505 16.510 2500.955 16.810 ;
        RECT 2283.505 16.495 2283.835 16.510 ;
        RECT 2500.625 16.495 2500.955 16.510 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2297.770 244.020 2298.090 244.080 ;
        RECT 2304.210 244.020 2304.530 244.080 ;
        RECT 2297.770 243.880 2304.530 244.020 ;
        RECT 2297.770 243.820 2298.090 243.880 ;
        RECT 2304.210 243.820 2304.530 243.880 ;
        RECT 2304.210 18.940 2304.530 19.000 ;
        RECT 2518.110 18.940 2518.430 19.000 ;
        RECT 2304.210 18.800 2518.430 18.940 ;
        RECT 2304.210 18.740 2304.530 18.800 ;
        RECT 2518.110 18.740 2518.430 18.800 ;
      LAYER via ;
        RECT 2297.800 243.820 2298.060 244.080 ;
        RECT 2304.240 243.820 2304.500 244.080 ;
        RECT 2304.240 18.740 2304.500 19.000 ;
        RECT 2518.140 18.740 2518.400 19.000 ;
      LAYER met2 ;
        RECT 2297.750 260.000 2298.030 264.000 ;
        RECT 2297.860 244.110 2298.000 260.000 ;
        RECT 2297.800 243.790 2298.060 244.110 ;
        RECT 2304.240 243.790 2304.500 244.110 ;
        RECT 2304.300 19.030 2304.440 243.790 ;
        RECT 2304.240 18.710 2304.500 19.030 ;
        RECT 2518.140 18.710 2518.400 19.030 ;
        RECT 2518.200 2.400 2518.340 18.710 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2344.765 17.765 2346.775 17.935 ;
      LAYER mcon ;
        RECT 2346.605 17.765 2346.775 17.935 ;
      LAYER met1 ;
        RECT 2311.570 244.020 2311.890 244.080 ;
        RECT 2318.010 244.020 2318.330 244.080 ;
        RECT 2311.570 243.880 2318.330 244.020 ;
        RECT 2311.570 243.820 2311.890 243.880 ;
        RECT 2318.010 243.820 2318.330 243.880 ;
        RECT 2318.010 17.920 2318.330 17.980 ;
        RECT 2344.705 17.920 2344.995 17.965 ;
        RECT 2318.010 17.780 2344.995 17.920 ;
        RECT 2318.010 17.720 2318.330 17.780 ;
        RECT 2344.705 17.735 2344.995 17.780 ;
        RECT 2346.545 17.920 2346.835 17.965 ;
        RECT 2536.050 17.920 2536.370 17.980 ;
        RECT 2346.545 17.780 2536.370 17.920 ;
        RECT 2346.545 17.735 2346.835 17.780 ;
        RECT 2536.050 17.720 2536.370 17.780 ;
      LAYER via ;
        RECT 2311.600 243.820 2311.860 244.080 ;
        RECT 2318.040 243.820 2318.300 244.080 ;
        RECT 2318.040 17.720 2318.300 17.980 ;
        RECT 2536.080 17.720 2536.340 17.980 ;
      LAYER met2 ;
        RECT 2311.550 260.000 2311.830 264.000 ;
        RECT 2311.660 244.110 2311.800 260.000 ;
        RECT 2311.600 243.790 2311.860 244.110 ;
        RECT 2318.040 243.790 2318.300 244.110 ;
        RECT 2318.100 18.010 2318.240 243.790 ;
        RECT 2318.040 17.690 2318.300 18.010 ;
        RECT 2536.080 17.690 2536.340 18.010 ;
        RECT 2536.140 2.400 2536.280 17.690 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2325.830 246.740 2326.150 246.800 ;
        RECT 2553.530 246.740 2553.850 246.800 ;
        RECT 2325.830 246.600 2553.850 246.740 ;
        RECT 2325.830 246.540 2326.150 246.600 ;
        RECT 2553.530 246.540 2553.850 246.600 ;
      LAYER via ;
        RECT 2325.860 246.540 2326.120 246.800 ;
        RECT 2553.560 246.540 2553.820 246.800 ;
      LAYER met2 ;
        RECT 2325.810 260.000 2326.090 264.000 ;
        RECT 2325.920 246.830 2326.060 260.000 ;
        RECT 2325.860 246.510 2326.120 246.830 ;
        RECT 2553.560 246.510 2553.820 246.830 ;
        RECT 2553.620 17.410 2553.760 246.510 ;
        RECT 2553.620 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2340.090 244.020 2340.410 244.080 ;
        RECT 2345.610 244.020 2345.930 244.080 ;
        RECT 2340.090 243.880 2345.930 244.020 ;
        RECT 2340.090 243.820 2340.410 243.880 ;
        RECT 2345.610 243.820 2345.930 243.880 ;
        RECT 2345.150 17.920 2345.470 17.980 ;
        RECT 2345.150 17.780 2346.300 17.920 ;
        RECT 2345.150 17.720 2345.470 17.780 ;
        RECT 2346.160 17.580 2346.300 17.780 ;
        RECT 2571.930 17.580 2572.250 17.640 ;
        RECT 2346.160 17.440 2572.250 17.580 ;
        RECT 2571.930 17.380 2572.250 17.440 ;
      LAYER via ;
        RECT 2340.120 243.820 2340.380 244.080 ;
        RECT 2345.640 243.820 2345.900 244.080 ;
        RECT 2345.180 17.720 2345.440 17.980 ;
        RECT 2571.960 17.380 2572.220 17.640 ;
      LAYER met2 ;
        RECT 2340.070 260.000 2340.350 264.000 ;
        RECT 2340.180 244.110 2340.320 260.000 ;
        RECT 2340.120 243.790 2340.380 244.110 ;
        RECT 2345.640 243.790 2345.900 244.110 ;
        RECT 2345.700 26.250 2345.840 243.790 ;
        RECT 2345.240 26.110 2345.840 26.250 ;
        RECT 2345.240 18.010 2345.380 26.110 ;
        RECT 2345.180 17.690 2345.440 18.010 ;
        RECT 2571.960 17.350 2572.220 17.670 ;
        RECT 2572.020 2.400 2572.160 17.350 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2353.890 244.020 2354.210 244.080 ;
        RECT 2359.410 244.020 2359.730 244.080 ;
        RECT 2353.890 243.880 2359.730 244.020 ;
        RECT 2353.890 243.820 2354.210 243.880 ;
        RECT 2359.410 243.820 2359.730 243.880 ;
        RECT 2359.410 18.260 2359.730 18.320 ;
        RECT 2589.410 18.260 2589.730 18.320 ;
        RECT 2359.410 18.120 2589.730 18.260 ;
        RECT 2359.410 18.060 2359.730 18.120 ;
        RECT 2589.410 18.060 2589.730 18.120 ;
      LAYER via ;
        RECT 2353.920 243.820 2354.180 244.080 ;
        RECT 2359.440 243.820 2359.700 244.080 ;
        RECT 2359.440 18.060 2359.700 18.320 ;
        RECT 2589.440 18.060 2589.700 18.320 ;
      LAYER met2 ;
        RECT 2353.870 260.000 2354.150 264.000 ;
        RECT 2353.980 244.110 2354.120 260.000 ;
        RECT 2353.920 243.790 2354.180 244.110 ;
        RECT 2359.440 243.790 2359.700 244.110 ;
        RECT 2359.500 18.350 2359.640 243.790 ;
        RECT 2359.440 18.030 2359.700 18.350 ;
        RECT 2589.440 18.030 2589.700 18.350 ;
        RECT 2589.500 2.400 2589.640 18.030 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 245.040 827.930 245.100 ;
        RECT 960.090 245.040 960.410 245.100 ;
        RECT 827.610 244.900 960.410 245.040 ;
        RECT 827.610 244.840 827.930 244.900 ;
        RECT 960.090 244.840 960.410 244.900 ;
        RECT 823.470 15.540 823.790 15.600 ;
        RECT 827.610 15.540 827.930 15.600 ;
        RECT 823.470 15.400 827.930 15.540 ;
        RECT 823.470 15.340 823.790 15.400 ;
        RECT 827.610 15.340 827.930 15.400 ;
      LAYER via ;
        RECT 827.640 244.840 827.900 245.100 ;
        RECT 960.120 244.840 960.380 245.100 ;
        RECT 823.500 15.340 823.760 15.600 ;
        RECT 827.640 15.340 827.900 15.600 ;
      LAYER met2 ;
        RECT 960.070 260.000 960.350 264.000 ;
        RECT 960.180 245.130 960.320 260.000 ;
        RECT 827.640 244.810 827.900 245.130 ;
        RECT 960.120 244.810 960.380 245.130 ;
        RECT 827.700 15.630 827.840 244.810 ;
        RECT 823.500 15.310 823.760 15.630 ;
        RECT 827.640 15.310 827.900 15.630 ;
        RECT 823.560 2.400 823.700 15.310 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2368.150 244.020 2368.470 244.080 ;
        RECT 2373.210 244.020 2373.530 244.080 ;
        RECT 2368.150 243.880 2373.530 244.020 ;
        RECT 2368.150 243.820 2368.470 243.880 ;
        RECT 2373.210 243.820 2373.530 243.880 ;
        RECT 2373.210 17.240 2373.530 17.300 ;
        RECT 2606.890 17.240 2607.210 17.300 ;
        RECT 2373.210 17.100 2607.210 17.240 ;
        RECT 2373.210 17.040 2373.530 17.100 ;
        RECT 2606.890 17.040 2607.210 17.100 ;
      LAYER via ;
        RECT 2368.180 243.820 2368.440 244.080 ;
        RECT 2373.240 243.820 2373.500 244.080 ;
        RECT 2373.240 17.040 2373.500 17.300 ;
        RECT 2606.920 17.040 2607.180 17.300 ;
      LAYER met2 ;
        RECT 2368.130 260.000 2368.410 264.000 ;
        RECT 2368.240 244.110 2368.380 260.000 ;
        RECT 2368.180 243.790 2368.440 244.110 ;
        RECT 2373.240 243.790 2373.500 244.110 ;
        RECT 2373.300 17.330 2373.440 243.790 ;
        RECT 2373.240 17.010 2373.500 17.330 ;
        RECT 2606.920 17.010 2607.180 17.330 ;
        RECT 2606.980 16.730 2607.120 17.010 ;
        RECT 2606.980 16.590 2607.580 16.730 ;
        RECT 2607.440 2.400 2607.580 16.590 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2382.410 246.400 2382.730 246.460 ;
        RECT 2622.070 246.400 2622.390 246.460 ;
        RECT 2382.410 246.260 2622.390 246.400 ;
        RECT 2382.410 246.200 2382.730 246.260 ;
        RECT 2622.070 246.200 2622.390 246.260 ;
      LAYER via ;
        RECT 2382.440 246.200 2382.700 246.460 ;
        RECT 2622.100 246.200 2622.360 246.460 ;
      LAYER met2 ;
        RECT 2382.390 260.000 2382.670 264.000 ;
        RECT 2382.500 246.490 2382.640 260.000 ;
        RECT 2382.440 246.170 2382.700 246.490 ;
        RECT 2622.100 246.170 2622.360 246.490 ;
        RECT 2622.160 16.730 2622.300 246.170 ;
        RECT 2622.160 16.590 2625.520 16.730 ;
        RECT 2625.380 2.400 2625.520 16.590 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2396.210 244.020 2396.530 244.080 ;
        RECT 2400.810 244.020 2401.130 244.080 ;
        RECT 2396.210 243.880 2401.130 244.020 ;
        RECT 2396.210 243.820 2396.530 243.880 ;
        RECT 2400.810 243.820 2401.130 243.880 ;
        RECT 2400.810 16.220 2401.130 16.280 ;
        RECT 2643.230 16.220 2643.550 16.280 ;
        RECT 2400.810 16.080 2643.550 16.220 ;
        RECT 2400.810 16.020 2401.130 16.080 ;
        RECT 2643.230 16.020 2643.550 16.080 ;
      LAYER via ;
        RECT 2396.240 243.820 2396.500 244.080 ;
        RECT 2400.840 243.820 2401.100 244.080 ;
        RECT 2400.840 16.020 2401.100 16.280 ;
        RECT 2643.260 16.020 2643.520 16.280 ;
      LAYER met2 ;
        RECT 2396.190 260.000 2396.470 264.000 ;
        RECT 2396.300 244.110 2396.440 260.000 ;
        RECT 2396.240 243.790 2396.500 244.110 ;
        RECT 2400.840 243.790 2401.100 244.110 ;
        RECT 2400.900 16.310 2401.040 243.790 ;
        RECT 2400.840 15.990 2401.100 16.310 ;
        RECT 2643.260 15.990 2643.520 16.310 ;
        RECT 2643.320 2.400 2643.460 15.990 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2410.470 246.060 2410.790 246.120 ;
        RECT 2656.570 246.060 2656.890 246.120 ;
        RECT 2410.470 245.920 2656.890 246.060 ;
        RECT 2410.470 245.860 2410.790 245.920 ;
        RECT 2656.570 245.860 2656.890 245.920 ;
      LAYER via ;
        RECT 2410.500 245.860 2410.760 246.120 ;
        RECT 2656.600 245.860 2656.860 246.120 ;
      LAYER met2 ;
        RECT 2410.450 260.000 2410.730 264.000 ;
        RECT 2410.560 246.150 2410.700 260.000 ;
        RECT 2410.500 245.830 2410.760 246.150 ;
        RECT 2656.600 245.830 2656.860 246.150 ;
        RECT 2656.660 17.410 2656.800 245.830 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2424.270 244.020 2424.590 244.080 ;
        RECT 2428.410 244.020 2428.730 244.080 ;
        RECT 2424.270 243.880 2428.730 244.020 ;
        RECT 2424.270 243.820 2424.590 243.880 ;
        RECT 2428.410 243.820 2428.730 243.880 ;
        RECT 2428.410 16.560 2428.730 16.620 ;
        RECT 2678.650 16.560 2678.970 16.620 ;
        RECT 2428.410 16.420 2678.970 16.560 ;
        RECT 2428.410 16.360 2428.730 16.420 ;
        RECT 2678.650 16.360 2678.970 16.420 ;
      LAYER via ;
        RECT 2424.300 243.820 2424.560 244.080 ;
        RECT 2428.440 243.820 2428.700 244.080 ;
        RECT 2428.440 16.360 2428.700 16.620 ;
        RECT 2678.680 16.360 2678.940 16.620 ;
      LAYER met2 ;
        RECT 2424.250 260.000 2424.530 264.000 ;
        RECT 2424.360 244.110 2424.500 260.000 ;
        RECT 2424.300 243.790 2424.560 244.110 ;
        RECT 2428.440 243.790 2428.700 244.110 ;
        RECT 2428.500 16.650 2428.640 243.790 ;
        RECT 2428.440 16.330 2428.700 16.650 ;
        RECT 2678.680 16.330 2678.940 16.650 ;
        RECT 2678.740 2.400 2678.880 16.330 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2438.530 245.720 2438.850 245.780 ;
        RECT 2691.070 245.720 2691.390 245.780 ;
        RECT 2438.530 245.580 2691.390 245.720 ;
        RECT 2438.530 245.520 2438.850 245.580 ;
        RECT 2691.070 245.520 2691.390 245.580 ;
      LAYER via ;
        RECT 2438.560 245.520 2438.820 245.780 ;
        RECT 2691.100 245.520 2691.360 245.780 ;
      LAYER met2 ;
        RECT 2438.510 260.000 2438.790 264.000 ;
        RECT 2438.620 245.810 2438.760 260.000 ;
        RECT 2438.560 245.490 2438.820 245.810 ;
        RECT 2691.100 245.490 2691.360 245.810 ;
        RECT 2691.160 17.410 2691.300 245.490 ;
        RECT 2691.160 17.270 2696.820 17.410 ;
        RECT 2696.680 2.400 2696.820 17.270 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2477.245 16.745 2477.415 19.635 ;
      LAYER mcon ;
        RECT 2477.245 19.465 2477.415 19.635 ;
      LAYER met1 ;
        RECT 2456.010 19.620 2456.330 19.680 ;
        RECT 2477.185 19.620 2477.475 19.665 ;
        RECT 2456.010 19.480 2477.475 19.620 ;
        RECT 2456.010 19.420 2456.330 19.480 ;
        RECT 2477.185 19.435 2477.475 19.480 ;
        RECT 2477.185 16.900 2477.475 16.945 ;
        RECT 2714.530 16.900 2714.850 16.960 ;
        RECT 2477.185 16.760 2714.850 16.900 ;
        RECT 2477.185 16.715 2477.475 16.760 ;
        RECT 2714.530 16.700 2714.850 16.760 ;
      LAYER via ;
        RECT 2456.040 19.420 2456.300 19.680 ;
        RECT 2714.560 16.700 2714.820 16.960 ;
      LAYER met2 ;
        RECT 2452.770 260.170 2453.050 264.000 ;
        RECT 2452.770 260.030 2456.240 260.170 ;
        RECT 2452.770 260.000 2453.050 260.030 ;
        RECT 2456.100 19.710 2456.240 260.030 ;
        RECT 2456.040 19.390 2456.300 19.710 ;
        RECT 2714.560 16.670 2714.820 16.990 ;
        RECT 2714.620 2.400 2714.760 16.670 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2466.590 245.380 2466.910 245.440 ;
        RECT 2732.470 245.380 2732.790 245.440 ;
        RECT 2466.590 245.240 2732.790 245.380 ;
        RECT 2466.590 245.180 2466.910 245.240 ;
        RECT 2732.470 245.180 2732.790 245.240 ;
      LAYER via ;
        RECT 2466.620 245.180 2466.880 245.440 ;
        RECT 2732.500 245.180 2732.760 245.440 ;
      LAYER met2 ;
        RECT 2466.570 260.000 2466.850 264.000 ;
        RECT 2466.680 245.470 2466.820 260.000 ;
        RECT 2466.620 245.150 2466.880 245.470 ;
        RECT 2732.500 245.150 2732.760 245.470 ;
        RECT 2732.560 2.400 2732.700 245.150 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2483.610 20.640 2483.930 20.700 ;
        RECT 2750.410 20.640 2750.730 20.700 ;
        RECT 2483.610 20.500 2750.730 20.640 ;
        RECT 2483.610 20.440 2483.930 20.500 ;
        RECT 2750.410 20.440 2750.730 20.500 ;
      LAYER via ;
        RECT 2483.640 20.440 2483.900 20.700 ;
        RECT 2750.440 20.440 2750.700 20.700 ;
      LAYER met2 ;
        RECT 2480.830 260.170 2481.110 264.000 ;
        RECT 2480.830 260.030 2483.840 260.170 ;
        RECT 2480.830 260.000 2481.110 260.030 ;
        RECT 2483.700 20.730 2483.840 260.030 ;
        RECT 2483.640 20.410 2483.900 20.730 ;
        RECT 2750.440 20.410 2750.700 20.730 ;
        RECT 2750.500 2.400 2750.640 20.410 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2494.650 245.040 2494.970 245.100 ;
        RECT 2766.970 245.040 2767.290 245.100 ;
        RECT 2494.650 244.900 2767.290 245.040 ;
        RECT 2494.650 244.840 2494.970 244.900 ;
        RECT 2766.970 244.840 2767.290 244.900 ;
      LAYER via ;
        RECT 2494.680 244.840 2494.940 245.100 ;
        RECT 2767.000 244.840 2767.260 245.100 ;
      LAYER met2 ;
        RECT 2494.630 260.000 2494.910 264.000 ;
        RECT 2494.740 245.130 2494.880 260.000 ;
        RECT 2494.680 244.810 2494.940 245.130 ;
        RECT 2767.000 244.810 2767.260 245.130 ;
        RECT 2767.060 17.410 2767.200 244.810 ;
        RECT 2767.060 17.270 2768.120 17.410 ;
        RECT 2767.980 2.400 2768.120 17.270 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 17.580 841.270 17.640 ;
        RECT 972.970 17.580 973.290 17.640 ;
        RECT 840.950 17.440 973.290 17.580 ;
        RECT 840.950 17.380 841.270 17.440 ;
        RECT 972.970 17.380 973.290 17.440 ;
      LAYER via ;
        RECT 840.980 17.380 841.240 17.640 ;
        RECT 973.000 17.380 973.260 17.640 ;
      LAYER met2 ;
        RECT 973.870 260.170 974.150 264.000 ;
        RECT 973.060 260.030 974.150 260.170 ;
        RECT 973.060 17.670 973.200 260.030 ;
        RECT 973.870 260.000 974.150 260.030 ;
        RECT 840.980 17.350 841.240 17.670 ;
        RECT 973.000 17.350 973.260 17.670 ;
        RECT 841.040 2.400 841.180 17.350 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2511.210 20.300 2511.530 20.360 ;
        RECT 2785.830 20.300 2786.150 20.360 ;
        RECT 2511.210 20.160 2786.150 20.300 ;
        RECT 2511.210 20.100 2511.530 20.160 ;
        RECT 2785.830 20.100 2786.150 20.160 ;
      LAYER via ;
        RECT 2511.240 20.100 2511.500 20.360 ;
        RECT 2785.860 20.100 2786.120 20.360 ;
      LAYER met2 ;
        RECT 2508.890 260.170 2509.170 264.000 ;
        RECT 2508.890 260.030 2511.440 260.170 ;
        RECT 2508.890 260.000 2509.170 260.030 ;
        RECT 2511.300 20.390 2511.440 260.030 ;
        RECT 2511.240 20.070 2511.500 20.390 ;
        RECT 2785.860 20.070 2786.120 20.390 ;
        RECT 2785.920 2.400 2786.060 20.070 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2525.010 19.960 2525.330 20.020 ;
        RECT 2803.770 19.960 2804.090 20.020 ;
        RECT 2525.010 19.820 2804.090 19.960 ;
        RECT 2525.010 19.760 2525.330 19.820 ;
        RECT 2803.770 19.760 2804.090 19.820 ;
      LAYER via ;
        RECT 2525.040 19.760 2525.300 20.020 ;
        RECT 2803.800 19.760 2804.060 20.020 ;
      LAYER met2 ;
        RECT 2523.150 260.170 2523.430 264.000 ;
        RECT 2523.150 260.030 2525.240 260.170 ;
        RECT 2523.150 260.000 2523.430 260.030 ;
        RECT 2525.100 20.050 2525.240 260.030 ;
        RECT 2525.040 19.730 2525.300 20.050 ;
        RECT 2803.800 19.730 2804.060 20.050 ;
        RECT 2803.860 2.400 2804.000 19.730 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2538.810 19.620 2539.130 19.680 ;
        RECT 2821.710 19.620 2822.030 19.680 ;
        RECT 2538.810 19.480 2822.030 19.620 ;
        RECT 2538.810 19.420 2539.130 19.480 ;
        RECT 2821.710 19.420 2822.030 19.480 ;
      LAYER via ;
        RECT 2538.840 19.420 2539.100 19.680 ;
        RECT 2821.740 19.420 2822.000 19.680 ;
      LAYER met2 ;
        RECT 2536.950 260.170 2537.230 264.000 ;
        RECT 2536.950 260.030 2539.040 260.170 ;
        RECT 2536.950 260.000 2537.230 260.030 ;
        RECT 2538.900 19.710 2539.040 260.030 ;
        RECT 2538.840 19.390 2539.100 19.710 ;
        RECT 2821.740 19.390 2822.000 19.710 ;
        RECT 2821.800 2.400 2821.940 19.390 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2552.610 19.280 2552.930 19.340 ;
        RECT 2839.190 19.280 2839.510 19.340 ;
        RECT 2552.610 19.140 2839.510 19.280 ;
        RECT 2552.610 19.080 2552.930 19.140 ;
        RECT 2839.190 19.080 2839.510 19.140 ;
      LAYER via ;
        RECT 2552.640 19.080 2552.900 19.340 ;
        RECT 2839.220 19.080 2839.480 19.340 ;
      LAYER met2 ;
        RECT 2551.210 260.170 2551.490 264.000 ;
        RECT 2551.210 260.030 2552.840 260.170 ;
        RECT 2551.210 260.000 2551.490 260.030 ;
        RECT 2552.700 19.370 2552.840 260.030 ;
        RECT 2552.640 19.050 2552.900 19.370 ;
        RECT 2839.220 19.050 2839.480 19.370 ;
        RECT 2839.280 2.400 2839.420 19.050 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2565.490 17.920 2565.810 17.980 ;
        RECT 2857.130 17.920 2857.450 17.980 ;
        RECT 2565.490 17.780 2857.450 17.920 ;
        RECT 2565.490 17.720 2565.810 17.780 ;
        RECT 2857.130 17.720 2857.450 17.780 ;
      LAYER via ;
        RECT 2565.520 17.720 2565.780 17.980 ;
        RECT 2857.160 17.720 2857.420 17.980 ;
      LAYER met2 ;
        RECT 2565.010 260.170 2565.290 264.000 ;
        RECT 2565.010 260.030 2566.640 260.170 ;
        RECT 2565.010 260.000 2565.290 260.030 ;
        RECT 2566.500 59.570 2566.640 260.030 ;
        RECT 2565.580 59.430 2566.640 59.570 ;
        RECT 2565.580 18.010 2565.720 59.430 ;
        RECT 2565.520 17.690 2565.780 18.010 ;
        RECT 2857.160 17.690 2857.420 18.010 ;
        RECT 2857.220 2.400 2857.360 17.690 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2875.070 17.920 2875.390 17.980 ;
        RECT 2857.680 17.780 2875.390 17.920 ;
        RECT 2579.750 17.580 2580.070 17.640 ;
        RECT 2857.680 17.580 2857.820 17.780 ;
        RECT 2875.070 17.720 2875.390 17.780 ;
        RECT 2579.750 17.440 2857.820 17.580 ;
        RECT 2579.750 17.380 2580.070 17.440 ;
      LAYER via ;
        RECT 2579.780 17.380 2580.040 17.640 ;
        RECT 2875.100 17.720 2875.360 17.980 ;
      LAYER met2 ;
        RECT 2579.270 260.170 2579.550 264.000 ;
        RECT 2579.270 260.030 2579.980 260.170 ;
        RECT 2579.270 260.000 2579.550 260.030 ;
        RECT 2579.840 17.670 2579.980 260.030 ;
        RECT 2875.100 17.690 2875.360 18.010 ;
        RECT 2579.780 17.350 2580.040 17.670 ;
        RECT 2875.160 2.400 2875.300 17.690 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2593.530 260.000 2593.810 264.000 ;
        RECT 2593.640 16.845 2593.780 260.000 ;
        RECT 2593.570 16.475 2593.850 16.845 ;
        RECT 2893.030 16.475 2893.310 16.845 ;
        RECT 2893.100 2.400 2893.240 16.475 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 2593.570 16.520 2593.850 16.800 ;
        RECT 2893.030 16.520 2893.310 16.800 ;
      LAYER met3 ;
        RECT 2593.545 16.810 2593.875 16.825 ;
        RECT 2893.005 16.810 2893.335 16.825 ;
        RECT 2593.545 16.510 2893.335 16.810 ;
        RECT 2593.545 16.495 2593.875 16.510 ;
        RECT 2893.005 16.495 2893.335 16.510 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.330 260.170 2607.610 264.000 ;
        RECT 2607.330 260.030 2608.040 260.170 ;
        RECT 2607.330 260.000 2607.610 260.030 ;
        RECT 2607.900 18.205 2608.040 260.030 ;
        RECT 2607.830 17.835 2608.110 18.205 ;
        RECT 2910.970 17.835 2911.250 18.205 ;
        RECT 2911.040 2.400 2911.180 17.835 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 2607.830 17.880 2608.110 18.160 ;
        RECT 2910.970 17.880 2911.250 18.160 ;
      LAYER met3 ;
        RECT 2607.805 18.170 2608.135 18.185 ;
        RECT 2910.945 18.170 2911.275 18.185 ;
        RECT 2607.805 17.870 2911.275 18.170 ;
        RECT 2607.805 17.855 2608.135 17.870 ;
        RECT 2910.945 17.855 2911.275 17.870 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 246.060 862.430 246.120 ;
        RECT 988.150 246.060 988.470 246.120 ;
        RECT 862.110 245.920 988.470 246.060 ;
        RECT 862.110 245.860 862.430 245.920 ;
        RECT 988.150 245.860 988.470 245.920 ;
        RECT 858.890 17.920 859.210 17.980 ;
        RECT 862.110 17.920 862.430 17.980 ;
        RECT 858.890 17.780 862.430 17.920 ;
        RECT 858.890 17.720 859.210 17.780 ;
        RECT 862.110 17.720 862.430 17.780 ;
      LAYER via ;
        RECT 862.140 245.860 862.400 246.120 ;
        RECT 988.180 245.860 988.440 246.120 ;
        RECT 858.920 17.720 859.180 17.980 ;
        RECT 862.140 17.720 862.400 17.980 ;
      LAYER met2 ;
        RECT 988.130 260.000 988.410 264.000 ;
        RECT 988.240 246.150 988.380 260.000 ;
        RECT 862.140 245.830 862.400 246.150 ;
        RECT 988.180 245.830 988.440 246.150 ;
        RECT 862.200 18.010 862.340 245.830 ;
        RECT 858.920 17.690 859.180 18.010 ;
        RECT 862.140 17.690 862.400 18.010 ;
        RECT 858.980 2.400 859.120 17.690 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.830 16.900 877.150 16.960 ;
        RECT 1000.570 16.900 1000.890 16.960 ;
        RECT 876.830 16.760 1000.890 16.900 ;
        RECT 876.830 16.700 877.150 16.760 ;
        RECT 1000.570 16.700 1000.890 16.760 ;
      LAYER via ;
        RECT 876.860 16.700 877.120 16.960 ;
        RECT 1000.600 16.700 1000.860 16.960 ;
      LAYER met2 ;
        RECT 1002.390 260.170 1002.670 264.000 ;
        RECT 1000.660 260.030 1002.670 260.170 ;
        RECT 1000.660 16.990 1000.800 260.030 ;
        RECT 1002.390 260.000 1002.670 260.030 ;
        RECT 876.860 16.670 877.120 16.990 ;
        RECT 1000.600 16.670 1000.860 16.990 ;
        RECT 876.920 2.400 877.060 16.670 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 246.400 896.930 246.460 ;
        RECT 1016.210 246.400 1016.530 246.460 ;
        RECT 896.610 246.260 1016.530 246.400 ;
        RECT 896.610 246.200 896.930 246.260 ;
        RECT 1016.210 246.200 1016.530 246.260 ;
      LAYER via ;
        RECT 896.640 246.200 896.900 246.460 ;
        RECT 1016.240 246.200 1016.500 246.460 ;
      LAYER met2 ;
        RECT 1016.190 260.000 1016.470 264.000 ;
        RECT 1016.300 246.490 1016.440 260.000 ;
        RECT 896.640 246.170 896.900 246.490 ;
        RECT 1016.240 246.170 1016.500 246.490 ;
        RECT 896.700 17.410 896.840 246.170 ;
        RECT 894.860 17.270 896.840 17.410 ;
        RECT 894.860 2.400 895.000 17.270 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 18.940 913.030 19.000 ;
        RECT 1028.170 18.940 1028.490 19.000 ;
        RECT 912.710 18.800 1028.490 18.940 ;
        RECT 912.710 18.740 913.030 18.800 ;
        RECT 1028.170 18.740 1028.490 18.800 ;
      LAYER via ;
        RECT 912.740 18.740 913.000 19.000 ;
        RECT 1028.200 18.740 1028.460 19.000 ;
      LAYER met2 ;
        RECT 1030.450 260.170 1030.730 264.000 ;
        RECT 1028.260 260.030 1030.730 260.170 ;
        RECT 1028.260 19.030 1028.400 260.030 ;
        RECT 1030.450 260.000 1030.730 260.030 ;
        RECT 912.740 18.710 913.000 19.030 ;
        RECT 1028.200 18.710 1028.460 19.030 ;
        RECT 912.800 2.400 912.940 18.710 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 246.740 931.430 246.800 ;
        RECT 1044.270 246.740 1044.590 246.800 ;
        RECT 931.110 246.600 1044.590 246.740 ;
        RECT 931.110 246.540 931.430 246.600 ;
        RECT 1044.270 246.540 1044.590 246.600 ;
      LAYER via ;
        RECT 931.140 246.540 931.400 246.800 ;
        RECT 1044.300 246.540 1044.560 246.800 ;
      LAYER met2 ;
        RECT 1044.250 260.000 1044.530 264.000 ;
        RECT 1044.360 246.830 1044.500 260.000 ;
        RECT 931.140 246.510 931.400 246.830 ;
        RECT 1044.300 246.510 1044.560 246.830 ;
        RECT 931.200 3.130 931.340 246.510 ;
        RECT 930.280 2.990 931.340 3.130 ;
        RECT 930.280 2.400 930.420 2.990 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 17.240 948.450 17.300 ;
        RECT 1055.770 17.240 1056.090 17.300 ;
        RECT 948.130 17.100 1056.090 17.240 ;
        RECT 948.130 17.040 948.450 17.100 ;
        RECT 1055.770 17.040 1056.090 17.100 ;
      LAYER via ;
        RECT 948.160 17.040 948.420 17.300 ;
        RECT 1055.800 17.040 1056.060 17.300 ;
      LAYER met2 ;
        RECT 1058.510 260.170 1058.790 264.000 ;
        RECT 1055.860 260.030 1058.790 260.170 ;
        RECT 1055.860 17.330 1056.000 260.030 ;
        RECT 1058.510 260.000 1058.790 260.030 ;
        RECT 948.160 17.010 948.420 17.330 ;
        RECT 1055.800 17.010 1056.060 17.330 ;
        RECT 948.220 2.400 948.360 17.010 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.070 16.220 966.390 16.280 ;
        RECT 1070.030 16.220 1070.350 16.280 ;
        RECT 966.070 16.080 1070.350 16.220 ;
        RECT 966.070 16.020 966.390 16.080 ;
        RECT 1070.030 16.020 1070.350 16.080 ;
      LAYER via ;
        RECT 966.100 16.020 966.360 16.280 ;
        RECT 1070.060 16.020 1070.320 16.280 ;
      LAYER met2 ;
        RECT 1072.770 260.170 1073.050 264.000 ;
        RECT 1070.120 260.030 1073.050 260.170 ;
        RECT 1070.120 16.310 1070.260 260.030 ;
        RECT 1072.770 260.000 1073.050 260.030 ;
        RECT 966.100 15.990 966.360 16.310 ;
        RECT 1070.060 15.990 1070.320 16.310 ;
        RECT 966.160 2.400 966.300 15.990 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 984.010 20.300 984.330 20.360 ;
        RECT 1083.370 20.300 1083.690 20.360 ;
        RECT 984.010 20.160 1083.690 20.300 ;
        RECT 984.010 20.100 984.330 20.160 ;
        RECT 1083.370 20.100 1083.690 20.160 ;
      LAYER via ;
        RECT 984.040 20.100 984.300 20.360 ;
        RECT 1083.400 20.100 1083.660 20.360 ;
      LAYER met2 ;
        RECT 1086.570 260.170 1086.850 264.000 ;
        RECT 1083.460 260.030 1086.850 260.170 ;
        RECT 1083.460 20.390 1083.600 260.030 ;
        RECT 1086.570 260.000 1086.850 260.030 ;
        RECT 984.040 20.070 984.300 20.390 ;
        RECT 1083.400 20.070 1083.660 20.390 ;
        RECT 984.100 2.400 984.240 20.070 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 113.800 669.230 113.860 ;
        RECT 828.070 113.800 828.390 113.860 ;
        RECT 668.910 113.660 828.390 113.800 ;
        RECT 668.910 113.600 669.230 113.660 ;
        RECT 828.070 113.600 828.390 113.660 ;
        RECT 662.930 17.920 663.250 17.980 ;
        RECT 668.910 17.920 669.230 17.980 ;
        RECT 662.930 17.780 669.230 17.920 ;
        RECT 662.930 17.720 663.250 17.780 ;
        RECT 668.910 17.720 669.230 17.780 ;
      LAYER via ;
        RECT 668.940 113.600 669.200 113.860 ;
        RECT 828.100 113.600 828.360 113.860 ;
        RECT 662.960 17.720 663.220 17.980 ;
        RECT 668.940 17.720 669.200 17.980 ;
      LAYER met2 ;
        RECT 833.110 260.170 833.390 264.000 ;
        RECT 829.540 260.030 833.390 260.170 ;
        RECT 829.540 230.250 829.680 260.030 ;
        RECT 833.110 260.000 833.390 260.030 ;
        RECT 828.160 230.110 829.680 230.250 ;
        RECT 828.160 113.890 828.300 230.110 ;
        RECT 668.940 113.570 669.200 113.890 ;
        RECT 828.100 113.570 828.360 113.890 ;
        RECT 669.000 18.010 669.140 113.570 ;
        RECT 662.960 17.690 663.220 18.010 ;
        RECT 668.940 17.690 669.200 18.010 ;
        RECT 663.020 2.400 663.160 17.690 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.950 16.900 1002.270 16.960 ;
        RECT 1097.630 16.900 1097.950 16.960 ;
        RECT 1001.950 16.760 1097.950 16.900 ;
        RECT 1001.950 16.700 1002.270 16.760 ;
        RECT 1097.630 16.700 1097.950 16.760 ;
      LAYER via ;
        RECT 1001.980 16.700 1002.240 16.960 ;
        RECT 1097.660 16.700 1097.920 16.960 ;
      LAYER met2 ;
        RECT 1100.830 260.170 1101.110 264.000 ;
        RECT 1097.720 260.030 1101.110 260.170 ;
        RECT 1097.720 16.990 1097.860 260.030 ;
        RECT 1100.830 260.000 1101.110 260.030 ;
        RECT 1001.980 16.670 1002.240 16.990 ;
        RECT 1097.660 16.670 1097.920 16.990 ;
        RECT 1002.040 2.400 1002.180 16.670 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1019.430 18.600 1019.750 18.660 ;
        RECT 1019.430 18.460 1042.200 18.600 ;
        RECT 1019.430 18.400 1019.750 18.460 ;
        RECT 1042.060 17.920 1042.200 18.460 ;
        RECT 1110.970 17.920 1111.290 17.980 ;
        RECT 1042.060 17.780 1111.290 17.920 ;
        RECT 1110.970 17.720 1111.290 17.780 ;
      LAYER via ;
        RECT 1019.460 18.400 1019.720 18.660 ;
        RECT 1111.000 17.720 1111.260 17.980 ;
      LAYER met2 ;
        RECT 1114.630 260.170 1114.910 264.000 ;
        RECT 1111.060 260.030 1114.910 260.170 ;
        RECT 1019.460 18.370 1019.720 18.690 ;
        RECT 1019.520 2.400 1019.660 18.370 ;
        RECT 1111.060 18.010 1111.200 260.030 ;
        RECT 1114.630 260.000 1114.910 260.030 ;
        RECT 1111.000 17.690 1111.260 18.010 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 246.060 1041.830 246.120 ;
        RECT 1128.910 246.060 1129.230 246.120 ;
        RECT 1041.510 245.920 1129.230 246.060 ;
        RECT 1041.510 245.860 1041.830 245.920 ;
        RECT 1128.910 245.860 1129.230 245.920 ;
        RECT 1037.370 17.920 1037.690 17.980 ;
        RECT 1041.510 17.920 1041.830 17.980 ;
        RECT 1037.370 17.780 1041.830 17.920 ;
        RECT 1037.370 17.720 1037.690 17.780 ;
        RECT 1041.510 17.720 1041.830 17.780 ;
      LAYER via ;
        RECT 1041.540 245.860 1041.800 246.120 ;
        RECT 1128.940 245.860 1129.200 246.120 ;
        RECT 1037.400 17.720 1037.660 17.980 ;
        RECT 1041.540 17.720 1041.800 17.980 ;
      LAYER met2 ;
        RECT 1128.890 260.000 1129.170 264.000 ;
        RECT 1129.000 246.150 1129.140 260.000 ;
        RECT 1041.540 245.830 1041.800 246.150 ;
        RECT 1128.940 245.830 1129.200 246.150 ;
        RECT 1041.600 18.010 1041.740 245.830 ;
        RECT 1037.400 17.690 1037.660 18.010 ;
        RECT 1041.540 17.690 1041.800 18.010 ;
        RECT 1037.460 2.400 1037.600 17.690 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1105.065 18.785 1105.235 19.975 ;
      LAYER mcon ;
        RECT 1105.065 19.805 1105.235 19.975 ;
      LAYER met1 ;
        RECT 1105.005 19.960 1105.295 20.005 ;
        RECT 1138.570 19.960 1138.890 20.020 ;
        RECT 1105.005 19.820 1138.890 19.960 ;
        RECT 1105.005 19.775 1105.295 19.820 ;
        RECT 1138.570 19.760 1138.890 19.820 ;
        RECT 1055.310 18.940 1055.630 19.000 ;
        RECT 1105.005 18.940 1105.295 18.985 ;
        RECT 1055.310 18.800 1105.295 18.940 ;
        RECT 1055.310 18.740 1055.630 18.800 ;
        RECT 1105.005 18.755 1105.295 18.800 ;
      LAYER via ;
        RECT 1138.600 19.760 1138.860 20.020 ;
        RECT 1055.340 18.740 1055.600 19.000 ;
      LAYER met2 ;
        RECT 1143.150 260.170 1143.430 264.000 ;
        RECT 1138.660 260.030 1143.430 260.170 ;
        RECT 1138.660 20.050 1138.800 260.030 ;
        RECT 1143.150 260.000 1143.430 260.030 ;
        RECT 1138.600 19.730 1138.860 20.050 ;
        RECT 1055.340 18.710 1055.600 19.030 ;
        RECT 1055.400 2.400 1055.540 18.710 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 246.400 1076.330 246.460 ;
        RECT 1156.970 246.400 1157.290 246.460 ;
        RECT 1076.010 246.260 1157.290 246.400 ;
        RECT 1076.010 246.200 1076.330 246.260 ;
        RECT 1156.970 246.200 1157.290 246.260 ;
        RECT 1073.250 17.580 1073.570 17.640 ;
        RECT 1076.010 17.580 1076.330 17.640 ;
        RECT 1073.250 17.440 1076.330 17.580 ;
        RECT 1073.250 17.380 1073.570 17.440 ;
        RECT 1076.010 17.380 1076.330 17.440 ;
      LAYER via ;
        RECT 1076.040 246.200 1076.300 246.460 ;
        RECT 1157.000 246.200 1157.260 246.460 ;
        RECT 1073.280 17.380 1073.540 17.640 ;
        RECT 1076.040 17.380 1076.300 17.640 ;
      LAYER met2 ;
        RECT 1156.950 260.000 1157.230 264.000 ;
        RECT 1157.060 246.490 1157.200 260.000 ;
        RECT 1076.040 246.170 1076.300 246.490 ;
        RECT 1157.000 246.170 1157.260 246.490 ;
        RECT 1076.100 17.670 1076.240 246.170 ;
        RECT 1073.280 17.350 1073.540 17.670 ;
        RECT 1076.040 17.350 1076.300 17.670 ;
        RECT 1073.340 2.400 1073.480 17.350 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 247.420 1097.030 247.480 ;
        RECT 1171.230 247.420 1171.550 247.480 ;
        RECT 1096.710 247.280 1171.550 247.420 ;
        RECT 1096.710 247.220 1097.030 247.280 ;
        RECT 1171.230 247.220 1171.550 247.280 ;
        RECT 1091.190 20.300 1091.510 20.360 ;
        RECT 1096.710 20.300 1097.030 20.360 ;
        RECT 1091.190 20.160 1097.030 20.300 ;
        RECT 1091.190 20.100 1091.510 20.160 ;
        RECT 1096.710 20.100 1097.030 20.160 ;
      LAYER via ;
        RECT 1096.740 247.220 1097.000 247.480 ;
        RECT 1171.260 247.220 1171.520 247.480 ;
        RECT 1091.220 20.100 1091.480 20.360 ;
        RECT 1096.740 20.100 1097.000 20.360 ;
      LAYER met2 ;
        RECT 1171.210 260.000 1171.490 264.000 ;
        RECT 1171.320 247.510 1171.460 260.000 ;
        RECT 1096.740 247.190 1097.000 247.510 ;
        RECT 1171.260 247.190 1171.520 247.510 ;
        RECT 1096.800 20.390 1096.940 247.190 ;
        RECT 1091.220 20.070 1091.480 20.390 ;
        RECT 1096.740 20.070 1097.000 20.390 ;
        RECT 1091.280 17.410 1091.420 20.070 ;
        RECT 1090.820 17.270 1091.420 17.410 ;
        RECT 1090.820 2.400 1090.960 17.270 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.510 245.040 1110.830 245.100 ;
        RECT 1185.030 245.040 1185.350 245.100 ;
        RECT 1110.510 244.900 1185.350 245.040 ;
        RECT 1110.510 244.840 1110.830 244.900 ;
        RECT 1185.030 244.840 1185.350 244.900 ;
      LAYER via ;
        RECT 1110.540 244.840 1110.800 245.100 ;
        RECT 1185.060 244.840 1185.320 245.100 ;
      LAYER met2 ;
        RECT 1185.010 260.000 1185.290 264.000 ;
        RECT 1185.120 245.130 1185.260 260.000 ;
        RECT 1110.540 244.810 1110.800 245.130 ;
        RECT 1185.060 244.810 1185.320 245.130 ;
        RECT 1110.600 3.130 1110.740 244.810 ;
        RECT 1108.760 2.990 1110.740 3.130 ;
        RECT 1108.760 2.400 1108.900 2.990 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 245.720 1131.530 245.780 ;
        RECT 1199.290 245.720 1199.610 245.780 ;
        RECT 1131.210 245.580 1199.610 245.720 ;
        RECT 1131.210 245.520 1131.530 245.580 ;
        RECT 1199.290 245.520 1199.610 245.580 ;
        RECT 1126.610 17.920 1126.930 17.980 ;
        RECT 1131.210 17.920 1131.530 17.980 ;
        RECT 1126.610 17.780 1131.530 17.920 ;
        RECT 1126.610 17.720 1126.930 17.780 ;
        RECT 1131.210 17.720 1131.530 17.780 ;
      LAYER via ;
        RECT 1131.240 245.520 1131.500 245.780 ;
        RECT 1199.320 245.520 1199.580 245.780 ;
        RECT 1126.640 17.720 1126.900 17.980 ;
        RECT 1131.240 17.720 1131.500 17.980 ;
      LAYER met2 ;
        RECT 1199.270 260.000 1199.550 264.000 ;
        RECT 1199.380 245.810 1199.520 260.000 ;
        RECT 1131.240 245.490 1131.500 245.810 ;
        RECT 1199.320 245.490 1199.580 245.810 ;
        RECT 1131.300 18.010 1131.440 245.490 ;
        RECT 1126.640 17.690 1126.900 18.010 ;
        RECT 1131.240 17.690 1131.500 18.010 ;
        RECT 1126.700 2.400 1126.840 17.690 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 248.440 1162.810 248.500 ;
        RECT 1213.550 248.440 1213.870 248.500 ;
        RECT 1162.490 248.300 1213.870 248.440 ;
        RECT 1162.490 248.240 1162.810 248.300 ;
        RECT 1213.550 248.240 1213.870 248.300 ;
        RECT 1144.550 18.940 1144.870 19.000 ;
        RECT 1162.490 18.940 1162.810 19.000 ;
        RECT 1144.550 18.800 1162.810 18.940 ;
        RECT 1144.550 18.740 1144.870 18.800 ;
        RECT 1162.490 18.740 1162.810 18.800 ;
      LAYER via ;
        RECT 1162.520 248.240 1162.780 248.500 ;
        RECT 1213.580 248.240 1213.840 248.500 ;
        RECT 1144.580 18.740 1144.840 19.000 ;
        RECT 1162.520 18.740 1162.780 19.000 ;
      LAYER met2 ;
        RECT 1213.530 260.000 1213.810 264.000 ;
        RECT 1213.640 248.530 1213.780 260.000 ;
        RECT 1162.520 248.210 1162.780 248.530 ;
        RECT 1213.580 248.210 1213.840 248.530 ;
        RECT 1162.580 19.030 1162.720 248.210 ;
        RECT 1144.580 18.710 1144.840 19.030 ;
        RECT 1162.520 18.710 1162.780 19.030 ;
        RECT 1144.640 2.400 1144.780 18.710 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 246.400 1166.030 246.460 ;
        RECT 1227.350 246.400 1227.670 246.460 ;
        RECT 1165.710 246.260 1227.670 246.400 ;
        RECT 1165.710 246.200 1166.030 246.260 ;
        RECT 1227.350 246.200 1227.670 246.260 ;
        RECT 1162.490 17.580 1162.810 17.640 ;
        RECT 1165.710 17.580 1166.030 17.640 ;
        RECT 1162.490 17.440 1166.030 17.580 ;
        RECT 1162.490 17.380 1162.810 17.440 ;
        RECT 1165.710 17.380 1166.030 17.440 ;
      LAYER via ;
        RECT 1165.740 246.200 1166.000 246.460 ;
        RECT 1227.380 246.200 1227.640 246.460 ;
        RECT 1162.520 17.380 1162.780 17.640 ;
        RECT 1165.740 17.380 1166.000 17.640 ;
      LAYER met2 ;
        RECT 1227.330 260.000 1227.610 264.000 ;
        RECT 1227.440 246.490 1227.580 260.000 ;
        RECT 1165.740 246.170 1166.000 246.490 ;
        RECT 1227.380 246.170 1227.640 246.490 ;
        RECT 1165.800 17.670 1165.940 246.170 ;
        RECT 1162.520 17.350 1162.780 17.670 ;
        RECT 1165.740 17.350 1166.000 17.670 ;
        RECT 1162.580 2.400 1162.720 17.350 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 843.785 193.205 843.955 241.315 ;
      LAYER mcon ;
        RECT 843.785 241.145 843.955 241.315 ;
      LAYER met1 ;
        RECT 843.710 241.300 844.030 241.360 ;
        RECT 843.515 241.160 844.030 241.300 ;
        RECT 843.710 241.100 844.030 241.160 ;
        RECT 843.725 193.360 844.015 193.405 ;
        RECT 844.170 193.360 844.490 193.420 ;
        RECT 843.725 193.220 844.490 193.360 ;
        RECT 843.725 193.175 844.015 193.220 ;
        RECT 844.170 193.160 844.490 193.220 ;
        RECT 682.710 120.600 683.030 120.660 ;
        RECT 844.170 120.600 844.490 120.660 ;
        RECT 682.710 120.460 844.490 120.600 ;
        RECT 682.710 120.400 683.030 120.460 ;
        RECT 844.170 120.400 844.490 120.460 ;
        RECT 680.410 17.920 680.730 17.980 ;
        RECT 682.710 17.920 683.030 17.980 ;
        RECT 680.410 17.780 683.030 17.920 ;
        RECT 680.410 17.720 680.730 17.780 ;
        RECT 682.710 17.720 683.030 17.780 ;
      LAYER via ;
        RECT 843.740 241.100 844.000 241.360 ;
        RECT 844.200 193.160 844.460 193.420 ;
        RECT 682.740 120.400 683.000 120.660 ;
        RECT 844.200 120.400 844.460 120.660 ;
        RECT 680.440 17.720 680.700 17.980 ;
        RECT 682.740 17.720 683.000 17.980 ;
      LAYER met2 ;
        RECT 847.370 260.850 847.650 264.000 ;
        RECT 843.800 260.710 847.650 260.850 ;
        RECT 843.800 241.390 843.940 260.710 ;
        RECT 847.370 260.000 847.650 260.710 ;
        RECT 843.740 241.070 844.000 241.390 ;
        RECT 844.200 193.130 844.460 193.450 ;
        RECT 844.260 120.690 844.400 193.130 ;
        RECT 682.740 120.370 683.000 120.690 ;
        RECT 844.200 120.370 844.460 120.690 ;
        RECT 682.800 18.010 682.940 120.370 ;
        RECT 680.440 17.690 680.700 18.010 ;
        RECT 682.740 17.690 683.000 18.010 ;
        RECT 680.500 2.400 680.640 17.690 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 247.760 1186.270 247.820 ;
        RECT 1240.230 247.760 1240.550 247.820 ;
        RECT 1185.950 247.620 1240.550 247.760 ;
        RECT 1185.950 247.560 1186.270 247.620 ;
        RECT 1240.230 247.560 1240.550 247.620 ;
        RECT 1179.970 17.920 1180.290 17.980 ;
        RECT 1185.950 17.920 1186.270 17.980 ;
        RECT 1179.970 17.780 1186.270 17.920 ;
        RECT 1179.970 17.720 1180.290 17.780 ;
        RECT 1185.950 17.720 1186.270 17.780 ;
      LAYER via ;
        RECT 1185.980 247.560 1186.240 247.820 ;
        RECT 1240.260 247.560 1240.520 247.820 ;
        RECT 1180.000 17.720 1180.260 17.980 ;
        RECT 1185.980 17.720 1186.240 17.980 ;
      LAYER met2 ;
        RECT 1241.590 260.170 1241.870 264.000 ;
        RECT 1240.320 260.030 1241.870 260.170 ;
        RECT 1240.320 247.850 1240.460 260.030 ;
        RECT 1241.590 260.000 1241.870 260.030 ;
        RECT 1185.980 247.530 1186.240 247.850 ;
        RECT 1240.260 247.530 1240.520 247.850 ;
        RECT 1186.040 18.010 1186.180 247.530 ;
        RECT 1180.000 17.690 1180.260 18.010 ;
        RECT 1185.980 17.690 1186.240 18.010 ;
        RECT 1180.060 2.400 1180.200 17.690 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 245.040 1200.530 245.100 ;
        RECT 1255.870 245.040 1256.190 245.100 ;
        RECT 1200.210 244.900 1256.190 245.040 ;
        RECT 1200.210 244.840 1200.530 244.900 ;
        RECT 1255.870 244.840 1256.190 244.900 ;
        RECT 1197.910 17.580 1198.230 17.640 ;
        RECT 1200.210 17.580 1200.530 17.640 ;
        RECT 1197.910 17.440 1200.530 17.580 ;
        RECT 1197.910 17.380 1198.230 17.440 ;
        RECT 1200.210 17.380 1200.530 17.440 ;
      LAYER via ;
        RECT 1200.240 244.840 1200.500 245.100 ;
        RECT 1255.900 244.840 1256.160 245.100 ;
        RECT 1197.940 17.380 1198.200 17.640 ;
        RECT 1200.240 17.380 1200.500 17.640 ;
      LAYER met2 ;
        RECT 1255.850 260.000 1256.130 264.000 ;
        RECT 1255.960 245.130 1256.100 260.000 ;
        RECT 1200.240 244.810 1200.500 245.130 ;
        RECT 1255.900 244.810 1256.160 245.130 ;
        RECT 1200.300 17.670 1200.440 244.810 ;
        RECT 1197.940 17.350 1198.200 17.670 ;
        RECT 1200.240 17.350 1200.500 17.670 ;
        RECT 1198.000 2.400 1198.140 17.350 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 245.720 1221.230 245.780 ;
        RECT 1269.670 245.720 1269.990 245.780 ;
        RECT 1220.910 245.580 1269.990 245.720 ;
        RECT 1220.910 245.520 1221.230 245.580 ;
        RECT 1269.670 245.520 1269.990 245.580 ;
        RECT 1215.850 17.580 1216.170 17.640 ;
        RECT 1220.910 17.580 1221.230 17.640 ;
        RECT 1215.850 17.440 1221.230 17.580 ;
        RECT 1215.850 17.380 1216.170 17.440 ;
        RECT 1220.910 17.380 1221.230 17.440 ;
      LAYER via ;
        RECT 1220.940 245.520 1221.200 245.780 ;
        RECT 1269.700 245.520 1269.960 245.780 ;
        RECT 1215.880 17.380 1216.140 17.640 ;
        RECT 1220.940 17.380 1221.200 17.640 ;
      LAYER met2 ;
        RECT 1269.650 260.000 1269.930 264.000 ;
        RECT 1269.760 245.810 1269.900 260.000 ;
        RECT 1220.940 245.490 1221.200 245.810 ;
        RECT 1269.700 245.490 1269.960 245.810 ;
        RECT 1221.000 17.670 1221.140 245.490 ;
        RECT 1215.880 17.350 1216.140 17.670 ;
        RECT 1220.940 17.350 1221.200 17.670 ;
        RECT 1215.940 2.400 1216.080 17.350 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.710 246.400 1235.030 246.460 ;
        RECT 1283.930 246.400 1284.250 246.460 ;
        RECT 1234.710 246.260 1284.250 246.400 ;
        RECT 1234.710 246.200 1235.030 246.260 ;
        RECT 1283.930 246.200 1284.250 246.260 ;
      LAYER via ;
        RECT 1234.740 246.200 1235.000 246.460 ;
        RECT 1283.960 246.200 1284.220 246.460 ;
      LAYER met2 ;
        RECT 1283.910 260.000 1284.190 264.000 ;
        RECT 1284.020 246.490 1284.160 260.000 ;
        RECT 1234.740 246.170 1235.000 246.490 ;
        RECT 1283.960 246.170 1284.220 246.490 ;
        RECT 1234.800 16.730 1234.940 246.170 ;
        RECT 1233.880 16.590 1234.940 16.730 ;
        RECT 1233.880 2.400 1234.020 16.590 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 246.740 1255.730 246.800 ;
        RECT 1297.730 246.740 1298.050 246.800 ;
        RECT 1255.410 246.600 1298.050 246.740 ;
        RECT 1255.410 246.540 1255.730 246.600 ;
        RECT 1297.730 246.540 1298.050 246.600 ;
        RECT 1251.730 17.580 1252.050 17.640 ;
        RECT 1255.410 17.580 1255.730 17.640 ;
        RECT 1251.730 17.440 1255.730 17.580 ;
        RECT 1251.730 17.380 1252.050 17.440 ;
        RECT 1255.410 17.380 1255.730 17.440 ;
      LAYER via ;
        RECT 1255.440 246.540 1255.700 246.800 ;
        RECT 1297.760 246.540 1298.020 246.800 ;
        RECT 1251.760 17.380 1252.020 17.640 ;
        RECT 1255.440 17.380 1255.700 17.640 ;
      LAYER met2 ;
        RECT 1297.710 260.000 1297.990 264.000 ;
        RECT 1297.820 246.830 1297.960 260.000 ;
        RECT 1255.440 246.510 1255.700 246.830 ;
        RECT 1297.760 246.510 1298.020 246.830 ;
        RECT 1255.500 17.670 1255.640 246.510 ;
        RECT 1251.760 17.350 1252.020 17.670 ;
        RECT 1255.440 17.350 1255.700 17.670 ;
        RECT 1251.820 2.400 1251.960 17.350 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1286.690 248.100 1287.010 248.160 ;
        RECT 1311.990 248.100 1312.310 248.160 ;
        RECT 1286.690 247.960 1312.310 248.100 ;
        RECT 1286.690 247.900 1287.010 247.960 ;
        RECT 1311.990 247.900 1312.310 247.960 ;
        RECT 1269.210 16.560 1269.530 16.620 ;
        RECT 1286.690 16.560 1287.010 16.620 ;
        RECT 1269.210 16.420 1287.010 16.560 ;
        RECT 1269.210 16.360 1269.530 16.420 ;
        RECT 1286.690 16.360 1287.010 16.420 ;
      LAYER via ;
        RECT 1286.720 247.900 1286.980 248.160 ;
        RECT 1312.020 247.900 1312.280 248.160 ;
        RECT 1269.240 16.360 1269.500 16.620 ;
        RECT 1286.720 16.360 1286.980 16.620 ;
      LAYER met2 ;
        RECT 1311.970 260.000 1312.250 264.000 ;
        RECT 1312.080 248.190 1312.220 260.000 ;
        RECT 1286.720 247.870 1286.980 248.190 ;
        RECT 1312.020 247.870 1312.280 248.190 ;
        RECT 1286.780 16.650 1286.920 247.870 ;
        RECT 1269.240 16.330 1269.500 16.650 ;
        RECT 1286.720 16.330 1286.980 16.650 ;
        RECT 1269.300 2.400 1269.440 16.330 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 245.720 1290.230 245.780 ;
        RECT 1326.250 245.720 1326.570 245.780 ;
        RECT 1289.910 245.580 1326.570 245.720 ;
        RECT 1289.910 245.520 1290.230 245.580 ;
        RECT 1326.250 245.520 1326.570 245.580 ;
        RECT 1287.150 17.580 1287.470 17.640 ;
        RECT 1289.910 17.580 1290.230 17.640 ;
        RECT 1287.150 17.440 1290.230 17.580 ;
        RECT 1287.150 17.380 1287.470 17.440 ;
        RECT 1289.910 17.380 1290.230 17.440 ;
      LAYER via ;
        RECT 1289.940 245.520 1290.200 245.780 ;
        RECT 1326.280 245.520 1326.540 245.780 ;
        RECT 1287.180 17.380 1287.440 17.640 ;
        RECT 1289.940 17.380 1290.200 17.640 ;
      LAYER met2 ;
        RECT 1326.230 260.000 1326.510 264.000 ;
        RECT 1326.340 245.810 1326.480 260.000 ;
        RECT 1289.940 245.490 1290.200 245.810 ;
        RECT 1326.280 245.490 1326.540 245.810 ;
        RECT 1290.000 17.670 1290.140 245.490 ;
        RECT 1287.180 17.350 1287.440 17.670 ;
        RECT 1289.940 17.350 1290.200 17.670 ;
        RECT 1287.240 2.400 1287.380 17.350 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 248.440 1310.930 248.500 ;
        RECT 1340.050 248.440 1340.370 248.500 ;
        RECT 1310.610 248.300 1340.370 248.440 ;
        RECT 1310.610 248.240 1310.930 248.300 ;
        RECT 1340.050 248.240 1340.370 248.300 ;
        RECT 1305.090 16.220 1305.410 16.280 ;
        RECT 1310.610 16.220 1310.930 16.280 ;
        RECT 1305.090 16.080 1310.930 16.220 ;
        RECT 1305.090 16.020 1305.410 16.080 ;
        RECT 1310.610 16.020 1310.930 16.080 ;
      LAYER via ;
        RECT 1310.640 248.240 1310.900 248.500 ;
        RECT 1340.080 248.240 1340.340 248.500 ;
        RECT 1305.120 16.020 1305.380 16.280 ;
        RECT 1310.640 16.020 1310.900 16.280 ;
      LAYER met2 ;
        RECT 1340.030 260.000 1340.310 264.000 ;
        RECT 1340.140 248.530 1340.280 260.000 ;
        RECT 1310.640 248.210 1310.900 248.530 ;
        RECT 1340.080 248.210 1340.340 248.530 ;
        RECT 1310.700 16.310 1310.840 248.210 ;
        RECT 1305.120 15.990 1305.380 16.310 ;
        RECT 1310.640 15.990 1310.900 16.310 ;
        RECT 1305.180 2.400 1305.320 15.990 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 245.380 1324.730 245.440 ;
        RECT 1354.310 245.380 1354.630 245.440 ;
        RECT 1324.410 245.240 1354.630 245.380 ;
        RECT 1324.410 245.180 1324.730 245.240 ;
        RECT 1354.310 245.180 1354.630 245.240 ;
      LAYER via ;
        RECT 1324.440 245.180 1324.700 245.440 ;
        RECT 1354.340 245.180 1354.600 245.440 ;
      LAYER met2 ;
        RECT 1354.290 260.000 1354.570 264.000 ;
        RECT 1354.400 245.470 1354.540 260.000 ;
        RECT 1324.440 245.150 1324.700 245.470 ;
        RECT 1354.340 245.150 1354.600 245.470 ;
        RECT 1324.500 17.410 1324.640 245.150 ;
        RECT 1323.120 17.270 1324.640 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 243.680 1345.430 243.740 ;
        RECT 1368.110 243.680 1368.430 243.740 ;
        RECT 1345.110 243.540 1368.430 243.680 ;
        RECT 1345.110 243.480 1345.430 243.540 ;
        RECT 1368.110 243.480 1368.430 243.540 ;
        RECT 1340.510 17.580 1340.830 17.640 ;
        RECT 1345.110 17.580 1345.430 17.640 ;
        RECT 1340.510 17.440 1345.430 17.580 ;
        RECT 1340.510 17.380 1340.830 17.440 ;
        RECT 1345.110 17.380 1345.430 17.440 ;
      LAYER via ;
        RECT 1345.140 243.480 1345.400 243.740 ;
        RECT 1368.140 243.480 1368.400 243.740 ;
        RECT 1340.540 17.380 1340.800 17.640 ;
        RECT 1345.140 17.380 1345.400 17.640 ;
      LAYER met2 ;
        RECT 1368.090 260.000 1368.370 264.000 ;
        RECT 1368.200 243.770 1368.340 260.000 ;
        RECT 1345.140 243.450 1345.400 243.770 ;
        RECT 1368.140 243.450 1368.400 243.770 ;
        RECT 1345.200 17.670 1345.340 243.450 ;
        RECT 1340.540 17.350 1340.800 17.670 ;
        RECT 1345.140 17.350 1345.400 17.670 ;
        RECT 1340.600 2.400 1340.740 17.350 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 127.740 703.730 127.800 ;
        RECT 855.670 127.740 855.990 127.800 ;
        RECT 703.410 127.600 855.990 127.740 ;
        RECT 703.410 127.540 703.730 127.600 ;
        RECT 855.670 127.540 855.990 127.600 ;
        RECT 698.350 17.920 698.670 17.980 ;
        RECT 703.410 17.920 703.730 17.980 ;
        RECT 698.350 17.780 703.730 17.920 ;
        RECT 698.350 17.720 698.670 17.780 ;
        RECT 703.410 17.720 703.730 17.780 ;
      LAYER via ;
        RECT 703.440 127.540 703.700 127.800 ;
        RECT 855.700 127.540 855.960 127.800 ;
        RECT 698.380 17.720 698.640 17.980 ;
        RECT 703.440 17.720 703.700 17.980 ;
      LAYER met2 ;
        RECT 861.170 260.170 861.450 264.000 ;
        RECT 859.440 260.030 861.450 260.170 ;
        RECT 859.440 222.770 859.580 260.030 ;
        RECT 861.170 260.000 861.450 260.030 ;
        RECT 855.760 222.630 859.580 222.770 ;
        RECT 855.760 127.830 855.900 222.630 ;
        RECT 703.440 127.510 703.700 127.830 ;
        RECT 855.700 127.510 855.960 127.830 ;
        RECT 703.500 18.010 703.640 127.510 ;
        RECT 698.380 17.690 698.640 18.010 ;
        RECT 703.440 17.690 703.700 18.010 ;
        RECT 698.440 2.400 698.580 17.690 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.910 244.360 1359.230 244.420 ;
        RECT 1382.370 244.360 1382.690 244.420 ;
        RECT 1358.910 244.220 1382.690 244.360 ;
        RECT 1358.910 244.160 1359.230 244.220 ;
        RECT 1382.370 244.160 1382.690 244.220 ;
      LAYER via ;
        RECT 1358.940 244.160 1359.200 244.420 ;
        RECT 1382.400 244.160 1382.660 244.420 ;
      LAYER met2 ;
        RECT 1382.350 260.000 1382.630 264.000 ;
        RECT 1382.460 244.450 1382.600 260.000 ;
        RECT 1358.940 244.130 1359.200 244.450 ;
        RECT 1382.400 244.130 1382.660 244.450 ;
        RECT 1359.000 17.410 1359.140 244.130 ;
        RECT 1358.540 17.270 1359.140 17.410 ;
        RECT 1358.540 2.400 1358.680 17.270 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.610 248.440 1379.930 248.500 ;
        RECT 1396.630 248.440 1396.950 248.500 ;
        RECT 1379.610 248.300 1396.950 248.440 ;
        RECT 1379.610 248.240 1379.930 248.300 ;
        RECT 1396.630 248.240 1396.950 248.300 ;
        RECT 1376.390 17.580 1376.710 17.640 ;
        RECT 1379.610 17.580 1379.930 17.640 ;
        RECT 1376.390 17.440 1379.930 17.580 ;
        RECT 1376.390 17.380 1376.710 17.440 ;
        RECT 1379.610 17.380 1379.930 17.440 ;
      LAYER via ;
        RECT 1379.640 248.240 1379.900 248.500 ;
        RECT 1396.660 248.240 1396.920 248.500 ;
        RECT 1376.420 17.380 1376.680 17.640 ;
        RECT 1379.640 17.380 1379.900 17.640 ;
      LAYER met2 ;
        RECT 1396.610 260.000 1396.890 264.000 ;
        RECT 1396.720 248.530 1396.860 260.000 ;
        RECT 1379.640 248.210 1379.900 248.530 ;
        RECT 1396.660 248.210 1396.920 248.530 ;
        RECT 1379.700 17.670 1379.840 248.210 ;
        RECT 1376.420 17.350 1376.680 17.670 ;
        RECT 1379.640 17.350 1379.900 17.670 ;
        RECT 1376.480 2.400 1376.620 17.350 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 243.680 1400.630 243.740 ;
        RECT 1410.430 243.680 1410.750 243.740 ;
        RECT 1400.310 243.540 1410.750 243.680 ;
        RECT 1400.310 243.480 1400.630 243.540 ;
        RECT 1410.430 243.480 1410.750 243.540 ;
        RECT 1399.390 24.720 1399.710 24.780 ;
        RECT 1400.310 24.720 1400.630 24.780 ;
        RECT 1399.390 24.580 1400.630 24.720 ;
        RECT 1399.390 24.520 1399.710 24.580 ;
        RECT 1400.310 24.520 1400.630 24.580 ;
        RECT 1394.330 20.640 1394.650 20.700 ;
        RECT 1399.390 20.640 1399.710 20.700 ;
        RECT 1394.330 20.500 1399.710 20.640 ;
        RECT 1394.330 20.440 1394.650 20.500 ;
        RECT 1399.390 20.440 1399.710 20.500 ;
      LAYER via ;
        RECT 1400.340 243.480 1400.600 243.740 ;
        RECT 1410.460 243.480 1410.720 243.740 ;
        RECT 1399.420 24.520 1399.680 24.780 ;
        RECT 1400.340 24.520 1400.600 24.780 ;
        RECT 1394.360 20.440 1394.620 20.700 ;
        RECT 1399.420 20.440 1399.680 20.700 ;
      LAYER met2 ;
        RECT 1410.410 260.000 1410.690 264.000 ;
        RECT 1410.520 243.770 1410.660 260.000 ;
        RECT 1400.340 243.450 1400.600 243.770 ;
        RECT 1410.460 243.450 1410.720 243.770 ;
        RECT 1400.400 24.810 1400.540 243.450 ;
        RECT 1399.420 24.490 1399.680 24.810 ;
        RECT 1400.340 24.490 1400.600 24.810 ;
        RECT 1399.480 20.730 1399.620 24.490 ;
        RECT 1394.360 20.410 1394.620 20.730 ;
        RECT 1399.420 20.410 1399.680 20.730 ;
        RECT 1394.420 2.400 1394.560 20.410 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1412.270 15.880 1412.590 15.940 ;
        RECT 1421.470 15.880 1421.790 15.940 ;
        RECT 1412.270 15.740 1421.790 15.880 ;
        RECT 1412.270 15.680 1412.590 15.740 ;
        RECT 1421.470 15.680 1421.790 15.740 ;
      LAYER via ;
        RECT 1412.300 15.680 1412.560 15.940 ;
        RECT 1421.500 15.680 1421.760 15.940 ;
      LAYER met2 ;
        RECT 1424.670 260.170 1424.950 264.000 ;
        RECT 1421.560 260.030 1424.950 260.170 ;
        RECT 1421.560 15.970 1421.700 260.030 ;
        RECT 1424.670 260.000 1424.950 260.030 ;
        RECT 1412.300 15.650 1412.560 15.970 ;
        RECT 1421.500 15.650 1421.760 15.970 ;
        RECT 1412.360 2.400 1412.500 15.650 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 241.640 1435.130 241.700 ;
        RECT 1438.490 241.640 1438.810 241.700 ;
        RECT 1434.810 241.500 1438.810 241.640 ;
        RECT 1434.810 241.440 1435.130 241.500 ;
        RECT 1438.490 241.440 1438.810 241.500 ;
        RECT 1429.750 18.260 1430.070 18.320 ;
        RECT 1434.810 18.260 1435.130 18.320 ;
        RECT 1429.750 18.120 1435.130 18.260 ;
        RECT 1429.750 18.060 1430.070 18.120 ;
        RECT 1434.810 18.060 1435.130 18.120 ;
      LAYER via ;
        RECT 1434.840 241.440 1435.100 241.700 ;
        RECT 1438.520 241.440 1438.780 241.700 ;
        RECT 1429.780 18.060 1430.040 18.320 ;
        RECT 1434.840 18.060 1435.100 18.320 ;
      LAYER met2 ;
        RECT 1438.470 260.000 1438.750 264.000 ;
        RECT 1438.580 241.730 1438.720 260.000 ;
        RECT 1434.840 241.410 1435.100 241.730 ;
        RECT 1438.520 241.410 1438.780 241.730 ;
        RECT 1434.900 18.350 1435.040 241.410 ;
        RECT 1429.780 18.030 1430.040 18.350 ;
        RECT 1434.840 18.030 1435.100 18.350 ;
        RECT 1429.840 2.400 1429.980 18.030 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1447.690 20.640 1448.010 20.700 ;
        RECT 1449.530 20.640 1449.850 20.700 ;
        RECT 1447.690 20.500 1449.850 20.640 ;
        RECT 1447.690 20.440 1448.010 20.500 ;
        RECT 1449.530 20.440 1449.850 20.500 ;
      LAYER via ;
        RECT 1447.720 20.440 1447.980 20.700 ;
        RECT 1449.560 20.440 1449.820 20.700 ;
      LAYER met2 ;
        RECT 1452.730 260.170 1453.010 264.000 ;
        RECT 1449.620 260.030 1453.010 260.170 ;
        RECT 1449.620 20.730 1449.760 260.030 ;
        RECT 1452.730 260.000 1453.010 260.030 ;
        RECT 1447.720 20.410 1447.980 20.730 ;
        RECT 1449.560 20.410 1449.820 20.730 ;
        RECT 1447.780 2.400 1447.920 20.410 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.870 20.640 1463.190 20.700 ;
        RECT 1465.630 20.640 1465.950 20.700 ;
        RECT 1462.870 20.500 1465.950 20.640 ;
        RECT 1462.870 20.440 1463.190 20.500 ;
        RECT 1465.630 20.440 1465.950 20.500 ;
      LAYER via ;
        RECT 1462.900 20.440 1463.160 20.700 ;
        RECT 1465.660 20.440 1465.920 20.700 ;
      LAYER met2 ;
        RECT 1466.990 260.170 1467.270 264.000 ;
        RECT 1462.960 260.030 1467.270 260.170 ;
        RECT 1462.960 20.730 1463.100 260.030 ;
        RECT 1466.990 260.000 1467.270 260.030 ;
        RECT 1462.900 20.410 1463.160 20.730 ;
        RECT 1465.660 20.410 1465.920 20.730 ;
        RECT 1465.720 2.400 1465.860 20.410 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.110 244.020 1483.430 244.080 ;
        RECT 1484.490 244.020 1484.810 244.080 ;
        RECT 1483.110 243.880 1484.810 244.020 ;
        RECT 1483.110 243.820 1483.430 243.880 ;
        RECT 1484.490 243.820 1484.810 243.880 ;
        RECT 1484.490 206.960 1484.810 207.020 ;
        RECT 1485.410 206.960 1485.730 207.020 ;
        RECT 1484.490 206.820 1485.730 206.960 ;
        RECT 1484.490 206.760 1484.810 206.820 ;
        RECT 1485.410 206.760 1485.730 206.820 ;
        RECT 1484.950 145.080 1485.270 145.140 ;
        RECT 1485.410 145.080 1485.730 145.140 ;
        RECT 1484.950 144.940 1485.730 145.080 ;
        RECT 1484.950 144.880 1485.270 144.940 ;
        RECT 1485.410 144.880 1485.730 144.940 ;
        RECT 1484.950 137.940 1485.270 138.000 ;
        RECT 1485.410 137.940 1485.730 138.000 ;
        RECT 1484.950 137.800 1485.730 137.940 ;
        RECT 1484.950 137.740 1485.270 137.800 ;
        RECT 1485.410 137.740 1485.730 137.800 ;
        RECT 1483.570 22.000 1483.890 22.060 ;
        RECT 1485.410 22.000 1485.730 22.060 ;
        RECT 1483.570 21.860 1485.730 22.000 ;
        RECT 1483.570 21.800 1483.890 21.860 ;
        RECT 1485.410 21.800 1485.730 21.860 ;
      LAYER via ;
        RECT 1483.140 243.820 1483.400 244.080 ;
        RECT 1484.520 243.820 1484.780 244.080 ;
        RECT 1484.520 206.760 1484.780 207.020 ;
        RECT 1485.440 206.760 1485.700 207.020 ;
        RECT 1484.980 144.880 1485.240 145.140 ;
        RECT 1485.440 144.880 1485.700 145.140 ;
        RECT 1484.980 137.740 1485.240 138.000 ;
        RECT 1485.440 137.740 1485.700 138.000 ;
        RECT 1483.600 21.800 1483.860 22.060 ;
        RECT 1485.440 21.800 1485.700 22.060 ;
      LAYER met2 ;
        RECT 1480.790 260.850 1481.070 264.000 ;
        RECT 1480.790 260.710 1483.340 260.850 ;
        RECT 1480.790 260.000 1481.070 260.710 ;
        RECT 1483.200 244.110 1483.340 260.710 ;
        RECT 1483.140 243.790 1483.400 244.110 ;
        RECT 1484.520 243.790 1484.780 244.110 ;
        RECT 1484.580 207.050 1484.720 243.790 ;
        RECT 1484.520 206.730 1484.780 207.050 ;
        RECT 1485.440 206.730 1485.700 207.050 ;
        RECT 1485.500 145.170 1485.640 206.730 ;
        RECT 1484.980 144.850 1485.240 145.170 ;
        RECT 1485.440 144.850 1485.700 145.170 ;
        RECT 1485.040 138.030 1485.180 144.850 ;
        RECT 1484.980 137.710 1485.240 138.030 ;
        RECT 1485.440 137.710 1485.700 138.030 ;
        RECT 1485.500 22.090 1485.640 137.710 ;
        RECT 1483.600 21.770 1483.860 22.090 ;
        RECT 1485.440 21.770 1485.700 22.090 ;
        RECT 1483.660 2.400 1483.800 21.770 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.910 20.640 1497.230 20.700 ;
        RECT 1501.510 20.640 1501.830 20.700 ;
        RECT 1496.910 20.500 1501.830 20.640 ;
        RECT 1496.910 20.440 1497.230 20.500 ;
        RECT 1501.510 20.440 1501.830 20.500 ;
      LAYER via ;
        RECT 1496.940 20.440 1497.200 20.700 ;
        RECT 1501.540 20.440 1501.800 20.700 ;
      LAYER met2 ;
        RECT 1495.050 260.170 1495.330 264.000 ;
        RECT 1495.050 260.030 1497.140 260.170 ;
        RECT 1495.050 260.000 1495.330 260.030 ;
        RECT 1497.000 20.730 1497.140 260.030 ;
        RECT 1496.940 20.410 1497.200 20.730 ;
        RECT 1501.540 20.410 1501.800 20.730 ;
        RECT 1501.600 2.400 1501.740 20.410 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.250 17.920 1510.570 17.980 ;
        RECT 1518.990 17.920 1519.310 17.980 ;
        RECT 1510.250 17.780 1519.310 17.920 ;
        RECT 1510.250 17.720 1510.570 17.780 ;
        RECT 1518.990 17.720 1519.310 17.780 ;
      LAYER via ;
        RECT 1510.280 17.720 1510.540 17.980 ;
        RECT 1519.020 17.720 1519.280 17.980 ;
      LAYER met2 ;
        RECT 1509.310 260.170 1509.590 264.000 ;
        RECT 1509.310 260.030 1510.480 260.170 ;
        RECT 1509.310 260.000 1509.590 260.030 ;
        RECT 1510.340 18.010 1510.480 260.030 ;
        RECT 1510.280 17.690 1510.540 18.010 ;
        RECT 1519.020 17.690 1519.280 18.010 ;
        RECT 1519.080 2.400 1519.220 17.690 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.470 231.100 869.790 231.160 ;
        RECT 874.070 231.100 874.390 231.160 ;
        RECT 869.470 230.960 874.390 231.100 ;
        RECT 869.470 230.900 869.790 230.960 ;
        RECT 874.070 230.900 874.390 230.960 ;
        RECT 869.470 18.260 869.790 18.320 ;
        RECT 718.220 18.120 745.960 18.260 ;
        RECT 716.290 17.920 716.610 17.980 ;
        RECT 718.220 17.920 718.360 18.120 ;
        RECT 716.290 17.780 718.360 17.920 ;
        RECT 716.290 17.720 716.610 17.780 ;
        RECT 745.820 17.580 745.960 18.120 ;
        RECT 858.520 18.120 869.790 18.260 ;
        RECT 858.520 17.920 858.660 18.120 ;
        RECT 869.470 18.060 869.790 18.120 ;
        RECT 786.760 17.780 858.660 17.920 ;
        RECT 786.760 17.580 786.900 17.780 ;
        RECT 745.820 17.440 786.900 17.580 ;
      LAYER via ;
        RECT 869.500 230.900 869.760 231.160 ;
        RECT 874.100 230.900 874.360 231.160 ;
        RECT 716.320 17.720 716.580 17.980 ;
        RECT 869.500 18.060 869.760 18.320 ;
      LAYER met2 ;
        RECT 875.430 260.170 875.710 264.000 ;
        RECT 874.160 260.030 875.710 260.170 ;
        RECT 874.160 231.190 874.300 260.030 ;
        RECT 875.430 260.000 875.710 260.030 ;
        RECT 869.500 230.870 869.760 231.190 ;
        RECT 874.100 230.870 874.360 231.190 ;
        RECT 869.560 18.350 869.700 230.870 ;
        RECT 869.500 18.030 869.760 18.350 ;
        RECT 716.320 17.690 716.580 18.010 ;
        RECT 716.380 2.400 716.520 17.690 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.050 20.300 1524.370 20.360 ;
        RECT 1536.930 20.300 1537.250 20.360 ;
        RECT 1524.050 20.160 1537.250 20.300 ;
        RECT 1524.050 20.100 1524.370 20.160 ;
        RECT 1536.930 20.100 1537.250 20.160 ;
      LAYER via ;
        RECT 1524.080 20.100 1524.340 20.360 ;
        RECT 1536.960 20.100 1537.220 20.360 ;
      LAYER met2 ;
        RECT 1523.110 260.170 1523.390 264.000 ;
        RECT 1523.110 260.030 1524.280 260.170 ;
        RECT 1523.110 260.000 1523.390 260.030 ;
        RECT 1524.140 20.390 1524.280 260.030 ;
        RECT 1524.080 20.070 1524.340 20.390 ;
        RECT 1536.960 20.070 1537.220 20.390 ;
        RECT 1537.020 2.400 1537.160 20.070 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.310 17.240 1538.630 17.300 ;
        RECT 1554.870 17.240 1555.190 17.300 ;
        RECT 1538.310 17.100 1555.190 17.240 ;
        RECT 1538.310 17.040 1538.630 17.100 ;
        RECT 1554.870 17.040 1555.190 17.100 ;
      LAYER via ;
        RECT 1538.340 17.040 1538.600 17.300 ;
        RECT 1554.900 17.040 1555.160 17.300 ;
      LAYER met2 ;
        RECT 1537.370 260.170 1537.650 264.000 ;
        RECT 1537.370 260.030 1538.540 260.170 ;
        RECT 1537.370 260.000 1537.650 260.030 ;
        RECT 1538.400 17.330 1538.540 260.030 ;
        RECT 1538.340 17.010 1538.600 17.330 ;
        RECT 1554.900 17.010 1555.160 17.330 ;
        RECT 1554.960 2.400 1555.100 17.010 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1551.650 16.900 1551.970 16.960 ;
        RECT 1572.810 16.900 1573.130 16.960 ;
        RECT 1551.650 16.760 1573.130 16.900 ;
        RECT 1551.650 16.700 1551.970 16.760 ;
        RECT 1572.810 16.700 1573.130 16.760 ;
      LAYER via ;
        RECT 1551.680 16.700 1551.940 16.960 ;
        RECT 1572.840 16.700 1573.100 16.960 ;
      LAYER met2 ;
        RECT 1551.170 260.170 1551.450 264.000 ;
        RECT 1551.170 260.030 1551.880 260.170 ;
        RECT 1551.170 260.000 1551.450 260.030 ;
        RECT 1551.740 16.990 1551.880 260.030 ;
        RECT 1551.680 16.670 1551.940 16.990 ;
        RECT 1572.840 16.670 1573.100 16.990 ;
        RECT 1572.900 2.400 1573.040 16.670 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.450 18.600 1565.770 18.660 ;
        RECT 1590.290 18.600 1590.610 18.660 ;
        RECT 1565.450 18.460 1590.610 18.600 ;
        RECT 1565.450 18.400 1565.770 18.460 ;
        RECT 1590.290 18.400 1590.610 18.460 ;
      LAYER via ;
        RECT 1565.480 18.400 1565.740 18.660 ;
        RECT 1590.320 18.400 1590.580 18.660 ;
      LAYER met2 ;
        RECT 1565.430 260.000 1565.710 264.000 ;
        RECT 1565.540 18.690 1565.680 260.000 ;
        RECT 1565.480 18.370 1565.740 18.690 ;
        RECT 1590.320 18.370 1590.580 18.690 ;
        RECT 1590.380 2.400 1590.520 18.370 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.250 17.240 1579.570 17.300 ;
        RECT 1608.230 17.240 1608.550 17.300 ;
        RECT 1579.250 17.100 1608.550 17.240 ;
        RECT 1579.250 17.040 1579.570 17.100 ;
        RECT 1608.230 17.040 1608.550 17.100 ;
      LAYER via ;
        RECT 1579.280 17.040 1579.540 17.300 ;
        RECT 1608.260 17.040 1608.520 17.300 ;
      LAYER met2 ;
        RECT 1579.690 260.170 1579.970 264.000 ;
        RECT 1579.340 260.030 1579.970 260.170 ;
        RECT 1579.340 17.330 1579.480 260.030 ;
        RECT 1579.690 260.000 1579.970 260.030 ;
        RECT 1579.280 17.010 1579.540 17.330 ;
        RECT 1608.260 17.010 1608.520 17.330 ;
        RECT 1608.320 2.400 1608.460 17.010 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 17.580 1593.830 17.640 ;
        RECT 1626.170 17.580 1626.490 17.640 ;
        RECT 1593.510 17.440 1626.490 17.580 ;
        RECT 1593.510 17.380 1593.830 17.440 ;
        RECT 1626.170 17.380 1626.490 17.440 ;
      LAYER via ;
        RECT 1593.540 17.380 1593.800 17.640 ;
        RECT 1626.200 17.380 1626.460 17.640 ;
      LAYER met2 ;
        RECT 1593.490 260.000 1593.770 264.000 ;
        RECT 1593.600 17.670 1593.740 260.000 ;
        RECT 1593.540 17.350 1593.800 17.670 ;
        RECT 1626.200 17.350 1626.460 17.670 ;
        RECT 1626.260 2.400 1626.400 17.350 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1607.770 244.020 1608.090 244.080 ;
        RECT 1613.750 244.020 1614.070 244.080 ;
        RECT 1607.770 243.880 1614.070 244.020 ;
        RECT 1607.770 243.820 1608.090 243.880 ;
        RECT 1613.750 243.820 1614.070 243.880 ;
        RECT 1613.750 17.920 1614.070 17.980 ;
        RECT 1644.110 17.920 1644.430 17.980 ;
        RECT 1613.750 17.780 1644.430 17.920 ;
        RECT 1613.750 17.720 1614.070 17.780 ;
        RECT 1644.110 17.720 1644.430 17.780 ;
      LAYER via ;
        RECT 1607.800 243.820 1608.060 244.080 ;
        RECT 1613.780 243.820 1614.040 244.080 ;
        RECT 1613.780 17.720 1614.040 17.980 ;
        RECT 1644.140 17.720 1644.400 17.980 ;
      LAYER met2 ;
        RECT 1607.750 260.000 1608.030 264.000 ;
        RECT 1607.860 244.110 1608.000 260.000 ;
        RECT 1607.800 243.790 1608.060 244.110 ;
        RECT 1613.780 243.790 1614.040 244.110 ;
        RECT 1613.840 18.010 1613.980 243.790 ;
        RECT 1613.780 17.690 1614.040 18.010 ;
        RECT 1644.140 17.690 1644.400 18.010 ;
        RECT 1644.200 2.400 1644.340 17.690 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1621.570 248.440 1621.890 248.500 ;
        RECT 1631.690 248.440 1632.010 248.500 ;
        RECT 1621.570 248.300 1632.010 248.440 ;
        RECT 1621.570 248.240 1621.890 248.300 ;
        RECT 1631.690 248.240 1632.010 248.300 ;
        RECT 1631.690 17.580 1632.010 17.640 ;
        RECT 1662.050 17.580 1662.370 17.640 ;
        RECT 1631.690 17.440 1662.370 17.580 ;
        RECT 1631.690 17.380 1632.010 17.440 ;
        RECT 1662.050 17.380 1662.370 17.440 ;
      LAYER via ;
        RECT 1621.600 248.240 1621.860 248.500 ;
        RECT 1631.720 248.240 1631.980 248.500 ;
        RECT 1631.720 17.380 1631.980 17.640 ;
        RECT 1662.080 17.380 1662.340 17.640 ;
      LAYER met2 ;
        RECT 1621.550 260.000 1621.830 264.000 ;
        RECT 1621.660 248.530 1621.800 260.000 ;
        RECT 1621.600 248.210 1621.860 248.530 ;
        RECT 1631.720 248.210 1631.980 248.530 ;
        RECT 1631.780 17.670 1631.920 248.210 ;
        RECT 1631.720 17.350 1631.980 17.670 ;
        RECT 1662.080 17.350 1662.340 17.670 ;
        RECT 1662.140 2.400 1662.280 17.350 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1635.830 244.020 1636.150 244.080 ;
        RECT 1641.810 244.020 1642.130 244.080 ;
        RECT 1635.830 243.880 1642.130 244.020 ;
        RECT 1635.830 243.820 1636.150 243.880 ;
        RECT 1641.810 243.820 1642.130 243.880 ;
        RECT 1641.810 19.280 1642.130 19.340 ;
        RECT 1679.530 19.280 1679.850 19.340 ;
        RECT 1641.810 19.140 1679.850 19.280 ;
        RECT 1641.810 19.080 1642.130 19.140 ;
        RECT 1679.530 19.080 1679.850 19.140 ;
      LAYER via ;
        RECT 1635.860 243.820 1636.120 244.080 ;
        RECT 1641.840 243.820 1642.100 244.080 ;
        RECT 1641.840 19.080 1642.100 19.340 ;
        RECT 1679.560 19.080 1679.820 19.340 ;
      LAYER met2 ;
        RECT 1635.810 260.000 1636.090 264.000 ;
        RECT 1635.920 244.110 1636.060 260.000 ;
        RECT 1635.860 243.790 1636.120 244.110 ;
        RECT 1641.840 243.790 1642.100 244.110 ;
        RECT 1641.900 19.370 1642.040 243.790 ;
        RECT 1641.840 19.050 1642.100 19.370 ;
        RECT 1679.560 19.050 1679.820 19.370 ;
        RECT 1679.620 2.400 1679.760 19.050 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1650.090 244.020 1650.410 244.080 ;
        RECT 1655.610 244.020 1655.930 244.080 ;
        RECT 1650.090 243.880 1655.930 244.020 ;
        RECT 1650.090 243.820 1650.410 243.880 ;
        RECT 1655.610 243.820 1655.930 243.880 ;
        RECT 1655.610 20.300 1655.930 20.360 ;
        RECT 1697.470 20.300 1697.790 20.360 ;
        RECT 1655.610 20.160 1697.790 20.300 ;
        RECT 1655.610 20.100 1655.930 20.160 ;
        RECT 1697.470 20.100 1697.790 20.160 ;
      LAYER via ;
        RECT 1650.120 243.820 1650.380 244.080 ;
        RECT 1655.640 243.820 1655.900 244.080 ;
        RECT 1655.640 20.100 1655.900 20.360 ;
        RECT 1697.500 20.100 1697.760 20.360 ;
      LAYER met2 ;
        RECT 1650.070 260.000 1650.350 264.000 ;
        RECT 1650.180 244.110 1650.320 260.000 ;
        RECT 1650.120 243.790 1650.380 244.110 ;
        RECT 1655.640 243.790 1655.900 244.110 ;
        RECT 1655.700 20.390 1655.840 243.790 ;
        RECT 1655.640 20.070 1655.900 20.390 ;
        RECT 1697.500 20.070 1697.760 20.390 ;
        RECT 1697.560 2.400 1697.700 20.070 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 883.270 234.500 883.590 234.560 ;
        RECT 887.870 234.500 888.190 234.560 ;
        RECT 883.270 234.360 888.190 234.500 ;
        RECT 883.270 234.300 883.590 234.360 ;
        RECT 887.870 234.300 888.190 234.360 ;
        RECT 734.230 18.600 734.550 18.660 ;
        RECT 883.270 18.600 883.590 18.660 ;
        RECT 734.230 18.460 883.590 18.600 ;
        RECT 734.230 18.400 734.550 18.460 ;
        RECT 883.270 18.400 883.590 18.460 ;
      LAYER via ;
        RECT 883.300 234.300 883.560 234.560 ;
        RECT 887.900 234.300 888.160 234.560 ;
        RECT 734.260 18.400 734.520 18.660 ;
        RECT 883.300 18.400 883.560 18.660 ;
      LAYER met2 ;
        RECT 889.690 260.170 889.970 264.000 ;
        RECT 887.960 260.030 889.970 260.170 ;
        RECT 887.960 234.590 888.100 260.030 ;
        RECT 889.690 260.000 889.970 260.030 ;
        RECT 883.300 234.270 883.560 234.590 ;
        RECT 887.900 234.270 888.160 234.590 ;
        RECT 883.360 18.690 883.500 234.270 ;
        RECT 734.260 18.370 734.520 18.690 ;
        RECT 883.300 18.370 883.560 18.690 ;
        RECT 734.320 2.400 734.460 18.370 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1663.890 244.020 1664.210 244.080 ;
        RECT 1669.410 244.020 1669.730 244.080 ;
        RECT 1663.890 243.880 1669.730 244.020 ;
        RECT 1663.890 243.820 1664.210 243.880 ;
        RECT 1669.410 243.820 1669.730 243.880 ;
        RECT 1669.410 16.900 1669.730 16.960 ;
        RECT 1715.410 16.900 1715.730 16.960 ;
        RECT 1669.410 16.760 1715.730 16.900 ;
        RECT 1669.410 16.700 1669.730 16.760 ;
        RECT 1715.410 16.700 1715.730 16.760 ;
      LAYER via ;
        RECT 1663.920 243.820 1664.180 244.080 ;
        RECT 1669.440 243.820 1669.700 244.080 ;
        RECT 1669.440 16.700 1669.700 16.960 ;
        RECT 1715.440 16.700 1715.700 16.960 ;
      LAYER met2 ;
        RECT 1663.870 260.000 1664.150 264.000 ;
        RECT 1663.980 244.110 1664.120 260.000 ;
        RECT 1663.920 243.790 1664.180 244.110 ;
        RECT 1669.440 243.790 1669.700 244.110 ;
        RECT 1669.500 16.990 1669.640 243.790 ;
        RECT 1669.440 16.670 1669.700 16.990 ;
        RECT 1715.440 16.670 1715.700 16.990 ;
        RECT 1715.500 2.400 1715.640 16.670 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1678.150 244.020 1678.470 244.080 ;
        RECT 1683.210 244.020 1683.530 244.080 ;
        RECT 1678.150 243.880 1683.530 244.020 ;
        RECT 1678.150 243.820 1678.470 243.880 ;
        RECT 1683.210 243.820 1683.530 243.880 ;
        RECT 1683.210 19.280 1683.530 19.340 ;
        RECT 1733.350 19.280 1733.670 19.340 ;
        RECT 1683.210 19.140 1733.670 19.280 ;
        RECT 1683.210 19.080 1683.530 19.140 ;
        RECT 1733.350 19.080 1733.670 19.140 ;
      LAYER via ;
        RECT 1678.180 243.820 1678.440 244.080 ;
        RECT 1683.240 243.820 1683.500 244.080 ;
        RECT 1683.240 19.080 1683.500 19.340 ;
        RECT 1733.380 19.080 1733.640 19.340 ;
      LAYER met2 ;
        RECT 1678.130 260.000 1678.410 264.000 ;
        RECT 1678.240 244.110 1678.380 260.000 ;
        RECT 1678.180 243.790 1678.440 244.110 ;
        RECT 1683.240 243.790 1683.500 244.110 ;
        RECT 1683.300 19.370 1683.440 243.790 ;
        RECT 1683.240 19.050 1683.500 19.370 ;
        RECT 1733.380 19.050 1733.640 19.370 ;
        RECT 1733.440 2.400 1733.580 19.050 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1692.410 244.020 1692.730 244.080 ;
        RECT 1697.010 244.020 1697.330 244.080 ;
        RECT 1692.410 243.880 1697.330 244.020 ;
        RECT 1692.410 243.820 1692.730 243.880 ;
        RECT 1697.010 243.820 1697.330 243.880 ;
        RECT 1697.010 18.940 1697.330 19.000 ;
        RECT 1751.290 18.940 1751.610 19.000 ;
        RECT 1697.010 18.800 1751.610 18.940 ;
        RECT 1697.010 18.740 1697.330 18.800 ;
        RECT 1751.290 18.740 1751.610 18.800 ;
      LAYER via ;
        RECT 1692.440 243.820 1692.700 244.080 ;
        RECT 1697.040 243.820 1697.300 244.080 ;
        RECT 1697.040 18.740 1697.300 19.000 ;
        RECT 1751.320 18.740 1751.580 19.000 ;
      LAYER met2 ;
        RECT 1692.390 260.000 1692.670 264.000 ;
        RECT 1692.500 244.110 1692.640 260.000 ;
        RECT 1692.440 243.790 1692.700 244.110 ;
        RECT 1697.040 243.790 1697.300 244.110 ;
        RECT 1697.100 19.030 1697.240 243.790 ;
        RECT 1697.040 18.710 1697.300 19.030 ;
        RECT 1751.320 18.710 1751.580 19.030 ;
        RECT 1751.380 2.400 1751.520 18.710 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1706.210 244.020 1706.530 244.080 ;
        RECT 1710.810 244.020 1711.130 244.080 ;
        RECT 1706.210 243.880 1711.130 244.020 ;
        RECT 1706.210 243.820 1706.530 243.880 ;
        RECT 1710.810 243.820 1711.130 243.880 ;
        RECT 1710.810 20.300 1711.130 20.360 ;
        RECT 1768.770 20.300 1769.090 20.360 ;
        RECT 1710.810 20.160 1769.090 20.300 ;
        RECT 1710.810 20.100 1711.130 20.160 ;
        RECT 1768.770 20.100 1769.090 20.160 ;
      LAYER via ;
        RECT 1706.240 243.820 1706.500 244.080 ;
        RECT 1710.840 243.820 1711.100 244.080 ;
        RECT 1710.840 20.100 1711.100 20.360 ;
        RECT 1768.800 20.100 1769.060 20.360 ;
      LAYER met2 ;
        RECT 1706.190 260.000 1706.470 264.000 ;
        RECT 1706.300 244.110 1706.440 260.000 ;
        RECT 1706.240 243.790 1706.500 244.110 ;
        RECT 1710.840 243.790 1711.100 244.110 ;
        RECT 1710.900 20.390 1711.040 243.790 ;
        RECT 1710.840 20.070 1711.100 20.390 ;
        RECT 1768.800 20.070 1769.060 20.390 ;
        RECT 1768.860 2.400 1769.000 20.070 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1720.470 244.020 1720.790 244.080 ;
        RECT 1724.610 244.020 1724.930 244.080 ;
        RECT 1720.470 243.880 1724.930 244.020 ;
        RECT 1720.470 243.820 1720.790 243.880 ;
        RECT 1724.610 243.820 1724.930 243.880 ;
        RECT 1724.610 16.220 1724.930 16.280 ;
        RECT 1786.710 16.220 1787.030 16.280 ;
        RECT 1724.610 16.080 1787.030 16.220 ;
        RECT 1724.610 16.020 1724.930 16.080 ;
        RECT 1786.710 16.020 1787.030 16.080 ;
      LAYER via ;
        RECT 1720.500 243.820 1720.760 244.080 ;
        RECT 1724.640 243.820 1724.900 244.080 ;
        RECT 1724.640 16.020 1724.900 16.280 ;
        RECT 1786.740 16.020 1787.000 16.280 ;
      LAYER met2 ;
        RECT 1720.450 260.000 1720.730 264.000 ;
        RECT 1720.560 244.110 1720.700 260.000 ;
        RECT 1720.500 243.790 1720.760 244.110 ;
        RECT 1724.640 243.790 1724.900 244.110 ;
        RECT 1724.700 16.310 1724.840 243.790 ;
        RECT 1724.640 15.990 1724.900 16.310 ;
        RECT 1786.740 15.990 1787.000 16.310 ;
        RECT 1786.800 2.400 1786.940 15.990 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1734.270 242.660 1734.590 242.720 ;
        RECT 1738.410 242.660 1738.730 242.720 ;
        RECT 1734.270 242.520 1738.730 242.660 ;
        RECT 1734.270 242.460 1734.590 242.520 ;
        RECT 1738.410 242.460 1738.730 242.520 ;
        RECT 1738.410 19.620 1738.730 19.680 ;
        RECT 1804.650 19.620 1804.970 19.680 ;
        RECT 1738.410 19.480 1804.970 19.620 ;
        RECT 1738.410 19.420 1738.730 19.480 ;
        RECT 1804.650 19.420 1804.970 19.480 ;
      LAYER via ;
        RECT 1734.300 242.460 1734.560 242.720 ;
        RECT 1738.440 242.460 1738.700 242.720 ;
        RECT 1738.440 19.420 1738.700 19.680 ;
        RECT 1804.680 19.420 1804.940 19.680 ;
      LAYER met2 ;
        RECT 1734.250 260.000 1734.530 264.000 ;
        RECT 1734.360 242.750 1734.500 260.000 ;
        RECT 1734.300 242.430 1734.560 242.750 ;
        RECT 1738.440 242.430 1738.700 242.750 ;
        RECT 1738.500 19.710 1738.640 242.430 ;
        RECT 1738.440 19.390 1738.700 19.710 ;
        RECT 1804.680 19.390 1804.940 19.710 ;
        RECT 1804.740 2.400 1804.880 19.390 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1752.210 20.640 1752.530 20.700 ;
        RECT 1822.590 20.640 1822.910 20.700 ;
        RECT 1752.210 20.500 1822.910 20.640 ;
        RECT 1752.210 20.440 1752.530 20.500 ;
        RECT 1822.590 20.440 1822.910 20.500 ;
      LAYER via ;
        RECT 1752.240 20.440 1752.500 20.700 ;
        RECT 1822.620 20.440 1822.880 20.700 ;
      LAYER met2 ;
        RECT 1748.510 260.170 1748.790 264.000 ;
        RECT 1748.510 260.030 1752.440 260.170 ;
        RECT 1748.510 260.000 1748.790 260.030 ;
        RECT 1752.300 20.730 1752.440 260.030 ;
        RECT 1752.240 20.410 1752.500 20.730 ;
        RECT 1822.620 20.410 1822.880 20.730 ;
        RECT 1822.680 2.400 1822.820 20.410 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.010 16.560 1766.330 16.620 ;
        RECT 1840.070 16.560 1840.390 16.620 ;
        RECT 1766.010 16.420 1840.390 16.560 ;
        RECT 1766.010 16.360 1766.330 16.420 ;
        RECT 1840.070 16.360 1840.390 16.420 ;
      LAYER via ;
        RECT 1766.040 16.360 1766.300 16.620 ;
        RECT 1840.100 16.360 1840.360 16.620 ;
      LAYER met2 ;
        RECT 1762.770 260.170 1763.050 264.000 ;
        RECT 1762.770 260.030 1766.240 260.170 ;
        RECT 1762.770 260.000 1763.050 260.030 ;
        RECT 1766.100 16.650 1766.240 260.030 ;
        RECT 1766.040 16.330 1766.300 16.650 ;
        RECT 1840.100 16.330 1840.360 16.650 ;
        RECT 1840.160 2.400 1840.300 16.330 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1779.810 18.260 1780.130 18.320 ;
        RECT 1858.010 18.260 1858.330 18.320 ;
        RECT 1779.810 18.120 1858.330 18.260 ;
        RECT 1779.810 18.060 1780.130 18.120 ;
        RECT 1858.010 18.060 1858.330 18.120 ;
      LAYER via ;
        RECT 1779.840 18.060 1780.100 18.320 ;
        RECT 1858.040 18.060 1858.300 18.320 ;
      LAYER met2 ;
        RECT 1776.570 260.170 1776.850 264.000 ;
        RECT 1776.570 260.030 1780.040 260.170 ;
        RECT 1776.570 260.000 1776.850 260.030 ;
        RECT 1779.900 18.350 1780.040 260.030 ;
        RECT 1779.840 18.030 1780.100 18.350 ;
        RECT 1858.040 18.030 1858.300 18.350 ;
        RECT 1858.100 2.400 1858.240 18.030 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 16.900 1793.930 16.960 ;
        RECT 1875.950 16.900 1876.270 16.960 ;
        RECT 1793.610 16.760 1876.270 16.900 ;
        RECT 1793.610 16.700 1793.930 16.760 ;
        RECT 1875.950 16.700 1876.270 16.760 ;
      LAYER via ;
        RECT 1793.640 16.700 1793.900 16.960 ;
        RECT 1875.980 16.700 1876.240 16.960 ;
      LAYER met2 ;
        RECT 1790.830 260.170 1791.110 264.000 ;
        RECT 1790.830 260.030 1793.840 260.170 ;
        RECT 1790.830 260.000 1791.110 260.030 ;
        RECT 1793.700 16.990 1793.840 260.030 ;
        RECT 1793.640 16.670 1793.900 16.990 ;
        RECT 1875.980 16.670 1876.240 16.990 ;
        RECT 1876.040 2.400 1876.180 16.670 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 897.070 244.020 897.390 244.080 ;
        RECT 901.670 244.020 901.990 244.080 ;
        RECT 897.070 243.880 901.990 244.020 ;
        RECT 897.070 243.820 897.390 243.880 ;
        RECT 901.670 243.820 901.990 243.880 ;
        RECT 752.170 19.620 752.490 19.680 ;
        RECT 897.070 19.620 897.390 19.680 ;
        RECT 752.170 19.480 897.390 19.620 ;
        RECT 752.170 19.420 752.490 19.480 ;
        RECT 897.070 19.420 897.390 19.480 ;
      LAYER via ;
        RECT 897.100 243.820 897.360 244.080 ;
        RECT 901.700 243.820 901.960 244.080 ;
        RECT 752.200 19.420 752.460 19.680 ;
        RECT 897.100 19.420 897.360 19.680 ;
      LAYER met2 ;
        RECT 903.490 260.170 903.770 264.000 ;
        RECT 901.760 260.030 903.770 260.170 ;
        RECT 901.760 244.110 901.900 260.030 ;
        RECT 903.490 260.000 903.770 260.030 ;
        RECT 897.100 243.790 897.360 244.110 ;
        RECT 901.700 243.790 901.960 244.110 ;
        RECT 897.160 19.710 897.300 243.790 ;
        RECT 752.200 19.390 752.460 19.710 ;
        RECT 897.100 19.390 897.360 19.710 ;
        RECT 752.260 2.400 752.400 19.390 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.410 19.960 1807.730 20.020 ;
        RECT 1893.890 19.960 1894.210 20.020 ;
        RECT 1807.410 19.820 1894.210 19.960 ;
        RECT 1807.410 19.760 1807.730 19.820 ;
        RECT 1893.890 19.760 1894.210 19.820 ;
      LAYER via ;
        RECT 1807.440 19.760 1807.700 20.020 ;
        RECT 1893.920 19.760 1894.180 20.020 ;
      LAYER met2 ;
        RECT 1804.630 260.170 1804.910 264.000 ;
        RECT 1804.630 260.030 1807.640 260.170 ;
        RECT 1804.630 260.000 1804.910 260.030 ;
        RECT 1807.500 20.050 1807.640 260.030 ;
        RECT 1807.440 19.730 1807.700 20.050 ;
        RECT 1893.920 19.730 1894.180 20.050 ;
        RECT 1893.980 2.400 1894.120 19.730 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 19.620 1821.530 19.680 ;
        RECT 1911.830 19.620 1912.150 19.680 ;
        RECT 1821.210 19.480 1912.150 19.620 ;
        RECT 1821.210 19.420 1821.530 19.480 ;
        RECT 1911.830 19.420 1912.150 19.480 ;
      LAYER via ;
        RECT 1821.240 19.420 1821.500 19.680 ;
        RECT 1911.860 19.420 1912.120 19.680 ;
      LAYER met2 ;
        RECT 1818.890 260.170 1819.170 264.000 ;
        RECT 1818.890 260.030 1821.440 260.170 ;
        RECT 1818.890 260.000 1819.170 260.030 ;
        RECT 1821.300 19.710 1821.440 260.030 ;
        RECT 1821.240 19.390 1821.500 19.710 ;
        RECT 1911.860 19.390 1912.120 19.710 ;
        RECT 1911.920 2.400 1912.060 19.390 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1835.010 20.640 1835.330 20.700 ;
        RECT 1929.310 20.640 1929.630 20.700 ;
        RECT 1835.010 20.500 1929.630 20.640 ;
        RECT 1835.010 20.440 1835.330 20.500 ;
        RECT 1929.310 20.440 1929.630 20.500 ;
      LAYER via ;
        RECT 1835.040 20.440 1835.300 20.700 ;
        RECT 1929.340 20.440 1929.600 20.700 ;
      LAYER met2 ;
        RECT 1833.150 260.170 1833.430 264.000 ;
        RECT 1833.150 260.030 1835.240 260.170 ;
        RECT 1833.150 260.000 1833.430 260.030 ;
        RECT 1835.100 20.730 1835.240 260.030 ;
        RECT 1835.040 20.410 1835.300 20.730 ;
        RECT 1929.340 20.410 1929.600 20.730 ;
        RECT 1929.400 2.400 1929.540 20.410 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.810 17.920 1849.130 17.980 ;
        RECT 1947.250 17.920 1947.570 17.980 ;
        RECT 1848.810 17.780 1947.570 17.920 ;
        RECT 1848.810 17.720 1849.130 17.780 ;
        RECT 1947.250 17.720 1947.570 17.780 ;
      LAYER via ;
        RECT 1848.840 17.720 1849.100 17.980 ;
        RECT 1947.280 17.720 1947.540 17.980 ;
      LAYER met2 ;
        RECT 1846.950 260.170 1847.230 264.000 ;
        RECT 1846.950 260.030 1849.040 260.170 ;
        RECT 1846.950 260.000 1847.230 260.030 ;
        RECT 1848.900 18.010 1849.040 260.030 ;
        RECT 1848.840 17.690 1849.100 18.010 ;
        RECT 1947.280 17.690 1947.540 18.010 ;
        RECT 1947.340 2.400 1947.480 17.690 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 20.300 1862.930 20.360 ;
        RECT 1965.190 20.300 1965.510 20.360 ;
        RECT 1862.610 20.160 1965.510 20.300 ;
        RECT 1862.610 20.100 1862.930 20.160 ;
        RECT 1965.190 20.100 1965.510 20.160 ;
      LAYER via ;
        RECT 1862.640 20.100 1862.900 20.360 ;
        RECT 1965.220 20.100 1965.480 20.360 ;
      LAYER met2 ;
        RECT 1861.210 260.170 1861.490 264.000 ;
        RECT 1861.210 260.030 1862.840 260.170 ;
        RECT 1861.210 260.000 1861.490 260.030 ;
        RECT 1862.700 20.390 1862.840 260.030 ;
        RECT 1862.640 20.070 1862.900 20.390 ;
        RECT 1965.220 20.070 1965.480 20.390 ;
        RECT 1965.280 2.400 1965.420 20.070 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1875.950 17.580 1876.270 17.640 ;
        RECT 1983.130 17.580 1983.450 17.640 ;
        RECT 1875.950 17.440 1983.450 17.580 ;
        RECT 1875.950 17.380 1876.270 17.440 ;
        RECT 1983.130 17.380 1983.450 17.440 ;
      LAYER via ;
        RECT 1875.980 17.380 1876.240 17.640 ;
        RECT 1983.160 17.380 1983.420 17.640 ;
      LAYER met2 ;
        RECT 1875.010 260.170 1875.290 264.000 ;
        RECT 1875.010 260.030 1876.180 260.170 ;
        RECT 1875.010 260.000 1875.290 260.030 ;
        RECT 1876.040 17.670 1876.180 260.030 ;
        RECT 1875.980 17.350 1876.240 17.670 ;
        RECT 1983.160 17.350 1983.420 17.670 ;
        RECT 1983.220 2.400 1983.360 17.350 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1889.750 18.260 1890.070 18.320 ;
        RECT 2001.070 18.260 2001.390 18.320 ;
        RECT 1889.750 18.120 2001.390 18.260 ;
        RECT 1889.750 18.060 1890.070 18.120 ;
        RECT 2001.070 18.060 2001.390 18.120 ;
      LAYER via ;
        RECT 1889.780 18.060 1890.040 18.320 ;
        RECT 2001.100 18.060 2001.360 18.320 ;
      LAYER met2 ;
        RECT 1889.270 260.170 1889.550 264.000 ;
        RECT 1889.270 260.030 1889.980 260.170 ;
        RECT 1889.270 260.000 1889.550 260.030 ;
        RECT 1889.840 18.350 1889.980 260.030 ;
        RECT 1889.780 18.030 1890.040 18.350 ;
        RECT 2001.100 18.030 2001.360 18.350 ;
        RECT 2001.160 2.400 2001.300 18.030 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1903.550 17.240 1903.870 17.300 ;
        RECT 2018.550 17.240 2018.870 17.300 ;
        RECT 1903.550 17.100 2018.870 17.240 ;
        RECT 1903.550 17.040 1903.870 17.100 ;
        RECT 2018.550 17.040 2018.870 17.100 ;
      LAYER via ;
        RECT 1903.580 17.040 1903.840 17.300 ;
        RECT 2018.580 17.040 2018.840 17.300 ;
      LAYER met2 ;
        RECT 1903.530 260.000 1903.810 264.000 ;
        RECT 1903.640 17.330 1903.780 260.000 ;
        RECT 1903.580 17.010 1903.840 17.330 ;
        RECT 2018.580 17.010 2018.840 17.330 ;
        RECT 2018.640 2.400 2018.780 17.010 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 18.600 1918.130 18.660 ;
        RECT 2036.490 18.600 2036.810 18.660 ;
        RECT 1917.810 18.460 2036.810 18.600 ;
        RECT 1917.810 18.400 1918.130 18.460 ;
        RECT 2036.490 18.400 2036.810 18.460 ;
      LAYER via ;
        RECT 1917.840 18.400 1918.100 18.660 ;
        RECT 2036.520 18.400 2036.780 18.660 ;
      LAYER met2 ;
        RECT 1917.330 260.170 1917.610 264.000 ;
        RECT 1917.330 260.030 1918.040 260.170 ;
        RECT 1917.330 260.000 1917.610 260.030 ;
        RECT 1917.900 18.690 1918.040 260.030 ;
        RECT 1917.840 18.370 1918.100 18.690 ;
        RECT 2036.520 18.370 2036.780 18.690 ;
        RECT 2036.580 2.400 2036.720 18.370 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.610 19.620 1931.930 19.680 ;
        RECT 2054.430 19.620 2054.750 19.680 ;
        RECT 1931.610 19.480 2054.750 19.620 ;
        RECT 1931.610 19.420 1931.930 19.480 ;
        RECT 2054.430 19.420 2054.750 19.480 ;
      LAYER via ;
        RECT 1931.640 19.420 1931.900 19.680 ;
        RECT 2054.460 19.420 2054.720 19.680 ;
      LAYER met2 ;
        RECT 1931.590 260.000 1931.870 264.000 ;
        RECT 1931.700 19.710 1931.840 260.000 ;
        RECT 1931.640 19.390 1931.900 19.710 ;
        RECT 2054.460 19.390 2054.720 19.710 ;
        RECT 2054.520 2.400 2054.660 19.390 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 769.650 19.280 769.970 19.340 ;
        RECT 917.770 19.280 918.090 19.340 ;
        RECT 769.650 19.140 918.090 19.280 ;
        RECT 769.650 19.080 769.970 19.140 ;
        RECT 917.770 19.080 918.090 19.140 ;
      LAYER via ;
        RECT 769.680 19.080 769.940 19.340 ;
        RECT 917.800 19.080 918.060 19.340 ;
      LAYER met2 ;
        RECT 917.750 260.000 918.030 264.000 ;
        RECT 917.860 19.370 918.000 260.000 ;
        RECT 769.680 19.050 769.940 19.370 ;
        RECT 917.800 19.050 918.060 19.370 ;
        RECT 769.740 2.400 769.880 19.050 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1945.870 244.020 1946.190 244.080 ;
        RECT 1952.310 244.020 1952.630 244.080 ;
        RECT 1945.870 243.880 1952.630 244.020 ;
        RECT 1945.870 243.820 1946.190 243.880 ;
        RECT 1952.310 243.820 1952.630 243.880 ;
        RECT 1952.310 18.940 1952.630 19.000 ;
        RECT 2072.370 18.940 2072.690 19.000 ;
        RECT 1952.310 18.800 2072.690 18.940 ;
        RECT 1952.310 18.740 1952.630 18.800 ;
        RECT 2072.370 18.740 2072.690 18.800 ;
      LAYER via ;
        RECT 1945.900 243.820 1946.160 244.080 ;
        RECT 1952.340 243.820 1952.600 244.080 ;
        RECT 1952.340 18.740 1952.600 19.000 ;
        RECT 2072.400 18.740 2072.660 19.000 ;
      LAYER met2 ;
        RECT 1945.850 260.000 1946.130 264.000 ;
        RECT 1945.960 244.110 1946.100 260.000 ;
        RECT 1945.900 243.790 1946.160 244.110 ;
        RECT 1952.340 243.790 1952.600 244.110 ;
        RECT 1952.400 19.030 1952.540 243.790 ;
        RECT 1952.340 18.710 1952.600 19.030 ;
        RECT 2072.400 18.710 2072.660 19.030 ;
        RECT 2072.460 2.400 2072.600 18.710 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1959.670 244.020 1959.990 244.080 ;
        RECT 1966.110 244.020 1966.430 244.080 ;
        RECT 1959.670 243.880 1966.430 244.020 ;
        RECT 1959.670 243.820 1959.990 243.880 ;
        RECT 1966.110 243.820 1966.430 243.880 ;
        RECT 1966.110 20.300 1966.430 20.360 ;
        RECT 2089.850 20.300 2090.170 20.360 ;
        RECT 1966.110 20.160 2090.170 20.300 ;
        RECT 1966.110 20.100 1966.430 20.160 ;
        RECT 2089.850 20.100 2090.170 20.160 ;
      LAYER via ;
        RECT 1959.700 243.820 1959.960 244.080 ;
        RECT 1966.140 243.820 1966.400 244.080 ;
        RECT 1966.140 20.100 1966.400 20.360 ;
        RECT 2089.880 20.100 2090.140 20.360 ;
      LAYER met2 ;
        RECT 1959.650 260.000 1959.930 264.000 ;
        RECT 1959.760 244.110 1959.900 260.000 ;
        RECT 1959.700 243.790 1959.960 244.110 ;
        RECT 1966.140 243.790 1966.400 244.110 ;
        RECT 1966.200 20.390 1966.340 243.790 ;
        RECT 1966.140 20.070 1966.400 20.390 ;
        RECT 2089.880 20.070 2090.140 20.390 ;
        RECT 2089.940 2.400 2090.080 20.070 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.930 244.020 1974.250 244.080 ;
        RECT 1979.910 244.020 1980.230 244.080 ;
        RECT 1973.930 243.880 1980.230 244.020 ;
        RECT 1973.930 243.820 1974.250 243.880 ;
        RECT 1979.910 243.820 1980.230 243.880 ;
        RECT 1979.910 17.920 1980.230 17.980 ;
        RECT 2107.790 17.920 2108.110 17.980 ;
        RECT 1979.910 17.780 2108.110 17.920 ;
        RECT 1979.910 17.720 1980.230 17.780 ;
        RECT 2107.790 17.720 2108.110 17.780 ;
      LAYER via ;
        RECT 1973.960 243.820 1974.220 244.080 ;
        RECT 1979.940 243.820 1980.200 244.080 ;
        RECT 1979.940 17.720 1980.200 17.980 ;
        RECT 2107.820 17.720 2108.080 17.980 ;
      LAYER met2 ;
        RECT 1973.910 260.000 1974.190 264.000 ;
        RECT 1974.020 244.110 1974.160 260.000 ;
        RECT 1973.960 243.790 1974.220 244.110 ;
        RECT 1979.940 243.790 1980.200 244.110 ;
        RECT 1980.000 18.010 1980.140 243.790 ;
        RECT 1979.940 17.690 1980.200 18.010 ;
        RECT 2107.820 17.690 2108.080 18.010 ;
        RECT 2107.880 2.400 2108.020 17.690 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1987.730 244.020 1988.050 244.080 ;
        RECT 1993.710 244.020 1994.030 244.080 ;
        RECT 1987.730 243.880 1994.030 244.020 ;
        RECT 1987.730 243.820 1988.050 243.880 ;
        RECT 1993.710 243.820 1994.030 243.880 ;
        RECT 1993.710 17.580 1994.030 17.640 ;
        RECT 2125.730 17.580 2126.050 17.640 ;
        RECT 1993.710 17.440 2126.050 17.580 ;
        RECT 1993.710 17.380 1994.030 17.440 ;
        RECT 2125.730 17.380 2126.050 17.440 ;
      LAYER via ;
        RECT 1987.760 243.820 1988.020 244.080 ;
        RECT 1993.740 243.820 1994.000 244.080 ;
        RECT 1993.740 17.380 1994.000 17.640 ;
        RECT 2125.760 17.380 2126.020 17.640 ;
      LAYER met2 ;
        RECT 1987.710 260.000 1987.990 264.000 ;
        RECT 1987.820 244.110 1987.960 260.000 ;
        RECT 1987.760 243.790 1988.020 244.110 ;
        RECT 1993.740 243.790 1994.000 244.110 ;
        RECT 1993.800 17.670 1993.940 243.790 ;
        RECT 1993.740 17.350 1994.000 17.670 ;
        RECT 2125.760 17.350 2126.020 17.670 ;
        RECT 2125.820 2.400 2125.960 17.350 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2001.990 244.020 2002.310 244.080 ;
        RECT 2007.510 244.020 2007.830 244.080 ;
        RECT 2001.990 243.880 2007.830 244.020 ;
        RECT 2001.990 243.820 2002.310 243.880 ;
        RECT 2007.510 243.820 2007.830 243.880 ;
        RECT 2007.510 18.260 2007.830 18.320 ;
        RECT 2143.670 18.260 2143.990 18.320 ;
        RECT 2007.510 18.120 2143.990 18.260 ;
        RECT 2007.510 18.060 2007.830 18.120 ;
        RECT 2143.670 18.060 2143.990 18.120 ;
      LAYER via ;
        RECT 2002.020 243.820 2002.280 244.080 ;
        RECT 2007.540 243.820 2007.800 244.080 ;
        RECT 2007.540 18.060 2007.800 18.320 ;
        RECT 2143.700 18.060 2143.960 18.320 ;
      LAYER met2 ;
        RECT 2001.970 260.000 2002.250 264.000 ;
        RECT 2002.080 244.110 2002.220 260.000 ;
        RECT 2002.020 243.790 2002.280 244.110 ;
        RECT 2007.540 243.790 2007.800 244.110 ;
        RECT 2007.600 18.350 2007.740 243.790 ;
        RECT 2007.540 18.030 2007.800 18.350 ;
        RECT 2143.700 18.030 2143.960 18.350 ;
        RECT 2143.760 2.400 2143.900 18.030 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2016.250 244.020 2016.570 244.080 ;
        RECT 2021.310 244.020 2021.630 244.080 ;
        RECT 2016.250 243.880 2021.630 244.020 ;
        RECT 2016.250 243.820 2016.570 243.880 ;
        RECT 2021.310 243.820 2021.630 243.880 ;
        RECT 2021.310 17.240 2021.630 17.300 ;
        RECT 2161.610 17.240 2161.930 17.300 ;
        RECT 2021.310 17.100 2161.930 17.240 ;
        RECT 2021.310 17.040 2021.630 17.100 ;
        RECT 2161.610 17.040 2161.930 17.100 ;
      LAYER via ;
        RECT 2016.280 243.820 2016.540 244.080 ;
        RECT 2021.340 243.820 2021.600 244.080 ;
        RECT 2021.340 17.040 2021.600 17.300 ;
        RECT 2161.640 17.040 2161.900 17.300 ;
      LAYER met2 ;
        RECT 2016.230 260.000 2016.510 264.000 ;
        RECT 2016.340 244.110 2016.480 260.000 ;
        RECT 2016.280 243.790 2016.540 244.110 ;
        RECT 2021.340 243.790 2021.600 244.110 ;
        RECT 2021.400 17.330 2021.540 243.790 ;
        RECT 2021.340 17.010 2021.600 17.330 ;
        RECT 2161.640 17.010 2161.900 17.330 ;
        RECT 2161.700 2.400 2161.840 17.010 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2030.050 245.040 2030.370 245.100 ;
        RECT 2173.570 245.040 2173.890 245.100 ;
        RECT 2030.050 244.900 2173.890 245.040 ;
        RECT 2030.050 244.840 2030.370 244.900 ;
        RECT 2173.570 244.840 2173.890 244.900 ;
        RECT 2173.570 2.960 2173.890 3.020 ;
        RECT 2179.090 2.960 2179.410 3.020 ;
        RECT 2173.570 2.820 2179.410 2.960 ;
        RECT 2173.570 2.760 2173.890 2.820 ;
        RECT 2179.090 2.760 2179.410 2.820 ;
      LAYER via ;
        RECT 2030.080 244.840 2030.340 245.100 ;
        RECT 2173.600 244.840 2173.860 245.100 ;
        RECT 2173.600 2.760 2173.860 3.020 ;
        RECT 2179.120 2.760 2179.380 3.020 ;
      LAYER met2 ;
        RECT 2030.030 260.000 2030.310 264.000 ;
        RECT 2030.140 245.130 2030.280 260.000 ;
        RECT 2030.080 244.810 2030.340 245.130 ;
        RECT 2173.600 244.810 2173.860 245.130 ;
        RECT 2173.660 3.050 2173.800 244.810 ;
        RECT 2173.600 2.730 2173.860 3.050 ;
        RECT 2179.120 2.730 2179.380 3.050 ;
        RECT 2179.180 2.400 2179.320 2.730 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2044.310 244.020 2044.630 244.080 ;
        RECT 2048.910 244.020 2049.230 244.080 ;
        RECT 2044.310 243.880 2049.230 244.020 ;
        RECT 2044.310 243.820 2044.630 243.880 ;
        RECT 2048.910 243.820 2049.230 243.880 ;
        RECT 2048.910 19.960 2049.230 20.020 ;
        RECT 2197.030 19.960 2197.350 20.020 ;
        RECT 2048.910 19.820 2197.350 19.960 ;
        RECT 2048.910 19.760 2049.230 19.820 ;
        RECT 2197.030 19.760 2197.350 19.820 ;
      LAYER via ;
        RECT 2044.340 243.820 2044.600 244.080 ;
        RECT 2048.940 243.820 2049.200 244.080 ;
        RECT 2048.940 19.760 2049.200 20.020 ;
        RECT 2197.060 19.760 2197.320 20.020 ;
      LAYER met2 ;
        RECT 2044.290 260.000 2044.570 264.000 ;
        RECT 2044.400 244.110 2044.540 260.000 ;
        RECT 2044.340 243.790 2044.600 244.110 ;
        RECT 2048.940 243.790 2049.200 244.110 ;
        RECT 2049.000 20.050 2049.140 243.790 ;
        RECT 2048.940 19.730 2049.200 20.050 ;
        RECT 2197.060 19.730 2197.320 20.050 ;
        RECT 2197.120 2.400 2197.260 19.730 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2058.110 244.020 2058.430 244.080 ;
        RECT 2062.710 244.020 2063.030 244.080 ;
        RECT 2058.110 243.880 2063.030 244.020 ;
        RECT 2058.110 243.820 2058.430 243.880 ;
        RECT 2062.710 243.820 2063.030 243.880 ;
        RECT 2062.710 19.620 2063.030 19.680 ;
        RECT 2214.970 19.620 2215.290 19.680 ;
        RECT 2062.710 19.480 2215.290 19.620 ;
        RECT 2062.710 19.420 2063.030 19.480 ;
        RECT 2214.970 19.420 2215.290 19.480 ;
      LAYER via ;
        RECT 2058.140 243.820 2058.400 244.080 ;
        RECT 2062.740 243.820 2063.000 244.080 ;
        RECT 2062.740 19.420 2063.000 19.680 ;
        RECT 2215.000 19.420 2215.260 19.680 ;
      LAYER met2 ;
        RECT 2058.090 260.000 2058.370 264.000 ;
        RECT 2058.200 244.110 2058.340 260.000 ;
        RECT 2058.140 243.790 2058.400 244.110 ;
        RECT 2062.740 243.790 2063.000 244.110 ;
        RECT 2062.800 19.710 2062.940 243.790 ;
        RECT 2062.740 19.390 2063.000 19.710 ;
        RECT 2215.000 19.390 2215.260 19.710 ;
        RECT 2215.060 2.400 2215.200 19.390 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2072.370 244.020 2072.690 244.080 ;
        RECT 2076.510 244.020 2076.830 244.080 ;
        RECT 2072.370 243.880 2076.830 244.020 ;
        RECT 2072.370 243.820 2072.690 243.880 ;
        RECT 2076.510 243.820 2076.830 243.880 ;
        RECT 2076.510 19.280 2076.830 19.340 ;
        RECT 2232.910 19.280 2233.230 19.340 ;
        RECT 2076.510 19.140 2233.230 19.280 ;
        RECT 2076.510 19.080 2076.830 19.140 ;
        RECT 2232.910 19.080 2233.230 19.140 ;
      LAYER via ;
        RECT 2072.400 243.820 2072.660 244.080 ;
        RECT 2076.540 243.820 2076.800 244.080 ;
        RECT 2076.540 19.080 2076.800 19.340 ;
        RECT 2232.940 19.080 2233.200 19.340 ;
      LAYER met2 ;
        RECT 2072.350 260.000 2072.630 264.000 ;
        RECT 2072.460 244.110 2072.600 260.000 ;
        RECT 2072.400 243.790 2072.660 244.110 ;
        RECT 2076.540 243.790 2076.800 244.110 ;
        RECT 2076.600 19.370 2076.740 243.790 ;
        RECT 2076.540 19.050 2076.800 19.370 ;
        RECT 2232.940 19.050 2233.200 19.370 ;
        RECT 2233.000 2.400 2233.140 19.050 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 245.380 793.430 245.440 ;
        RECT 931.570 245.380 931.890 245.440 ;
        RECT 793.110 245.240 931.890 245.380 ;
        RECT 793.110 245.180 793.430 245.240 ;
        RECT 931.570 245.180 931.890 245.240 ;
        RECT 787.590 17.240 787.910 17.300 ;
        RECT 793.110 17.240 793.430 17.300 ;
        RECT 787.590 17.100 793.430 17.240 ;
        RECT 787.590 17.040 787.910 17.100 ;
        RECT 793.110 17.040 793.430 17.100 ;
      LAYER via ;
        RECT 793.140 245.180 793.400 245.440 ;
        RECT 931.600 245.180 931.860 245.440 ;
        RECT 787.620 17.040 787.880 17.300 ;
        RECT 793.140 17.040 793.400 17.300 ;
      LAYER met2 ;
        RECT 931.550 260.000 931.830 264.000 ;
        RECT 931.660 245.470 931.800 260.000 ;
        RECT 793.140 245.150 793.400 245.470 ;
        RECT 931.600 245.150 931.860 245.470 ;
        RECT 793.200 17.330 793.340 245.150 ;
        RECT 787.620 17.010 787.880 17.330 ;
        RECT 793.140 17.010 793.400 17.330 ;
        RECT 787.680 2.400 787.820 17.010 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2086.630 242.320 2086.950 242.380 ;
        RECT 2090.310 242.320 2090.630 242.380 ;
        RECT 2086.630 242.180 2090.630 242.320 ;
        RECT 2086.630 242.120 2086.950 242.180 ;
        RECT 2090.310 242.120 2090.630 242.180 ;
        RECT 2090.310 18.600 2090.630 18.660 ;
        RECT 2250.850 18.600 2251.170 18.660 ;
        RECT 2090.310 18.460 2251.170 18.600 ;
        RECT 2090.310 18.400 2090.630 18.460 ;
        RECT 2250.850 18.400 2251.170 18.460 ;
      LAYER via ;
        RECT 2086.660 242.120 2086.920 242.380 ;
        RECT 2090.340 242.120 2090.600 242.380 ;
        RECT 2090.340 18.400 2090.600 18.660 ;
        RECT 2250.880 18.400 2251.140 18.660 ;
      LAYER met2 ;
        RECT 2086.610 260.000 2086.890 264.000 ;
        RECT 2086.720 242.410 2086.860 260.000 ;
        RECT 2086.660 242.090 2086.920 242.410 ;
        RECT 2090.340 242.090 2090.600 242.410 ;
        RECT 2090.400 18.690 2090.540 242.090 ;
        RECT 2090.340 18.370 2090.600 18.690 ;
        RECT 2250.880 18.370 2251.140 18.690 ;
        RECT 2250.940 2.400 2251.080 18.370 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2100.430 244.020 2100.750 244.080 ;
        RECT 2104.110 244.020 2104.430 244.080 ;
        RECT 2100.430 243.880 2104.430 244.020 ;
        RECT 2100.430 243.820 2100.750 243.880 ;
        RECT 2104.110 243.820 2104.430 243.880 ;
        RECT 2104.110 15.880 2104.430 15.940 ;
        RECT 2268.330 15.880 2268.650 15.940 ;
        RECT 2104.110 15.740 2268.650 15.880 ;
        RECT 2104.110 15.680 2104.430 15.740 ;
        RECT 2268.330 15.680 2268.650 15.740 ;
      LAYER via ;
        RECT 2100.460 243.820 2100.720 244.080 ;
        RECT 2104.140 243.820 2104.400 244.080 ;
        RECT 2104.140 15.680 2104.400 15.940 ;
        RECT 2268.360 15.680 2268.620 15.940 ;
      LAYER met2 ;
        RECT 2100.410 260.000 2100.690 264.000 ;
        RECT 2100.520 244.110 2100.660 260.000 ;
        RECT 2100.460 243.790 2100.720 244.110 ;
        RECT 2104.140 243.790 2104.400 244.110 ;
        RECT 2104.200 15.970 2104.340 243.790 ;
        RECT 2104.140 15.650 2104.400 15.970 ;
        RECT 2268.360 15.650 2268.620 15.970 ;
        RECT 2268.420 2.400 2268.560 15.650 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.910 18.940 2118.230 19.000 ;
        RECT 2286.270 18.940 2286.590 19.000 ;
        RECT 2117.910 18.800 2286.590 18.940 ;
        RECT 2117.910 18.740 2118.230 18.800 ;
        RECT 2286.270 18.740 2286.590 18.800 ;
      LAYER via ;
        RECT 2117.940 18.740 2118.200 19.000 ;
        RECT 2286.300 18.740 2286.560 19.000 ;
      LAYER met2 ;
        RECT 2114.670 260.170 2114.950 264.000 ;
        RECT 2114.670 260.030 2118.140 260.170 ;
        RECT 2114.670 260.000 2114.950 260.030 ;
        RECT 2118.000 19.030 2118.140 260.030 ;
        RECT 2117.940 18.710 2118.200 19.030 ;
        RECT 2286.300 18.710 2286.560 19.030 ;
        RECT 2286.360 2.400 2286.500 18.710 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 17.920 2132.030 17.980 ;
        RECT 2304.210 17.920 2304.530 17.980 ;
        RECT 2131.710 17.780 2304.530 17.920 ;
        RECT 2131.710 17.720 2132.030 17.780 ;
        RECT 2304.210 17.720 2304.530 17.780 ;
      LAYER via ;
        RECT 2131.740 17.720 2132.000 17.980 ;
        RECT 2304.240 17.720 2304.500 17.980 ;
      LAYER met2 ;
        RECT 2128.470 260.170 2128.750 264.000 ;
        RECT 2128.470 260.030 2131.940 260.170 ;
        RECT 2128.470 260.000 2128.750 260.030 ;
        RECT 2131.800 18.010 2131.940 260.030 ;
        RECT 2131.740 17.690 2132.000 18.010 ;
        RECT 2304.240 17.690 2304.500 18.010 ;
        RECT 2304.300 2.400 2304.440 17.690 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.510 16.220 2145.830 16.280 ;
        RECT 2322.150 16.220 2322.470 16.280 ;
        RECT 2145.510 16.080 2322.470 16.220 ;
        RECT 2145.510 16.020 2145.830 16.080 ;
        RECT 2322.150 16.020 2322.470 16.080 ;
      LAYER via ;
        RECT 2145.540 16.020 2145.800 16.280 ;
        RECT 2322.180 16.020 2322.440 16.280 ;
      LAYER met2 ;
        RECT 2142.730 260.170 2143.010 264.000 ;
        RECT 2142.730 260.030 2145.740 260.170 ;
        RECT 2142.730 260.000 2143.010 260.030 ;
        RECT 2145.600 16.310 2145.740 260.030 ;
        RECT 2145.540 15.990 2145.800 16.310 ;
        RECT 2322.180 15.990 2322.440 16.310 ;
        RECT 2322.240 2.400 2322.380 15.990 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2159.310 17.580 2159.630 17.640 ;
        RECT 2339.170 17.580 2339.490 17.640 ;
        RECT 2159.310 17.440 2339.490 17.580 ;
        RECT 2159.310 17.380 2159.630 17.440 ;
        RECT 2339.170 17.380 2339.490 17.440 ;
      LAYER via ;
        RECT 2159.340 17.380 2159.600 17.640 ;
        RECT 2339.200 17.380 2339.460 17.640 ;
      LAYER met2 ;
        RECT 2156.990 260.170 2157.270 264.000 ;
        RECT 2156.990 260.030 2159.540 260.170 ;
        RECT 2156.990 260.000 2157.270 260.030 ;
        RECT 2159.400 17.670 2159.540 260.030 ;
        RECT 2159.340 17.350 2159.600 17.670 ;
        RECT 2339.200 17.350 2339.460 17.670 ;
        RECT 2339.260 16.730 2339.400 17.350 ;
        RECT 2339.260 16.590 2339.860 16.730 ;
        RECT 2339.720 2.400 2339.860 16.590 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2173.110 18.260 2173.430 18.320 ;
        RECT 2357.570 18.260 2357.890 18.320 ;
        RECT 2173.110 18.120 2357.890 18.260 ;
        RECT 2173.110 18.060 2173.430 18.120 ;
        RECT 2357.570 18.060 2357.890 18.120 ;
      LAYER via ;
        RECT 2173.140 18.060 2173.400 18.320 ;
        RECT 2357.600 18.060 2357.860 18.320 ;
      LAYER met2 ;
        RECT 2170.790 260.170 2171.070 264.000 ;
        RECT 2170.790 260.030 2173.340 260.170 ;
        RECT 2170.790 260.000 2171.070 260.030 ;
        RECT 2173.200 18.350 2173.340 260.030 ;
        RECT 2173.140 18.030 2173.400 18.350 ;
        RECT 2357.600 18.030 2357.860 18.350 ;
        RECT 2357.660 2.400 2357.800 18.030 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 16.900 2187.230 16.960 ;
        RECT 2375.510 16.900 2375.830 16.960 ;
        RECT 2186.910 16.760 2375.830 16.900 ;
        RECT 2186.910 16.700 2187.230 16.760 ;
        RECT 2375.510 16.700 2375.830 16.760 ;
      LAYER via ;
        RECT 2186.940 16.700 2187.200 16.960 ;
        RECT 2375.540 16.700 2375.800 16.960 ;
      LAYER met2 ;
        RECT 2185.050 260.170 2185.330 264.000 ;
        RECT 2185.050 260.030 2187.140 260.170 ;
        RECT 2185.050 260.000 2185.330 260.030 ;
        RECT 2187.000 16.990 2187.140 260.030 ;
        RECT 2186.940 16.670 2187.200 16.990 ;
        RECT 2375.540 16.670 2375.800 16.990 ;
        RECT 2375.600 2.400 2375.740 16.670 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2200.250 20.300 2200.570 20.360 ;
        RECT 2393.450 20.300 2393.770 20.360 ;
        RECT 2200.250 20.160 2393.770 20.300 ;
        RECT 2200.250 20.100 2200.570 20.160 ;
        RECT 2393.450 20.100 2393.770 20.160 ;
      LAYER via ;
        RECT 2200.280 20.100 2200.540 20.360 ;
        RECT 2393.480 20.100 2393.740 20.360 ;
      LAYER met2 ;
        RECT 2199.310 260.170 2199.590 264.000 ;
        RECT 2199.310 260.030 2200.480 260.170 ;
        RECT 2199.310 260.000 2199.590 260.030 ;
        RECT 2200.340 20.390 2200.480 260.030 ;
        RECT 2200.280 20.070 2200.540 20.390 ;
        RECT 2393.480 20.070 2393.740 20.390 ;
        RECT 2393.540 2.400 2393.680 20.070 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2213.110 260.170 2213.390 264.000 ;
        RECT 2213.110 260.030 2214.740 260.170 ;
        RECT 2213.110 260.000 2213.390 260.030 ;
        RECT 2214.600 17.525 2214.740 260.030 ;
        RECT 2214.530 17.155 2214.810 17.525 ;
        RECT 2411.410 17.155 2411.690 17.525 ;
        RECT 2411.480 2.400 2411.620 17.155 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 2214.530 17.200 2214.810 17.480 ;
        RECT 2411.410 17.200 2411.690 17.480 ;
      LAYER met3 ;
        RECT 2214.505 17.490 2214.835 17.505 ;
        RECT 2411.385 17.490 2411.715 17.505 ;
        RECT 2214.505 17.190 2411.715 17.490 ;
        RECT 2214.505 17.175 2214.835 17.190 ;
        RECT 2411.385 17.175 2411.715 17.190 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 805.530 17.240 805.850 17.300 ;
        RECT 945.370 17.240 945.690 17.300 ;
        RECT 805.530 17.100 945.690 17.240 ;
        RECT 805.530 17.040 805.850 17.100 ;
        RECT 945.370 17.040 945.690 17.100 ;
      LAYER via ;
        RECT 805.560 17.040 805.820 17.300 ;
        RECT 945.400 17.040 945.660 17.300 ;
      LAYER met2 ;
        RECT 945.810 260.170 946.090 264.000 ;
        RECT 945.460 260.030 946.090 260.170 ;
        RECT 945.460 17.330 945.600 260.030 ;
        RECT 945.810 260.000 946.090 260.030 ;
        RECT 805.560 17.010 805.820 17.330 ;
        RECT 945.400 17.010 945.660 17.330 ;
        RECT 805.620 2.400 805.760 17.010 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 306.890 241.640 307.210 241.700 ;
        RECT 312.410 241.640 312.730 241.700 ;
        RECT 306.890 241.500 312.730 241.640 ;
        RECT 306.890 241.440 307.210 241.500 ;
        RECT 312.410 241.440 312.730 241.500 ;
        RECT 2.830 30.840 3.150 30.900 ;
        RECT 306.890 30.840 307.210 30.900 ;
        RECT 2.830 30.700 307.210 30.840 ;
        RECT 2.830 30.640 3.150 30.700 ;
        RECT 306.890 30.640 307.210 30.700 ;
      LAYER via ;
        RECT 306.920 241.440 307.180 241.700 ;
        RECT 312.440 241.440 312.700 241.700 ;
        RECT 2.860 30.640 3.120 30.900 ;
        RECT 306.920 30.640 307.180 30.900 ;
      LAYER met2 ;
        RECT 312.390 260.000 312.670 264.000 ;
        RECT 312.500 241.730 312.640 260.000 ;
        RECT 306.920 241.410 307.180 241.730 ;
        RECT 312.440 241.410 312.700 241.730 ;
        RECT 306.980 30.930 307.120 241.410 ;
        RECT 2.860 30.610 3.120 30.930 ;
        RECT 306.920 30.610 307.180 30.930 ;
        RECT 2.920 2.400 3.060 30.610 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 311.565 96.645 311.735 144.755 ;
      LAYER mcon ;
        RECT 311.565 144.585 311.735 144.755 ;
      LAYER met1 ;
        RECT 311.950 206.960 312.270 207.020 ;
        RECT 315.630 206.960 315.950 207.020 ;
        RECT 311.950 206.820 315.950 206.960 ;
        RECT 311.950 206.760 312.270 206.820 ;
        RECT 315.630 206.760 315.950 206.820 ;
        RECT 311.490 144.740 311.810 144.800 ;
        RECT 311.295 144.600 311.810 144.740 ;
        RECT 311.490 144.540 311.810 144.600 ;
        RECT 311.505 96.800 311.795 96.845 ;
        RECT 312.410 96.800 312.730 96.860 ;
        RECT 311.505 96.660 312.730 96.800 ;
        RECT 311.505 96.615 311.795 96.660 ;
        RECT 312.410 96.600 312.730 96.660 ;
        RECT 8.350 37.980 8.670 38.040 ;
        RECT 312.410 37.980 312.730 38.040 ;
        RECT 8.350 37.840 312.730 37.980 ;
        RECT 8.350 37.780 8.670 37.840 ;
        RECT 312.410 37.780 312.730 37.840 ;
      LAYER via ;
        RECT 311.980 206.760 312.240 207.020 ;
        RECT 315.660 206.760 315.920 207.020 ;
        RECT 311.520 144.540 311.780 144.800 ;
        RECT 312.440 96.600 312.700 96.860 ;
        RECT 8.380 37.780 8.640 38.040 ;
        RECT 312.440 37.780 312.700 38.040 ;
      LAYER met2 ;
        RECT 316.990 260.170 317.270 264.000 ;
        RECT 315.720 260.030 317.270 260.170 ;
        RECT 315.720 207.050 315.860 260.030 ;
        RECT 316.990 260.000 317.270 260.030 ;
        RECT 311.980 206.730 312.240 207.050 ;
        RECT 315.660 206.730 315.920 207.050 ;
        RECT 312.040 158.850 312.180 206.730 ;
        RECT 311.120 158.710 312.180 158.850 ;
        RECT 311.120 158.170 311.260 158.710 ;
        RECT 311.120 158.030 311.720 158.170 ;
        RECT 311.580 144.830 311.720 158.030 ;
        RECT 311.520 144.510 311.780 144.830 ;
        RECT 312.440 96.570 312.700 96.890 ;
        RECT 312.500 38.070 312.640 96.570 ;
        RECT 8.380 37.750 8.640 38.070 ;
        RECT 312.440 37.750 312.700 38.070 ;
        RECT 8.440 2.400 8.580 37.750 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 51.580 20.630 51.640 ;
        RECT 317.470 51.580 317.790 51.640 ;
        RECT 20.310 51.440 317.790 51.580 ;
        RECT 20.310 51.380 20.630 51.440 ;
        RECT 317.470 51.380 317.790 51.440 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 20.310 17.580 20.630 17.640 ;
        RECT 14.330 17.440 20.630 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 20.310 17.380 20.630 17.440 ;
      LAYER via ;
        RECT 20.340 51.380 20.600 51.640 ;
        RECT 317.500 51.380 317.760 51.640 ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 20.340 17.380 20.600 17.640 ;
      LAYER met2 ;
        RECT 321.590 260.170 321.870 264.000 ;
        RECT 317.560 260.030 321.870 260.170 ;
        RECT 317.560 51.670 317.700 260.030 ;
        RECT 321.590 260.000 321.870 260.030 ;
        RECT 20.340 51.350 20.600 51.670 ;
        RECT 317.500 51.350 317.760 51.670 ;
        RECT 20.400 17.670 20.540 51.350 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 20.340 17.350 20.600 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.150 58.720 45.470 58.780 ;
        RECT 338.170 58.720 338.490 58.780 ;
        RECT 45.150 58.580 338.490 58.720 ;
        RECT 45.150 58.520 45.470 58.580 ;
        RECT 338.170 58.520 338.490 58.580 ;
        RECT 38.250 17.580 38.570 17.640 ;
        RECT 45.150 17.580 45.470 17.640 ;
        RECT 38.250 17.440 45.470 17.580 ;
        RECT 38.250 17.380 38.570 17.440 ;
        RECT 45.150 17.380 45.470 17.440 ;
      LAYER via ;
        RECT 45.180 58.520 45.440 58.780 ;
        RECT 338.200 58.520 338.460 58.780 ;
        RECT 38.280 17.380 38.540 17.640 ;
        RECT 45.180 17.380 45.440 17.640 ;
      LAYER met2 ;
        RECT 340.450 260.170 340.730 264.000 ;
        RECT 338.260 260.030 340.730 260.170 ;
        RECT 338.260 58.810 338.400 260.030 ;
        RECT 340.450 260.000 340.730 260.030 ;
        RECT 45.180 58.490 45.440 58.810 ;
        RECT 338.200 58.490 338.460 58.810 ;
        RECT 45.240 17.670 45.380 58.490 ;
        RECT 38.280 17.350 38.540 17.670 ;
        RECT 45.180 17.350 45.440 17.670 ;
        RECT 38.340 2.400 38.480 17.350 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.650 24.720 240.970 24.780 ;
        RECT 496.870 24.720 497.190 24.780 ;
        RECT 240.650 24.580 497.190 24.720 ;
        RECT 240.650 24.520 240.970 24.580 ;
        RECT 496.870 24.520 497.190 24.580 ;
      LAYER via ;
        RECT 240.680 24.520 240.940 24.780 ;
        RECT 496.900 24.520 497.160 24.780 ;
      LAYER met2 ;
        RECT 500.070 260.170 500.350 264.000 ;
        RECT 496.960 260.030 500.350 260.170 ;
        RECT 496.960 24.810 497.100 260.030 ;
        RECT 500.070 260.000 500.350 260.030 ;
        RECT 240.680 24.490 240.940 24.810 ;
        RECT 496.900 24.490 497.160 24.810 ;
        RECT 240.740 2.400 240.880 24.490 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 25.060 258.450 25.120 ;
        RECT 510.670 25.060 510.990 25.120 ;
        RECT 258.130 24.920 510.990 25.060 ;
        RECT 258.130 24.860 258.450 24.920 ;
        RECT 510.670 24.860 510.990 24.920 ;
      LAYER via ;
        RECT 258.160 24.860 258.420 25.120 ;
        RECT 510.700 24.860 510.960 25.120 ;
      LAYER met2 ;
        RECT 513.870 260.170 514.150 264.000 ;
        RECT 510.760 260.030 514.150 260.170 ;
        RECT 510.760 25.150 510.900 260.030 ;
        RECT 513.870 260.000 514.150 260.030 ;
        RECT 258.160 24.830 258.420 25.150 ;
        RECT 510.700 24.830 510.960 25.150 ;
        RECT 258.220 2.400 258.360 24.830 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 25.740 276.390 25.800 ;
        RECT 524.470 25.740 524.790 25.800 ;
        RECT 276.070 25.600 524.790 25.740 ;
        RECT 276.070 25.540 276.390 25.600 ;
        RECT 524.470 25.540 524.790 25.600 ;
      LAYER via ;
        RECT 276.100 25.540 276.360 25.800 ;
        RECT 524.500 25.540 524.760 25.800 ;
      LAYER met2 ;
        RECT 528.130 260.170 528.410 264.000 ;
        RECT 524.560 260.030 528.410 260.170 ;
        RECT 524.560 25.830 524.700 260.030 ;
        RECT 528.130 260.000 528.410 260.030 ;
        RECT 276.100 25.510 276.360 25.830 ;
        RECT 524.500 25.510 524.760 25.830 ;
        RECT 276.160 2.400 276.300 25.510 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 25.400 294.330 25.460 ;
        RECT 538.270 25.400 538.590 25.460 ;
        RECT 294.010 25.260 538.590 25.400 ;
        RECT 294.010 25.200 294.330 25.260 ;
        RECT 538.270 25.200 538.590 25.260 ;
      LAYER via ;
        RECT 294.040 25.200 294.300 25.460 ;
        RECT 538.300 25.200 538.560 25.460 ;
      LAYER met2 ;
        RECT 542.390 260.170 542.670 264.000 ;
        RECT 538.360 260.030 542.670 260.170 ;
        RECT 538.360 25.490 538.500 260.030 ;
        RECT 542.390 260.000 542.670 260.030 ;
        RECT 294.040 25.170 294.300 25.490 ;
        RECT 538.300 25.170 538.560 25.490 ;
        RECT 294.100 2.400 294.240 25.170 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 30.840 312.270 30.900 ;
        RECT 552.070 30.840 552.390 30.900 ;
        RECT 311.950 30.700 552.390 30.840 ;
        RECT 311.950 30.640 312.270 30.700 ;
        RECT 552.070 30.640 552.390 30.700 ;
      LAYER via ;
        RECT 311.980 30.640 312.240 30.900 ;
        RECT 552.100 30.640 552.360 30.900 ;
      LAYER met2 ;
        RECT 556.190 260.170 556.470 264.000 ;
        RECT 552.160 260.030 556.470 260.170 ;
        RECT 552.160 30.930 552.300 260.030 ;
        RECT 556.190 260.000 556.470 260.030 ;
        RECT 311.980 30.610 312.240 30.930 ;
        RECT 552.100 30.610 552.360 30.930 ;
        RECT 312.040 2.400 312.180 30.610 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 37.980 330.210 38.040 ;
        RECT 566.330 37.980 566.650 38.040 ;
        RECT 329.890 37.840 566.650 37.980 ;
        RECT 329.890 37.780 330.210 37.840 ;
        RECT 566.330 37.780 566.650 37.840 ;
      LAYER via ;
        RECT 329.920 37.780 330.180 38.040 ;
        RECT 566.360 37.780 566.620 38.040 ;
      LAYER met2 ;
        RECT 570.450 260.170 570.730 264.000 ;
        RECT 566.420 260.030 570.730 260.170 ;
        RECT 566.420 38.070 566.560 260.030 ;
        RECT 570.450 260.000 570.730 260.030 ;
        RECT 329.920 37.750 330.180 38.070 ;
        RECT 566.360 37.750 566.620 38.070 ;
        RECT 329.980 2.400 330.120 37.750 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.510 237.900 351.830 237.960 ;
        RECT 584.270 237.900 584.590 237.960 ;
        RECT 351.510 237.760 584.590 237.900 ;
        RECT 351.510 237.700 351.830 237.760 ;
        RECT 584.270 237.700 584.590 237.760 ;
        RECT 347.370 17.580 347.690 17.640 ;
        RECT 351.510 17.580 351.830 17.640 ;
        RECT 347.370 17.440 351.830 17.580 ;
        RECT 347.370 17.380 347.690 17.440 ;
        RECT 351.510 17.380 351.830 17.440 ;
      LAYER via ;
        RECT 351.540 237.700 351.800 237.960 ;
        RECT 584.300 237.700 584.560 237.960 ;
        RECT 347.400 17.380 347.660 17.640 ;
        RECT 351.540 17.380 351.800 17.640 ;
      LAYER met2 ;
        RECT 584.250 260.000 584.530 264.000 ;
        RECT 584.360 237.990 584.500 260.000 ;
        RECT 351.540 237.670 351.800 237.990 ;
        RECT 584.300 237.670 584.560 237.990 ;
        RECT 351.600 17.670 351.740 237.670 ;
        RECT 347.400 17.350 347.660 17.670 ;
        RECT 351.540 17.350 351.800 17.670 ;
        RECT 347.460 2.400 347.600 17.350 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.930 231.440 594.250 231.500 ;
        RECT 597.150 231.440 597.470 231.500 ;
        RECT 593.930 231.300 597.470 231.440 ;
        RECT 593.930 231.240 594.250 231.300 ;
        RECT 597.150 231.240 597.470 231.300 ;
        RECT 365.310 24.040 365.630 24.100 ;
        RECT 593.930 24.040 594.250 24.100 ;
        RECT 365.310 23.900 594.250 24.040 ;
        RECT 365.310 23.840 365.630 23.900 ;
        RECT 593.930 23.840 594.250 23.900 ;
      LAYER via ;
        RECT 593.960 231.240 594.220 231.500 ;
        RECT 597.180 231.240 597.440 231.500 ;
        RECT 365.340 23.840 365.600 24.100 ;
        RECT 593.960 23.840 594.220 24.100 ;
      LAYER met2 ;
        RECT 598.510 260.170 598.790 264.000 ;
        RECT 597.240 260.030 598.790 260.170 ;
        RECT 597.240 231.530 597.380 260.030 ;
        RECT 598.510 260.000 598.790 260.030 ;
        RECT 593.960 231.210 594.220 231.530 ;
        RECT 597.180 231.210 597.440 231.530 ;
        RECT 594.020 24.130 594.160 231.210 ;
        RECT 365.340 23.810 365.600 24.130 ;
        RECT 593.960 23.810 594.220 24.130 ;
        RECT 365.400 2.400 365.540 23.810 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.590 241.640 603.910 241.700 ;
        RECT 612.790 241.640 613.110 241.700 ;
        RECT 603.590 241.500 613.110 241.640 ;
        RECT 603.590 241.440 603.910 241.500 ;
        RECT 612.790 241.440 613.110 241.500 ;
        RECT 383.250 44.780 383.570 44.840 ;
        RECT 603.590 44.780 603.910 44.840 ;
        RECT 383.250 44.640 603.910 44.780 ;
        RECT 383.250 44.580 383.570 44.640 ;
        RECT 603.590 44.580 603.910 44.640 ;
      LAYER via ;
        RECT 603.620 241.440 603.880 241.700 ;
        RECT 612.820 241.440 613.080 241.700 ;
        RECT 383.280 44.580 383.540 44.840 ;
        RECT 603.620 44.580 603.880 44.840 ;
      LAYER met2 ;
        RECT 612.770 260.000 613.050 264.000 ;
        RECT 612.880 241.730 613.020 260.000 ;
        RECT 603.620 241.410 603.880 241.730 ;
        RECT 612.820 241.410 613.080 241.730 ;
        RECT 603.680 44.870 603.820 241.410 ;
        RECT 383.280 44.550 383.540 44.870 ;
        RECT 603.620 44.550 603.880 44.870 ;
        RECT 383.340 2.400 383.480 44.550 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 621.605 144.925 621.775 193.035 ;
      LAYER mcon ;
        RECT 621.605 192.865 621.775 193.035 ;
      LAYER met1 ;
        RECT 621.070 206.960 621.390 207.020 ;
        RECT 621.990 206.960 622.310 207.020 ;
        RECT 621.070 206.820 622.310 206.960 ;
        RECT 621.070 206.760 621.390 206.820 ;
        RECT 621.990 206.760 622.310 206.820 ;
        RECT 621.545 193.020 621.835 193.065 ;
        RECT 621.990 193.020 622.310 193.080 ;
        RECT 621.545 192.880 622.310 193.020 ;
        RECT 621.545 192.835 621.835 192.880 ;
        RECT 621.990 192.820 622.310 192.880 ;
        RECT 621.530 145.080 621.850 145.140 ;
        RECT 621.335 144.940 621.850 145.080 ;
        RECT 621.530 144.880 621.850 144.940 ;
        RECT 621.530 110.540 621.850 110.800 ;
        RECT 621.620 110.120 621.760 110.540 ;
        RECT 621.530 109.860 621.850 110.120 ;
        RECT 401.190 51.580 401.510 51.640 ;
        RECT 621.990 51.580 622.310 51.640 ;
        RECT 401.190 51.440 622.310 51.580 ;
        RECT 401.190 51.380 401.510 51.440 ;
        RECT 621.990 51.380 622.310 51.440 ;
      LAYER via ;
        RECT 621.100 206.760 621.360 207.020 ;
        RECT 622.020 206.760 622.280 207.020 ;
        RECT 622.020 192.820 622.280 193.080 ;
        RECT 621.560 144.880 621.820 145.140 ;
        RECT 621.560 110.540 621.820 110.800 ;
        RECT 621.560 109.860 621.820 110.120 ;
        RECT 401.220 51.380 401.480 51.640 ;
        RECT 622.020 51.380 622.280 51.640 ;
      LAYER met2 ;
        RECT 626.570 260.170 626.850 264.000 ;
        RECT 624.380 260.030 626.850 260.170 ;
        RECT 624.380 230.250 624.520 260.030 ;
        RECT 626.570 260.000 626.850 260.030 ;
        RECT 621.160 230.110 624.520 230.250 ;
        RECT 621.160 207.050 621.300 230.110 ;
        RECT 621.100 206.730 621.360 207.050 ;
        RECT 622.020 206.730 622.280 207.050 ;
        RECT 622.080 193.110 622.220 206.730 ;
        RECT 622.020 192.790 622.280 193.110 ;
        RECT 621.560 144.850 621.820 145.170 ;
        RECT 621.620 110.830 621.760 144.850 ;
        RECT 621.560 110.510 621.820 110.830 ;
        RECT 621.560 109.830 621.820 110.150 ;
        RECT 621.620 62.290 621.760 109.830 ;
        RECT 621.620 62.150 622.220 62.290 ;
        RECT 622.080 51.670 622.220 62.150 ;
        RECT 401.220 51.350 401.480 51.670 ;
        RECT 622.020 51.350 622.280 51.670 ;
        RECT 401.280 2.400 401.420 51.350 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 24.040 62.490 24.100 ;
        RECT 358.870 24.040 359.190 24.100 ;
        RECT 62.170 23.900 359.190 24.040 ;
        RECT 62.170 23.840 62.490 23.900 ;
        RECT 358.870 23.840 359.190 23.900 ;
      LAYER via ;
        RECT 62.200 23.840 62.460 24.100 ;
        RECT 358.900 23.840 359.160 24.100 ;
      LAYER met2 ;
        RECT 359.310 260.170 359.590 264.000 ;
        RECT 358.960 260.030 359.590 260.170 ;
        RECT 358.960 24.130 359.100 260.030 ;
        RECT 359.310 260.000 359.590 260.030 ;
        RECT 62.200 23.810 62.460 24.130 ;
        RECT 358.900 23.810 359.160 24.130 ;
        RECT 62.260 2.400 62.400 23.810 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 631.190 241.640 631.510 241.700 ;
        RECT 640.850 241.640 641.170 241.700 ;
        RECT 631.190 241.500 641.170 241.640 ;
        RECT 631.190 241.440 631.510 241.500 ;
        RECT 640.850 241.440 641.170 241.500 ;
        RECT 420.510 58.720 420.830 58.780 ;
        RECT 631.190 58.720 631.510 58.780 ;
        RECT 420.510 58.580 631.510 58.720 ;
        RECT 420.510 58.520 420.830 58.580 ;
        RECT 631.190 58.520 631.510 58.580 ;
        RECT 419.130 2.960 419.450 3.020 ;
        RECT 420.510 2.960 420.830 3.020 ;
        RECT 419.130 2.820 420.830 2.960 ;
        RECT 419.130 2.760 419.450 2.820 ;
        RECT 420.510 2.760 420.830 2.820 ;
      LAYER via ;
        RECT 631.220 241.440 631.480 241.700 ;
        RECT 640.880 241.440 641.140 241.700 ;
        RECT 420.540 58.520 420.800 58.780 ;
        RECT 631.220 58.520 631.480 58.780 ;
        RECT 419.160 2.760 419.420 3.020 ;
        RECT 420.540 2.760 420.800 3.020 ;
      LAYER met2 ;
        RECT 640.830 260.000 641.110 264.000 ;
        RECT 640.940 241.730 641.080 260.000 ;
        RECT 631.220 241.410 631.480 241.730 ;
        RECT 640.880 241.410 641.140 241.730 ;
        RECT 631.280 58.810 631.420 241.410 ;
        RECT 420.540 58.490 420.800 58.810 ;
        RECT 631.220 58.490 631.480 58.810 ;
        RECT 420.600 3.050 420.740 58.490 ;
        RECT 419.160 2.730 419.420 3.050 ;
        RECT 420.540 2.730 420.800 3.050 ;
        RECT 419.220 2.400 419.360 2.730 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 231.100 441.530 231.160 ;
        RECT 654.650 231.100 654.970 231.160 ;
        RECT 441.210 230.960 654.970 231.100 ;
        RECT 441.210 230.900 441.530 230.960 ;
        RECT 654.650 230.900 654.970 230.960 ;
        RECT 436.610 14.520 436.930 14.580 ;
        RECT 441.210 14.520 441.530 14.580 ;
        RECT 436.610 14.380 441.530 14.520 ;
        RECT 436.610 14.320 436.930 14.380 ;
        RECT 441.210 14.320 441.530 14.380 ;
      LAYER via ;
        RECT 441.240 230.900 441.500 231.160 ;
        RECT 654.680 230.900 654.940 231.160 ;
        RECT 436.640 14.320 436.900 14.580 ;
        RECT 441.240 14.320 441.500 14.580 ;
      LAYER met2 ;
        RECT 654.630 260.000 654.910 264.000 ;
        RECT 654.740 231.190 654.880 260.000 ;
        RECT 441.240 230.870 441.500 231.190 ;
        RECT 654.680 230.870 654.940 231.190 ;
        RECT 441.300 14.610 441.440 230.870 ;
        RECT 436.640 14.290 436.900 14.610 ;
        RECT 441.240 14.290 441.500 14.610 ;
        RECT 436.700 2.400 436.840 14.290 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 664.310 193.360 664.630 193.420 ;
        RECT 667.070 193.360 667.390 193.420 ;
        RECT 664.310 193.220 667.390 193.360 ;
        RECT 664.310 193.160 664.630 193.220 ;
        RECT 667.070 193.160 667.390 193.220 ;
        RECT 455.010 113.800 455.330 113.860 ;
        RECT 664.310 113.800 664.630 113.860 ;
        RECT 455.010 113.660 664.630 113.800 ;
        RECT 455.010 113.600 455.330 113.660 ;
        RECT 664.310 113.600 664.630 113.660 ;
      LAYER via ;
        RECT 664.340 193.160 664.600 193.420 ;
        RECT 667.100 193.160 667.360 193.420 ;
        RECT 455.040 113.600 455.300 113.860 ;
        RECT 664.340 113.600 664.600 113.860 ;
      LAYER met2 ;
        RECT 668.890 260.170 669.170 264.000 ;
        RECT 667.160 260.030 669.170 260.170 ;
        RECT 667.160 193.450 667.300 260.030 ;
        RECT 668.890 260.000 669.170 260.030 ;
        RECT 664.340 193.130 664.600 193.450 ;
        RECT 667.100 193.130 667.360 193.450 ;
        RECT 664.400 113.890 664.540 193.130 ;
        RECT 455.040 113.570 455.300 113.890 ;
        RECT 664.340 113.570 664.600 113.890 ;
        RECT 455.100 2.960 455.240 113.570 ;
        RECT 454.640 2.820 455.240 2.960 ;
        RECT 454.640 2.400 454.780 2.820 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.710 65.520 476.030 65.580 ;
        RECT 683.170 65.520 683.490 65.580 ;
        RECT 475.710 65.380 683.490 65.520 ;
        RECT 475.710 65.320 476.030 65.380 ;
        RECT 683.170 65.320 683.490 65.380 ;
        RECT 472.490 14.520 472.810 14.580 ;
        RECT 475.710 14.520 476.030 14.580 ;
        RECT 472.490 14.380 476.030 14.520 ;
        RECT 472.490 14.320 472.810 14.380 ;
        RECT 475.710 14.320 476.030 14.380 ;
      LAYER via ;
        RECT 475.740 65.320 476.000 65.580 ;
        RECT 683.200 65.320 683.460 65.580 ;
        RECT 472.520 14.320 472.780 14.580 ;
        RECT 475.740 14.320 476.000 14.580 ;
      LAYER met2 ;
        RECT 683.150 260.000 683.430 264.000 ;
        RECT 683.260 65.610 683.400 260.000 ;
        RECT 475.740 65.290 476.000 65.610 ;
        RECT 683.200 65.290 683.460 65.610 ;
        RECT 475.800 14.610 475.940 65.290 ;
        RECT 472.520 14.290 472.780 14.610 ;
        RECT 475.740 14.290 476.000 14.610 ;
        RECT 472.580 2.400 472.720 14.290 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 72.320 496.730 72.380 ;
        RECT 697.430 72.320 697.750 72.380 ;
        RECT 496.410 72.180 697.750 72.320 ;
        RECT 496.410 72.120 496.730 72.180 ;
        RECT 697.430 72.120 697.750 72.180 ;
        RECT 490.430 16.900 490.750 16.960 ;
        RECT 496.410 16.900 496.730 16.960 ;
        RECT 490.430 16.760 496.730 16.900 ;
        RECT 490.430 16.700 490.750 16.760 ;
        RECT 496.410 16.700 496.730 16.760 ;
      LAYER via ;
        RECT 496.440 72.120 496.700 72.380 ;
        RECT 697.460 72.120 697.720 72.380 ;
        RECT 490.460 16.700 490.720 16.960 ;
        RECT 496.440 16.700 496.700 16.960 ;
      LAYER met2 ;
        RECT 696.950 260.170 697.230 264.000 ;
        RECT 696.950 260.030 697.660 260.170 ;
        RECT 696.950 260.000 697.230 260.030 ;
        RECT 697.520 72.410 697.660 260.030 ;
        RECT 496.440 72.090 496.700 72.410 ;
        RECT 697.460 72.090 697.720 72.410 ;
        RECT 496.500 16.990 496.640 72.090 ;
        RECT 490.460 16.670 490.720 16.990 ;
        RECT 496.440 16.670 496.700 16.990 ;
        RECT 490.520 2.400 490.660 16.670 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 79.460 510.530 79.520 ;
        RECT 711.230 79.460 711.550 79.520 ;
        RECT 510.210 79.320 711.550 79.460 ;
        RECT 510.210 79.260 510.530 79.320 ;
        RECT 711.230 79.260 711.550 79.320 ;
        RECT 507.910 16.900 508.230 16.960 ;
        RECT 510.210 16.900 510.530 16.960 ;
        RECT 507.910 16.760 510.530 16.900 ;
        RECT 507.910 16.700 508.230 16.760 ;
        RECT 510.210 16.700 510.530 16.760 ;
      LAYER via ;
        RECT 510.240 79.260 510.500 79.520 ;
        RECT 711.260 79.260 711.520 79.520 ;
        RECT 507.940 16.700 508.200 16.960 ;
        RECT 510.240 16.700 510.500 16.960 ;
      LAYER met2 ;
        RECT 711.210 260.000 711.490 264.000 ;
        RECT 711.320 79.550 711.460 260.000 ;
        RECT 510.240 79.230 510.500 79.550 ;
        RECT 711.260 79.230 711.520 79.550 ;
        RECT 510.300 16.990 510.440 79.230 ;
        RECT 507.940 16.670 508.200 16.990 ;
        RECT 510.240 16.670 510.500 16.990 ;
        RECT 508.000 2.400 508.140 16.670 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.910 210.360 531.230 210.420 ;
        RECT 725.030 210.360 725.350 210.420 ;
        RECT 530.910 210.220 725.350 210.360 ;
        RECT 530.910 210.160 531.230 210.220 ;
        RECT 725.030 210.160 725.350 210.220 ;
        RECT 525.850 16.900 526.170 16.960 ;
        RECT 530.910 16.900 531.230 16.960 ;
        RECT 525.850 16.760 531.230 16.900 ;
        RECT 525.850 16.700 526.170 16.760 ;
        RECT 530.910 16.700 531.230 16.760 ;
      LAYER via ;
        RECT 530.940 210.160 531.200 210.420 ;
        RECT 725.060 210.160 725.320 210.420 ;
        RECT 525.880 16.700 526.140 16.960 ;
        RECT 530.940 16.700 531.200 16.960 ;
      LAYER met2 ;
        RECT 725.010 260.000 725.290 264.000 ;
        RECT 725.120 210.450 725.260 260.000 ;
        RECT 530.940 210.130 531.200 210.450 ;
        RECT 725.060 210.130 725.320 210.450 ;
        RECT 531.000 16.990 531.140 210.130 ;
        RECT 525.880 16.670 526.140 16.990 ;
        RECT 530.940 16.670 531.200 16.990 ;
        RECT 525.940 2.400 526.080 16.670 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 734.690 244.020 735.010 244.080 ;
        RECT 739.290 244.020 739.610 244.080 ;
        RECT 734.690 243.880 739.610 244.020 ;
        RECT 734.690 243.820 735.010 243.880 ;
        RECT 739.290 243.820 739.610 243.880 ;
        RECT 544.710 107.000 545.030 107.060 ;
        RECT 734.690 107.000 735.010 107.060 ;
        RECT 544.710 106.860 735.010 107.000 ;
        RECT 544.710 106.800 545.030 106.860 ;
        RECT 734.690 106.800 735.010 106.860 ;
      LAYER via ;
        RECT 734.720 243.820 734.980 244.080 ;
        RECT 739.320 243.820 739.580 244.080 ;
        RECT 544.740 106.800 545.000 107.060 ;
        RECT 734.720 106.800 734.980 107.060 ;
      LAYER met2 ;
        RECT 739.270 260.000 739.550 264.000 ;
        RECT 739.380 244.110 739.520 260.000 ;
        RECT 734.720 243.790 734.980 244.110 ;
        RECT 739.320 243.790 739.580 244.110 ;
        RECT 734.780 107.090 734.920 243.790 ;
        RECT 544.740 106.770 545.000 107.090 ;
        RECT 734.720 106.770 734.980 107.090 ;
        RECT 544.800 3.130 544.940 106.770 ;
        RECT 543.880 2.990 544.940 3.130 ;
        RECT 543.880 2.400 544.020 2.990 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 30.840 562.050 30.900 ;
        RECT 752.630 30.840 752.950 30.900 ;
        RECT 561.730 30.700 752.950 30.840 ;
        RECT 561.730 30.640 562.050 30.700 ;
        RECT 752.630 30.640 752.950 30.700 ;
      LAYER via ;
        RECT 561.760 30.640 562.020 30.900 ;
        RECT 752.660 30.640 752.920 30.900 ;
      LAYER met2 ;
        RECT 753.530 260.170 753.810 264.000 ;
        RECT 752.720 260.030 753.810 260.170 ;
        RECT 752.720 30.930 752.860 260.030 ;
        RECT 753.530 260.000 753.810 260.030 ;
        RECT 561.760 30.610 562.020 30.930 ;
        RECT 752.660 30.610 752.920 30.930 ;
        RECT 561.820 2.400 561.960 30.610 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 37.980 579.990 38.040 ;
        RECT 766.430 37.980 766.750 38.040 ;
        RECT 579.670 37.840 766.750 37.980 ;
        RECT 579.670 37.780 579.990 37.840 ;
        RECT 766.430 37.780 766.750 37.840 ;
      LAYER via ;
        RECT 579.700 37.780 579.960 38.040 ;
        RECT 766.460 37.780 766.720 38.040 ;
      LAYER met2 ;
        RECT 767.330 260.170 767.610 264.000 ;
        RECT 766.520 260.030 767.610 260.170 ;
        RECT 766.520 38.070 766.660 260.030 ;
        RECT 767.330 260.000 767.610 260.030 ;
        RECT 579.700 37.750 579.960 38.070 ;
        RECT 766.460 37.750 766.720 38.070 ;
        RECT 579.760 2.400 579.900 37.750 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 373.665 96.645 373.835 111.775 ;
      LAYER mcon ;
        RECT 373.665 111.605 373.835 111.775 ;
      LAYER met1 ;
        RECT 373.590 193.360 373.910 193.420 ;
        RECT 374.510 193.360 374.830 193.420 ;
        RECT 373.590 193.220 374.830 193.360 ;
        RECT 373.590 193.160 373.910 193.220 ;
        RECT 374.510 193.160 374.830 193.220 ;
        RECT 373.590 111.760 373.910 111.820 ;
        RECT 373.395 111.620 373.910 111.760 ;
        RECT 373.590 111.560 373.910 111.620 ;
        RECT 373.590 96.800 373.910 96.860 ;
        RECT 373.395 96.660 373.910 96.800 ;
        RECT 373.590 96.600 373.910 96.660 ;
        RECT 86.550 24.380 86.870 24.440 ;
        RECT 373.590 24.380 373.910 24.440 ;
        RECT 86.550 24.240 373.910 24.380 ;
        RECT 86.550 24.180 86.870 24.240 ;
        RECT 373.590 24.180 373.910 24.240 ;
      LAYER via ;
        RECT 373.620 193.160 373.880 193.420 ;
        RECT 374.540 193.160 374.800 193.420 ;
        RECT 373.620 111.560 373.880 111.820 ;
        RECT 373.620 96.600 373.880 96.860 ;
        RECT 86.580 24.180 86.840 24.440 ;
        RECT 373.620 24.180 373.880 24.440 ;
      LAYER met2 ;
        RECT 377.710 260.850 377.990 264.000 ;
        RECT 375.060 260.710 377.990 260.850 ;
        RECT 375.060 256.090 375.200 260.710 ;
        RECT 377.710 260.000 377.990 260.710 ;
        RECT 374.600 255.950 375.200 256.090 ;
        RECT 374.600 193.450 374.740 255.950 ;
        RECT 373.620 193.130 373.880 193.450 ;
        RECT 374.540 193.130 374.800 193.450 ;
        RECT 373.680 111.850 373.820 193.130 ;
        RECT 373.620 111.530 373.880 111.850 ;
        RECT 373.620 96.570 373.880 96.890 ;
        RECT 373.680 24.470 373.820 96.570 ;
        RECT 86.580 24.150 86.840 24.470 ;
        RECT 373.620 24.150 373.880 24.470 ;
        RECT 86.640 12.650 86.780 24.150 ;
        RECT 86.180 12.510 86.780 12.650 ;
        RECT 86.180 2.400 86.320 12.510 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 45.120 597.470 45.180 ;
        RECT 780.230 45.120 780.550 45.180 ;
        RECT 597.150 44.980 780.550 45.120 ;
        RECT 597.150 44.920 597.470 44.980 ;
        RECT 780.230 44.920 780.550 44.980 ;
      LAYER via ;
        RECT 597.180 44.920 597.440 45.180 ;
        RECT 780.260 44.920 780.520 45.180 ;
      LAYER met2 ;
        RECT 781.590 260.170 781.870 264.000 ;
        RECT 780.320 260.030 781.870 260.170 ;
        RECT 780.320 45.210 780.460 260.030 ;
        RECT 781.590 260.000 781.870 260.030 ;
        RECT 597.180 44.890 597.440 45.210 ;
        RECT 780.260 44.890 780.520 45.210 ;
        RECT 597.240 2.400 597.380 44.890 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 134.540 620.930 134.600 ;
        RECT 793.570 134.540 793.890 134.600 ;
        RECT 620.610 134.400 793.890 134.540 ;
        RECT 620.610 134.340 620.930 134.400 ;
        RECT 793.570 134.340 793.890 134.400 ;
        RECT 615.090 17.920 615.410 17.980 ;
        RECT 620.610 17.920 620.930 17.980 ;
        RECT 615.090 17.780 620.930 17.920 ;
        RECT 615.090 17.720 615.410 17.780 ;
        RECT 620.610 17.720 620.930 17.780 ;
      LAYER via ;
        RECT 620.640 134.340 620.900 134.600 ;
        RECT 793.600 134.340 793.860 134.600 ;
        RECT 615.120 17.720 615.380 17.980 ;
        RECT 620.640 17.720 620.900 17.980 ;
      LAYER met2 ;
        RECT 795.850 260.170 796.130 264.000 ;
        RECT 793.660 260.030 796.130 260.170 ;
        RECT 793.660 134.630 793.800 260.030 ;
        RECT 795.850 260.000 796.130 260.030 ;
        RECT 620.640 134.310 620.900 134.630 ;
        RECT 793.600 134.310 793.860 134.630 ;
        RECT 620.700 18.010 620.840 134.310 ;
        RECT 615.120 17.690 615.380 18.010 ;
        RECT 620.640 17.690 620.900 18.010 ;
        RECT 615.180 2.400 615.320 17.690 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 231.100 110.330 231.160 ;
        RECT 110.010 230.960 370.140 231.100 ;
        RECT 110.010 230.900 110.330 230.960 ;
        RECT 370.000 230.760 370.140 230.960 ;
        RECT 394.750 230.760 395.070 230.820 ;
        RECT 370.000 230.620 395.070 230.760 ;
        RECT 394.750 230.560 395.070 230.620 ;
      LAYER via ;
        RECT 110.040 230.900 110.300 231.160 ;
        RECT 394.780 230.560 395.040 230.820 ;
      LAYER met2 ;
        RECT 396.570 260.170 396.850 264.000 ;
        RECT 394.840 260.030 396.850 260.170 ;
        RECT 110.040 230.870 110.300 231.190 ;
        RECT 110.100 17.410 110.240 230.870 ;
        RECT 394.840 230.850 394.980 260.030 ;
        RECT 396.570 260.000 396.850 260.030 ;
        RECT 394.780 230.530 395.040 230.850 ;
        RECT 109.640 17.270 110.240 17.410 ;
        RECT 109.640 2.400 109.780 17.270 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 137.610 224.300 137.930 224.360 ;
        RECT 414.530 224.300 414.850 224.360 ;
        RECT 137.610 224.160 414.850 224.300 ;
        RECT 137.610 224.100 137.930 224.160 ;
        RECT 414.530 224.100 414.850 224.160 ;
        RECT 133.470 16.900 133.790 16.960 ;
        RECT 137.610 16.900 137.930 16.960 ;
        RECT 133.470 16.760 137.930 16.900 ;
        RECT 133.470 16.700 133.790 16.760 ;
        RECT 137.610 16.700 137.930 16.760 ;
      LAYER via ;
        RECT 137.640 224.100 137.900 224.360 ;
        RECT 414.560 224.100 414.820 224.360 ;
        RECT 133.500 16.700 133.760 16.960 ;
        RECT 137.640 16.700 137.900 16.960 ;
      LAYER met2 ;
        RECT 415.430 260.170 415.710 264.000 ;
        RECT 414.620 260.030 415.710 260.170 ;
        RECT 414.620 224.390 414.760 260.030 ;
        RECT 415.430 260.000 415.710 260.030 ;
        RECT 137.640 224.070 137.900 224.390 ;
        RECT 414.560 224.070 414.820 224.390 ;
        RECT 137.700 16.990 137.840 224.070 ;
        RECT 133.500 16.670 133.760 16.990 ;
        RECT 137.640 16.670 137.900 16.990 ;
        RECT 133.560 2.400 133.700 16.670 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 65.520 151.730 65.580 ;
        RECT 427.870 65.520 428.190 65.580 ;
        RECT 151.410 65.380 428.190 65.520 ;
        RECT 151.410 65.320 151.730 65.380 ;
        RECT 427.870 65.320 428.190 65.380 ;
      LAYER via ;
        RECT 151.440 65.320 151.700 65.580 ;
        RECT 427.900 65.320 428.160 65.580 ;
      LAYER met2 ;
        RECT 429.690 260.170 429.970 264.000 ;
        RECT 427.960 260.030 429.970 260.170 ;
        RECT 427.960 65.610 428.100 260.030 ;
        RECT 429.690 260.000 429.970 260.030 ;
        RECT 151.440 65.290 151.700 65.610 ;
        RECT 427.900 65.290 428.160 65.610 ;
        RECT 151.500 2.400 151.640 65.290 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 217.160 172.430 217.220 ;
        RECT 442.130 217.160 442.450 217.220 ;
        RECT 172.110 217.020 442.450 217.160 ;
        RECT 172.110 216.960 172.430 217.020 ;
        RECT 442.130 216.960 442.450 217.020 ;
        RECT 169.350 16.900 169.670 16.960 ;
        RECT 172.110 16.900 172.430 16.960 ;
        RECT 169.350 16.760 172.430 16.900 ;
        RECT 169.350 16.700 169.670 16.760 ;
        RECT 172.110 16.700 172.430 16.760 ;
      LAYER via ;
        RECT 172.140 216.960 172.400 217.220 ;
        RECT 442.160 216.960 442.420 217.220 ;
        RECT 169.380 16.700 169.640 16.960 ;
        RECT 172.140 16.700 172.400 16.960 ;
      LAYER met2 ;
        RECT 443.490 260.170 443.770 264.000 ;
        RECT 442.220 260.030 443.770 260.170 ;
        RECT 442.220 217.250 442.360 260.030 ;
        RECT 443.490 260.000 443.770 260.030 ;
        RECT 172.140 216.930 172.400 217.250 ;
        RECT 442.160 216.930 442.420 217.250 ;
        RECT 172.200 16.990 172.340 216.930 ;
        RECT 169.380 16.670 169.640 16.990 ;
        RECT 172.140 16.670 172.400 16.990 ;
        RECT 169.440 2.400 169.580 16.670 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 72.320 192.670 72.380 ;
        RECT 455.470 72.320 455.790 72.380 ;
        RECT 192.350 72.180 455.790 72.320 ;
        RECT 192.350 72.120 192.670 72.180 ;
        RECT 455.470 72.120 455.790 72.180 ;
        RECT 186.830 16.900 187.150 16.960 ;
        RECT 192.350 16.900 192.670 16.960 ;
        RECT 186.830 16.760 192.670 16.900 ;
        RECT 186.830 16.700 187.150 16.760 ;
        RECT 192.350 16.700 192.670 16.760 ;
      LAYER via ;
        RECT 192.380 72.120 192.640 72.380 ;
        RECT 455.500 72.120 455.760 72.380 ;
        RECT 186.860 16.700 187.120 16.960 ;
        RECT 192.380 16.700 192.640 16.960 ;
      LAYER met2 ;
        RECT 457.750 260.170 458.030 264.000 ;
        RECT 455.560 260.030 458.030 260.170 ;
        RECT 455.560 72.410 455.700 260.030 ;
        RECT 457.750 260.000 458.030 260.030 ;
        RECT 192.380 72.090 192.640 72.410 ;
        RECT 455.500 72.090 455.760 72.410 ;
        RECT 192.440 16.990 192.580 72.090 ;
        RECT 186.860 16.670 187.120 16.990 ;
        RECT 192.380 16.670 192.640 16.990 ;
        RECT 186.920 2.400 187.060 16.670 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 206.610 79.460 206.930 79.520 ;
        RECT 469.270 79.460 469.590 79.520 ;
        RECT 206.610 79.320 469.590 79.460 ;
        RECT 206.610 79.260 206.930 79.320 ;
        RECT 469.270 79.260 469.590 79.320 ;
      LAYER via ;
        RECT 206.640 79.260 206.900 79.520 ;
        RECT 469.300 79.260 469.560 79.520 ;
      LAYER met2 ;
        RECT 471.550 260.170 471.830 264.000 ;
        RECT 469.360 260.030 471.830 260.170 ;
        RECT 469.360 79.550 469.500 260.030 ;
        RECT 471.550 260.000 471.830 260.030 ;
        RECT 206.640 79.230 206.900 79.550 ;
        RECT 469.300 79.230 469.560 79.550 ;
        RECT 206.700 17.410 206.840 79.230 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 86.260 227.630 86.320 ;
        RECT 483.070 86.260 483.390 86.320 ;
        RECT 227.310 86.120 483.390 86.260 ;
        RECT 227.310 86.060 227.630 86.120 ;
        RECT 483.070 86.060 483.390 86.120 ;
        RECT 222.710 16.560 223.030 16.620 ;
        RECT 227.310 16.560 227.630 16.620 ;
        RECT 222.710 16.420 227.630 16.560 ;
        RECT 222.710 16.360 223.030 16.420 ;
        RECT 227.310 16.360 227.630 16.420 ;
      LAYER via ;
        RECT 227.340 86.060 227.600 86.320 ;
        RECT 483.100 86.060 483.360 86.320 ;
        RECT 222.740 16.360 223.000 16.620 ;
        RECT 227.340 16.360 227.600 16.620 ;
      LAYER met2 ;
        RECT 485.810 260.170 486.090 264.000 ;
        RECT 483.160 260.030 486.090 260.170 ;
        RECT 483.160 86.350 483.300 260.030 ;
        RECT 485.810 260.000 486.090 260.030 ;
        RECT 227.340 86.030 227.600 86.350 ;
        RECT 483.100 86.030 483.360 86.350 ;
        RECT 227.400 16.650 227.540 86.030 ;
        RECT 222.740 16.330 223.000 16.650 ;
        RECT 227.340 16.330 227.600 16.650 ;
        RECT 222.800 2.400 222.940 16.330 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.590 237.900 51.910 237.960 ;
        RECT 326.210 237.900 326.530 237.960 ;
        RECT 51.590 237.760 326.530 237.900 ;
        RECT 51.590 237.700 51.910 237.760 ;
        RECT 326.210 237.700 326.530 237.760 ;
        RECT 51.590 18.260 51.910 18.320 ;
        RECT 37.880 18.120 51.910 18.260 ;
        RECT 37.880 17.580 38.020 18.120 ;
        RECT 51.590 18.060 51.910 18.120 ;
        RECT 20.860 17.440 38.020 17.580 ;
        RECT 20.310 16.900 20.630 16.960 ;
        RECT 20.860 16.900 21.000 17.440 ;
        RECT 20.310 16.760 21.000 16.900 ;
        RECT 20.310 16.700 20.630 16.760 ;
      LAYER via ;
        RECT 51.620 237.700 51.880 237.960 ;
        RECT 326.240 237.700 326.500 237.960 ;
        RECT 51.620 18.060 51.880 18.320 ;
        RECT 20.340 16.700 20.600 16.960 ;
      LAYER met2 ;
        RECT 326.190 260.000 326.470 264.000 ;
        RECT 326.300 237.990 326.440 260.000 ;
        RECT 51.620 237.670 51.880 237.990 ;
        RECT 326.240 237.670 326.500 237.990 ;
        RECT 51.680 18.350 51.820 237.670 ;
        RECT 51.620 18.030 51.880 18.350 ;
        RECT 20.340 16.670 20.600 16.990 ;
        RECT 20.400 2.400 20.540 16.670 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 52.050 93.060 52.370 93.120 ;
        RECT 345.530 93.060 345.850 93.120 ;
        RECT 52.050 92.920 345.850 93.060 ;
        RECT 52.050 92.860 52.370 92.920 ;
        RECT 345.530 92.860 345.850 92.920 ;
        RECT 44.230 14.860 44.550 14.920 ;
        RECT 52.050 14.860 52.370 14.920 ;
        RECT 44.230 14.720 52.370 14.860 ;
        RECT 44.230 14.660 44.550 14.720 ;
        RECT 52.050 14.660 52.370 14.720 ;
      LAYER via ;
        RECT 52.080 92.860 52.340 93.120 ;
        RECT 345.560 92.860 345.820 93.120 ;
        RECT 44.260 14.660 44.520 14.920 ;
        RECT 52.080 14.660 52.340 14.920 ;
      LAYER met2 ;
        RECT 345.050 260.170 345.330 264.000 ;
        RECT 345.050 260.030 345.760 260.170 ;
        RECT 345.050 260.000 345.330 260.030 ;
        RECT 345.620 93.150 345.760 260.030 ;
        RECT 52.080 92.830 52.340 93.150 ;
        RECT 345.560 92.830 345.820 93.150 ;
        RECT 52.140 14.950 52.280 92.830 ;
        RECT 44.260 14.630 44.520 14.950 ;
        RECT 52.080 14.630 52.340 14.950 ;
        RECT 44.320 2.400 44.460 14.630 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 203.560 248.330 203.620 ;
        RECT 504.230 203.560 504.550 203.620 ;
        RECT 248.010 203.420 504.550 203.560 ;
        RECT 248.010 203.360 248.330 203.420 ;
        RECT 504.230 203.360 504.550 203.420 ;
      LAYER via ;
        RECT 248.040 203.360 248.300 203.620 ;
        RECT 504.260 203.360 504.520 203.620 ;
      LAYER met2 ;
        RECT 504.670 260.170 504.950 264.000 ;
        RECT 504.320 260.030 504.950 260.170 ;
        RECT 504.320 203.650 504.460 260.030 ;
        RECT 504.670 260.000 504.950 260.030 ;
        RECT 248.040 203.330 248.300 203.650 ;
        RECT 504.260 203.330 504.520 203.650 ;
        RECT 248.100 17.410 248.240 203.330 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 196.760 269.030 196.820 ;
        RECT 518.030 196.760 518.350 196.820 ;
        RECT 268.710 196.620 518.350 196.760 ;
        RECT 268.710 196.560 269.030 196.620 ;
        RECT 518.030 196.560 518.350 196.620 ;
        RECT 264.110 16.900 264.430 16.960 ;
        RECT 268.710 16.900 269.030 16.960 ;
        RECT 264.110 16.760 269.030 16.900 ;
        RECT 264.110 16.700 264.430 16.760 ;
        RECT 268.710 16.700 269.030 16.760 ;
      LAYER via ;
        RECT 268.740 196.560 269.000 196.820 ;
        RECT 518.060 196.560 518.320 196.820 ;
        RECT 264.140 16.700 264.400 16.960 ;
        RECT 268.740 16.700 269.000 16.960 ;
      LAYER met2 ;
        RECT 518.470 260.170 518.750 264.000 ;
        RECT 518.120 260.030 518.750 260.170 ;
        RECT 518.120 196.850 518.260 260.030 ;
        RECT 518.470 260.000 518.750 260.030 ;
        RECT 268.740 196.530 269.000 196.850 ;
        RECT 518.060 196.530 518.320 196.850 ;
        RECT 268.800 16.990 268.940 196.530 ;
        RECT 264.140 16.670 264.400 16.990 ;
        RECT 268.740 16.670 269.000 16.990 ;
        RECT 264.200 2.400 264.340 16.670 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 189.620 282.370 189.680 ;
        RECT 531.830 189.620 532.150 189.680 ;
        RECT 282.050 189.480 532.150 189.620 ;
        RECT 282.050 189.420 282.370 189.480 ;
        RECT 531.830 189.420 532.150 189.480 ;
      LAYER via ;
        RECT 282.080 189.420 282.340 189.680 ;
        RECT 531.860 189.420 532.120 189.680 ;
      LAYER met2 ;
        RECT 532.730 260.170 533.010 264.000 ;
        RECT 531.920 260.030 533.010 260.170 ;
        RECT 531.920 189.710 532.060 260.030 ;
        RECT 532.730 260.000 533.010 260.030 ;
        RECT 282.080 189.390 282.340 189.710 ;
        RECT 531.860 189.390 532.120 189.710 ;
        RECT 282.140 2.400 282.280 189.390 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 541.490 244.020 541.810 244.080 ;
        RECT 547.010 244.020 547.330 244.080 ;
        RECT 541.490 243.880 547.330 244.020 ;
        RECT 541.490 243.820 541.810 243.880 ;
        RECT 547.010 243.820 547.330 243.880 ;
        RECT 303.210 107.000 303.530 107.060 ;
        RECT 541.490 107.000 541.810 107.060 ;
        RECT 303.210 106.860 541.810 107.000 ;
        RECT 303.210 106.800 303.530 106.860 ;
        RECT 541.490 106.800 541.810 106.860 ;
        RECT 299.990 17.240 300.310 17.300 ;
        RECT 303.210 17.240 303.530 17.300 ;
        RECT 299.990 17.100 303.530 17.240 ;
        RECT 299.990 17.040 300.310 17.100 ;
        RECT 303.210 17.040 303.530 17.100 ;
      LAYER via ;
        RECT 541.520 243.820 541.780 244.080 ;
        RECT 547.040 243.820 547.300 244.080 ;
        RECT 303.240 106.800 303.500 107.060 ;
        RECT 541.520 106.800 541.780 107.060 ;
        RECT 300.020 17.040 300.280 17.300 ;
        RECT 303.240 17.040 303.500 17.300 ;
      LAYER met2 ;
        RECT 546.990 260.000 547.270 264.000 ;
        RECT 547.100 244.110 547.240 260.000 ;
        RECT 541.520 243.790 541.780 244.110 ;
        RECT 547.040 243.790 547.300 244.110 ;
        RECT 541.580 107.090 541.720 243.790 ;
        RECT 303.240 106.770 303.500 107.090 ;
        RECT 541.520 106.770 541.780 107.090 ;
        RECT 303.300 17.330 303.440 106.770 ;
        RECT 300.020 17.010 300.280 17.330 ;
        RECT 303.240 17.010 303.500 17.330 ;
        RECT 300.080 2.400 300.220 17.010 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 555.290 241.640 555.610 241.700 ;
        RECT 560.810 241.640 561.130 241.700 ;
        RECT 555.290 241.500 561.130 241.640 ;
        RECT 555.290 241.440 555.610 241.500 ;
        RECT 560.810 241.440 561.130 241.500 ;
        RECT 323.450 99.860 323.770 99.920 ;
        RECT 555.290 99.860 555.610 99.920 ;
        RECT 323.450 99.720 555.610 99.860 ;
        RECT 323.450 99.660 323.770 99.720 ;
        RECT 555.290 99.660 555.610 99.720 ;
        RECT 317.930 17.920 318.250 17.980 ;
        RECT 323.450 17.920 323.770 17.980 ;
        RECT 317.930 17.780 323.770 17.920 ;
        RECT 317.930 17.720 318.250 17.780 ;
        RECT 323.450 17.720 323.770 17.780 ;
      LAYER via ;
        RECT 555.320 241.440 555.580 241.700 ;
        RECT 560.840 241.440 561.100 241.700 ;
        RECT 323.480 99.660 323.740 99.920 ;
        RECT 555.320 99.660 555.580 99.920 ;
        RECT 317.960 17.720 318.220 17.980 ;
        RECT 323.480 17.720 323.740 17.980 ;
      LAYER met2 ;
        RECT 560.790 260.000 561.070 264.000 ;
        RECT 560.900 241.730 561.040 260.000 ;
        RECT 555.320 241.410 555.580 241.730 ;
        RECT 560.840 241.410 561.100 241.730 ;
        RECT 555.380 99.950 555.520 241.410 ;
        RECT 323.480 99.630 323.740 99.950 ;
        RECT 555.320 99.630 555.580 99.950 ;
        RECT 323.540 18.010 323.680 99.630 ;
        RECT 317.960 17.690 318.220 18.010 ;
        RECT 323.480 17.690 323.740 18.010 ;
        RECT 318.020 2.400 318.160 17.690 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 337.710 120.600 338.030 120.660 ;
        RECT 572.770 120.600 573.090 120.660 ;
        RECT 337.710 120.460 573.090 120.600 ;
        RECT 337.710 120.400 338.030 120.460 ;
        RECT 572.770 120.400 573.090 120.460 ;
      LAYER via ;
        RECT 337.740 120.400 338.000 120.660 ;
        RECT 572.800 120.400 573.060 120.660 ;
      LAYER met2 ;
        RECT 575.050 260.170 575.330 264.000 ;
        RECT 572.860 260.030 575.330 260.170 ;
        RECT 572.860 120.690 573.000 260.030 ;
        RECT 575.050 260.000 575.330 260.030 ;
        RECT 337.740 120.370 338.000 120.690 ;
        RECT 572.800 120.370 573.060 120.690 ;
        RECT 337.800 3.130 337.940 120.370 ;
        RECT 335.960 2.990 337.940 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 93.060 358.730 93.120 ;
        RECT 586.570 93.060 586.890 93.120 ;
        RECT 358.410 92.920 586.890 93.060 ;
        RECT 358.410 92.860 358.730 92.920 ;
        RECT 586.570 92.860 586.890 92.920 ;
        RECT 353.350 18.260 353.670 18.320 ;
        RECT 358.410 18.260 358.730 18.320 ;
        RECT 353.350 18.120 358.730 18.260 ;
        RECT 353.350 18.060 353.670 18.120 ;
        RECT 358.410 18.060 358.730 18.120 ;
      LAYER via ;
        RECT 358.440 92.860 358.700 93.120 ;
        RECT 586.600 92.860 586.860 93.120 ;
        RECT 353.380 18.060 353.640 18.320 ;
        RECT 358.440 18.060 358.700 18.320 ;
      LAYER met2 ;
        RECT 589.310 260.170 589.590 264.000 ;
        RECT 586.660 260.030 589.590 260.170 ;
        RECT 586.660 93.150 586.800 260.030 ;
        RECT 589.310 260.000 589.590 260.030 ;
        RECT 358.440 92.830 358.700 93.150 ;
        RECT 586.600 92.830 586.860 93.150 ;
        RECT 358.500 18.350 358.640 92.830 ;
        RECT 353.380 18.030 353.640 18.350 ;
        RECT 358.440 18.030 358.700 18.350 ;
        RECT 353.440 2.400 353.580 18.030 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 127.740 372.530 127.800 ;
        RECT 600.370 127.740 600.690 127.800 ;
        RECT 372.210 127.600 600.690 127.740 ;
        RECT 372.210 127.540 372.530 127.600 ;
        RECT 600.370 127.540 600.690 127.600 ;
        RECT 371.290 2.960 371.610 3.020 ;
        RECT 372.210 2.960 372.530 3.020 ;
        RECT 371.290 2.820 372.530 2.960 ;
        RECT 371.290 2.760 371.610 2.820 ;
        RECT 372.210 2.760 372.530 2.820 ;
      LAYER via ;
        RECT 372.240 127.540 372.500 127.800 ;
        RECT 600.400 127.540 600.660 127.800 ;
        RECT 371.320 2.760 371.580 3.020 ;
        RECT 372.240 2.760 372.500 3.020 ;
      LAYER met2 ;
        RECT 603.110 260.170 603.390 264.000 ;
        RECT 600.460 260.030 603.390 260.170 ;
        RECT 600.460 127.830 600.600 260.030 ;
        RECT 603.110 260.000 603.390 260.030 ;
        RECT 372.240 127.510 372.500 127.830 ;
        RECT 600.400 127.510 600.660 127.830 ;
        RECT 372.300 3.050 372.440 127.510 ;
        RECT 371.320 2.730 371.580 3.050 ;
        RECT 372.240 2.730 372.500 3.050 ;
        RECT 371.380 2.400 371.520 2.730 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 134.540 393.230 134.600 ;
        RECT 614.170 134.540 614.490 134.600 ;
        RECT 392.910 134.400 614.490 134.540 ;
        RECT 392.910 134.340 393.230 134.400 ;
        RECT 614.170 134.340 614.490 134.400 ;
        RECT 389.230 18.260 389.550 18.320 ;
        RECT 392.910 18.260 393.230 18.320 ;
        RECT 389.230 18.120 393.230 18.260 ;
        RECT 389.230 18.060 389.550 18.120 ;
        RECT 392.910 18.060 393.230 18.120 ;
      LAYER via ;
        RECT 392.940 134.340 393.200 134.600 ;
        RECT 614.200 134.340 614.460 134.600 ;
        RECT 389.260 18.060 389.520 18.320 ;
        RECT 392.940 18.060 393.200 18.320 ;
      LAYER met2 ;
        RECT 617.370 260.170 617.650 264.000 ;
        RECT 614.260 260.030 617.650 260.170 ;
        RECT 614.260 134.630 614.400 260.030 ;
        RECT 617.370 260.000 617.650 260.030 ;
        RECT 392.940 134.310 393.200 134.630 ;
        RECT 614.200 134.310 614.460 134.630 ;
        RECT 393.000 18.350 393.140 134.310 ;
        RECT 389.260 18.030 389.520 18.350 ;
        RECT 392.940 18.030 393.200 18.350 ;
        RECT 389.320 2.400 389.460 18.030 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 141.340 413.930 141.400 ;
        RECT 627.970 141.340 628.290 141.400 ;
        RECT 413.610 141.200 628.290 141.340 ;
        RECT 413.610 141.140 413.930 141.200 ;
        RECT 627.970 141.140 628.290 141.200 ;
        RECT 407.170 15.540 407.490 15.600 ;
        RECT 413.610 15.540 413.930 15.600 ;
        RECT 407.170 15.400 413.930 15.540 ;
        RECT 407.170 15.340 407.490 15.400 ;
        RECT 413.610 15.340 413.930 15.400 ;
      LAYER via ;
        RECT 413.640 141.140 413.900 141.400 ;
        RECT 628.000 141.140 628.260 141.400 ;
        RECT 407.200 15.340 407.460 15.600 ;
        RECT 413.640 15.340 413.900 15.600 ;
      LAYER met2 ;
        RECT 631.170 260.170 631.450 264.000 ;
        RECT 628.060 260.030 631.450 260.170 ;
        RECT 628.060 141.430 628.200 260.030 ;
        RECT 631.170 260.000 631.450 260.030 ;
        RECT 413.640 141.110 413.900 141.430 ;
        RECT 628.000 141.110 628.260 141.430 ;
        RECT 413.700 15.630 413.840 141.110 ;
        RECT 407.200 15.310 407.460 15.630 ;
        RECT 413.640 15.310 413.900 15.630 ;
        RECT 407.260 2.400 407.400 15.310 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 72.290 182.820 72.610 182.880 ;
        RECT 360.250 182.820 360.570 182.880 ;
        RECT 72.290 182.680 360.570 182.820 ;
        RECT 72.290 182.620 72.610 182.680 ;
        RECT 360.250 182.620 360.570 182.680 ;
        RECT 68.150 17.580 68.470 17.640 ;
        RECT 72.290 17.580 72.610 17.640 ;
        RECT 68.150 17.440 72.610 17.580 ;
        RECT 68.150 17.380 68.470 17.440 ;
        RECT 72.290 17.380 72.610 17.440 ;
      LAYER via ;
        RECT 72.320 182.620 72.580 182.880 ;
        RECT 360.280 182.620 360.540 182.880 ;
        RECT 68.180 17.380 68.440 17.640 ;
        RECT 72.320 17.380 72.580 17.640 ;
      LAYER met2 ;
        RECT 363.910 260.170 364.190 264.000 ;
        RECT 360.340 260.030 364.190 260.170 ;
        RECT 360.340 182.910 360.480 260.030 ;
        RECT 363.910 260.000 364.190 260.030 ;
        RECT 72.320 182.590 72.580 182.910 ;
        RECT 360.280 182.590 360.540 182.910 ;
        RECT 72.380 17.670 72.520 182.590 ;
        RECT 68.180 17.350 68.440 17.670 ;
        RECT 72.320 17.350 72.580 17.670 ;
        RECT 68.240 2.400 68.380 17.350 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 148.480 427.730 148.540 ;
        RECT 641.770 148.480 642.090 148.540 ;
        RECT 427.410 148.340 642.090 148.480 ;
        RECT 427.410 148.280 427.730 148.340 ;
        RECT 641.770 148.280 642.090 148.340 ;
        RECT 424.650 19.280 424.970 19.340 ;
        RECT 427.410 19.280 427.730 19.340 ;
        RECT 424.650 19.140 427.730 19.280 ;
        RECT 424.650 19.080 424.970 19.140 ;
        RECT 427.410 19.080 427.730 19.140 ;
      LAYER via ;
        RECT 427.440 148.280 427.700 148.540 ;
        RECT 641.800 148.280 642.060 148.540 ;
        RECT 424.680 19.080 424.940 19.340 ;
        RECT 427.440 19.080 427.700 19.340 ;
      LAYER met2 ;
        RECT 645.430 260.170 645.710 264.000 ;
        RECT 641.860 260.030 645.710 260.170 ;
        RECT 641.860 148.570 642.000 260.030 ;
        RECT 645.430 260.000 645.710 260.030 ;
        RECT 427.440 148.250 427.700 148.570 ;
        RECT 641.800 148.250 642.060 148.570 ;
        RECT 427.500 19.370 427.640 148.250 ;
        RECT 424.680 19.050 424.940 19.370 ;
        RECT 427.440 19.050 427.700 19.370 ;
        RECT 424.740 2.400 424.880 19.050 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 155.280 448.430 155.340 ;
        RECT 655.570 155.280 655.890 155.340 ;
        RECT 448.110 155.140 655.890 155.280 ;
        RECT 448.110 155.080 448.430 155.140 ;
        RECT 655.570 155.080 655.890 155.140 ;
        RECT 442.590 19.280 442.910 19.340 ;
        RECT 448.110 19.280 448.430 19.340 ;
        RECT 442.590 19.140 448.430 19.280 ;
        RECT 442.590 19.080 442.910 19.140 ;
        RECT 448.110 19.080 448.430 19.140 ;
      LAYER via ;
        RECT 448.140 155.080 448.400 155.340 ;
        RECT 655.600 155.080 655.860 155.340 ;
        RECT 442.620 19.080 442.880 19.340 ;
        RECT 448.140 19.080 448.400 19.340 ;
      LAYER met2 ;
        RECT 659.690 260.170 659.970 264.000 ;
        RECT 655.660 260.030 659.970 260.170 ;
        RECT 655.660 155.370 655.800 260.030 ;
        RECT 659.690 260.000 659.970 260.030 ;
        RECT 448.140 155.050 448.400 155.370 ;
        RECT 655.600 155.050 655.860 155.370 ;
        RECT 448.200 19.370 448.340 155.050 ;
        RECT 442.620 19.050 442.880 19.370 ;
        RECT 448.140 19.050 448.400 19.370 ;
        RECT 442.680 2.400 442.820 19.050 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 224.300 462.230 224.360 ;
        RECT 669.370 224.300 669.690 224.360 ;
        RECT 461.910 224.160 669.690 224.300 ;
        RECT 461.910 224.100 462.230 224.160 ;
        RECT 669.370 224.100 669.690 224.160 ;
      LAYER via ;
        RECT 461.940 224.100 462.200 224.360 ;
        RECT 669.400 224.100 669.660 224.360 ;
      LAYER met2 ;
        RECT 673.490 260.170 673.770 264.000 ;
        RECT 669.460 260.030 673.770 260.170 ;
        RECT 669.460 224.390 669.600 260.030 ;
        RECT 673.490 260.000 673.770 260.030 ;
        RECT 461.940 224.070 462.200 224.390 ;
        RECT 669.400 224.070 669.660 224.390 ;
        RECT 462.000 3.130 462.140 224.070 ;
        RECT 461.080 2.990 462.140 3.130 ;
        RECT 461.080 2.960 461.220 2.990 ;
        RECT 460.620 2.820 461.220 2.960 ;
        RECT 460.620 2.400 460.760 2.820 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 162.080 482.930 162.140 ;
        RECT 683.630 162.080 683.950 162.140 ;
        RECT 482.610 161.940 683.950 162.080 ;
        RECT 482.610 161.880 482.930 161.940 ;
        RECT 683.630 161.880 683.950 161.940 ;
        RECT 478.470 16.900 478.790 16.960 ;
        RECT 482.610 16.900 482.930 16.960 ;
        RECT 478.470 16.760 482.930 16.900 ;
        RECT 478.470 16.700 478.790 16.760 ;
        RECT 482.610 16.700 482.930 16.760 ;
      LAYER via ;
        RECT 482.640 161.880 482.900 162.140 ;
        RECT 683.660 161.880 683.920 162.140 ;
        RECT 478.500 16.700 478.760 16.960 ;
        RECT 482.640 16.700 482.900 16.960 ;
      LAYER met2 ;
        RECT 687.750 260.170 688.030 264.000 ;
        RECT 683.720 260.030 688.030 260.170 ;
        RECT 683.720 162.170 683.860 260.030 ;
        RECT 687.750 260.000 688.030 260.030 ;
        RECT 482.640 161.850 482.900 162.170 ;
        RECT 683.660 161.850 683.920 162.170 ;
        RECT 482.700 16.990 482.840 161.850 ;
        RECT 478.500 16.670 478.760 16.990 ;
        RECT 482.640 16.670 482.900 16.990 ;
        RECT 478.560 2.400 478.700 16.670 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.970 244.020 697.290 244.080 ;
        RECT 700.190 244.020 700.510 244.080 ;
        RECT 696.970 243.880 700.510 244.020 ;
        RECT 696.970 243.820 697.290 243.880 ;
        RECT 700.190 243.820 700.510 243.880 ;
        RECT 495.950 19.280 496.270 19.340 ;
        RECT 696.970 19.280 697.290 19.340 ;
        RECT 495.950 19.140 697.290 19.280 ;
        RECT 495.950 19.080 496.270 19.140 ;
        RECT 696.970 19.080 697.290 19.140 ;
      LAYER via ;
        RECT 697.000 243.820 697.260 244.080 ;
        RECT 700.220 243.820 700.480 244.080 ;
        RECT 495.980 19.080 496.240 19.340 ;
        RECT 697.000 19.080 697.260 19.340 ;
      LAYER met2 ;
        RECT 701.550 260.170 701.830 264.000 ;
        RECT 700.280 260.030 701.830 260.170 ;
        RECT 700.280 244.110 700.420 260.030 ;
        RECT 701.550 260.000 701.830 260.030 ;
        RECT 697.000 243.790 697.260 244.110 ;
        RECT 700.220 243.790 700.480 244.110 ;
        RECT 697.060 19.370 697.200 243.790 ;
        RECT 495.980 19.050 496.240 19.370 ;
        RECT 697.000 19.050 697.260 19.370 ;
        RECT 496.040 9.930 496.180 19.050 ;
        RECT 496.040 9.790 496.640 9.930 ;
        RECT 496.500 2.400 496.640 9.790 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 245.380 517.430 245.440 ;
        RECT 715.830 245.380 716.150 245.440 ;
        RECT 517.110 245.240 716.150 245.380 ;
        RECT 517.110 245.180 517.430 245.240 ;
        RECT 715.830 245.180 716.150 245.240 ;
        RECT 513.890 16.900 514.210 16.960 ;
        RECT 517.110 16.900 517.430 16.960 ;
        RECT 513.890 16.760 517.430 16.900 ;
        RECT 513.890 16.700 514.210 16.760 ;
        RECT 517.110 16.700 517.430 16.760 ;
      LAYER via ;
        RECT 517.140 245.180 517.400 245.440 ;
        RECT 715.860 245.180 716.120 245.440 ;
        RECT 513.920 16.700 514.180 16.960 ;
        RECT 517.140 16.700 517.400 16.960 ;
      LAYER met2 ;
        RECT 715.810 260.000 716.090 264.000 ;
        RECT 715.920 245.470 716.060 260.000 ;
        RECT 517.140 245.150 517.400 245.470 ;
        RECT 715.860 245.150 716.120 245.470 ;
        RECT 517.200 16.990 517.340 245.150 ;
        RECT 513.920 16.670 514.180 16.990 ;
        RECT 517.140 16.670 517.400 16.990 ;
        RECT 513.980 2.400 514.120 16.670 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.570 244.020 724.890 244.080 ;
        RECT 728.710 244.020 729.030 244.080 ;
        RECT 724.570 243.880 729.030 244.020 ;
        RECT 724.570 243.820 724.890 243.880 ;
        RECT 728.710 243.820 729.030 243.880 ;
        RECT 531.830 20.640 532.150 20.700 ;
        RECT 724.570 20.640 724.890 20.700 ;
        RECT 531.830 20.500 724.890 20.640 ;
        RECT 531.830 20.440 532.150 20.500 ;
        RECT 724.570 20.440 724.890 20.500 ;
      LAYER via ;
        RECT 724.600 243.820 724.860 244.080 ;
        RECT 728.740 243.820 729.000 244.080 ;
        RECT 531.860 20.440 532.120 20.700 ;
        RECT 724.600 20.440 724.860 20.700 ;
      LAYER met2 ;
        RECT 730.070 260.170 730.350 264.000 ;
        RECT 728.800 260.030 730.350 260.170 ;
        RECT 728.800 244.110 728.940 260.030 ;
        RECT 730.070 260.000 730.350 260.030 ;
        RECT 724.600 243.790 724.860 244.110 ;
        RECT 728.740 243.790 729.000 244.110 ;
        RECT 724.660 20.730 724.800 243.790 ;
        RECT 531.860 20.410 532.120 20.730 ;
        RECT 724.600 20.410 724.860 20.730 ;
        RECT 531.920 2.400 532.060 20.410 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 738.905 48.365 739.075 96.475 ;
      LAYER mcon ;
        RECT 738.905 96.305 739.075 96.475 ;
      LAYER met1 ;
        RECT 738.830 255.240 739.150 255.300 ;
        RECT 740.210 255.240 740.530 255.300 ;
        RECT 738.830 255.100 740.530 255.240 ;
        RECT 738.830 255.040 739.150 255.100 ;
        RECT 740.210 255.040 740.530 255.100 ;
        RECT 738.845 96.460 739.135 96.505 ;
        RECT 739.290 96.460 739.610 96.520 ;
        RECT 738.845 96.320 739.610 96.460 ;
        RECT 738.845 96.275 739.135 96.320 ;
        RECT 739.290 96.260 739.610 96.320 ;
        RECT 738.830 48.520 739.150 48.580 ;
        RECT 738.635 48.380 739.150 48.520 ;
        RECT 738.830 48.320 739.150 48.380 ;
        RECT 549.770 20.300 550.090 20.360 ;
        RECT 738.830 20.300 739.150 20.360 ;
        RECT 549.770 20.160 739.150 20.300 ;
        RECT 549.770 20.100 550.090 20.160 ;
        RECT 738.830 20.100 739.150 20.160 ;
      LAYER via ;
        RECT 738.860 255.040 739.120 255.300 ;
        RECT 740.240 255.040 740.500 255.300 ;
        RECT 739.320 96.260 739.580 96.520 ;
        RECT 738.860 48.320 739.120 48.580 ;
        RECT 549.800 20.100 550.060 20.360 ;
        RECT 738.860 20.100 739.120 20.360 ;
      LAYER met2 ;
        RECT 743.870 260.170 744.150 264.000 ;
        RECT 740.300 260.030 744.150 260.170 ;
        RECT 740.300 255.330 740.440 260.030 ;
        RECT 743.870 260.000 744.150 260.030 ;
        RECT 738.860 255.010 739.120 255.330 ;
        RECT 740.240 255.010 740.500 255.330 ;
        RECT 738.920 158.850 739.060 255.010 ;
        RECT 738.920 158.710 739.520 158.850 ;
        RECT 739.380 96.550 739.520 158.710 ;
        RECT 739.320 96.230 739.580 96.550 ;
        RECT 738.860 48.290 739.120 48.610 ;
        RECT 738.920 20.390 739.060 48.290 ;
        RECT 549.800 20.070 550.060 20.390 ;
        RECT 738.860 20.070 739.120 20.390 ;
        RECT 549.860 2.400 550.000 20.070 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 754.085 48.365 754.255 110.755 ;
      LAYER mcon ;
        RECT 754.085 110.585 754.255 110.755 ;
      LAYER met1 ;
        RECT 754.010 131.480 754.330 131.540 ;
        RECT 754.470 131.480 754.790 131.540 ;
        RECT 754.010 131.340 754.790 131.480 ;
        RECT 754.010 131.280 754.330 131.340 ;
        RECT 754.470 131.280 754.790 131.340 ;
        RECT 753.090 110.740 753.410 110.800 ;
        RECT 754.025 110.740 754.315 110.785 ;
        RECT 753.090 110.600 754.315 110.740 ;
        RECT 753.090 110.540 753.410 110.600 ;
        RECT 754.025 110.555 754.315 110.600 ;
        RECT 754.010 48.520 754.330 48.580 ;
        RECT 753.815 48.380 754.330 48.520 ;
        RECT 754.010 48.320 754.330 48.380 ;
        RECT 567.710 16.900 568.030 16.960 ;
        RECT 754.010 16.900 754.330 16.960 ;
        RECT 567.710 16.760 754.330 16.900 ;
        RECT 567.710 16.700 568.030 16.760 ;
        RECT 754.010 16.700 754.330 16.760 ;
      LAYER via ;
        RECT 754.040 131.280 754.300 131.540 ;
        RECT 754.500 131.280 754.760 131.540 ;
        RECT 753.120 110.540 753.380 110.800 ;
        RECT 754.040 48.320 754.300 48.580 ;
        RECT 567.740 16.700 568.000 16.960 ;
        RECT 754.040 16.700 754.300 16.960 ;
      LAYER met2 ;
        RECT 758.130 260.850 758.410 264.000 ;
        RECT 754.560 260.710 758.410 260.850 ;
        RECT 754.560 131.570 754.700 260.710 ;
        RECT 758.130 260.000 758.410 260.710 ;
        RECT 754.040 131.250 754.300 131.570 ;
        RECT 754.500 131.250 754.760 131.570 ;
        RECT 754.100 130.970 754.240 131.250 ;
        RECT 753.180 130.830 754.240 130.970 ;
        RECT 753.180 110.830 753.320 130.830 ;
        RECT 753.120 110.510 753.380 110.830 ;
        RECT 754.040 48.290 754.300 48.610 ;
        RECT 754.100 16.990 754.240 48.290 ;
        RECT 567.740 16.670 568.000 16.990 ;
        RECT 754.040 16.670 754.300 16.990 ;
        RECT 567.800 2.400 567.940 16.670 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 765.970 231.440 766.290 231.500 ;
        RECT 771.030 231.440 771.350 231.500 ;
        RECT 765.970 231.300 771.350 231.440 ;
        RECT 765.970 231.240 766.290 231.300 ;
        RECT 771.030 231.240 771.350 231.300 ;
        RECT 585.650 16.560 585.970 16.620 ;
        RECT 765.970 16.560 766.290 16.620 ;
        RECT 585.650 16.420 766.290 16.560 ;
        RECT 585.650 16.360 585.970 16.420 ;
        RECT 765.970 16.360 766.290 16.420 ;
      LAYER via ;
        RECT 766.000 231.240 766.260 231.500 ;
        RECT 771.060 231.240 771.320 231.500 ;
        RECT 585.680 16.360 585.940 16.620 ;
        RECT 766.000 16.360 766.260 16.620 ;
      LAYER met2 ;
        RECT 772.390 260.170 772.670 264.000 ;
        RECT 771.120 260.030 772.670 260.170 ;
        RECT 771.120 231.530 771.260 260.030 ;
        RECT 772.390 260.000 772.670 260.030 ;
        RECT 766.000 231.210 766.260 231.530 ;
        RECT 771.060 231.210 771.320 231.530 ;
        RECT 766.060 16.650 766.200 231.210 ;
        RECT 585.680 16.330 585.940 16.650 ;
        RECT 766.000 16.330 766.260 16.650 ;
        RECT 585.740 2.400 585.880 16.330 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 99.890 176.020 100.210 176.080 ;
        RECT 379.570 176.020 379.890 176.080 ;
        RECT 99.890 175.880 379.890 176.020 ;
        RECT 99.890 175.820 100.210 175.880 ;
        RECT 379.570 175.820 379.890 175.880 ;
        RECT 91.610 16.900 91.930 16.960 ;
        RECT 99.890 16.900 100.210 16.960 ;
        RECT 91.610 16.760 100.210 16.900 ;
        RECT 91.610 16.700 91.930 16.760 ;
        RECT 99.890 16.700 100.210 16.760 ;
      LAYER via ;
        RECT 99.920 175.820 100.180 176.080 ;
        RECT 379.600 175.820 379.860 176.080 ;
        RECT 91.640 16.700 91.900 16.960 ;
        RECT 99.920 16.700 100.180 16.960 ;
      LAYER met2 ;
        RECT 382.770 260.170 383.050 264.000 ;
        RECT 379.660 260.030 383.050 260.170 ;
        RECT 379.660 176.110 379.800 260.030 ;
        RECT 382.770 260.000 383.050 260.030 ;
        RECT 99.920 175.790 100.180 176.110 ;
        RECT 379.600 175.790 379.860 176.110 ;
        RECT 99.980 16.990 100.120 175.790 ;
        RECT 91.640 16.670 91.900 16.990 ;
        RECT 99.920 16.670 100.180 16.990 ;
        RECT 91.700 2.400 91.840 16.670 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.770 231.440 780.090 231.500 ;
        RECT 784.830 231.440 785.150 231.500 ;
        RECT 779.770 231.300 785.150 231.440 ;
        RECT 779.770 231.240 780.090 231.300 ;
        RECT 784.830 231.240 785.150 231.300 ;
        RECT 603.130 16.220 603.450 16.280 ;
        RECT 779.770 16.220 780.090 16.280 ;
        RECT 603.130 16.080 780.090 16.220 ;
        RECT 603.130 16.020 603.450 16.080 ;
        RECT 779.770 16.020 780.090 16.080 ;
      LAYER via ;
        RECT 779.800 231.240 780.060 231.500 ;
        RECT 784.860 231.240 785.120 231.500 ;
        RECT 603.160 16.020 603.420 16.280 ;
        RECT 779.800 16.020 780.060 16.280 ;
      LAYER met2 ;
        RECT 786.190 260.170 786.470 264.000 ;
        RECT 784.920 260.030 786.470 260.170 ;
        RECT 784.920 231.530 785.060 260.030 ;
        RECT 786.190 260.000 786.470 260.030 ;
        RECT 779.800 231.210 780.060 231.530 ;
        RECT 784.860 231.210 785.120 231.530 ;
        RECT 779.860 16.310 780.000 231.210 ;
        RECT 603.160 15.990 603.420 16.310 ;
        RECT 779.800 15.990 780.060 16.310 ;
        RECT 603.220 2.400 603.360 15.990 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.510 245.040 627.830 245.100 ;
        RECT 800.470 245.040 800.790 245.100 ;
        RECT 627.510 244.900 800.790 245.040 ;
        RECT 627.510 244.840 627.830 244.900 ;
        RECT 800.470 244.840 800.790 244.900 ;
        RECT 621.070 17.920 621.390 17.980 ;
        RECT 627.510 17.920 627.830 17.980 ;
        RECT 621.070 17.780 627.830 17.920 ;
        RECT 621.070 17.720 621.390 17.780 ;
        RECT 627.510 17.720 627.830 17.780 ;
      LAYER via ;
        RECT 627.540 244.840 627.800 245.100 ;
        RECT 800.500 244.840 800.760 245.100 ;
        RECT 621.100 17.720 621.360 17.980 ;
        RECT 627.540 17.720 627.800 17.980 ;
      LAYER met2 ;
        RECT 800.450 260.000 800.730 264.000 ;
        RECT 800.560 245.130 800.700 260.000 ;
        RECT 627.540 244.810 627.800 245.130 ;
        RECT 800.500 244.810 800.760 245.130 ;
        RECT 627.600 18.010 627.740 244.810 ;
        RECT 621.100 17.690 621.360 18.010 ;
        RECT 627.540 17.690 627.800 18.010 ;
        RECT 621.160 2.400 621.300 17.690 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 396.590 244.020 396.910 244.080 ;
        RECT 401.190 244.020 401.510 244.080 ;
        RECT 396.590 243.880 401.510 244.020 ;
        RECT 396.590 243.820 396.910 243.880 ;
        RECT 401.190 243.820 401.510 243.880 ;
        RECT 116.910 113.800 117.230 113.860 ;
        RECT 396.590 113.800 396.910 113.860 ;
        RECT 116.910 113.660 396.910 113.800 ;
        RECT 116.910 113.600 117.230 113.660 ;
        RECT 396.590 113.600 396.910 113.660 ;
      LAYER via ;
        RECT 396.620 243.820 396.880 244.080 ;
        RECT 401.220 243.820 401.480 244.080 ;
        RECT 116.940 113.600 117.200 113.860 ;
        RECT 396.620 113.600 396.880 113.860 ;
      LAYER met2 ;
        RECT 401.170 260.000 401.450 264.000 ;
        RECT 401.280 244.110 401.420 260.000 ;
        RECT 396.620 243.790 396.880 244.110 ;
        RECT 401.220 243.790 401.480 244.110 ;
        RECT 396.680 113.890 396.820 243.790 ;
        RECT 116.940 113.570 117.200 113.890 ;
        RECT 396.620 113.570 396.880 113.890 ;
        RECT 117.000 17.410 117.140 113.570 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 414.070 193.360 414.390 193.420 ;
        RECT 418.670 193.360 418.990 193.420 ;
        RECT 414.070 193.220 418.990 193.360 ;
        RECT 414.070 193.160 414.390 193.220 ;
        RECT 418.670 193.160 418.990 193.220 ;
        RECT 144.510 168.880 144.830 168.940 ;
        RECT 414.070 168.880 414.390 168.940 ;
        RECT 144.510 168.740 414.390 168.880 ;
        RECT 144.510 168.680 144.830 168.740 ;
        RECT 414.070 168.680 414.390 168.740 ;
        RECT 139.450 16.900 139.770 16.960 ;
        RECT 144.510 16.900 144.830 16.960 ;
        RECT 139.450 16.760 144.830 16.900 ;
        RECT 139.450 16.700 139.770 16.760 ;
        RECT 144.510 16.700 144.830 16.760 ;
      LAYER via ;
        RECT 414.100 193.160 414.360 193.420 ;
        RECT 418.700 193.160 418.960 193.420 ;
        RECT 144.540 168.680 144.800 168.940 ;
        RECT 414.100 168.680 414.360 168.940 ;
        RECT 139.480 16.700 139.740 16.960 ;
        RECT 144.540 16.700 144.800 16.960 ;
      LAYER met2 ;
        RECT 420.030 260.170 420.310 264.000 ;
        RECT 418.760 260.030 420.310 260.170 ;
        RECT 418.760 193.450 418.900 260.030 ;
        RECT 420.030 260.000 420.310 260.030 ;
        RECT 414.100 193.130 414.360 193.450 ;
        RECT 418.700 193.130 418.960 193.450 ;
        RECT 414.160 168.970 414.300 193.130 ;
        RECT 144.540 168.650 144.800 168.970 ;
        RECT 414.100 168.650 414.360 168.970 ;
        RECT 144.600 16.990 144.740 168.650 ;
        RECT 139.480 16.670 139.740 16.990 ;
        RECT 144.540 16.670 144.800 16.990 ;
        RECT 139.540 2.400 139.680 16.670 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 428.865 193.205 429.035 217.515 ;
      LAYER mcon ;
        RECT 428.865 217.345 429.035 217.515 ;
      LAYER met1 ;
        RECT 428.805 217.500 429.095 217.545 ;
        RECT 432.470 217.500 432.790 217.560 ;
        RECT 428.805 217.360 432.790 217.500 ;
        RECT 428.805 217.315 429.095 217.360 ;
        RECT 432.470 217.300 432.790 217.360 ;
        RECT 428.790 193.360 429.110 193.420 ;
        RECT 428.595 193.220 429.110 193.360 ;
        RECT 428.790 193.160 429.110 193.220 ;
        RECT 158.310 162.080 158.630 162.140 ;
        RECT 428.790 162.080 429.110 162.140 ;
        RECT 158.310 161.940 429.110 162.080 ;
        RECT 158.310 161.880 158.630 161.940 ;
        RECT 428.790 161.880 429.110 161.940 ;
      LAYER via ;
        RECT 432.500 217.300 432.760 217.560 ;
        RECT 428.820 193.160 429.080 193.420 ;
        RECT 158.340 161.880 158.600 162.140 ;
        RECT 428.820 161.880 429.080 162.140 ;
      LAYER met2 ;
        RECT 434.290 260.170 434.570 264.000 ;
        RECT 432.560 260.030 434.570 260.170 ;
        RECT 432.560 217.590 432.700 260.030 ;
        RECT 434.290 260.000 434.570 260.030 ;
        RECT 432.500 217.270 432.760 217.590 ;
        RECT 428.820 193.130 429.080 193.450 ;
        RECT 428.880 162.170 429.020 193.130 ;
        RECT 158.340 161.850 158.600 162.170 ;
        RECT 428.820 161.850 429.080 162.170 ;
        RECT 158.400 17.410 158.540 161.850 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 179.010 155.280 179.330 155.340 ;
        RECT 441.670 155.280 441.990 155.340 ;
        RECT 179.010 155.140 441.990 155.280 ;
        RECT 179.010 155.080 179.330 155.140 ;
        RECT 441.670 155.080 441.990 155.140 ;
        RECT 174.870 16.900 175.190 16.960 ;
        RECT 179.010 16.900 179.330 16.960 ;
        RECT 174.870 16.760 179.330 16.900 ;
        RECT 174.870 16.700 175.190 16.760 ;
        RECT 179.010 16.700 179.330 16.760 ;
      LAYER via ;
        RECT 179.040 155.080 179.300 155.340 ;
        RECT 441.700 155.080 441.960 155.340 ;
        RECT 174.900 16.700 175.160 16.960 ;
        RECT 179.040 16.700 179.300 16.960 ;
      LAYER met2 ;
        RECT 448.090 260.170 448.370 264.000 ;
        RECT 446.360 260.030 448.370 260.170 ;
        RECT 446.360 214.610 446.500 260.030 ;
        RECT 448.090 260.000 448.370 260.030 ;
        RECT 441.760 214.470 446.500 214.610 ;
        RECT 441.760 155.370 441.900 214.470 ;
        RECT 179.040 155.050 179.300 155.370 ;
        RECT 441.700 155.050 441.960 155.370 ;
        RECT 179.100 16.990 179.240 155.050 ;
        RECT 174.900 16.670 175.160 16.990 ;
        RECT 179.040 16.670 179.300 16.990 ;
        RECT 174.960 2.400 175.100 16.670 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 148.140 193.130 148.200 ;
        RECT 462.830 148.140 463.150 148.200 ;
        RECT 192.810 148.000 463.150 148.140 ;
        RECT 192.810 147.940 193.130 148.000 ;
        RECT 462.830 147.940 463.150 148.000 ;
      LAYER via ;
        RECT 192.840 147.940 193.100 148.200 ;
        RECT 462.860 147.940 463.120 148.200 ;
      LAYER met2 ;
        RECT 462.350 260.170 462.630 264.000 ;
        RECT 462.350 260.030 463.060 260.170 ;
        RECT 462.350 260.000 462.630 260.030 ;
        RECT 462.920 148.230 463.060 260.030 ;
        RECT 192.840 147.910 193.100 148.230 ;
        RECT 462.860 147.910 463.120 148.230 ;
        RECT 192.900 2.400 193.040 147.910 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 210.360 213.830 210.420 ;
        RECT 476.630 210.360 476.950 210.420 ;
        RECT 213.510 210.220 476.950 210.360 ;
        RECT 213.510 210.160 213.830 210.220 ;
        RECT 476.630 210.160 476.950 210.220 ;
        RECT 210.750 16.900 211.070 16.960 ;
        RECT 213.510 16.900 213.830 16.960 ;
        RECT 210.750 16.760 213.830 16.900 ;
        RECT 210.750 16.700 211.070 16.760 ;
        RECT 213.510 16.700 213.830 16.760 ;
      LAYER via ;
        RECT 213.540 210.160 213.800 210.420 ;
        RECT 476.660 210.160 476.920 210.420 ;
        RECT 210.780 16.700 211.040 16.960 ;
        RECT 213.540 16.700 213.800 16.960 ;
      LAYER met2 ;
        RECT 476.610 260.000 476.890 264.000 ;
        RECT 476.720 210.450 476.860 260.000 ;
        RECT 213.540 210.130 213.800 210.450 ;
        RECT 476.660 210.130 476.920 210.450 ;
        RECT 213.600 16.990 213.740 210.130 ;
        RECT 210.780 16.670 211.040 16.990 ;
        RECT 213.540 16.670 213.800 16.990 ;
        RECT 210.840 2.400 210.980 16.670 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 228.690 20.640 229.010 20.700 ;
        RECT 489.970 20.640 490.290 20.700 ;
        RECT 228.690 20.500 490.290 20.640 ;
        RECT 228.690 20.440 229.010 20.500 ;
        RECT 489.970 20.440 490.290 20.500 ;
      LAYER via ;
        RECT 228.720 20.440 228.980 20.700 ;
        RECT 490.000 20.440 490.260 20.700 ;
      LAYER met2 ;
        RECT 490.410 260.170 490.690 264.000 ;
        RECT 490.060 260.030 490.690 260.170 ;
        RECT 490.060 20.730 490.200 260.030 ;
        RECT 490.410 260.000 490.690 260.030 ;
        RECT 228.720 20.410 228.980 20.730 ;
        RECT 490.000 20.410 490.260 20.730 ;
        RECT 228.780 2.400 228.920 20.410 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 65.390 245.720 65.710 245.780 ;
        RECT 349.670 245.720 349.990 245.780 ;
        RECT 65.390 245.580 349.990 245.720 ;
        RECT 65.390 245.520 65.710 245.580 ;
        RECT 349.670 245.520 349.990 245.580 ;
        RECT 50.210 16.220 50.530 16.280 ;
        RECT 65.390 16.220 65.710 16.280 ;
        RECT 50.210 16.080 65.710 16.220 ;
        RECT 50.210 16.020 50.530 16.080 ;
        RECT 65.390 16.020 65.710 16.080 ;
      LAYER via ;
        RECT 65.420 245.520 65.680 245.780 ;
        RECT 349.700 245.520 349.960 245.780 ;
        RECT 50.240 16.020 50.500 16.280 ;
        RECT 65.420 16.020 65.680 16.280 ;
      LAYER met2 ;
        RECT 349.650 260.000 349.930 264.000 ;
        RECT 349.760 245.810 349.900 260.000 ;
        RECT 65.420 245.490 65.680 245.810 ;
        RECT 349.700 245.490 349.960 245.810 ;
        RECT 65.480 16.310 65.620 245.490 ;
        RECT 50.240 15.990 50.500 16.310 ;
        RECT 65.420 15.990 65.680 16.310 ;
        RECT 50.300 2.400 50.440 15.990 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 246.060 255.230 246.120 ;
        RECT 509.290 246.060 509.610 246.120 ;
        RECT 254.910 245.920 509.610 246.060 ;
        RECT 254.910 245.860 255.230 245.920 ;
        RECT 509.290 245.860 509.610 245.920 ;
        RECT 252.610 16.900 252.930 16.960 ;
        RECT 254.910 16.900 255.230 16.960 ;
        RECT 252.610 16.760 255.230 16.900 ;
        RECT 252.610 16.700 252.930 16.760 ;
        RECT 254.910 16.700 255.230 16.760 ;
      LAYER via ;
        RECT 254.940 245.860 255.200 246.120 ;
        RECT 509.320 245.860 509.580 246.120 ;
        RECT 252.640 16.700 252.900 16.960 ;
        RECT 254.940 16.700 255.200 16.960 ;
      LAYER met2 ;
        RECT 509.270 260.000 509.550 264.000 ;
        RECT 509.380 246.150 509.520 260.000 ;
        RECT 254.940 245.830 255.200 246.150 ;
        RECT 509.320 245.830 509.580 246.150 ;
        RECT 255.000 16.990 255.140 245.830 ;
        RECT 252.640 16.670 252.900 16.990 ;
        RECT 254.940 16.670 255.200 16.990 ;
        RECT 252.700 2.400 252.840 16.670 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 517.570 244.020 517.890 244.080 ;
        RECT 521.710 244.020 522.030 244.080 ;
        RECT 517.570 243.880 522.030 244.020 ;
        RECT 517.570 243.820 517.890 243.880 ;
        RECT 521.710 243.820 522.030 243.880 ;
        RECT 270.090 16.560 270.410 16.620 ;
        RECT 517.570 16.560 517.890 16.620 ;
        RECT 270.090 16.420 517.890 16.560 ;
        RECT 270.090 16.360 270.410 16.420 ;
        RECT 517.570 16.360 517.890 16.420 ;
      LAYER via ;
        RECT 517.600 243.820 517.860 244.080 ;
        RECT 521.740 243.820 522.000 244.080 ;
        RECT 270.120 16.360 270.380 16.620 ;
        RECT 517.600 16.360 517.860 16.620 ;
      LAYER met2 ;
        RECT 523.530 260.170 523.810 264.000 ;
        RECT 521.800 260.030 523.810 260.170 ;
        RECT 521.800 244.110 521.940 260.030 ;
        RECT 523.530 260.000 523.810 260.030 ;
        RECT 517.600 243.790 517.860 244.110 ;
        RECT 521.740 243.790 522.000 244.110 ;
        RECT 517.660 16.650 517.800 243.790 ;
        RECT 270.120 16.330 270.380 16.650 ;
        RECT 517.600 16.330 517.860 16.650 ;
        RECT 270.180 2.400 270.320 16.330 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 246.400 289.730 246.460 ;
        RECT 537.350 246.400 537.670 246.460 ;
        RECT 289.410 246.260 537.670 246.400 ;
        RECT 289.410 246.200 289.730 246.260 ;
        RECT 537.350 246.200 537.670 246.260 ;
      LAYER via ;
        RECT 289.440 246.200 289.700 246.460 ;
        RECT 537.380 246.200 537.640 246.460 ;
      LAYER met2 ;
        RECT 537.330 260.000 537.610 264.000 ;
        RECT 537.440 246.490 537.580 260.000 ;
        RECT 289.440 246.170 289.700 246.490 ;
        RECT 537.380 246.170 537.640 246.490 ;
        RECT 289.500 17.410 289.640 246.170 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 547.085 144.925 547.255 193.035 ;
      LAYER mcon ;
        RECT 547.085 192.865 547.255 193.035 ;
      LAYER met1 ;
        RECT 547.010 193.020 547.330 193.080 ;
        RECT 546.815 192.880 547.330 193.020 ;
        RECT 547.010 192.820 547.330 192.880 ;
        RECT 547.025 145.080 547.315 145.125 ;
        RECT 547.470 145.080 547.790 145.140 ;
        RECT 547.025 144.940 547.790 145.080 ;
        RECT 547.025 144.895 547.315 144.940 ;
        RECT 547.470 144.880 547.790 144.940 ;
        RECT 546.550 96.800 546.870 96.860 ;
        RECT 547.010 96.800 547.330 96.860 ;
        RECT 546.550 96.660 547.330 96.800 ;
        RECT 546.550 96.600 546.870 96.660 ;
        RECT 547.010 96.600 547.330 96.660 ;
        RECT 305.970 16.220 306.290 16.280 ;
        RECT 547.010 16.220 547.330 16.280 ;
        RECT 305.970 16.080 547.330 16.220 ;
        RECT 305.970 16.020 306.290 16.080 ;
        RECT 547.010 16.020 547.330 16.080 ;
      LAYER via ;
        RECT 547.040 192.820 547.300 193.080 ;
        RECT 547.500 144.880 547.760 145.140 ;
        RECT 546.580 96.600 546.840 96.860 ;
        RECT 547.040 96.600 547.300 96.860 ;
        RECT 306.000 16.020 306.260 16.280 ;
        RECT 547.040 16.020 547.300 16.280 ;
      LAYER met2 ;
        RECT 551.590 260.170 551.870 264.000 ;
        RECT 550.320 260.030 551.870 260.170 ;
        RECT 550.320 194.325 550.460 260.030 ;
        RECT 551.590 260.000 551.870 260.030 ;
        RECT 550.250 193.955 550.530 194.325 ;
        RECT 546.570 193.530 546.850 193.645 ;
        RECT 546.570 193.390 547.240 193.530 ;
        RECT 546.570 193.275 546.850 193.390 ;
        RECT 547.100 193.110 547.240 193.390 ;
        RECT 547.040 192.790 547.300 193.110 ;
        RECT 547.500 144.850 547.760 145.170 ;
        RECT 547.560 111.250 547.700 144.850 ;
        RECT 547.100 111.110 547.700 111.250 ;
        RECT 547.100 96.890 547.240 111.110 ;
        RECT 546.580 96.570 546.840 96.890 ;
        RECT 547.040 96.570 547.300 96.890 ;
        RECT 546.640 62.290 546.780 96.570 ;
        RECT 546.640 62.150 547.240 62.290 ;
        RECT 547.100 16.310 547.240 62.150 ;
        RECT 306.000 15.990 306.260 16.310 ;
        RECT 547.040 15.990 547.300 16.310 ;
        RECT 306.060 2.400 306.200 15.990 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 550.250 194.000 550.530 194.280 ;
        RECT 546.570 193.320 546.850 193.600 ;
      LAYER met3 ;
        RECT 550.225 194.290 550.555 194.305 ;
        RECT 545.870 193.990 550.555 194.290 ;
        RECT 545.870 193.610 546.170 193.990 ;
        RECT 550.225 193.975 550.555 193.990 ;
        RECT 546.545 193.610 546.875 193.625 ;
        RECT 545.870 193.310 546.875 193.610 ;
        RECT 546.545 193.295 546.875 193.310 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 246.740 324.230 246.800 ;
        RECT 565.870 246.740 566.190 246.800 ;
        RECT 323.910 246.600 566.190 246.740 ;
        RECT 323.910 246.540 324.230 246.600 ;
        RECT 565.870 246.540 566.190 246.600 ;
      LAYER via ;
        RECT 323.940 246.540 324.200 246.800 ;
        RECT 565.900 246.540 566.160 246.800 ;
      LAYER met2 ;
        RECT 565.850 260.000 566.130 264.000 ;
        RECT 565.960 246.830 566.100 260.000 ;
        RECT 323.940 246.510 324.200 246.830 ;
        RECT 565.900 246.510 566.160 246.830 ;
        RECT 324.000 2.400 324.140 246.510 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 17.240 341.710 17.300 ;
        RECT 580.590 17.240 580.910 17.300 ;
        RECT 341.390 17.100 580.910 17.240 ;
        RECT 341.390 17.040 341.710 17.100 ;
        RECT 580.590 17.040 580.910 17.100 ;
      LAYER via ;
        RECT 341.420 17.040 341.680 17.300 ;
        RECT 580.620 17.040 580.880 17.300 ;
      LAYER met2 ;
        RECT 579.650 260.170 579.930 264.000 ;
        RECT 579.650 260.030 580.820 260.170 ;
        RECT 579.650 260.000 579.930 260.030 ;
        RECT 580.680 17.330 580.820 260.030 ;
        RECT 341.420 17.010 341.680 17.330 ;
        RECT 580.620 17.010 580.880 17.330 ;
        RECT 341.480 2.400 341.620 17.010 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 15.880 359.650 15.940 ;
        RECT 359.330 15.740 567.020 15.880 ;
        RECT 359.330 15.680 359.650 15.740 ;
        RECT 566.880 15.540 567.020 15.740 ;
        RECT 594.390 15.540 594.710 15.600 ;
        RECT 566.880 15.400 594.710 15.540 ;
        RECT 594.390 15.340 594.710 15.400 ;
      LAYER via ;
        RECT 359.360 15.680 359.620 15.940 ;
        RECT 594.420 15.340 594.680 15.600 ;
      LAYER met2 ;
        RECT 593.910 260.170 594.190 264.000 ;
        RECT 593.910 260.030 594.620 260.170 ;
        RECT 593.910 260.000 594.190 260.030 ;
        RECT 359.360 15.650 359.620 15.970 ;
        RECT 359.420 2.400 359.560 15.650 ;
        RECT 594.480 15.630 594.620 260.030 ;
        RECT 594.420 15.310 594.680 15.630 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 569.165 15.725 569.335 17.595 ;
      LAYER mcon ;
        RECT 569.165 17.425 569.335 17.595 ;
      LAYER met1 ;
        RECT 377.270 17.920 377.590 17.980 ;
        RECT 377.270 17.780 448.340 17.920 ;
        RECT 377.270 17.720 377.590 17.780 ;
        RECT 448.200 17.580 448.340 17.780 ;
        RECT 569.105 17.580 569.395 17.625 ;
        RECT 448.200 17.440 569.395 17.580 ;
        RECT 569.105 17.395 569.395 17.440 ;
        RECT 569.105 15.880 569.395 15.925 ;
        RECT 607.730 15.880 608.050 15.940 ;
        RECT 569.105 15.740 608.050 15.880 ;
        RECT 569.105 15.695 569.395 15.740 ;
        RECT 607.730 15.680 608.050 15.740 ;
      LAYER via ;
        RECT 377.300 17.720 377.560 17.980 ;
        RECT 607.760 15.680 608.020 15.940 ;
      LAYER met2 ;
        RECT 607.710 260.000 607.990 264.000 ;
        RECT 377.300 17.690 377.560 18.010 ;
        RECT 377.360 2.400 377.500 17.690 ;
        RECT 607.820 15.970 607.960 260.000 ;
        RECT 607.760 15.650 608.020 15.970 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 245.040 400.130 245.100 ;
        RECT 621.990 245.040 622.310 245.100 ;
        RECT 399.810 244.900 622.310 245.040 ;
        RECT 399.810 244.840 400.130 244.900 ;
        RECT 621.990 244.840 622.310 244.900 ;
        RECT 395.210 4.320 395.530 4.380 ;
        RECT 399.810 4.320 400.130 4.380 ;
        RECT 395.210 4.180 400.130 4.320 ;
        RECT 395.210 4.120 395.530 4.180 ;
        RECT 399.810 4.120 400.130 4.180 ;
      LAYER via ;
        RECT 399.840 244.840 400.100 245.100 ;
        RECT 622.020 244.840 622.280 245.100 ;
        RECT 395.240 4.120 395.500 4.380 ;
        RECT 399.840 4.120 400.100 4.380 ;
      LAYER met2 ;
        RECT 621.970 260.000 622.250 264.000 ;
        RECT 622.080 245.130 622.220 260.000 ;
        RECT 399.840 244.810 400.100 245.130 ;
        RECT 622.020 244.810 622.280 245.130 ;
        RECT 399.900 4.410 400.040 244.810 ;
        RECT 395.240 4.090 395.500 4.410 ;
        RECT 399.840 4.090 400.100 4.410 ;
        RECT 395.300 2.400 395.440 4.090 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 636.230 260.170 636.510 264.000 ;
        RECT 635.420 260.030 636.510 260.170 ;
        RECT 635.420 16.845 635.560 260.030 ;
        RECT 636.230 260.000 636.510 260.030 ;
        RECT 413.170 16.475 413.450 16.845 ;
        RECT 635.350 16.475 635.630 16.845 ;
        RECT 413.240 2.400 413.380 16.475 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 413.170 16.520 413.450 16.800 ;
        RECT 635.350 16.520 635.630 16.800 ;
      LAYER met3 ;
        RECT 413.145 16.810 413.475 16.825 ;
        RECT 635.325 16.810 635.655 16.825 ;
        RECT 413.145 16.510 635.655 16.810 ;
        RECT 413.145 16.495 413.475 16.510 ;
        RECT 635.325 16.495 635.655 16.510 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 317.545 15.385 317.715 17.935 ;
      LAYER mcon ;
        RECT 317.545 17.765 317.715 17.935 ;
      LAYER met1 ;
        RECT 74.130 17.920 74.450 17.980 ;
        RECT 317.485 17.920 317.775 17.965 ;
        RECT 74.130 17.780 317.775 17.920 ;
        RECT 74.130 17.720 74.450 17.780 ;
        RECT 317.485 17.735 317.775 17.780 ;
        RECT 317.485 15.540 317.775 15.585 ;
        RECT 365.770 15.540 366.090 15.600 ;
        RECT 317.485 15.400 366.090 15.540 ;
        RECT 317.485 15.355 317.775 15.400 ;
        RECT 365.770 15.340 366.090 15.400 ;
      LAYER via ;
        RECT 74.160 17.720 74.420 17.980 ;
        RECT 365.800 15.340 366.060 15.600 ;
      LAYER met2 ;
        RECT 368.510 260.170 368.790 264.000 ;
        RECT 365.860 260.030 368.790 260.170 ;
        RECT 74.160 17.690 74.420 18.010 ;
        RECT 74.220 2.400 74.360 17.690 ;
        RECT 365.860 15.630 366.000 260.030 ;
        RECT 368.510 260.000 368.790 260.030 ;
        RECT 365.800 15.310 366.060 15.630 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.030 260.170 650.310 264.000 ;
        RECT 649.680 260.030 650.310 260.170 ;
        RECT 649.680 17.525 649.820 260.030 ;
        RECT 650.030 260.000 650.310 260.030 ;
        RECT 430.650 17.155 430.930 17.525 ;
        RECT 649.610 17.155 649.890 17.525 ;
        RECT 430.720 2.400 430.860 17.155 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 430.650 17.200 430.930 17.480 ;
        RECT 649.610 17.200 649.890 17.480 ;
      LAYER met3 ;
        RECT 430.625 17.490 430.955 17.505 ;
        RECT 649.585 17.490 649.915 17.505 ;
        RECT 430.625 17.190 649.915 17.490 ;
        RECT 430.625 17.175 430.955 17.190 ;
        RECT 649.585 17.175 649.915 17.190 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 608.725 15.725 608.895 17.935 ;
      LAYER mcon ;
        RECT 608.725 17.765 608.895 17.935 ;
      LAYER met1 ;
        RECT 448.570 17.920 448.890 17.980 ;
        RECT 608.665 17.920 608.955 17.965 ;
        RECT 448.570 17.780 608.955 17.920 ;
        RECT 448.570 17.720 448.890 17.780 ;
        RECT 608.665 17.735 608.955 17.780 ;
        RECT 608.665 15.880 608.955 15.925 ;
        RECT 662.470 15.880 662.790 15.940 ;
        RECT 608.665 15.740 662.790 15.880 ;
        RECT 608.665 15.695 608.955 15.740 ;
        RECT 662.470 15.680 662.790 15.740 ;
      LAYER via ;
        RECT 448.600 17.720 448.860 17.980 ;
        RECT 662.500 15.680 662.760 15.940 ;
      LAYER met2 ;
        RECT 664.290 260.170 664.570 264.000 ;
        RECT 662.560 260.030 664.570 260.170 ;
        RECT 448.600 17.690 448.860 18.010 ;
        RECT 448.660 2.400 448.800 17.690 ;
        RECT 662.560 15.970 662.700 260.030 ;
        RECT 664.290 260.000 664.570 260.030 ;
        RECT 662.500 15.650 662.760 15.970 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 18.260 466.830 18.320 ;
        RECT 676.270 18.260 676.590 18.320 ;
        RECT 466.510 18.120 676.590 18.260 ;
        RECT 466.510 18.060 466.830 18.120 ;
        RECT 676.270 18.060 676.590 18.120 ;
      LAYER via ;
        RECT 466.540 18.060 466.800 18.320 ;
        RECT 676.300 18.060 676.560 18.320 ;
      LAYER met2 ;
        RECT 678.090 260.170 678.370 264.000 ;
        RECT 676.360 260.030 678.370 260.170 ;
        RECT 676.360 18.350 676.500 260.030 ;
        RECT 678.090 260.000 678.370 260.030 ;
        RECT 466.540 18.030 466.800 18.350 ;
        RECT 676.300 18.030 676.560 18.350 ;
        RECT 466.600 2.400 466.740 18.030 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 18.940 484.770 19.000 ;
        RECT 690.070 18.940 690.390 19.000 ;
        RECT 484.450 18.800 690.390 18.940 ;
        RECT 484.450 18.740 484.770 18.800 ;
        RECT 690.070 18.740 690.390 18.800 ;
      LAYER via ;
        RECT 484.480 18.740 484.740 19.000 ;
        RECT 690.100 18.740 690.360 19.000 ;
      LAYER met2 ;
        RECT 692.350 260.170 692.630 264.000 ;
        RECT 690.160 260.030 692.630 260.170 ;
        RECT 690.160 19.030 690.300 260.030 ;
        RECT 692.350 260.000 692.630 260.030 ;
        RECT 484.480 18.710 484.740 19.030 ;
        RECT 690.100 18.710 690.360 19.030 ;
        RECT 484.540 2.400 484.680 18.710 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 502.390 18.600 502.710 18.660 ;
        RECT 703.870 18.600 704.190 18.660 ;
        RECT 502.390 18.460 704.190 18.600 ;
        RECT 502.390 18.400 502.710 18.460 ;
        RECT 703.870 18.400 704.190 18.460 ;
      LAYER via ;
        RECT 502.420 18.400 502.680 18.660 ;
        RECT 703.900 18.400 704.160 18.660 ;
      LAYER met2 ;
        RECT 706.610 260.170 706.890 264.000 ;
        RECT 703.960 260.030 706.890 260.170 ;
        RECT 703.960 18.690 704.100 260.030 ;
        RECT 706.610 260.000 706.890 260.030 ;
        RECT 502.420 18.370 502.680 18.690 ;
        RECT 703.900 18.370 704.160 18.690 ;
        RECT 502.480 2.400 502.620 18.370 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 19.620 520.190 19.680 ;
        RECT 519.870 19.480 704.560 19.620 ;
        RECT 519.870 19.420 520.190 19.480 ;
        RECT 704.420 18.260 704.560 19.480 ;
        RECT 717.670 18.260 717.990 18.320 ;
        RECT 704.420 18.120 717.990 18.260 ;
        RECT 717.670 18.060 717.990 18.120 ;
      LAYER via ;
        RECT 519.900 19.420 520.160 19.680 ;
        RECT 717.700 18.060 717.960 18.320 ;
      LAYER met2 ;
        RECT 720.410 260.170 720.690 264.000 ;
        RECT 717.760 260.030 720.690 260.170 ;
        RECT 519.900 19.390 520.160 19.710 ;
        RECT 519.960 2.400 520.100 19.390 ;
        RECT 717.760 18.350 717.900 260.030 ;
        RECT 720.410 260.000 720.690 260.030 ;
        RECT 717.700 18.030 717.960 18.350 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 245.720 538.130 245.780 ;
        RECT 734.690 245.720 735.010 245.780 ;
        RECT 537.810 245.580 735.010 245.720 ;
        RECT 537.810 245.520 538.130 245.580 ;
        RECT 734.690 245.520 735.010 245.580 ;
      LAYER via ;
        RECT 537.840 245.520 538.100 245.780 ;
        RECT 734.720 245.520 734.980 245.780 ;
      LAYER met2 ;
        RECT 734.670 260.000 734.950 264.000 ;
        RECT 734.780 245.810 734.920 260.000 ;
        RECT 537.840 245.490 538.100 245.810 ;
        RECT 734.720 245.490 734.980 245.810 ;
        RECT 537.900 2.400 538.040 245.490 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 19.960 556.070 20.020 ;
        RECT 745.270 19.960 745.590 20.020 ;
        RECT 555.750 19.820 745.590 19.960 ;
        RECT 555.750 19.760 556.070 19.820 ;
        RECT 745.270 19.760 745.590 19.820 ;
      LAYER via ;
        RECT 555.780 19.760 556.040 20.020 ;
        RECT 745.300 19.760 745.560 20.020 ;
      LAYER met2 ;
        RECT 748.470 260.170 748.750 264.000 ;
        RECT 745.360 260.030 748.750 260.170 ;
        RECT 745.360 20.050 745.500 260.030 ;
        RECT 748.470 260.000 748.750 260.030 ;
        RECT 555.780 19.730 556.040 20.050 ;
        RECT 745.300 19.730 745.560 20.050 ;
        RECT 555.840 2.400 555.980 19.730 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.210 246.060 579.530 246.120 ;
        RECT 762.750 246.060 763.070 246.120 ;
        RECT 579.210 245.920 763.070 246.060 ;
        RECT 579.210 245.860 579.530 245.920 ;
        RECT 762.750 245.860 763.070 245.920 ;
        RECT 573.690 16.220 574.010 16.280 ;
        RECT 579.210 16.220 579.530 16.280 ;
        RECT 573.690 16.080 579.530 16.220 ;
        RECT 573.690 16.020 574.010 16.080 ;
        RECT 579.210 16.020 579.530 16.080 ;
      LAYER via ;
        RECT 579.240 245.860 579.500 246.120 ;
        RECT 762.780 245.860 763.040 246.120 ;
        RECT 573.720 16.020 573.980 16.280 ;
        RECT 579.240 16.020 579.500 16.280 ;
      LAYER met2 ;
        RECT 762.730 260.000 763.010 264.000 ;
        RECT 762.840 246.150 762.980 260.000 ;
        RECT 579.240 245.830 579.500 246.150 ;
        RECT 762.780 245.830 763.040 246.150 ;
        RECT 579.300 16.310 579.440 245.830 ;
        RECT 573.720 15.990 573.980 16.310 ;
        RECT 579.240 15.990 579.500 16.310 ;
        RECT 573.780 2.400 573.920 15.990 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 739.365 17.085 739.535 18.955 ;
      LAYER mcon ;
        RECT 739.365 18.785 739.535 18.955 ;
      LAYER met1 ;
        RECT 739.305 18.940 739.595 18.985 ;
        RECT 773.330 18.940 773.650 19.000 ;
        RECT 739.305 18.800 773.650 18.940 ;
        RECT 739.305 18.755 739.595 18.800 ;
        RECT 773.330 18.740 773.650 18.800 ;
        RECT 591.170 17.240 591.490 17.300 ;
        RECT 739.305 17.240 739.595 17.285 ;
        RECT 591.170 17.100 739.595 17.240 ;
        RECT 591.170 17.040 591.490 17.100 ;
        RECT 739.305 17.055 739.595 17.100 ;
      LAYER via ;
        RECT 773.360 18.740 773.620 19.000 ;
        RECT 591.200 17.040 591.460 17.300 ;
      LAYER met2 ;
        RECT 776.990 260.170 777.270 264.000 ;
        RECT 773.420 260.030 777.270 260.170 ;
        RECT 773.420 19.030 773.560 260.030 ;
        RECT 776.990 260.000 777.270 260.030 ;
        RECT 773.360 18.710 773.620 19.030 ;
        RECT 591.200 17.010 591.460 17.330 ;
        RECT 591.260 2.400 591.400 17.010 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 387.370 260.000 387.650 264.000 ;
        RECT 387.480 16.845 387.620 260.000 ;
        RECT 97.610 16.475 97.890 16.845 ;
        RECT 387.410 16.475 387.690 16.845 ;
        RECT 97.680 2.400 97.820 16.475 ;
        RECT 97.470 -4.800 98.030 2.400 ;
      LAYER via2 ;
        RECT 97.610 16.520 97.890 16.800 ;
        RECT 387.410 16.520 387.690 16.800 ;
      LAYER met3 ;
        RECT 97.585 16.810 97.915 16.825 ;
        RECT 387.385 16.810 387.715 16.825 ;
        RECT 97.585 16.510 387.715 16.810 ;
        RECT 97.585 16.495 97.915 16.510 ;
        RECT 387.385 16.495 387.715 16.510 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 246.400 614.030 246.460 ;
        RECT 790.810 246.400 791.130 246.460 ;
        RECT 613.710 246.260 791.130 246.400 ;
        RECT 613.710 246.200 614.030 246.260 ;
        RECT 790.810 246.200 791.130 246.260 ;
        RECT 609.110 17.920 609.430 17.980 ;
        RECT 613.710 17.920 614.030 17.980 ;
        RECT 609.110 17.780 614.030 17.920 ;
        RECT 609.110 17.720 609.430 17.780 ;
        RECT 613.710 17.720 614.030 17.780 ;
      LAYER via ;
        RECT 613.740 246.200 614.000 246.460 ;
        RECT 790.840 246.200 791.100 246.460 ;
        RECT 609.140 17.720 609.400 17.980 ;
        RECT 613.740 17.720 614.000 17.980 ;
      LAYER met2 ;
        RECT 790.790 260.000 791.070 264.000 ;
        RECT 790.900 246.490 791.040 260.000 ;
        RECT 613.740 246.170 614.000 246.490 ;
        RECT 790.840 246.170 791.100 246.490 ;
        RECT 613.800 18.010 613.940 246.170 ;
        RECT 609.140 17.690 609.400 18.010 ;
        RECT 613.740 17.690 614.000 18.010 ;
        RECT 609.200 2.400 609.340 17.690 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 628.060 17.780 648.900 17.920 ;
        RECT 627.050 17.580 627.370 17.640 ;
        RECT 628.060 17.580 628.200 17.780 ;
        RECT 627.050 17.440 628.200 17.580 ;
        RECT 648.760 17.580 648.900 17.780 ;
        RECT 801.390 17.580 801.710 17.640 ;
        RECT 648.760 17.440 739.980 17.580 ;
        RECT 627.050 17.380 627.370 17.440 ;
        RECT 739.840 17.240 739.980 17.440 ;
        RECT 787.220 17.440 801.710 17.580 ;
        RECT 787.220 17.240 787.360 17.440 ;
        RECT 801.390 17.380 801.710 17.440 ;
        RECT 739.840 17.100 787.360 17.240 ;
      LAYER via ;
        RECT 627.080 17.380 627.340 17.640 ;
        RECT 801.420 17.380 801.680 17.640 ;
      LAYER met2 ;
        RECT 805.050 260.170 805.330 264.000 ;
        RECT 801.480 260.030 805.330 260.170 ;
        RECT 801.480 17.670 801.620 260.030 ;
        RECT 805.050 260.000 805.330 260.030 ;
        RECT 627.080 17.350 627.340 17.670 ;
        RECT 801.420 17.350 801.680 17.670 ;
        RECT 627.140 2.400 627.280 17.350 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 400.730 138.280 401.050 138.340 ;
        RECT 401.190 138.280 401.510 138.340 ;
        RECT 400.730 138.140 401.510 138.280 ;
        RECT 400.730 138.080 401.050 138.140 ;
        RECT 401.190 138.080 401.510 138.140 ;
        RECT 400.270 62.120 400.590 62.180 ;
        RECT 402.110 62.120 402.430 62.180 ;
        RECT 400.270 61.980 402.430 62.120 ;
        RECT 400.270 61.920 400.590 61.980 ;
        RECT 402.110 61.920 402.430 61.980 ;
        RECT 121.510 18.600 121.830 18.660 ;
        RECT 400.730 18.600 401.050 18.660 ;
        RECT 121.510 18.460 401.050 18.600 ;
        RECT 121.510 18.400 121.830 18.460 ;
        RECT 400.730 18.400 401.050 18.460 ;
      LAYER via ;
        RECT 400.760 138.080 401.020 138.340 ;
        RECT 401.220 138.080 401.480 138.340 ;
        RECT 400.300 61.920 400.560 62.180 ;
        RECT 402.140 61.920 402.400 62.180 ;
        RECT 121.540 18.400 121.800 18.660 ;
        RECT 400.760 18.400 401.020 18.660 ;
      LAYER met2 ;
        RECT 406.230 260.170 406.510 264.000 ;
        RECT 404.960 260.030 406.510 260.170 ;
        RECT 404.960 230.250 405.100 260.030 ;
        RECT 406.230 260.000 406.510 260.030 ;
        RECT 401.280 230.110 405.100 230.250 ;
        RECT 401.280 138.370 401.420 230.110 ;
        RECT 400.760 138.050 401.020 138.370 ;
        RECT 401.220 138.050 401.480 138.370 ;
        RECT 400.820 96.405 400.960 138.050 ;
        RECT 400.750 96.035 401.030 96.405 ;
        RECT 402.130 96.035 402.410 96.405 ;
        RECT 402.200 62.210 402.340 96.035 ;
        RECT 400.300 61.890 400.560 62.210 ;
        RECT 402.140 61.890 402.400 62.210 ;
        RECT 400.360 48.010 400.500 61.890 ;
        RECT 400.360 47.870 400.960 48.010 ;
        RECT 400.820 18.690 400.960 47.870 ;
        RECT 121.540 18.370 121.800 18.690 ;
        RECT 400.760 18.370 401.020 18.690 ;
        RECT 121.600 2.400 121.740 18.370 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 400.750 96.080 401.030 96.360 ;
        RECT 402.130 96.080 402.410 96.360 ;
      LAYER met3 ;
        RECT 400.725 96.370 401.055 96.385 ;
        RECT 402.105 96.370 402.435 96.385 ;
        RECT 400.725 96.070 402.435 96.370 ;
        RECT 400.725 96.055 401.055 96.070 ;
        RECT 402.105 96.055 402.435 96.070 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 18.940 145.750 19.000 ;
        RECT 420.970 18.940 421.290 19.000 ;
        RECT 145.430 18.800 421.290 18.940 ;
        RECT 145.430 18.740 145.750 18.800 ;
        RECT 420.970 18.740 421.290 18.800 ;
      LAYER via ;
        RECT 145.460 18.740 145.720 19.000 ;
        RECT 421.000 18.740 421.260 19.000 ;
      LAYER met2 ;
        RECT 424.630 260.170 424.910 264.000 ;
        RECT 421.060 260.030 424.910 260.170 ;
        RECT 421.060 19.030 421.200 260.030 ;
        RECT 424.630 260.000 424.910 260.030 ;
        RECT 145.460 18.710 145.720 19.030 ;
        RECT 421.000 18.710 421.260 19.030 ;
        RECT 145.520 2.400 145.660 18.710 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 19.280 163.690 19.340 ;
        RECT 163.370 19.140 421.660 19.280 ;
        RECT 163.370 19.080 163.690 19.140 ;
        RECT 421.520 18.940 421.660 19.140 ;
        RECT 434.770 18.940 435.090 19.000 ;
        RECT 421.520 18.800 435.090 18.940 ;
        RECT 434.770 18.740 435.090 18.800 ;
      LAYER via ;
        RECT 163.400 19.080 163.660 19.340 ;
        RECT 434.800 18.740 435.060 19.000 ;
      LAYER met2 ;
        RECT 438.890 260.170 439.170 264.000 ;
        RECT 434.860 260.030 439.170 260.170 ;
        RECT 163.400 19.050 163.660 19.370 ;
        RECT 163.460 2.400 163.600 19.050 ;
        RECT 434.860 19.030 435.000 260.030 ;
        RECT 438.890 260.000 439.170 260.030 ;
        RECT 434.800 18.710 435.060 19.030 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 19.960 181.170 20.020 ;
        RECT 448.570 19.960 448.890 20.020 ;
        RECT 180.850 19.820 448.890 19.960 ;
        RECT 180.850 19.760 181.170 19.820 ;
        RECT 448.570 19.760 448.890 19.820 ;
      LAYER via ;
        RECT 180.880 19.760 181.140 20.020 ;
        RECT 448.600 19.760 448.860 20.020 ;
      LAYER met2 ;
        RECT 453.150 260.170 453.430 264.000 ;
        RECT 448.660 260.030 453.430 260.170 ;
        RECT 448.660 20.050 448.800 260.030 ;
        RECT 453.150 260.000 453.430 260.030 ;
        RECT 180.880 19.730 181.140 20.050 ;
        RECT 448.600 19.730 448.860 20.050 ;
        RECT 180.940 2.400 181.080 19.730 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 462.370 244.020 462.690 244.080 ;
        RECT 465.590 244.020 465.910 244.080 ;
        RECT 462.370 243.880 465.910 244.020 ;
        RECT 462.370 243.820 462.690 243.880 ;
        RECT 465.590 243.820 465.910 243.880 ;
        RECT 198.790 19.620 199.110 19.680 ;
        RECT 462.370 19.620 462.690 19.680 ;
        RECT 198.790 19.480 462.690 19.620 ;
        RECT 198.790 19.420 199.110 19.480 ;
        RECT 462.370 19.420 462.690 19.480 ;
      LAYER via ;
        RECT 462.400 243.820 462.660 244.080 ;
        RECT 465.620 243.820 465.880 244.080 ;
        RECT 198.820 19.420 199.080 19.680 ;
        RECT 462.400 19.420 462.660 19.680 ;
      LAYER met2 ;
        RECT 466.950 260.170 467.230 264.000 ;
        RECT 465.680 260.030 467.230 260.170 ;
        RECT 465.680 244.110 465.820 260.030 ;
        RECT 466.950 260.000 467.230 260.030 ;
        RECT 462.400 243.790 462.660 244.110 ;
        RECT 465.620 243.790 465.880 244.110 ;
        RECT 462.460 19.710 462.600 243.790 ;
        RECT 198.820 19.390 199.080 19.710 ;
        RECT 462.400 19.390 462.660 19.710 ;
        RECT 198.880 2.400 199.020 19.390 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 476.170 244.020 476.490 244.080 ;
        RECT 479.390 244.020 479.710 244.080 ;
        RECT 476.170 243.880 479.710 244.020 ;
        RECT 476.170 243.820 476.490 243.880 ;
        RECT 479.390 243.820 479.710 243.880 ;
        RECT 216.730 20.300 217.050 20.360 ;
        RECT 216.730 20.160 463.060 20.300 ;
        RECT 216.730 20.100 217.050 20.160 ;
        RECT 462.920 19.280 463.060 20.160 ;
        RECT 476.170 19.280 476.490 19.340 ;
        RECT 462.920 19.140 476.490 19.280 ;
        RECT 476.170 19.080 476.490 19.140 ;
      LAYER via ;
        RECT 476.200 243.820 476.460 244.080 ;
        RECT 479.420 243.820 479.680 244.080 ;
        RECT 216.760 20.100 217.020 20.360 ;
        RECT 476.200 19.080 476.460 19.340 ;
      LAYER met2 ;
        RECT 481.210 260.170 481.490 264.000 ;
        RECT 479.480 260.030 481.490 260.170 ;
        RECT 479.480 244.110 479.620 260.030 ;
        RECT 481.210 260.000 481.490 260.030 ;
        RECT 476.200 243.790 476.460 244.110 ;
        RECT 479.420 243.790 479.680 244.110 ;
        RECT 216.760 20.070 217.020 20.390 ;
        RECT 216.820 2.400 216.960 20.070 ;
        RECT 476.260 19.370 476.400 243.790 ;
        RECT 476.200 19.050 476.460 19.370 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 478.085 16.745 478.255 18.615 ;
      LAYER mcon ;
        RECT 478.085 18.445 478.255 18.615 ;
      LAYER met1 ;
        RECT 490.430 179.760 490.750 179.820 ;
        RECT 491.350 179.760 491.670 179.820 ;
        RECT 490.430 179.620 491.670 179.760 ;
        RECT 490.430 179.560 490.750 179.620 ;
        RECT 491.350 179.560 491.670 179.620 ;
        RECT 490.430 83.200 490.750 83.260 ;
        RECT 491.350 83.200 491.670 83.260 ;
        RECT 490.430 83.060 491.670 83.200 ;
        RECT 490.430 83.000 490.750 83.060 ;
        RECT 491.350 83.000 491.670 83.060 ;
        RECT 478.025 18.600 478.315 18.645 ;
        RECT 491.350 18.600 491.670 18.660 ;
        RECT 478.025 18.460 491.670 18.600 ;
        RECT 478.025 18.415 478.315 18.460 ;
        RECT 491.350 18.400 491.670 18.460 ;
        RECT 478.025 16.900 478.315 16.945 ;
        RECT 269.260 16.760 478.315 16.900 ;
        RECT 234.670 16.560 234.990 16.620 ;
        RECT 269.260 16.560 269.400 16.760 ;
        RECT 478.025 16.715 478.315 16.760 ;
        RECT 234.670 16.420 269.400 16.560 ;
        RECT 234.670 16.360 234.990 16.420 ;
      LAYER via ;
        RECT 490.460 179.560 490.720 179.820 ;
        RECT 491.380 179.560 491.640 179.820 ;
        RECT 490.460 83.000 490.720 83.260 ;
        RECT 491.380 83.000 491.640 83.260 ;
        RECT 491.380 18.400 491.640 18.660 ;
        RECT 234.700 16.360 234.960 16.620 ;
      LAYER met2 ;
        RECT 495.010 260.170 495.290 264.000 ;
        RECT 491.440 260.030 495.290 260.170 ;
        RECT 491.440 179.850 491.580 260.030 ;
        RECT 495.010 260.000 495.290 260.030 ;
        RECT 490.460 179.530 490.720 179.850 ;
        RECT 491.380 179.530 491.640 179.850 ;
        RECT 490.520 130.970 490.660 179.530 ;
        RECT 490.520 130.830 491.580 130.970 ;
        RECT 491.440 83.290 491.580 130.830 ;
        RECT 490.460 82.970 490.720 83.290 ;
        RECT 491.380 82.970 491.640 83.290 ;
        RECT 490.520 34.410 490.660 82.970 ;
        RECT 490.520 34.270 491.580 34.410 ;
        RECT 491.440 18.690 491.580 34.270 ;
        RECT 491.380 18.370 491.640 18.690 ;
        RECT 234.700 16.330 234.960 16.650 ;
        RECT 234.760 2.400 234.900 16.330 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 352.430 17.920 352.750 17.980 ;
        RECT 56.190 17.780 72.980 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 72.840 17.580 72.980 17.780 ;
        RECT 327.680 17.780 352.750 17.920 ;
        RECT 327.680 17.580 327.820 17.780 ;
        RECT 352.430 17.720 352.750 17.780 ;
        RECT 72.840 17.440 327.820 17.580 ;
      LAYER via ;
        RECT 56.220 17.720 56.480 17.980 ;
        RECT 352.460 17.720 352.720 17.980 ;
      LAYER met2 ;
        RECT 354.250 260.170 354.530 264.000 ;
        RECT 352.520 260.030 354.530 260.170 ;
        RECT 352.520 18.010 352.660 260.030 ;
        RECT 354.250 260.000 354.530 260.030 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 352.460 17.690 352.720 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 245.040 86.410 245.100 ;
        RECT 373.130 245.040 373.450 245.100 ;
        RECT 86.090 244.900 373.450 245.040 ;
        RECT 86.090 244.840 86.410 244.900 ;
        RECT 373.130 244.840 373.450 244.900 ;
        RECT 80.110 15.880 80.430 15.940 ;
        RECT 86.090 15.880 86.410 15.940 ;
        RECT 80.110 15.740 86.410 15.880 ;
        RECT 80.110 15.680 80.430 15.740 ;
        RECT 86.090 15.680 86.410 15.740 ;
      LAYER via ;
        RECT 86.120 244.840 86.380 245.100 ;
        RECT 373.160 244.840 373.420 245.100 ;
        RECT 80.140 15.680 80.400 15.940 ;
        RECT 86.120 15.680 86.380 15.940 ;
      LAYER met2 ;
        RECT 373.110 260.000 373.390 264.000 ;
        RECT 373.220 245.130 373.360 260.000 ;
        RECT 86.120 244.810 86.380 245.130 ;
        RECT 373.160 244.810 373.420 245.130 ;
        RECT 86.180 15.970 86.320 244.810 ;
        RECT 80.140 15.650 80.400 15.970 ;
        RECT 86.120 15.650 86.380 15.970 ;
        RECT 80.200 2.400 80.340 15.650 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 386.930 231.100 387.250 231.160 ;
        RECT 390.150 231.100 390.470 231.160 ;
        RECT 386.930 230.960 390.470 231.100 ;
        RECT 386.930 230.900 387.250 230.960 ;
        RECT 390.150 230.900 390.470 230.960 ;
        RECT 103.570 18.260 103.890 18.320 ;
        RECT 386.930 18.260 387.250 18.320 ;
        RECT 103.570 18.120 353.120 18.260 ;
        RECT 103.570 18.060 103.890 18.120 ;
        RECT 352.980 17.920 353.120 18.120 ;
        RECT 358.960 18.120 387.250 18.260 ;
        RECT 358.960 17.920 359.100 18.120 ;
        RECT 386.930 18.060 387.250 18.120 ;
        RECT 352.980 17.780 359.100 17.920 ;
      LAYER via ;
        RECT 386.960 230.900 387.220 231.160 ;
        RECT 390.180 230.900 390.440 231.160 ;
        RECT 103.600 18.060 103.860 18.320 ;
        RECT 386.960 18.060 387.220 18.320 ;
      LAYER met2 ;
        RECT 391.970 260.170 392.250 264.000 ;
        RECT 390.240 260.030 392.250 260.170 ;
        RECT 390.240 231.190 390.380 260.030 ;
        RECT 391.970 260.000 392.250 260.030 ;
        RECT 386.960 230.870 387.220 231.190 ;
        RECT 390.180 230.870 390.440 231.190 ;
        RECT 387.020 18.350 387.160 230.870 ;
        RECT 103.600 18.030 103.860 18.350 ;
        RECT 386.960 18.030 387.220 18.350 ;
        RECT 103.660 2.400 103.800 18.030 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 410.830 260.170 411.110 264.000 ;
        RECT 407.720 260.030 411.110 260.170 ;
        RECT 407.720 17.525 407.860 260.030 ;
        RECT 410.830 260.000 411.110 260.030 ;
        RECT 127.510 17.155 127.790 17.525 ;
        RECT 407.650 17.155 407.930 17.525 ;
        RECT 127.580 2.400 127.720 17.155 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 127.510 17.200 127.790 17.480 ;
        RECT 407.650 17.200 407.930 17.480 ;
      LAYER met3 ;
        RECT 127.485 17.490 127.815 17.505 ;
        RECT 407.625 17.490 407.955 17.505 ;
        RECT 127.485 17.190 407.955 17.490 ;
        RECT 127.485 17.175 127.815 17.190 ;
        RECT 407.625 17.175 407.955 17.190 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 245.380 45.010 245.440 ;
        RECT 330.810 245.380 331.130 245.440 ;
        RECT 44.690 245.240 331.130 245.380 ;
        RECT 44.690 245.180 45.010 245.240 ;
        RECT 330.810 245.180 331.130 245.240 ;
        RECT 26.290 18.940 26.610 19.000 ;
        RECT 44.690 18.940 45.010 19.000 ;
        RECT 26.290 18.800 45.010 18.940 ;
        RECT 26.290 18.740 26.610 18.800 ;
        RECT 44.690 18.740 45.010 18.800 ;
      LAYER via ;
        RECT 44.720 245.180 44.980 245.440 ;
        RECT 330.840 245.180 331.100 245.440 ;
        RECT 26.320 18.740 26.580 19.000 ;
        RECT 44.720 18.740 44.980 19.000 ;
      LAYER met2 ;
        RECT 330.790 260.000 331.070 264.000 ;
        RECT 330.900 245.470 331.040 260.000 ;
        RECT 44.720 245.150 44.980 245.470 ;
        RECT 330.840 245.150 331.100 245.470 ;
        RECT 44.780 19.030 44.920 245.150 ;
        RECT 26.320 18.710 26.580 19.030 ;
        RECT 44.720 18.710 44.980 19.030 ;
        RECT 26.380 2.400 26.520 18.710 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 299.605 15.725 299.775 17.255 ;
      LAYER mcon ;
        RECT 299.605 17.085 299.775 17.255 ;
      LAYER met1 ;
        RECT 32.270 17.240 32.590 17.300 ;
        RECT 299.545 17.240 299.835 17.285 ;
        RECT 32.270 17.100 299.835 17.240 ;
        RECT 32.270 17.040 32.590 17.100 ;
        RECT 299.545 17.055 299.835 17.100 ;
        RECT 299.545 15.880 299.835 15.925 ;
        RECT 331.730 15.880 332.050 15.940 ;
        RECT 299.545 15.740 332.050 15.880 ;
        RECT 299.545 15.695 299.835 15.740 ;
        RECT 331.730 15.680 332.050 15.740 ;
      LAYER via ;
        RECT 32.300 17.040 32.560 17.300 ;
        RECT 331.760 15.680 332.020 15.940 ;
      LAYER met2 ;
        RECT 335.850 260.170 336.130 264.000 ;
        RECT 331.820 260.030 336.130 260.170 ;
        RECT 32.300 17.010 32.560 17.330 ;
        RECT 32.360 2.400 32.500 17.010 ;
        RECT 331.820 15.970 331.960 260.030 ;
        RECT 335.850 260.000 336.130 260.030 ;
        RECT 331.760 15.650 332.020 15.970 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 3260.000 367.020 3528.900 ;
        RECT 544.020 3260.000 547.020 3528.900 ;
        RECT 724.020 3260.000 727.020 3528.900 ;
        RECT 904.020 3260.000 907.020 3528.900 ;
        RECT 1084.020 3260.000 1087.020 3528.900 ;
        RECT 1264.020 3260.000 1267.020 3528.900 ;
        RECT 1444.020 3260.000 1447.020 3528.900 ;
        RECT 1624.020 3260.000 1627.020 3528.900 ;
        RECT 1804.020 3260.000 1807.020 3528.900 ;
        RECT 1984.020 3260.000 1987.020 3528.900 ;
        RECT 2164.020 3260.000 2167.020 3528.900 ;
        RECT 2344.020 3260.000 2347.020 3528.900 ;
        RECT 2524.020 3260.000 2527.020 3528.900 ;
        RECT 364.020 -9.220 367.020 260.000 ;
        RECT 544.020 -9.220 547.020 260.000 ;
        RECT 724.020 -9.220 727.020 260.000 ;
        RECT 904.020 -9.220 907.020 260.000 ;
        RECT 1084.020 -9.220 1087.020 260.000 ;
        RECT 1264.020 -9.220 1267.020 260.000 ;
        RECT 1444.020 -9.220 1447.020 260.000 ;
        RECT 1624.020 -9.220 1627.020 260.000 ;
        RECT 1804.020 -9.220 1807.020 260.000 ;
        RECT 1984.020 -9.220 1987.020 260.000 ;
        RECT 2164.020 -9.220 2167.020 260.000 ;
        RECT 2344.020 -9.220 2347.020 260.000 ;
        RECT 2524.020 -9.220 2527.020 260.000 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 3260.000 457.020 3528.900 ;
        RECT 634.020 3260.000 637.020 3528.900 ;
        RECT 814.020 3260.000 817.020 3528.900 ;
        RECT 994.020 3260.000 997.020 3528.900 ;
        RECT 1174.020 3260.000 1177.020 3528.900 ;
        RECT 1354.020 3260.000 1357.020 3528.900 ;
        RECT 1534.020 3260.000 1537.020 3528.900 ;
        RECT 1714.020 3260.000 1717.020 3528.900 ;
        RECT 1894.020 3260.000 1897.020 3528.900 ;
        RECT 2074.020 3260.000 2077.020 3528.900 ;
        RECT 2254.020 3260.000 2257.020 3528.900 ;
        RECT 2434.020 3260.000 2437.020 3528.900 ;
        RECT 454.020 -9.220 457.020 260.000 ;
        RECT 634.020 -9.220 637.020 260.000 ;
        RECT 814.020 -9.220 817.020 260.000 ;
        RECT 994.020 -9.220 997.020 260.000 ;
        RECT 1174.020 -9.220 1177.020 260.000 ;
        RECT 1354.020 -9.220 1357.020 260.000 ;
        RECT 1534.020 -9.220 1537.020 260.000 ;
        RECT 1714.020 -9.220 1717.020 260.000 ;
        RECT 1894.020 -9.220 1897.020 260.000 ;
        RECT 2074.020 -9.220 2077.020 260.000 ;
        RECT 2254.020 -9.220 2257.020 260.000 ;
        RECT 2434.020 -9.220 2437.020 260.000 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 3260.000 385.020 3538.100 ;
        RECT 562.020 3260.000 565.020 3538.100 ;
        RECT 742.020 3260.000 745.020 3538.100 ;
        RECT 922.020 3260.000 925.020 3538.100 ;
        RECT 1102.020 3260.000 1105.020 3538.100 ;
        RECT 1282.020 3260.000 1285.020 3538.100 ;
        RECT 1462.020 3260.000 1465.020 3538.100 ;
        RECT 1642.020 3260.000 1645.020 3538.100 ;
        RECT 1822.020 3260.000 1825.020 3538.100 ;
        RECT 2002.020 3260.000 2005.020 3538.100 ;
        RECT 2182.020 3260.000 2185.020 3538.100 ;
        RECT 2362.020 3260.000 2365.020 3538.100 ;
        RECT 2542.020 3260.000 2545.020 3538.100 ;
        RECT 382.020 -18.420 385.020 260.000 ;
        RECT 562.020 -18.420 565.020 260.000 ;
        RECT 742.020 -18.420 745.020 260.000 ;
        RECT 922.020 -18.420 925.020 260.000 ;
        RECT 1102.020 -18.420 1105.020 260.000 ;
        RECT 1282.020 -18.420 1285.020 260.000 ;
        RECT 1462.020 -18.420 1465.020 260.000 ;
        RECT 1642.020 -18.420 1645.020 260.000 ;
        RECT 1822.020 -18.420 1825.020 260.000 ;
        RECT 2002.020 -18.420 2005.020 260.000 ;
        RECT 2182.020 -18.420 2185.020 260.000 ;
        RECT 2362.020 -18.420 2365.020 260.000 ;
        RECT 2542.020 -18.420 2545.020 260.000 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 3260.000 475.020 3538.100 ;
        RECT 652.020 3260.000 655.020 3538.100 ;
        RECT 832.020 3260.000 835.020 3538.100 ;
        RECT 1012.020 3260.000 1015.020 3538.100 ;
        RECT 1192.020 3260.000 1195.020 3538.100 ;
        RECT 1372.020 3260.000 1375.020 3538.100 ;
        RECT 1552.020 3260.000 1555.020 3538.100 ;
        RECT 1732.020 3260.000 1735.020 3538.100 ;
        RECT 1912.020 3260.000 1915.020 3538.100 ;
        RECT 2092.020 3260.000 2095.020 3538.100 ;
        RECT 2272.020 3260.000 2275.020 3538.100 ;
        RECT 2452.020 3260.000 2455.020 3538.100 ;
        RECT 472.020 -18.420 475.020 260.000 ;
        RECT 652.020 -18.420 655.020 260.000 ;
        RECT 832.020 -18.420 835.020 260.000 ;
        RECT 1012.020 -18.420 1015.020 260.000 ;
        RECT 1192.020 -18.420 1195.020 260.000 ;
        RECT 1372.020 -18.420 1375.020 260.000 ;
        RECT 1552.020 -18.420 1555.020 260.000 ;
        RECT 1732.020 -18.420 1735.020 260.000 ;
        RECT 1912.020 -18.420 1915.020 260.000 ;
        RECT 2092.020 -18.420 2095.020 260.000 ;
        RECT 2272.020 -18.420 2275.020 260.000 ;
        RECT 2452.020 -18.420 2455.020 260.000 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 3260.000 403.020 3547.300 ;
        RECT 580.020 3260.000 583.020 3547.300 ;
        RECT 760.020 3260.000 763.020 3547.300 ;
        RECT 940.020 3260.000 943.020 3547.300 ;
        RECT 1120.020 3260.000 1123.020 3547.300 ;
        RECT 1300.020 3260.000 1303.020 3547.300 ;
        RECT 1480.020 3260.000 1483.020 3547.300 ;
        RECT 1660.020 3260.000 1663.020 3547.300 ;
        RECT 1840.020 3260.000 1843.020 3547.300 ;
        RECT 2020.020 3260.000 2023.020 3547.300 ;
        RECT 2200.020 3260.000 2203.020 3547.300 ;
        RECT 2380.020 3260.000 2383.020 3547.300 ;
        RECT 2560.020 3260.000 2563.020 3547.300 ;
        RECT 400.020 -27.620 403.020 260.000 ;
        RECT 580.020 -27.620 583.020 260.000 ;
        RECT 760.020 -27.620 763.020 260.000 ;
        RECT 940.020 -27.620 943.020 260.000 ;
        RECT 1120.020 -27.620 1123.020 260.000 ;
        RECT 1300.020 -27.620 1303.020 260.000 ;
        RECT 1480.020 -27.620 1483.020 260.000 ;
        RECT 1660.020 -27.620 1663.020 260.000 ;
        RECT 1840.020 -27.620 1843.020 260.000 ;
        RECT 2020.020 -27.620 2023.020 260.000 ;
        RECT 2200.020 -27.620 2203.020 260.000 ;
        RECT 2380.020 -27.620 2383.020 260.000 ;
        RECT 2560.020 -27.620 2563.020 260.000 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 3260.000 313.020 3547.300 ;
        RECT 490.020 3260.000 493.020 3547.300 ;
        RECT 670.020 3260.000 673.020 3547.300 ;
        RECT 850.020 3260.000 853.020 3547.300 ;
        RECT 1030.020 3260.000 1033.020 3547.300 ;
        RECT 1210.020 3260.000 1213.020 3547.300 ;
        RECT 1390.020 3260.000 1393.020 3547.300 ;
        RECT 1570.020 3260.000 1573.020 3547.300 ;
        RECT 1750.020 3260.000 1753.020 3547.300 ;
        RECT 1930.020 3260.000 1933.020 3547.300 ;
        RECT 2110.020 3260.000 2113.020 3547.300 ;
        RECT 2290.020 3260.000 2293.020 3547.300 ;
        RECT 2470.020 3260.000 2473.020 3547.300 ;
        RECT 310.020 -27.620 313.020 260.000 ;
        RECT 490.020 -27.620 493.020 260.000 ;
        RECT 670.020 -27.620 673.020 260.000 ;
        RECT 850.020 -27.620 853.020 260.000 ;
        RECT 1030.020 -27.620 1033.020 260.000 ;
        RECT 1210.020 -27.620 1213.020 260.000 ;
        RECT 1390.020 -27.620 1393.020 260.000 ;
        RECT 1570.020 -27.620 1573.020 260.000 ;
        RECT 1750.020 -27.620 1753.020 260.000 ;
        RECT 1930.020 -27.620 1933.020 260.000 ;
        RECT 2110.020 -27.620 2113.020 260.000 ;
        RECT 2290.020 -27.620 2293.020 260.000 ;
        RECT 2470.020 -27.620 2473.020 260.000 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 3260.000 421.020 3556.500 ;
        RECT 598.020 3260.000 601.020 3556.500 ;
        RECT 778.020 3260.000 781.020 3556.500 ;
        RECT 958.020 3260.000 961.020 3556.500 ;
        RECT 1138.020 3260.000 1141.020 3556.500 ;
        RECT 1318.020 3260.000 1321.020 3556.500 ;
        RECT 1498.020 3260.000 1501.020 3556.500 ;
        RECT 1678.020 3260.000 1681.020 3556.500 ;
        RECT 1858.020 3260.000 1861.020 3556.500 ;
        RECT 2038.020 3260.000 2041.020 3556.500 ;
        RECT 2218.020 3260.000 2221.020 3556.500 ;
        RECT 2398.020 3260.000 2401.020 3556.500 ;
        RECT 2578.020 3260.000 2581.020 3556.500 ;
        RECT 418.020 -36.820 421.020 260.000 ;
        RECT 598.020 -36.820 601.020 260.000 ;
        RECT 778.020 -36.820 781.020 260.000 ;
        RECT 958.020 -36.820 961.020 260.000 ;
        RECT 1138.020 -36.820 1141.020 260.000 ;
        RECT 1318.020 -36.820 1321.020 260.000 ;
        RECT 1498.020 -36.820 1501.020 260.000 ;
        RECT 1678.020 -36.820 1681.020 260.000 ;
        RECT 1858.020 -36.820 1861.020 260.000 ;
        RECT 2038.020 -36.820 2041.020 260.000 ;
        RECT 2218.020 -36.820 2221.020 260.000 ;
        RECT 2398.020 -36.820 2401.020 260.000 ;
        RECT 2578.020 -36.820 2581.020 260.000 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 3260.000 331.020 3556.500 ;
        RECT 508.020 3260.000 511.020 3556.500 ;
        RECT 688.020 3260.000 691.020 3556.500 ;
        RECT 868.020 3260.000 871.020 3556.500 ;
        RECT 1048.020 3260.000 1051.020 3556.500 ;
        RECT 1228.020 3260.000 1231.020 3556.500 ;
        RECT 1408.020 3260.000 1411.020 3556.500 ;
        RECT 1588.020 3260.000 1591.020 3556.500 ;
        RECT 1768.020 3260.000 1771.020 3556.500 ;
        RECT 1948.020 3260.000 1951.020 3556.500 ;
        RECT 2128.020 3260.000 2131.020 3556.500 ;
        RECT 2308.020 3260.000 2311.020 3556.500 ;
        RECT 2488.020 3260.000 2491.020 3556.500 ;
        RECT 328.020 -36.820 331.020 260.000 ;
        RECT 508.020 -36.820 511.020 260.000 ;
        RECT 688.020 -36.820 691.020 260.000 ;
        RECT 868.020 -36.820 871.020 260.000 ;
        RECT 1048.020 -36.820 1051.020 260.000 ;
        RECT 1228.020 -36.820 1231.020 260.000 ;
        RECT 1408.020 -36.820 1411.020 260.000 ;
        RECT 1588.020 -36.820 1591.020 260.000 ;
        RECT 1768.020 -36.820 1771.020 260.000 ;
        RECT 1948.020 -36.820 1951.020 260.000 ;
        RECT 2128.020 -36.820 2131.020 260.000 ;
        RECT 2308.020 -36.820 2311.020 260.000 ;
        RECT 2488.020 -36.820 2491.020 260.000 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 315.520 270.795 2604.480 3246.645 ;
      LAYER met1 ;
        RECT 312.370 269.900 2604.480 3246.800 ;
      LAYER met2 ;
        RECT 312.400 3255.720 352.130 3256.000 ;
        RECT 352.970 3255.720 437.230 3256.000 ;
        RECT 438.070 3255.720 522.330 3256.000 ;
        RECT 523.170 3255.720 607.430 3256.000 ;
        RECT 608.270 3255.720 692.530 3256.000 ;
        RECT 693.370 3255.720 777.630 3256.000 ;
        RECT 778.470 3255.720 863.190 3256.000 ;
        RECT 864.030 3255.720 948.290 3256.000 ;
        RECT 949.130 3255.720 1033.390 3256.000 ;
        RECT 1034.230 3255.720 1118.490 3256.000 ;
        RECT 1119.330 3255.720 1203.590 3256.000 ;
        RECT 1204.430 3255.720 1289.150 3256.000 ;
        RECT 1289.990 3255.720 1374.250 3256.000 ;
        RECT 1375.090 3255.720 1459.350 3256.000 ;
        RECT 1460.190 3255.720 1544.450 3256.000 ;
        RECT 1545.290 3255.720 1629.550 3256.000 ;
        RECT 1630.390 3255.720 1714.650 3256.000 ;
        RECT 1715.490 3255.720 1800.210 3256.000 ;
        RECT 1801.050 3255.720 1885.310 3256.000 ;
        RECT 1886.150 3255.720 1970.410 3256.000 ;
        RECT 1971.250 3255.720 2055.510 3256.000 ;
        RECT 2056.350 3255.720 2140.610 3256.000 ;
        RECT 2141.450 3255.720 2226.170 3256.000 ;
        RECT 2227.010 3255.720 2311.270 3256.000 ;
        RECT 2312.110 3255.720 2396.370 3256.000 ;
        RECT 2397.210 3255.720 2481.470 3256.000 ;
        RECT 2482.310 3255.720 2566.570 3256.000 ;
        RECT 2567.410 3255.720 2603.000 3256.000 ;
        RECT 312.400 264.280 2603.000 3255.720 ;
        RECT 312.950 264.000 316.710 264.280 ;
        RECT 317.550 264.000 321.310 264.280 ;
        RECT 322.150 264.000 325.910 264.280 ;
        RECT 326.750 264.000 330.510 264.280 ;
        RECT 331.350 264.000 335.570 264.280 ;
        RECT 336.410 264.000 340.170 264.280 ;
        RECT 341.010 264.000 344.770 264.280 ;
        RECT 345.610 264.000 349.370 264.280 ;
        RECT 350.210 264.000 353.970 264.280 ;
        RECT 354.810 264.000 359.030 264.280 ;
        RECT 359.870 264.000 363.630 264.280 ;
        RECT 364.470 264.000 368.230 264.280 ;
        RECT 369.070 264.000 372.830 264.280 ;
        RECT 373.670 264.000 377.430 264.280 ;
        RECT 378.270 264.000 382.490 264.280 ;
        RECT 383.330 264.000 387.090 264.280 ;
        RECT 387.930 264.000 391.690 264.280 ;
        RECT 392.530 264.000 396.290 264.280 ;
        RECT 397.130 264.000 400.890 264.280 ;
        RECT 401.730 264.000 405.950 264.280 ;
        RECT 406.790 264.000 410.550 264.280 ;
        RECT 411.390 264.000 415.150 264.280 ;
        RECT 415.990 264.000 419.750 264.280 ;
        RECT 420.590 264.000 424.350 264.280 ;
        RECT 425.190 264.000 429.410 264.280 ;
        RECT 430.250 264.000 434.010 264.280 ;
        RECT 434.850 264.000 438.610 264.280 ;
        RECT 439.450 264.000 443.210 264.280 ;
        RECT 444.050 264.000 447.810 264.280 ;
        RECT 448.650 264.000 452.870 264.280 ;
        RECT 453.710 264.000 457.470 264.280 ;
        RECT 458.310 264.000 462.070 264.280 ;
        RECT 462.910 264.000 466.670 264.280 ;
        RECT 467.510 264.000 471.270 264.280 ;
        RECT 472.110 264.000 476.330 264.280 ;
        RECT 477.170 264.000 480.930 264.280 ;
        RECT 481.770 264.000 485.530 264.280 ;
        RECT 486.370 264.000 490.130 264.280 ;
        RECT 490.970 264.000 494.730 264.280 ;
        RECT 495.570 264.000 499.790 264.280 ;
        RECT 500.630 264.000 504.390 264.280 ;
        RECT 505.230 264.000 508.990 264.280 ;
        RECT 509.830 264.000 513.590 264.280 ;
        RECT 514.430 264.000 518.190 264.280 ;
        RECT 519.030 264.000 523.250 264.280 ;
        RECT 524.090 264.000 527.850 264.280 ;
        RECT 528.690 264.000 532.450 264.280 ;
        RECT 533.290 264.000 537.050 264.280 ;
        RECT 537.890 264.000 542.110 264.280 ;
        RECT 542.950 264.000 546.710 264.280 ;
        RECT 547.550 264.000 551.310 264.280 ;
        RECT 552.150 264.000 555.910 264.280 ;
        RECT 556.750 264.000 560.510 264.280 ;
        RECT 561.350 264.000 565.570 264.280 ;
        RECT 566.410 264.000 570.170 264.280 ;
        RECT 571.010 264.000 574.770 264.280 ;
        RECT 575.610 264.000 579.370 264.280 ;
        RECT 580.210 264.000 583.970 264.280 ;
        RECT 584.810 264.000 589.030 264.280 ;
        RECT 589.870 264.000 593.630 264.280 ;
        RECT 594.470 264.000 598.230 264.280 ;
        RECT 599.070 264.000 602.830 264.280 ;
        RECT 603.670 264.000 607.430 264.280 ;
        RECT 608.270 264.000 612.490 264.280 ;
        RECT 613.330 264.000 617.090 264.280 ;
        RECT 617.930 264.000 621.690 264.280 ;
        RECT 622.530 264.000 626.290 264.280 ;
        RECT 627.130 264.000 630.890 264.280 ;
        RECT 631.730 264.000 635.950 264.280 ;
        RECT 636.790 264.000 640.550 264.280 ;
        RECT 641.390 264.000 645.150 264.280 ;
        RECT 645.990 264.000 649.750 264.280 ;
        RECT 650.590 264.000 654.350 264.280 ;
        RECT 655.190 264.000 659.410 264.280 ;
        RECT 660.250 264.000 664.010 264.280 ;
        RECT 664.850 264.000 668.610 264.280 ;
        RECT 669.450 264.000 673.210 264.280 ;
        RECT 674.050 264.000 677.810 264.280 ;
        RECT 678.650 264.000 682.870 264.280 ;
        RECT 683.710 264.000 687.470 264.280 ;
        RECT 688.310 264.000 692.070 264.280 ;
        RECT 692.910 264.000 696.670 264.280 ;
        RECT 697.510 264.000 701.270 264.280 ;
        RECT 702.110 264.000 706.330 264.280 ;
        RECT 707.170 264.000 710.930 264.280 ;
        RECT 711.770 264.000 715.530 264.280 ;
        RECT 716.370 264.000 720.130 264.280 ;
        RECT 720.970 264.000 724.730 264.280 ;
        RECT 725.570 264.000 729.790 264.280 ;
        RECT 730.630 264.000 734.390 264.280 ;
        RECT 735.230 264.000 738.990 264.280 ;
        RECT 739.830 264.000 743.590 264.280 ;
        RECT 744.430 264.000 748.190 264.280 ;
        RECT 749.030 264.000 753.250 264.280 ;
        RECT 754.090 264.000 757.850 264.280 ;
        RECT 758.690 264.000 762.450 264.280 ;
        RECT 763.290 264.000 767.050 264.280 ;
        RECT 767.890 264.000 772.110 264.280 ;
        RECT 772.950 264.000 776.710 264.280 ;
        RECT 777.550 264.000 781.310 264.280 ;
        RECT 782.150 264.000 785.910 264.280 ;
        RECT 786.750 264.000 790.510 264.280 ;
        RECT 791.350 264.000 795.570 264.280 ;
        RECT 796.410 264.000 800.170 264.280 ;
        RECT 801.010 264.000 804.770 264.280 ;
        RECT 805.610 264.000 809.370 264.280 ;
        RECT 810.210 264.000 813.970 264.280 ;
        RECT 814.810 264.000 819.030 264.280 ;
        RECT 819.870 264.000 823.630 264.280 ;
        RECT 824.470 264.000 828.230 264.280 ;
        RECT 829.070 264.000 832.830 264.280 ;
        RECT 833.670 264.000 837.430 264.280 ;
        RECT 838.270 264.000 842.490 264.280 ;
        RECT 843.330 264.000 847.090 264.280 ;
        RECT 847.930 264.000 851.690 264.280 ;
        RECT 852.530 264.000 856.290 264.280 ;
        RECT 857.130 264.000 860.890 264.280 ;
        RECT 861.730 264.000 865.950 264.280 ;
        RECT 866.790 264.000 870.550 264.280 ;
        RECT 871.390 264.000 875.150 264.280 ;
        RECT 875.990 264.000 879.750 264.280 ;
        RECT 880.590 264.000 884.350 264.280 ;
        RECT 885.190 264.000 889.410 264.280 ;
        RECT 890.250 264.000 894.010 264.280 ;
        RECT 894.850 264.000 898.610 264.280 ;
        RECT 899.450 264.000 903.210 264.280 ;
        RECT 904.050 264.000 907.810 264.280 ;
        RECT 908.650 264.000 912.870 264.280 ;
        RECT 913.710 264.000 917.470 264.280 ;
        RECT 918.310 264.000 922.070 264.280 ;
        RECT 922.910 264.000 926.670 264.280 ;
        RECT 927.510 264.000 931.270 264.280 ;
        RECT 932.110 264.000 936.330 264.280 ;
        RECT 937.170 264.000 940.930 264.280 ;
        RECT 941.770 264.000 945.530 264.280 ;
        RECT 946.370 264.000 950.130 264.280 ;
        RECT 950.970 264.000 954.730 264.280 ;
        RECT 955.570 264.000 959.790 264.280 ;
        RECT 960.630 264.000 964.390 264.280 ;
        RECT 965.230 264.000 968.990 264.280 ;
        RECT 969.830 264.000 973.590 264.280 ;
        RECT 974.430 264.000 978.190 264.280 ;
        RECT 979.030 264.000 983.250 264.280 ;
        RECT 984.090 264.000 987.850 264.280 ;
        RECT 988.690 264.000 992.450 264.280 ;
        RECT 993.290 264.000 997.050 264.280 ;
        RECT 997.890 264.000 1002.110 264.280 ;
        RECT 1002.950 264.000 1006.710 264.280 ;
        RECT 1007.550 264.000 1011.310 264.280 ;
        RECT 1012.150 264.000 1015.910 264.280 ;
        RECT 1016.750 264.000 1020.510 264.280 ;
        RECT 1021.350 264.000 1025.570 264.280 ;
        RECT 1026.410 264.000 1030.170 264.280 ;
        RECT 1031.010 264.000 1034.770 264.280 ;
        RECT 1035.610 264.000 1039.370 264.280 ;
        RECT 1040.210 264.000 1043.970 264.280 ;
        RECT 1044.810 264.000 1049.030 264.280 ;
        RECT 1049.870 264.000 1053.630 264.280 ;
        RECT 1054.470 264.000 1058.230 264.280 ;
        RECT 1059.070 264.000 1062.830 264.280 ;
        RECT 1063.670 264.000 1067.430 264.280 ;
        RECT 1068.270 264.000 1072.490 264.280 ;
        RECT 1073.330 264.000 1077.090 264.280 ;
        RECT 1077.930 264.000 1081.690 264.280 ;
        RECT 1082.530 264.000 1086.290 264.280 ;
        RECT 1087.130 264.000 1090.890 264.280 ;
        RECT 1091.730 264.000 1095.950 264.280 ;
        RECT 1096.790 264.000 1100.550 264.280 ;
        RECT 1101.390 264.000 1105.150 264.280 ;
        RECT 1105.990 264.000 1109.750 264.280 ;
        RECT 1110.590 264.000 1114.350 264.280 ;
        RECT 1115.190 264.000 1119.410 264.280 ;
        RECT 1120.250 264.000 1124.010 264.280 ;
        RECT 1124.850 264.000 1128.610 264.280 ;
        RECT 1129.450 264.000 1133.210 264.280 ;
        RECT 1134.050 264.000 1137.810 264.280 ;
        RECT 1138.650 264.000 1142.870 264.280 ;
        RECT 1143.710 264.000 1147.470 264.280 ;
        RECT 1148.310 264.000 1152.070 264.280 ;
        RECT 1152.910 264.000 1156.670 264.280 ;
        RECT 1157.510 264.000 1161.270 264.280 ;
        RECT 1162.110 264.000 1166.330 264.280 ;
        RECT 1167.170 264.000 1170.930 264.280 ;
        RECT 1171.770 264.000 1175.530 264.280 ;
        RECT 1176.370 264.000 1180.130 264.280 ;
        RECT 1180.970 264.000 1184.730 264.280 ;
        RECT 1185.570 264.000 1189.790 264.280 ;
        RECT 1190.630 264.000 1194.390 264.280 ;
        RECT 1195.230 264.000 1198.990 264.280 ;
        RECT 1199.830 264.000 1203.590 264.280 ;
        RECT 1204.430 264.000 1208.190 264.280 ;
        RECT 1209.030 264.000 1213.250 264.280 ;
        RECT 1214.090 264.000 1217.850 264.280 ;
        RECT 1218.690 264.000 1222.450 264.280 ;
        RECT 1223.290 264.000 1227.050 264.280 ;
        RECT 1227.890 264.000 1232.110 264.280 ;
        RECT 1232.950 264.000 1236.710 264.280 ;
        RECT 1237.550 264.000 1241.310 264.280 ;
        RECT 1242.150 264.000 1245.910 264.280 ;
        RECT 1246.750 264.000 1250.510 264.280 ;
        RECT 1251.350 264.000 1255.570 264.280 ;
        RECT 1256.410 264.000 1260.170 264.280 ;
        RECT 1261.010 264.000 1264.770 264.280 ;
        RECT 1265.610 264.000 1269.370 264.280 ;
        RECT 1270.210 264.000 1273.970 264.280 ;
        RECT 1274.810 264.000 1279.030 264.280 ;
        RECT 1279.870 264.000 1283.630 264.280 ;
        RECT 1284.470 264.000 1288.230 264.280 ;
        RECT 1289.070 264.000 1292.830 264.280 ;
        RECT 1293.670 264.000 1297.430 264.280 ;
        RECT 1298.270 264.000 1302.490 264.280 ;
        RECT 1303.330 264.000 1307.090 264.280 ;
        RECT 1307.930 264.000 1311.690 264.280 ;
        RECT 1312.530 264.000 1316.290 264.280 ;
        RECT 1317.130 264.000 1320.890 264.280 ;
        RECT 1321.730 264.000 1325.950 264.280 ;
        RECT 1326.790 264.000 1330.550 264.280 ;
        RECT 1331.390 264.000 1335.150 264.280 ;
        RECT 1335.990 264.000 1339.750 264.280 ;
        RECT 1340.590 264.000 1344.350 264.280 ;
        RECT 1345.190 264.000 1349.410 264.280 ;
        RECT 1350.250 264.000 1354.010 264.280 ;
        RECT 1354.850 264.000 1358.610 264.280 ;
        RECT 1359.450 264.000 1363.210 264.280 ;
        RECT 1364.050 264.000 1367.810 264.280 ;
        RECT 1368.650 264.000 1372.870 264.280 ;
        RECT 1373.710 264.000 1377.470 264.280 ;
        RECT 1378.310 264.000 1382.070 264.280 ;
        RECT 1382.910 264.000 1386.670 264.280 ;
        RECT 1387.510 264.000 1391.270 264.280 ;
        RECT 1392.110 264.000 1396.330 264.280 ;
        RECT 1397.170 264.000 1400.930 264.280 ;
        RECT 1401.770 264.000 1405.530 264.280 ;
        RECT 1406.370 264.000 1410.130 264.280 ;
        RECT 1410.970 264.000 1414.730 264.280 ;
        RECT 1415.570 264.000 1419.790 264.280 ;
        RECT 1420.630 264.000 1424.390 264.280 ;
        RECT 1425.230 264.000 1428.990 264.280 ;
        RECT 1429.830 264.000 1433.590 264.280 ;
        RECT 1434.430 264.000 1438.190 264.280 ;
        RECT 1439.030 264.000 1443.250 264.280 ;
        RECT 1444.090 264.000 1447.850 264.280 ;
        RECT 1448.690 264.000 1452.450 264.280 ;
        RECT 1453.290 264.000 1457.050 264.280 ;
        RECT 1457.890 264.000 1462.110 264.280 ;
        RECT 1462.950 264.000 1466.710 264.280 ;
        RECT 1467.550 264.000 1471.310 264.280 ;
        RECT 1472.150 264.000 1475.910 264.280 ;
        RECT 1476.750 264.000 1480.510 264.280 ;
        RECT 1481.350 264.000 1485.570 264.280 ;
        RECT 1486.410 264.000 1490.170 264.280 ;
        RECT 1491.010 264.000 1494.770 264.280 ;
        RECT 1495.610 264.000 1499.370 264.280 ;
        RECT 1500.210 264.000 1503.970 264.280 ;
        RECT 1504.810 264.000 1509.030 264.280 ;
        RECT 1509.870 264.000 1513.630 264.280 ;
        RECT 1514.470 264.000 1518.230 264.280 ;
        RECT 1519.070 264.000 1522.830 264.280 ;
        RECT 1523.670 264.000 1527.430 264.280 ;
        RECT 1528.270 264.000 1532.490 264.280 ;
        RECT 1533.330 264.000 1537.090 264.280 ;
        RECT 1537.930 264.000 1541.690 264.280 ;
        RECT 1542.530 264.000 1546.290 264.280 ;
        RECT 1547.130 264.000 1550.890 264.280 ;
        RECT 1551.730 264.000 1555.950 264.280 ;
        RECT 1556.790 264.000 1560.550 264.280 ;
        RECT 1561.390 264.000 1565.150 264.280 ;
        RECT 1565.990 264.000 1569.750 264.280 ;
        RECT 1570.590 264.000 1574.350 264.280 ;
        RECT 1575.190 264.000 1579.410 264.280 ;
        RECT 1580.250 264.000 1584.010 264.280 ;
        RECT 1584.850 264.000 1588.610 264.280 ;
        RECT 1589.450 264.000 1593.210 264.280 ;
        RECT 1594.050 264.000 1597.810 264.280 ;
        RECT 1598.650 264.000 1602.870 264.280 ;
        RECT 1603.710 264.000 1607.470 264.280 ;
        RECT 1608.310 264.000 1612.070 264.280 ;
        RECT 1612.910 264.000 1616.670 264.280 ;
        RECT 1617.510 264.000 1621.270 264.280 ;
        RECT 1622.110 264.000 1626.330 264.280 ;
        RECT 1627.170 264.000 1630.930 264.280 ;
        RECT 1631.770 264.000 1635.530 264.280 ;
        RECT 1636.370 264.000 1640.130 264.280 ;
        RECT 1640.970 264.000 1644.730 264.280 ;
        RECT 1645.570 264.000 1649.790 264.280 ;
        RECT 1650.630 264.000 1654.390 264.280 ;
        RECT 1655.230 264.000 1658.990 264.280 ;
        RECT 1659.830 264.000 1663.590 264.280 ;
        RECT 1664.430 264.000 1668.190 264.280 ;
        RECT 1669.030 264.000 1673.250 264.280 ;
        RECT 1674.090 264.000 1677.850 264.280 ;
        RECT 1678.690 264.000 1682.450 264.280 ;
        RECT 1683.290 264.000 1687.050 264.280 ;
        RECT 1687.890 264.000 1692.110 264.280 ;
        RECT 1692.950 264.000 1696.710 264.280 ;
        RECT 1697.550 264.000 1701.310 264.280 ;
        RECT 1702.150 264.000 1705.910 264.280 ;
        RECT 1706.750 264.000 1710.510 264.280 ;
        RECT 1711.350 264.000 1715.570 264.280 ;
        RECT 1716.410 264.000 1720.170 264.280 ;
        RECT 1721.010 264.000 1724.770 264.280 ;
        RECT 1725.610 264.000 1729.370 264.280 ;
        RECT 1730.210 264.000 1733.970 264.280 ;
        RECT 1734.810 264.000 1739.030 264.280 ;
        RECT 1739.870 264.000 1743.630 264.280 ;
        RECT 1744.470 264.000 1748.230 264.280 ;
        RECT 1749.070 264.000 1752.830 264.280 ;
        RECT 1753.670 264.000 1757.430 264.280 ;
        RECT 1758.270 264.000 1762.490 264.280 ;
        RECT 1763.330 264.000 1767.090 264.280 ;
        RECT 1767.930 264.000 1771.690 264.280 ;
        RECT 1772.530 264.000 1776.290 264.280 ;
        RECT 1777.130 264.000 1780.890 264.280 ;
        RECT 1781.730 264.000 1785.950 264.280 ;
        RECT 1786.790 264.000 1790.550 264.280 ;
        RECT 1791.390 264.000 1795.150 264.280 ;
        RECT 1795.990 264.000 1799.750 264.280 ;
        RECT 1800.590 264.000 1804.350 264.280 ;
        RECT 1805.190 264.000 1809.410 264.280 ;
        RECT 1810.250 264.000 1814.010 264.280 ;
        RECT 1814.850 264.000 1818.610 264.280 ;
        RECT 1819.450 264.000 1823.210 264.280 ;
        RECT 1824.050 264.000 1827.810 264.280 ;
        RECT 1828.650 264.000 1832.870 264.280 ;
        RECT 1833.710 264.000 1837.470 264.280 ;
        RECT 1838.310 264.000 1842.070 264.280 ;
        RECT 1842.910 264.000 1846.670 264.280 ;
        RECT 1847.510 264.000 1851.270 264.280 ;
        RECT 1852.110 264.000 1856.330 264.280 ;
        RECT 1857.170 264.000 1860.930 264.280 ;
        RECT 1861.770 264.000 1865.530 264.280 ;
        RECT 1866.370 264.000 1870.130 264.280 ;
        RECT 1870.970 264.000 1874.730 264.280 ;
        RECT 1875.570 264.000 1879.790 264.280 ;
        RECT 1880.630 264.000 1884.390 264.280 ;
        RECT 1885.230 264.000 1888.990 264.280 ;
        RECT 1889.830 264.000 1893.590 264.280 ;
        RECT 1894.430 264.000 1898.190 264.280 ;
        RECT 1899.030 264.000 1903.250 264.280 ;
        RECT 1904.090 264.000 1907.850 264.280 ;
        RECT 1908.690 264.000 1912.450 264.280 ;
        RECT 1913.290 264.000 1917.050 264.280 ;
        RECT 1917.890 264.000 1922.110 264.280 ;
        RECT 1922.950 264.000 1926.710 264.280 ;
        RECT 1927.550 264.000 1931.310 264.280 ;
        RECT 1932.150 264.000 1935.910 264.280 ;
        RECT 1936.750 264.000 1940.510 264.280 ;
        RECT 1941.350 264.000 1945.570 264.280 ;
        RECT 1946.410 264.000 1950.170 264.280 ;
        RECT 1951.010 264.000 1954.770 264.280 ;
        RECT 1955.610 264.000 1959.370 264.280 ;
        RECT 1960.210 264.000 1963.970 264.280 ;
        RECT 1964.810 264.000 1969.030 264.280 ;
        RECT 1969.870 264.000 1973.630 264.280 ;
        RECT 1974.470 264.000 1978.230 264.280 ;
        RECT 1979.070 264.000 1982.830 264.280 ;
        RECT 1983.670 264.000 1987.430 264.280 ;
        RECT 1988.270 264.000 1992.490 264.280 ;
        RECT 1993.330 264.000 1997.090 264.280 ;
        RECT 1997.930 264.000 2001.690 264.280 ;
        RECT 2002.530 264.000 2006.290 264.280 ;
        RECT 2007.130 264.000 2010.890 264.280 ;
        RECT 2011.730 264.000 2015.950 264.280 ;
        RECT 2016.790 264.000 2020.550 264.280 ;
        RECT 2021.390 264.000 2025.150 264.280 ;
        RECT 2025.990 264.000 2029.750 264.280 ;
        RECT 2030.590 264.000 2034.350 264.280 ;
        RECT 2035.190 264.000 2039.410 264.280 ;
        RECT 2040.250 264.000 2044.010 264.280 ;
        RECT 2044.850 264.000 2048.610 264.280 ;
        RECT 2049.450 264.000 2053.210 264.280 ;
        RECT 2054.050 264.000 2057.810 264.280 ;
        RECT 2058.650 264.000 2062.870 264.280 ;
        RECT 2063.710 264.000 2067.470 264.280 ;
        RECT 2068.310 264.000 2072.070 264.280 ;
        RECT 2072.910 264.000 2076.670 264.280 ;
        RECT 2077.510 264.000 2081.270 264.280 ;
        RECT 2082.110 264.000 2086.330 264.280 ;
        RECT 2087.170 264.000 2090.930 264.280 ;
        RECT 2091.770 264.000 2095.530 264.280 ;
        RECT 2096.370 264.000 2100.130 264.280 ;
        RECT 2100.970 264.000 2104.730 264.280 ;
        RECT 2105.570 264.000 2109.790 264.280 ;
        RECT 2110.630 264.000 2114.390 264.280 ;
        RECT 2115.230 264.000 2118.990 264.280 ;
        RECT 2119.830 264.000 2123.590 264.280 ;
        RECT 2124.430 264.000 2128.190 264.280 ;
        RECT 2129.030 264.000 2133.250 264.280 ;
        RECT 2134.090 264.000 2137.850 264.280 ;
        RECT 2138.690 264.000 2142.450 264.280 ;
        RECT 2143.290 264.000 2147.050 264.280 ;
        RECT 2147.890 264.000 2152.110 264.280 ;
        RECT 2152.950 264.000 2156.710 264.280 ;
        RECT 2157.550 264.000 2161.310 264.280 ;
        RECT 2162.150 264.000 2165.910 264.280 ;
        RECT 2166.750 264.000 2170.510 264.280 ;
        RECT 2171.350 264.000 2175.570 264.280 ;
        RECT 2176.410 264.000 2180.170 264.280 ;
        RECT 2181.010 264.000 2184.770 264.280 ;
        RECT 2185.610 264.000 2189.370 264.280 ;
        RECT 2190.210 264.000 2193.970 264.280 ;
        RECT 2194.810 264.000 2199.030 264.280 ;
        RECT 2199.870 264.000 2203.630 264.280 ;
        RECT 2204.470 264.000 2208.230 264.280 ;
        RECT 2209.070 264.000 2212.830 264.280 ;
        RECT 2213.670 264.000 2217.430 264.280 ;
        RECT 2218.270 264.000 2222.490 264.280 ;
        RECT 2223.330 264.000 2227.090 264.280 ;
        RECT 2227.930 264.000 2231.690 264.280 ;
        RECT 2232.530 264.000 2236.290 264.280 ;
        RECT 2237.130 264.000 2240.890 264.280 ;
        RECT 2241.730 264.000 2245.950 264.280 ;
        RECT 2246.790 264.000 2250.550 264.280 ;
        RECT 2251.390 264.000 2255.150 264.280 ;
        RECT 2255.990 264.000 2259.750 264.280 ;
        RECT 2260.590 264.000 2264.350 264.280 ;
        RECT 2265.190 264.000 2269.410 264.280 ;
        RECT 2270.250 264.000 2274.010 264.280 ;
        RECT 2274.850 264.000 2278.610 264.280 ;
        RECT 2279.450 264.000 2283.210 264.280 ;
        RECT 2284.050 264.000 2287.810 264.280 ;
        RECT 2288.650 264.000 2292.870 264.280 ;
        RECT 2293.710 264.000 2297.470 264.280 ;
        RECT 2298.310 264.000 2302.070 264.280 ;
        RECT 2302.910 264.000 2306.670 264.280 ;
        RECT 2307.510 264.000 2311.270 264.280 ;
        RECT 2312.110 264.000 2316.330 264.280 ;
        RECT 2317.170 264.000 2320.930 264.280 ;
        RECT 2321.770 264.000 2325.530 264.280 ;
        RECT 2326.370 264.000 2330.130 264.280 ;
        RECT 2330.970 264.000 2334.730 264.280 ;
        RECT 2335.570 264.000 2339.790 264.280 ;
        RECT 2340.630 264.000 2344.390 264.280 ;
        RECT 2345.230 264.000 2348.990 264.280 ;
        RECT 2349.830 264.000 2353.590 264.280 ;
        RECT 2354.430 264.000 2358.190 264.280 ;
        RECT 2359.030 264.000 2363.250 264.280 ;
        RECT 2364.090 264.000 2367.850 264.280 ;
        RECT 2368.690 264.000 2372.450 264.280 ;
        RECT 2373.290 264.000 2377.050 264.280 ;
        RECT 2377.890 264.000 2382.110 264.280 ;
        RECT 2382.950 264.000 2386.710 264.280 ;
        RECT 2387.550 264.000 2391.310 264.280 ;
        RECT 2392.150 264.000 2395.910 264.280 ;
        RECT 2396.750 264.000 2400.510 264.280 ;
        RECT 2401.350 264.000 2405.570 264.280 ;
        RECT 2406.410 264.000 2410.170 264.280 ;
        RECT 2411.010 264.000 2414.770 264.280 ;
        RECT 2415.610 264.000 2419.370 264.280 ;
        RECT 2420.210 264.000 2423.970 264.280 ;
        RECT 2424.810 264.000 2429.030 264.280 ;
        RECT 2429.870 264.000 2433.630 264.280 ;
        RECT 2434.470 264.000 2438.230 264.280 ;
        RECT 2439.070 264.000 2442.830 264.280 ;
        RECT 2443.670 264.000 2447.430 264.280 ;
        RECT 2448.270 264.000 2452.490 264.280 ;
        RECT 2453.330 264.000 2457.090 264.280 ;
        RECT 2457.930 264.000 2461.690 264.280 ;
        RECT 2462.530 264.000 2466.290 264.280 ;
        RECT 2467.130 264.000 2470.890 264.280 ;
        RECT 2471.730 264.000 2475.950 264.280 ;
        RECT 2476.790 264.000 2480.550 264.280 ;
        RECT 2481.390 264.000 2485.150 264.280 ;
        RECT 2485.990 264.000 2489.750 264.280 ;
        RECT 2490.590 264.000 2494.350 264.280 ;
        RECT 2495.190 264.000 2499.410 264.280 ;
        RECT 2500.250 264.000 2504.010 264.280 ;
        RECT 2504.850 264.000 2508.610 264.280 ;
        RECT 2509.450 264.000 2513.210 264.280 ;
        RECT 2514.050 264.000 2517.810 264.280 ;
        RECT 2518.650 264.000 2522.870 264.280 ;
        RECT 2523.710 264.000 2527.470 264.280 ;
        RECT 2528.310 264.000 2532.070 264.280 ;
        RECT 2532.910 264.000 2536.670 264.280 ;
        RECT 2537.510 264.000 2541.270 264.280 ;
        RECT 2542.110 264.000 2546.330 264.280 ;
        RECT 2547.170 264.000 2550.930 264.280 ;
        RECT 2551.770 264.000 2555.530 264.280 ;
        RECT 2556.370 264.000 2560.130 264.280 ;
        RECT 2560.970 264.000 2564.730 264.280 ;
        RECT 2565.570 264.000 2569.790 264.280 ;
        RECT 2570.630 264.000 2574.390 264.280 ;
        RECT 2575.230 264.000 2578.990 264.280 ;
        RECT 2579.830 264.000 2583.590 264.280 ;
        RECT 2584.430 264.000 2588.190 264.280 ;
        RECT 2589.030 264.000 2593.250 264.280 ;
        RECT 2594.090 264.000 2597.850 264.280 ;
        RECT 2598.690 264.000 2602.450 264.280 ;
      LAYER met3 ;
        RECT 314.000 3227.200 2606.010 3246.725 ;
        RECT 314.000 3225.800 2605.600 3227.200 ;
        RECT 314.000 3224.480 2606.010 3225.800 ;
        RECT 314.400 3223.080 2606.010 3224.480 ;
        RECT 314.000 3160.560 2606.010 3223.080 ;
        RECT 314.000 3159.160 2605.600 3160.560 ;
        RECT 314.000 3153.080 2606.010 3159.160 ;
        RECT 314.400 3151.680 2606.010 3153.080 ;
        RECT 314.000 3093.920 2606.010 3151.680 ;
        RECT 314.000 3092.520 2605.600 3093.920 ;
        RECT 314.000 3081.680 2606.010 3092.520 ;
        RECT 314.400 3080.280 2606.010 3081.680 ;
        RECT 314.000 3027.280 2606.010 3080.280 ;
        RECT 314.000 3025.880 2605.600 3027.280 ;
        RECT 314.000 3010.280 2606.010 3025.880 ;
        RECT 314.400 3008.880 2606.010 3010.280 ;
        RECT 314.000 2960.640 2606.010 3008.880 ;
        RECT 314.000 2959.240 2605.600 2960.640 ;
        RECT 314.000 2938.880 2606.010 2959.240 ;
        RECT 314.400 2937.480 2606.010 2938.880 ;
        RECT 314.000 2894.000 2606.010 2937.480 ;
        RECT 314.000 2892.600 2605.600 2894.000 ;
        RECT 314.000 2867.480 2606.010 2892.600 ;
        RECT 314.400 2866.080 2606.010 2867.480 ;
        RECT 314.000 2827.360 2606.010 2866.080 ;
        RECT 314.000 2825.960 2605.600 2827.360 ;
        RECT 314.000 2796.080 2606.010 2825.960 ;
        RECT 314.400 2794.680 2606.010 2796.080 ;
        RECT 314.000 2760.720 2606.010 2794.680 ;
        RECT 314.000 2759.320 2605.600 2760.720 ;
        RECT 314.000 2724.680 2606.010 2759.320 ;
        RECT 314.400 2723.280 2606.010 2724.680 ;
        RECT 314.000 2694.080 2606.010 2723.280 ;
        RECT 314.000 2692.680 2605.600 2694.080 ;
        RECT 314.000 2653.280 2606.010 2692.680 ;
        RECT 314.400 2651.880 2606.010 2653.280 ;
        RECT 314.000 2627.440 2606.010 2651.880 ;
        RECT 314.000 2626.040 2605.600 2627.440 ;
        RECT 314.000 2581.880 2606.010 2626.040 ;
        RECT 314.400 2580.480 2606.010 2581.880 ;
        RECT 314.000 2560.800 2606.010 2580.480 ;
        RECT 314.000 2559.400 2605.600 2560.800 ;
        RECT 314.000 2510.480 2606.010 2559.400 ;
        RECT 314.400 2509.080 2606.010 2510.480 ;
        RECT 314.000 2494.160 2606.010 2509.080 ;
        RECT 314.000 2492.760 2605.600 2494.160 ;
        RECT 314.000 2439.080 2606.010 2492.760 ;
        RECT 314.400 2437.680 2606.010 2439.080 ;
        RECT 314.000 2427.520 2606.010 2437.680 ;
        RECT 314.000 2426.120 2605.600 2427.520 ;
        RECT 314.000 2367.680 2606.010 2426.120 ;
        RECT 314.400 2366.280 2606.010 2367.680 ;
        RECT 314.000 2360.880 2606.010 2366.280 ;
        RECT 314.000 2359.480 2605.600 2360.880 ;
        RECT 314.000 2296.280 2606.010 2359.480 ;
        RECT 314.400 2294.880 2606.010 2296.280 ;
        RECT 314.000 2294.240 2606.010 2294.880 ;
        RECT 314.000 2292.840 2605.600 2294.240 ;
        RECT 314.000 2227.600 2606.010 2292.840 ;
        RECT 314.000 2226.200 2605.600 2227.600 ;
        RECT 314.000 2224.880 2606.010 2226.200 ;
        RECT 314.400 2223.480 2606.010 2224.880 ;
        RECT 314.000 2160.960 2606.010 2223.480 ;
        RECT 314.000 2159.560 2605.600 2160.960 ;
        RECT 314.000 2153.480 2606.010 2159.560 ;
        RECT 314.400 2152.080 2606.010 2153.480 ;
        RECT 314.000 2094.320 2606.010 2152.080 ;
        RECT 314.000 2092.920 2605.600 2094.320 ;
        RECT 314.000 2082.080 2606.010 2092.920 ;
        RECT 314.400 2080.680 2606.010 2082.080 ;
        RECT 314.000 2027.680 2606.010 2080.680 ;
        RECT 314.000 2026.280 2605.600 2027.680 ;
        RECT 314.000 2010.680 2606.010 2026.280 ;
        RECT 314.400 2009.280 2606.010 2010.680 ;
        RECT 314.000 1961.040 2606.010 2009.280 ;
        RECT 314.000 1959.640 2605.600 1961.040 ;
        RECT 314.000 1939.280 2606.010 1959.640 ;
        RECT 314.400 1937.880 2606.010 1939.280 ;
        RECT 314.000 1894.400 2606.010 1937.880 ;
        RECT 314.000 1893.000 2605.600 1894.400 ;
        RECT 314.000 1867.880 2606.010 1893.000 ;
        RECT 314.400 1866.480 2606.010 1867.880 ;
        RECT 314.000 1827.760 2606.010 1866.480 ;
        RECT 314.000 1826.360 2605.600 1827.760 ;
        RECT 314.000 1796.480 2606.010 1826.360 ;
        RECT 314.400 1795.080 2606.010 1796.480 ;
        RECT 314.000 1760.440 2606.010 1795.080 ;
        RECT 314.000 1759.040 2605.600 1760.440 ;
        RECT 314.000 1724.400 2606.010 1759.040 ;
        RECT 314.400 1723.000 2606.010 1724.400 ;
        RECT 314.000 1693.800 2606.010 1723.000 ;
        RECT 314.000 1692.400 2605.600 1693.800 ;
        RECT 314.000 1653.000 2606.010 1692.400 ;
        RECT 314.400 1651.600 2606.010 1653.000 ;
        RECT 314.000 1627.160 2606.010 1651.600 ;
        RECT 314.000 1625.760 2605.600 1627.160 ;
        RECT 314.000 1581.600 2606.010 1625.760 ;
        RECT 314.400 1580.200 2606.010 1581.600 ;
        RECT 314.000 1560.520 2606.010 1580.200 ;
        RECT 314.000 1559.120 2605.600 1560.520 ;
        RECT 314.000 1510.200 2606.010 1559.120 ;
        RECT 314.400 1508.800 2606.010 1510.200 ;
        RECT 314.000 1493.880 2606.010 1508.800 ;
        RECT 314.000 1492.480 2605.600 1493.880 ;
        RECT 314.000 1438.800 2606.010 1492.480 ;
        RECT 314.400 1437.400 2606.010 1438.800 ;
        RECT 314.000 1427.240 2606.010 1437.400 ;
        RECT 314.000 1425.840 2605.600 1427.240 ;
        RECT 314.000 1367.400 2606.010 1425.840 ;
        RECT 314.400 1366.000 2606.010 1367.400 ;
        RECT 314.000 1360.600 2606.010 1366.000 ;
        RECT 314.000 1359.200 2605.600 1360.600 ;
        RECT 314.000 1296.000 2606.010 1359.200 ;
        RECT 314.400 1294.600 2606.010 1296.000 ;
        RECT 314.000 1293.960 2606.010 1294.600 ;
        RECT 314.000 1292.560 2605.600 1293.960 ;
        RECT 314.000 1227.320 2606.010 1292.560 ;
        RECT 314.000 1225.920 2605.600 1227.320 ;
        RECT 314.000 1224.600 2606.010 1225.920 ;
        RECT 314.400 1223.200 2606.010 1224.600 ;
        RECT 314.000 1160.680 2606.010 1223.200 ;
        RECT 314.000 1159.280 2605.600 1160.680 ;
        RECT 314.000 1153.200 2606.010 1159.280 ;
        RECT 314.400 1151.800 2606.010 1153.200 ;
        RECT 314.000 1094.040 2606.010 1151.800 ;
        RECT 314.000 1092.640 2605.600 1094.040 ;
        RECT 314.000 1081.800 2606.010 1092.640 ;
        RECT 314.400 1080.400 2606.010 1081.800 ;
        RECT 314.000 1027.400 2606.010 1080.400 ;
        RECT 314.000 1026.000 2605.600 1027.400 ;
        RECT 314.000 1010.400 2606.010 1026.000 ;
        RECT 314.400 1009.000 2606.010 1010.400 ;
        RECT 314.000 960.760 2606.010 1009.000 ;
        RECT 314.000 959.360 2605.600 960.760 ;
        RECT 314.000 939.000 2606.010 959.360 ;
        RECT 314.400 937.600 2606.010 939.000 ;
        RECT 314.000 894.120 2606.010 937.600 ;
        RECT 314.000 892.720 2605.600 894.120 ;
        RECT 314.000 867.600 2606.010 892.720 ;
        RECT 314.400 866.200 2606.010 867.600 ;
        RECT 314.000 827.480 2606.010 866.200 ;
        RECT 314.000 826.080 2605.600 827.480 ;
        RECT 314.000 796.200 2606.010 826.080 ;
        RECT 314.400 794.800 2606.010 796.200 ;
        RECT 314.000 760.840 2606.010 794.800 ;
        RECT 314.000 759.440 2605.600 760.840 ;
        RECT 314.000 724.800 2606.010 759.440 ;
        RECT 314.400 723.400 2606.010 724.800 ;
        RECT 314.000 694.200 2606.010 723.400 ;
        RECT 314.000 692.800 2605.600 694.200 ;
        RECT 314.000 653.400 2606.010 692.800 ;
        RECT 314.400 652.000 2606.010 653.400 ;
        RECT 314.000 627.560 2606.010 652.000 ;
        RECT 314.000 626.160 2605.600 627.560 ;
        RECT 314.000 582.000 2606.010 626.160 ;
        RECT 314.400 580.600 2606.010 582.000 ;
        RECT 314.000 560.920 2606.010 580.600 ;
        RECT 314.000 559.520 2605.600 560.920 ;
        RECT 314.000 510.600 2606.010 559.520 ;
        RECT 314.400 509.200 2606.010 510.600 ;
        RECT 314.000 494.280 2606.010 509.200 ;
        RECT 314.000 492.880 2605.600 494.280 ;
        RECT 314.000 439.200 2606.010 492.880 ;
        RECT 314.400 437.800 2606.010 439.200 ;
        RECT 314.000 427.640 2606.010 437.800 ;
        RECT 314.000 426.240 2605.600 427.640 ;
        RECT 314.000 367.800 2606.010 426.240 ;
        RECT 314.400 366.400 2606.010 367.800 ;
        RECT 314.000 361.000 2606.010 366.400 ;
        RECT 314.000 359.600 2605.600 361.000 ;
        RECT 314.000 296.400 2606.010 359.600 ;
        RECT 314.400 295.000 2606.010 296.400 ;
        RECT 314.000 294.360 2606.010 295.000 ;
        RECT 314.000 292.960 2605.600 294.360 ;
        RECT 314.000 270.715 2606.010 292.960 ;
      LAYER met4 ;
        RECT 325.935 270.640 330.640 3246.800 ;
      LAYER met4 ;
        RECT 331.040 270.640 332.640 3246.800 ;
      LAYER met4 ;
        RECT 333.040 270.640 407.440 3246.800 ;
      LAYER met4 ;
        RECT 407.840 270.640 409.440 3246.800 ;
      LAYER met4 ;
        RECT 409.840 270.640 2590.385 3246.800 ;
  END
END user_project_wrapper
END LIBRARY

