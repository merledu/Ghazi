VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 379.110 36.620 379.430 36.680 ;
        RECT 400.730 36.620 401.050 36.680 ;
        RECT 379.110 36.480 401.050 36.620 ;
        RECT 379.110 36.420 379.430 36.480 ;
        RECT 400.730 36.420 401.050 36.480 ;
        RECT 414.070 36.620 414.390 36.680 ;
        RECT 461.450 36.620 461.770 36.680 ;
        RECT 414.070 36.480 461.770 36.620 ;
        RECT 414.070 36.420 414.390 36.480 ;
        RECT 461.450 36.420 461.770 36.480 ;
        RECT 800.470 36.620 800.790 36.680 ;
        RECT 847.850 36.620 848.170 36.680 ;
        RECT 800.470 36.480 848.170 36.620 ;
        RECT 800.470 36.420 800.790 36.480 ;
        RECT 847.850 36.420 848.170 36.480 ;
        RECT 2028.670 36.620 2028.990 36.680 ;
        RECT 2053.050 36.620 2053.370 36.680 ;
        RECT 2028.670 36.480 2053.370 36.620 ;
        RECT 2028.670 36.420 2028.990 36.480 ;
        RECT 2053.050 36.420 2053.370 36.480 ;
        RECT 2525.010 36.620 2525.330 36.680 ;
        RECT 2552.610 36.620 2552.930 36.680 ;
        RECT 2525.010 36.480 2552.930 36.620 ;
        RECT 2525.010 36.420 2525.330 36.480 ;
        RECT 2552.610 36.420 2552.930 36.480 ;
        RECT 2608.730 36.620 2609.050 36.680 ;
        RECT 2697.510 36.620 2697.830 36.680 ;
        RECT 2608.730 36.480 2697.830 36.620 ;
        RECT 2608.730 36.420 2609.050 36.480 ;
        RECT 2697.510 36.420 2697.830 36.480 ;
        RECT 2238.890 36.280 2239.210 36.340 ;
        RECT 2262.810 36.280 2263.130 36.340 ;
        RECT 2238.890 36.140 2263.130 36.280 ;
        RECT 2238.890 36.080 2239.210 36.140 ;
        RECT 2262.810 36.080 2263.130 36.140 ;
        RECT 2318.930 36.280 2319.250 36.340 ;
        RECT 2365.850 36.280 2366.170 36.340 ;
        RECT 2318.930 36.140 2366.170 36.280 ;
        RECT 2318.930 36.080 2319.250 36.140 ;
        RECT 2365.850 36.080 2366.170 36.140 ;
        RECT 753.550 35.940 753.870 36.000 ;
        RECT 787.130 35.940 787.450 36.000 ;
        RECT 753.550 35.800 787.450 35.940 ;
        RECT 753.550 35.740 753.870 35.800 ;
        RECT 787.130 35.740 787.450 35.800 ;
        RECT 868.550 35.940 868.870 36.000 ;
        RECT 872.690 35.940 873.010 36.000 ;
        RECT 868.550 35.800 873.010 35.940 ;
        RECT 868.550 35.740 868.870 35.800 ;
        RECT 872.690 35.740 873.010 35.800 ;
        RECT 1531.870 35.940 1532.190 36.000 ;
        RECT 1579.710 35.940 1580.030 36.000 ;
        RECT 1531.870 35.800 1580.030 35.940 ;
        RECT 1531.870 35.740 1532.190 35.800 ;
        RECT 1579.710 35.740 1580.030 35.800 ;
        RECT 511.130 35.600 511.450 35.660 ;
        RECT 558.050 35.600 558.370 35.660 ;
        RECT 511.130 35.460 558.370 35.600 ;
        RECT 511.130 35.400 511.450 35.460 ;
        RECT 558.050 35.400 558.370 35.460 ;
        RECT 2787.670 35.600 2787.990 35.660 ;
        RECT 2816.190 35.600 2816.510 35.660 ;
        RECT 2787.670 35.460 2816.510 35.600 ;
        RECT 2787.670 35.400 2787.990 35.460 ;
        RECT 2816.190 35.400 2816.510 35.460 ;
        RECT 607.270 35.260 607.590 35.320 ;
        RECT 655.110 35.260 655.430 35.320 ;
        RECT 607.270 35.120 655.430 35.260 ;
        RECT 607.270 35.060 607.590 35.120 ;
        RECT 655.110 35.060 655.430 35.120 ;
      LAYER via ;
        RECT 379.140 36.420 379.400 36.680 ;
        RECT 400.760 36.420 401.020 36.680 ;
        RECT 414.100 36.420 414.360 36.680 ;
        RECT 461.480 36.420 461.740 36.680 ;
        RECT 800.500 36.420 800.760 36.680 ;
        RECT 847.880 36.420 848.140 36.680 ;
        RECT 2028.700 36.420 2028.960 36.680 ;
        RECT 2053.080 36.420 2053.340 36.680 ;
        RECT 2525.040 36.420 2525.300 36.680 ;
        RECT 2552.640 36.420 2552.900 36.680 ;
        RECT 2608.760 36.420 2609.020 36.680 ;
        RECT 2697.540 36.420 2697.800 36.680 ;
        RECT 2238.920 36.080 2239.180 36.340 ;
        RECT 2262.840 36.080 2263.100 36.340 ;
        RECT 2318.960 36.080 2319.220 36.340 ;
        RECT 2365.880 36.080 2366.140 36.340 ;
        RECT 753.580 35.740 753.840 36.000 ;
        RECT 787.160 35.740 787.420 36.000 ;
        RECT 868.580 35.740 868.840 36.000 ;
        RECT 872.720 35.740 872.980 36.000 ;
        RECT 1531.900 35.740 1532.160 36.000 ;
        RECT 1579.740 35.740 1580.000 36.000 ;
        RECT 511.160 35.400 511.420 35.660 ;
        RECT 558.080 35.400 558.340 35.660 ;
        RECT 2787.700 35.400 2787.960 35.660 ;
        RECT 2816.220 35.400 2816.480 35.660 ;
        RECT 607.300 35.060 607.560 35.320 ;
        RECT 655.140 35.060 655.400 35.320 ;
      LAYER met2 ;
        RECT 296.790 3159.435 297.070 3159.805 ;
        RECT 296.860 3153.685 297.000 3159.435 ;
        RECT 296.790 3153.315 297.070 3153.685 ;
        RECT 1222.310 38.235 1222.590 38.605 ;
        RECT 1314.310 38.235 1314.590 38.605 ;
        RECT 606.370 36.875 606.650 37.245 ;
        RECT 717.230 36.875 717.510 37.245 ;
        RECT 379.140 36.565 379.400 36.710 ;
        RECT 400.760 36.565 401.020 36.710 ;
        RECT 414.100 36.565 414.360 36.710 ;
        RECT 461.480 36.565 461.740 36.710 ;
        RECT 379.130 36.195 379.410 36.565 ;
        RECT 400.750 36.195 401.030 36.565 ;
        RECT 414.090 36.195 414.370 36.565 ;
        RECT 461.470 36.195 461.750 36.565 ;
        RECT 495.970 36.450 496.250 36.565 ;
        RECT 496.890 36.450 497.170 36.565 ;
        RECT 495.970 36.310 497.170 36.450 ;
        RECT 495.970 36.195 496.250 36.310 ;
        RECT 496.890 36.195 497.170 36.310 ;
        RECT 511.150 35.515 511.430 35.885 ;
        RECT 558.070 35.515 558.350 35.885 ;
        RECT 511.160 35.370 511.420 35.515 ;
        RECT 558.080 35.370 558.340 35.515 ;
        RECT 606.440 35.205 606.580 36.875 ;
        RECT 717.300 35.885 717.440 36.875 ;
        RECT 800.500 36.565 800.760 36.710 ;
        RECT 847.880 36.565 848.140 36.710 ;
        RECT 787.150 36.195 787.430 36.565 ;
        RECT 800.490 36.195 800.770 36.565 ;
        RECT 847.870 36.195 848.150 36.565 ;
        RECT 868.570 36.195 868.850 36.565 ;
        RECT 787.220 36.030 787.360 36.195 ;
        RECT 868.640 36.030 868.780 36.195 ;
        RECT 655.130 35.515 655.410 35.885 ;
        RECT 717.230 35.515 717.510 35.885 ;
        RECT 753.580 35.710 753.840 36.030 ;
        RECT 787.160 35.710 787.420 36.030 ;
        RECT 868.580 35.710 868.840 36.030 ;
        RECT 872.720 35.710 872.980 36.030 ;
        RECT 1222.380 35.885 1222.520 38.235 ;
        RECT 1283.030 36.875 1283.310 37.245 ;
        RECT 1283.100 35.885 1283.240 36.875 ;
        RECT 1314.380 36.565 1314.520 38.235 ;
        RECT 1410.910 37.555 1411.190 37.925 ;
        RECT 2142.310 37.555 2142.590 37.925 ;
        RECT 2238.910 37.555 2239.190 37.925 ;
        RECT 1410.980 36.565 1411.120 37.555 ;
        RECT 2028.700 36.565 2028.960 36.710 ;
        RECT 2053.080 36.565 2053.340 36.710 ;
        RECT 1314.310 36.195 1314.590 36.565 ;
        RECT 1410.910 36.195 1411.190 36.565 ;
        RECT 1496.930 36.195 1497.210 36.565 ;
        RECT 1579.730 36.195 1580.010 36.565 ;
        RECT 1587.550 36.195 1587.830 36.565 ;
        RECT 2028.690 36.195 2028.970 36.565 ;
        RECT 2053.070 36.195 2053.350 36.565 ;
        RECT 655.200 35.350 655.340 35.515 ;
        RECT 607.300 35.205 607.560 35.350 ;
        RECT 606.370 34.835 606.650 35.205 ;
        RECT 607.290 34.835 607.570 35.205 ;
        RECT 655.140 35.030 655.400 35.350 ;
        RECT 753.640 35.205 753.780 35.710 ;
        RECT 872.780 35.205 872.920 35.710 ;
        RECT 1222.310 35.515 1222.590 35.885 ;
        RECT 1283.030 35.515 1283.310 35.885 ;
        RECT 1497.000 35.770 1497.140 36.195 ;
        RECT 1579.800 36.030 1579.940 36.195 ;
        RECT 1531.900 35.885 1532.160 36.030 ;
        RECT 1497.850 35.770 1498.130 35.885 ;
        RECT 1497.000 35.630 1498.130 35.770 ;
        RECT 1497.850 35.515 1498.130 35.630 ;
        RECT 1531.890 35.515 1532.170 35.885 ;
        RECT 1579.740 35.710 1580.000 36.030 ;
        RECT 1587.620 35.205 1587.760 36.195 ;
        RECT 2142.380 35.885 2142.520 37.555 ;
        RECT 2174.050 36.195 2174.330 36.565 ;
        RECT 2238.980 36.370 2239.120 37.555 ;
        RECT 2270.650 37.130 2270.930 37.245 ;
        RECT 2270.260 36.990 2270.930 37.130 ;
        RECT 2270.260 36.565 2270.400 36.990 ;
        RECT 2270.650 36.875 2270.930 36.990 ;
        RECT 2697.530 36.875 2697.810 37.245 ;
        RECT 2883.830 36.875 2884.110 37.245 ;
        RECT 2697.600 36.710 2697.740 36.875 ;
        RECT 2525.040 36.565 2525.300 36.710 ;
        RECT 2552.640 36.565 2552.900 36.710 ;
        RECT 2608.760 36.565 2609.020 36.710 ;
        RECT 2142.310 35.515 2142.590 35.885 ;
        RECT 2174.120 35.205 2174.260 36.195 ;
        RECT 2238.920 36.050 2239.180 36.370 ;
        RECT 2262.830 36.195 2263.110 36.565 ;
        RECT 2270.190 36.195 2270.470 36.565 ;
        RECT 2318.950 36.195 2319.230 36.565 ;
        RECT 2365.870 36.195 2366.150 36.565 ;
        RECT 2525.030 36.195 2525.310 36.565 ;
        RECT 2552.630 36.195 2552.910 36.565 ;
        RECT 2608.750 36.195 2609.030 36.565 ;
        RECT 2697.540 36.390 2697.800 36.710 ;
        RECT 2262.840 36.050 2263.100 36.195 ;
        RECT 2318.960 36.050 2319.220 36.195 ;
        RECT 2365.880 36.050 2366.140 36.195 ;
        RECT 2883.900 35.885 2884.040 36.875 ;
        RECT 2787.690 35.515 2787.970 35.885 ;
        RECT 2787.700 35.370 2787.960 35.515 ;
        RECT 2816.220 35.370 2816.480 35.690 ;
        RECT 2883.830 35.515 2884.110 35.885 ;
        RECT 2816.280 35.205 2816.420 35.370 ;
        RECT 753.570 34.835 753.850 35.205 ;
        RECT 872.710 34.835 872.990 35.205 ;
        RECT 1587.550 34.835 1587.830 35.205 ;
        RECT 2174.050 34.835 2174.330 35.205 ;
        RECT 2816.210 34.835 2816.490 35.205 ;
      LAYER via2 ;
        RECT 296.790 3159.480 297.070 3159.760 ;
        RECT 296.790 3153.360 297.070 3153.640 ;
        RECT 1222.310 38.280 1222.590 38.560 ;
        RECT 1314.310 38.280 1314.590 38.560 ;
        RECT 606.370 36.920 606.650 37.200 ;
        RECT 717.230 36.920 717.510 37.200 ;
        RECT 379.130 36.240 379.410 36.520 ;
        RECT 400.750 36.240 401.030 36.520 ;
        RECT 414.090 36.240 414.370 36.520 ;
        RECT 461.470 36.240 461.750 36.520 ;
        RECT 495.970 36.240 496.250 36.520 ;
        RECT 496.890 36.240 497.170 36.520 ;
        RECT 511.150 35.560 511.430 35.840 ;
        RECT 558.070 35.560 558.350 35.840 ;
        RECT 787.150 36.240 787.430 36.520 ;
        RECT 800.490 36.240 800.770 36.520 ;
        RECT 847.870 36.240 848.150 36.520 ;
        RECT 868.570 36.240 868.850 36.520 ;
        RECT 655.130 35.560 655.410 35.840 ;
        RECT 717.230 35.560 717.510 35.840 ;
        RECT 1283.030 36.920 1283.310 37.200 ;
        RECT 1410.910 37.600 1411.190 37.880 ;
        RECT 2142.310 37.600 2142.590 37.880 ;
        RECT 2238.910 37.600 2239.190 37.880 ;
        RECT 1314.310 36.240 1314.590 36.520 ;
        RECT 1410.910 36.240 1411.190 36.520 ;
        RECT 1496.930 36.240 1497.210 36.520 ;
        RECT 1579.730 36.240 1580.010 36.520 ;
        RECT 1587.550 36.240 1587.830 36.520 ;
        RECT 2028.690 36.240 2028.970 36.520 ;
        RECT 2053.070 36.240 2053.350 36.520 ;
        RECT 606.370 34.880 606.650 35.160 ;
        RECT 607.290 34.880 607.570 35.160 ;
        RECT 1222.310 35.560 1222.590 35.840 ;
        RECT 1283.030 35.560 1283.310 35.840 ;
        RECT 1497.850 35.560 1498.130 35.840 ;
        RECT 1531.890 35.560 1532.170 35.840 ;
        RECT 2174.050 36.240 2174.330 36.520 ;
        RECT 2270.650 36.920 2270.930 37.200 ;
        RECT 2697.530 36.920 2697.810 37.200 ;
        RECT 2883.830 36.920 2884.110 37.200 ;
        RECT 2142.310 35.560 2142.590 35.840 ;
        RECT 2262.830 36.240 2263.110 36.520 ;
        RECT 2270.190 36.240 2270.470 36.520 ;
        RECT 2318.950 36.240 2319.230 36.520 ;
        RECT 2365.870 36.240 2366.150 36.520 ;
        RECT 2525.030 36.240 2525.310 36.520 ;
        RECT 2552.630 36.240 2552.910 36.520 ;
        RECT 2608.750 36.240 2609.030 36.520 ;
        RECT 2787.690 35.560 2787.970 35.840 ;
        RECT 2883.830 35.560 2884.110 35.840 ;
        RECT 753.570 34.880 753.850 35.160 ;
        RECT 872.710 34.880 872.990 35.160 ;
        RECT 1587.550 34.880 1587.830 35.160 ;
        RECT 2174.050 34.880 2174.330 35.160 ;
        RECT 2816.210 34.880 2816.490 35.160 ;
      LAYER met3 ;
        RECT 296.765 3159.770 297.095 3159.785 ;
        RECT 310.000 3159.770 314.000 3160.160 ;
        RECT 296.765 3159.560 314.000 3159.770 ;
        RECT 296.765 3159.470 310.500 3159.560 ;
        RECT 296.765 3159.455 297.095 3159.470 ;
        RECT 261.550 3153.650 261.930 3153.660 ;
        RECT 296.765 3153.650 297.095 3153.665 ;
        RECT 261.550 3153.350 297.095 3153.650 ;
        RECT 261.550 3153.340 261.930 3153.350 ;
        RECT 296.765 3153.335 297.095 3153.350 ;
        RECT 2917.600 39.250 2924.800 39.700 ;
        RECT 2916.940 38.950 2924.800 39.250 ;
        RECT 1222.285 38.570 1222.615 38.585 ;
        RECT 1193.550 38.270 1222.615 38.570 ;
        RECT 663.590 37.890 663.970 37.900 ;
        RECT 663.590 37.590 669.450 37.890 ;
        RECT 663.590 37.580 663.970 37.590 ;
        RECT 558.710 37.210 559.090 37.220 ;
        RECT 606.345 37.210 606.675 37.225 ;
        RECT 558.710 36.910 606.675 37.210 ;
        RECT 669.150 37.210 669.450 37.590 ;
        RECT 717.205 37.210 717.535 37.225 ;
        RECT 1055.510 37.210 1055.890 37.220 ;
        RECT 1110.710 37.210 1111.090 37.220 ;
        RECT 1193.550 37.210 1193.850 38.270 ;
        RECT 1222.285 38.255 1222.615 38.270 ;
        RECT 1290.110 38.570 1290.490 38.580 ;
        RECT 1314.285 38.570 1314.615 38.585 ;
        RECT 1290.110 38.270 1314.615 38.570 ;
        RECT 1290.110 38.260 1290.490 38.270 ;
        RECT 1314.285 38.255 1314.615 38.270 ;
        RECT 1386.710 37.890 1387.090 37.900 ;
        RECT 1410.885 37.890 1411.215 37.905 ;
        RECT 1386.710 37.590 1411.215 37.890 ;
        RECT 1386.710 37.580 1387.090 37.590 ;
        RECT 1410.885 37.575 1411.215 37.590 ;
        RECT 2118.110 37.890 2118.490 37.900 ;
        RECT 2142.285 37.890 2142.615 37.905 ;
        RECT 2118.110 37.590 2142.615 37.890 ;
        RECT 2118.110 37.580 2118.490 37.590 ;
        RECT 2142.285 37.575 2142.615 37.590 ;
        RECT 2214.710 37.890 2215.090 37.900 ;
        RECT 2238.885 37.890 2239.215 37.905 ;
        RECT 2214.710 37.590 2239.215 37.890 ;
        RECT 2214.710 37.580 2215.090 37.590 ;
        RECT 2238.885 37.575 2239.215 37.590 ;
        RECT 2366.510 37.890 2366.890 37.900 ;
        RECT 2455.750 37.890 2456.130 37.900 ;
        RECT 2366.510 37.590 2456.130 37.890 ;
        RECT 2366.510 37.580 2366.890 37.590 ;
        RECT 2455.750 37.580 2456.130 37.590 ;
        RECT 669.150 36.910 717.535 37.210 ;
        RECT 558.710 36.900 559.090 36.910 ;
        RECT 606.345 36.895 606.675 36.910 ;
        RECT 717.205 36.895 717.535 36.910 ;
        RECT 903.750 36.910 951.890 37.210 ;
        RECT 261.550 36.530 261.930 36.540 ;
        RECT 379.105 36.530 379.435 36.545 ;
        RECT 261.550 36.230 379.435 36.530 ;
        RECT 261.550 36.220 261.930 36.230 ;
        RECT 379.105 36.215 379.435 36.230 ;
        RECT 400.725 36.530 401.055 36.545 ;
        RECT 414.065 36.530 414.395 36.545 ;
        RECT 400.725 36.230 414.395 36.530 ;
        RECT 400.725 36.215 401.055 36.230 ;
        RECT 414.065 36.215 414.395 36.230 ;
        RECT 461.445 36.530 461.775 36.545 ;
        RECT 495.945 36.530 496.275 36.545 ;
        RECT 461.445 36.230 496.275 36.530 ;
        RECT 461.445 36.215 461.775 36.230 ;
        RECT 495.945 36.215 496.275 36.230 ;
        RECT 496.865 36.530 497.195 36.545 ;
        RECT 787.125 36.530 787.455 36.545 ;
        RECT 800.465 36.530 800.795 36.545 ;
        RECT 496.865 36.230 510.290 36.530 ;
        RECT 496.865 36.215 497.195 36.230 ;
        RECT 509.990 35.850 510.290 36.230 ;
        RECT 787.125 36.230 800.795 36.530 ;
        RECT 787.125 36.215 787.455 36.230 ;
        RECT 800.465 36.215 800.795 36.230 ;
        RECT 847.845 36.530 848.175 36.545 ;
        RECT 868.545 36.530 868.875 36.545 ;
        RECT 847.845 36.230 868.875 36.530 ;
        RECT 847.845 36.215 848.175 36.230 ;
        RECT 868.545 36.215 868.875 36.230 ;
        RECT 511.125 35.850 511.455 35.865 ;
        RECT 509.990 35.550 511.455 35.850 ;
        RECT 511.125 35.535 511.455 35.550 ;
        RECT 558.045 35.850 558.375 35.865 ;
        RECT 558.710 35.850 559.090 35.860 ;
        RECT 558.045 35.550 559.090 35.850 ;
        RECT 558.045 35.535 558.375 35.550 ;
        RECT 558.710 35.540 559.090 35.550 ;
        RECT 655.105 35.850 655.435 35.865 ;
        RECT 662.670 35.850 663.050 35.860 ;
        RECT 655.105 35.550 663.050 35.850 ;
        RECT 655.105 35.535 655.435 35.550 ;
        RECT 662.670 35.540 663.050 35.550 ;
        RECT 717.205 35.850 717.535 35.865 ;
        RECT 717.205 35.550 718.210 35.850 ;
        RECT 717.205 35.535 717.535 35.550 ;
        RECT 606.345 35.170 606.675 35.185 ;
        RECT 607.265 35.170 607.595 35.185 ;
        RECT 606.345 34.870 607.595 35.170 ;
        RECT 717.910 35.170 718.210 35.550 ;
        RECT 753.545 35.170 753.875 35.185 ;
        RECT 717.910 34.870 753.875 35.170 ;
        RECT 606.345 34.855 606.675 34.870 ;
        RECT 607.265 34.855 607.595 34.870 ;
        RECT 753.545 34.855 753.875 34.870 ;
        RECT 872.685 35.170 873.015 35.185 ;
        RECT 903.750 35.170 904.050 36.910 ;
        RECT 951.590 35.850 951.890 36.910 ;
        RECT 1055.510 36.910 1103.690 37.210 ;
        RECT 1055.510 36.900 1055.890 36.910 ;
        RECT 1055.510 35.850 1055.890 35.860 ;
        RECT 951.590 35.550 1055.890 35.850 ;
        RECT 1055.510 35.540 1055.890 35.550 ;
        RECT 872.685 34.870 904.050 35.170 ;
        RECT 1103.390 35.170 1103.690 36.910 ;
        RECT 1110.710 36.910 1193.850 37.210 ;
        RECT 1234.910 37.210 1235.290 37.220 ;
        RECT 1283.005 37.210 1283.335 37.225 ;
        RECT 1234.910 36.910 1283.335 37.210 ;
        RECT 1110.710 36.900 1111.090 36.910 ;
        RECT 1234.910 36.900 1235.290 36.910 ;
        RECT 1283.005 36.895 1283.335 36.910 ;
        RECT 2270.625 37.210 2270.955 37.225 ;
        RECT 2697.505 37.210 2697.835 37.225 ;
        RECT 2835.710 37.210 2836.090 37.220 ;
        RECT 2883.805 37.210 2884.135 37.225 ;
        RECT 2270.625 36.910 2318.090 37.210 ;
        RECT 2697.100 36.910 2698.050 37.210 ;
        RECT 2270.625 36.895 2270.955 36.910 ;
        RECT 1290.110 36.220 1290.490 36.540 ;
        RECT 1314.285 36.530 1314.615 36.545 ;
        RECT 1386.710 36.530 1387.090 36.540 ;
        RECT 1314.285 36.230 1387.090 36.530 ;
        RECT 1222.285 35.850 1222.615 35.865 ;
        RECT 1234.910 35.850 1235.290 35.860 ;
        RECT 1222.285 35.550 1235.290 35.850 ;
        RECT 1222.285 35.535 1222.615 35.550 ;
        RECT 1234.910 35.540 1235.290 35.550 ;
        RECT 1283.005 35.850 1283.335 35.865 ;
        RECT 1290.150 35.850 1290.450 36.220 ;
        RECT 1314.285 36.215 1314.615 36.230 ;
        RECT 1386.710 36.220 1387.090 36.230 ;
        RECT 1410.885 36.530 1411.215 36.545 ;
        RECT 1442.830 36.530 1443.210 36.540 ;
        RECT 1496.905 36.530 1497.235 36.545 ;
        RECT 1410.885 36.230 1434.890 36.530 ;
        RECT 1410.885 36.215 1411.215 36.230 ;
        RECT 1283.005 35.550 1290.450 35.850 ;
        RECT 1434.590 35.850 1434.890 36.230 ;
        RECT 1442.830 36.230 1497.235 36.530 ;
        RECT 1442.830 36.220 1443.210 36.230 ;
        RECT 1496.905 36.215 1497.235 36.230 ;
        RECT 1579.705 36.530 1580.035 36.545 ;
        RECT 1587.525 36.530 1587.855 36.545 ;
        RECT 1981.030 36.530 1981.410 36.540 ;
        RECT 2028.665 36.530 2028.995 36.545 ;
        RECT 1579.705 36.230 1587.855 36.530 ;
        RECT 1579.705 36.215 1580.035 36.230 ;
        RECT 1587.525 36.215 1587.855 36.230 ;
        RECT 1731.750 36.230 1732.970 36.530 ;
        RECT 1441.910 35.850 1442.290 35.860 ;
        RECT 1434.590 35.550 1442.290 35.850 ;
        RECT 1283.005 35.535 1283.335 35.550 ;
        RECT 1441.910 35.540 1442.290 35.550 ;
        RECT 1497.825 35.850 1498.155 35.865 ;
        RECT 1531.865 35.850 1532.195 35.865 ;
        RECT 1497.825 35.550 1532.195 35.850 ;
        RECT 1497.825 35.535 1498.155 35.550 ;
        RECT 1531.865 35.535 1532.195 35.550 ;
        RECT 1110.710 35.170 1111.090 35.180 ;
        RECT 1103.390 34.870 1111.090 35.170 ;
        RECT 872.685 34.855 873.015 34.870 ;
        RECT 1110.710 34.860 1111.090 34.870 ;
        RECT 1587.525 35.170 1587.855 35.185 ;
        RECT 1731.750 35.170 1732.050 36.230 ;
        RECT 1732.670 35.850 1732.970 36.230 ;
        RECT 1981.030 36.230 2028.995 36.530 ;
        RECT 1981.030 36.220 1981.410 36.230 ;
        RECT 2028.665 36.215 2028.995 36.230 ;
        RECT 2053.045 36.530 2053.375 36.545 ;
        RECT 2118.110 36.530 2118.490 36.540 ;
        RECT 2053.045 36.230 2118.490 36.530 ;
        RECT 2053.045 36.215 2053.375 36.230 ;
        RECT 2118.110 36.220 2118.490 36.230 ;
        RECT 2174.025 36.530 2174.355 36.545 ;
        RECT 2214.710 36.530 2215.090 36.540 ;
        RECT 2174.025 36.230 2215.090 36.530 ;
        RECT 2174.025 36.215 2174.355 36.230 ;
        RECT 2214.710 36.220 2215.090 36.230 ;
        RECT 2262.805 36.530 2263.135 36.545 ;
        RECT 2270.165 36.530 2270.495 36.545 ;
        RECT 2262.805 36.230 2270.495 36.530 ;
        RECT 2317.790 36.530 2318.090 36.910 ;
        RECT 2697.505 36.895 2698.050 36.910 ;
        RECT 2835.710 36.910 2884.135 37.210 ;
        RECT 2835.710 36.900 2836.090 36.910 ;
        RECT 2883.805 36.895 2884.135 36.910 ;
        RECT 2318.925 36.530 2319.255 36.545 ;
        RECT 2317.790 36.230 2319.255 36.530 ;
        RECT 2262.805 36.215 2263.135 36.230 ;
        RECT 2270.165 36.215 2270.495 36.230 ;
        RECT 2318.925 36.215 2319.255 36.230 ;
        RECT 2365.845 36.530 2366.175 36.545 ;
        RECT 2366.510 36.530 2366.890 36.540 ;
        RECT 2365.845 36.230 2366.890 36.530 ;
        RECT 2365.845 36.215 2366.175 36.230 ;
        RECT 2366.510 36.220 2366.890 36.230 ;
        RECT 2456.670 36.530 2457.050 36.540 ;
        RECT 2525.005 36.530 2525.335 36.545 ;
        RECT 2456.670 36.230 2525.335 36.530 ;
        RECT 2456.670 36.220 2457.050 36.230 ;
        RECT 2525.005 36.215 2525.335 36.230 ;
        RECT 2552.605 36.530 2552.935 36.545 ;
        RECT 2608.725 36.530 2609.055 36.545 ;
        RECT 2552.605 36.230 2609.055 36.530 ;
        RECT 2552.605 36.215 2552.935 36.230 ;
        RECT 2608.725 36.215 2609.055 36.230 ;
        RECT 1786.910 35.850 1787.290 35.860 ;
        RECT 1980.110 35.850 1980.490 35.860 ;
        RECT 1732.670 35.550 1787.290 35.850 ;
        RECT 1786.910 35.540 1787.290 35.550 ;
        RECT 1834.790 35.550 1980.490 35.850 ;
        RECT 1587.525 34.870 1732.050 35.170 ;
        RECT 1787.830 35.170 1788.210 35.180 ;
        RECT 1834.790 35.170 1835.090 35.550 ;
        RECT 1980.110 35.540 1980.490 35.550 ;
        RECT 2142.285 35.850 2142.615 35.865 ;
        RECT 2697.750 35.850 2698.050 36.895 ;
        RECT 2916.940 36.530 2917.240 38.950 ;
        RECT 2917.600 38.500 2924.800 38.950 ;
        RECT 2897.390 36.230 2917.240 36.530 ;
        RECT 2787.665 35.850 2787.995 35.865 ;
        RECT 2142.285 35.550 2166.290 35.850 ;
        RECT 2697.750 35.550 2719.210 35.850 ;
        RECT 2142.285 35.535 2142.615 35.550 ;
        RECT 1787.830 34.870 1835.090 35.170 ;
        RECT 2165.990 35.170 2166.290 35.550 ;
        RECT 2174.025 35.170 2174.355 35.185 ;
        RECT 2165.990 34.870 2174.355 35.170 ;
        RECT 2718.910 35.170 2719.210 35.550 ;
        RECT 2745.590 35.550 2787.995 35.850 ;
        RECT 2745.590 35.170 2745.890 35.550 ;
        RECT 2787.665 35.535 2787.995 35.550 ;
        RECT 2883.805 35.850 2884.135 35.865 ;
        RECT 2897.390 35.850 2897.690 36.230 ;
        RECT 2883.805 35.550 2897.690 35.850 ;
        RECT 2883.805 35.535 2884.135 35.550 ;
        RECT 2718.910 34.870 2745.890 35.170 ;
        RECT 2816.185 35.170 2816.515 35.185 ;
        RECT 2835.710 35.170 2836.090 35.180 ;
        RECT 2816.185 34.870 2836.090 35.170 ;
        RECT 1587.525 34.855 1587.855 34.870 ;
        RECT 1787.830 34.860 1788.210 34.870 ;
        RECT 2174.025 34.855 2174.355 34.870 ;
        RECT 2816.185 34.855 2816.515 34.870 ;
        RECT 2835.710 34.860 2836.090 34.870 ;
      LAYER via3 ;
        RECT 261.580 3153.340 261.900 3153.660 ;
        RECT 663.620 37.580 663.940 37.900 ;
        RECT 558.740 36.900 559.060 37.220 ;
        RECT 261.580 36.220 261.900 36.540 ;
        RECT 558.740 35.540 559.060 35.860 ;
        RECT 662.700 35.540 663.020 35.860 ;
        RECT 1055.540 36.900 1055.860 37.220 ;
        RECT 1055.540 35.540 1055.860 35.860 ;
        RECT 1110.740 36.900 1111.060 37.220 ;
        RECT 1290.140 38.260 1290.460 38.580 ;
        RECT 1386.740 37.580 1387.060 37.900 ;
        RECT 2118.140 37.580 2118.460 37.900 ;
        RECT 2214.740 37.580 2215.060 37.900 ;
        RECT 2366.540 37.580 2366.860 37.900 ;
        RECT 2455.780 37.580 2456.100 37.900 ;
        RECT 1234.940 36.900 1235.260 37.220 ;
        RECT 1290.140 36.220 1290.460 36.540 ;
        RECT 1234.940 35.540 1235.260 35.860 ;
        RECT 1386.740 36.220 1387.060 36.540 ;
        RECT 1442.860 36.220 1443.180 36.540 ;
        RECT 1441.940 35.540 1442.260 35.860 ;
        RECT 1110.740 34.860 1111.060 35.180 ;
        RECT 1981.060 36.220 1981.380 36.540 ;
        RECT 2118.140 36.220 2118.460 36.540 ;
        RECT 2214.740 36.220 2215.060 36.540 ;
        RECT 2835.740 36.900 2836.060 37.220 ;
        RECT 2366.540 36.220 2366.860 36.540 ;
        RECT 2456.700 36.220 2457.020 36.540 ;
        RECT 1786.940 35.540 1787.260 35.860 ;
        RECT 1787.860 34.860 1788.180 35.180 ;
        RECT 1980.140 35.540 1980.460 35.860 ;
        RECT 2835.740 34.860 2836.060 35.180 ;
      LAYER met4 ;
        RECT 261.575 3153.335 261.905 3153.665 ;
        RECT 261.590 36.545 261.890 3153.335 ;
        RECT 1290.135 38.255 1290.465 38.585 ;
        RECT 663.615 37.575 663.945 37.905 ;
        RECT 558.735 36.895 559.065 37.225 ;
        RECT 261.575 36.215 261.905 36.545 ;
        RECT 558.750 35.865 559.050 36.895 ;
        RECT 558.735 35.535 559.065 35.865 ;
        RECT 662.695 35.850 663.025 35.865 ;
        RECT 663.630 35.850 663.930 37.575 ;
        RECT 1055.535 36.895 1055.865 37.225 ;
        RECT 1110.735 36.895 1111.065 37.225 ;
        RECT 1234.935 36.895 1235.265 37.225 ;
        RECT 1055.550 35.865 1055.850 36.895 ;
        RECT 662.695 35.550 663.930 35.850 ;
        RECT 662.695 35.535 663.025 35.550 ;
        RECT 1055.535 35.535 1055.865 35.865 ;
        RECT 1110.750 35.185 1111.050 36.895 ;
        RECT 1234.950 35.865 1235.250 36.895 ;
        RECT 1290.150 36.545 1290.450 38.255 ;
        RECT 1386.735 37.575 1387.065 37.905 ;
        RECT 2118.135 37.575 2118.465 37.905 ;
        RECT 2214.735 37.575 2215.065 37.905 ;
        RECT 2366.535 37.575 2366.865 37.905 ;
        RECT 2455.775 37.575 2456.105 37.905 ;
        RECT 1386.750 36.545 1387.050 37.575 ;
        RECT 2118.150 36.545 2118.450 37.575 ;
        RECT 2214.750 36.545 2215.050 37.575 ;
        RECT 2366.550 36.545 2366.850 37.575 ;
        RECT 1290.135 36.215 1290.465 36.545 ;
        RECT 1386.735 36.215 1387.065 36.545 ;
        RECT 1442.855 36.215 1443.185 36.545 ;
        RECT 1981.055 36.215 1981.385 36.545 ;
        RECT 2118.135 36.215 2118.465 36.545 ;
        RECT 2214.735 36.215 2215.065 36.545 ;
        RECT 2366.535 36.215 2366.865 36.545 ;
        RECT 1234.935 35.535 1235.265 35.865 ;
        RECT 1441.935 35.850 1442.265 35.865 ;
        RECT 1442.870 35.850 1443.170 36.215 ;
        RECT 1441.935 35.550 1443.170 35.850 ;
        RECT 1786.935 35.850 1787.265 35.865 ;
        RECT 1980.135 35.850 1980.465 35.865 ;
        RECT 1981.070 35.850 1981.370 36.215 ;
        RECT 1786.935 35.550 1788.170 35.850 ;
        RECT 1441.935 35.535 1442.265 35.550 ;
        RECT 1786.935 35.535 1787.265 35.550 ;
        RECT 1787.870 35.185 1788.170 35.550 ;
        RECT 1980.135 35.550 1981.370 35.850 ;
        RECT 2455.790 35.850 2456.090 37.575 ;
        RECT 2835.735 36.895 2836.065 37.225 ;
        RECT 2456.695 36.215 2457.025 36.545 ;
        RECT 2456.710 35.850 2457.010 36.215 ;
        RECT 2455.790 35.550 2457.010 35.850 ;
        RECT 1980.135 35.535 1980.465 35.550 ;
        RECT 2835.750 35.185 2836.050 36.895 ;
        RECT 1110.735 34.855 1111.065 35.185 ;
        RECT 1787.855 34.855 1788.185 35.185 ;
        RECT 2835.735 34.855 2836.065 35.185 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2680.490 2380.580 2680.810 2380.640 ;
        RECT 2900.830 2380.580 2901.150 2380.640 ;
        RECT 2680.490 2380.440 2901.150 2380.580 ;
        RECT 2680.490 2380.380 2680.810 2380.440 ;
        RECT 2900.830 2380.380 2901.150 2380.440 ;
        RECT 2615.170 1628.160 2615.490 1628.220 ;
        RECT 2680.490 1628.160 2680.810 1628.220 ;
        RECT 2615.170 1628.020 2680.810 1628.160 ;
        RECT 2615.170 1627.960 2615.490 1628.020 ;
        RECT 2680.490 1627.960 2680.810 1628.020 ;
      LAYER via ;
        RECT 2680.520 2380.380 2680.780 2380.640 ;
        RECT 2900.860 2380.380 2901.120 2380.640 ;
        RECT 2615.200 1627.960 2615.460 1628.220 ;
        RECT 2680.520 1627.960 2680.780 1628.220 ;
      LAYER met2 ;
        RECT 2900.850 2384.915 2901.130 2385.285 ;
        RECT 2900.920 2380.670 2901.060 2384.915 ;
        RECT 2680.520 2380.350 2680.780 2380.670 ;
        RECT 2900.860 2380.350 2901.120 2380.670 ;
        RECT 2615.190 1628.075 2615.470 1628.445 ;
        RECT 2680.580 1628.250 2680.720 2380.350 ;
        RECT 2615.200 1627.930 2615.460 1628.075 ;
        RECT 2680.520 1627.930 2680.780 1628.250 ;
      LAYER via2 ;
        RECT 2900.850 2384.960 2901.130 2385.240 ;
        RECT 2615.190 1628.120 2615.470 1628.400 ;
      LAYER met3 ;
        RECT 2900.825 2385.250 2901.155 2385.265 ;
        RECT 2917.600 2385.250 2924.800 2385.700 ;
        RECT 2900.825 2384.950 2924.800 2385.250 ;
        RECT 2900.825 2384.935 2901.155 2384.950 ;
        RECT 2917.600 2384.500 2924.800 2384.950 ;
        RECT 2606.000 1628.410 2610.000 1628.800 ;
        RECT 2615.165 1628.410 2615.495 1628.425 ;
        RECT 2606.000 1628.200 2615.495 1628.410 ;
        RECT 2609.580 1628.110 2615.495 1628.200 ;
        RECT 2615.165 1628.095 2615.495 1628.110 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2006.590 3264.920 2006.910 3264.980 ;
        RECT 2867.250 3264.920 2867.570 3264.980 ;
        RECT 2006.590 3264.780 2867.570 3264.920 ;
        RECT 2006.590 3264.720 2006.910 3264.780 ;
        RECT 2867.250 3264.720 2867.570 3264.780 ;
        RECT 2867.250 2621.980 2867.570 2622.040 ;
        RECT 2900.830 2621.980 2901.150 2622.040 ;
        RECT 2867.250 2621.840 2901.150 2621.980 ;
        RECT 2867.250 2621.780 2867.570 2621.840 ;
        RECT 2900.830 2621.780 2901.150 2621.840 ;
      LAYER via ;
        RECT 2006.620 3264.720 2006.880 3264.980 ;
        RECT 2867.280 3264.720 2867.540 3264.980 ;
        RECT 2867.280 2621.780 2867.540 2622.040 ;
        RECT 2900.860 2621.780 2901.120 2622.040 ;
      LAYER met2 ;
        RECT 2006.620 3264.690 2006.880 3265.010 ;
        RECT 2867.280 3264.690 2867.540 3265.010 ;
        RECT 2006.680 3260.000 2006.820 3264.690 ;
        RECT 2006.570 3256.000 2006.850 3260.000 ;
        RECT 2867.340 2622.070 2867.480 3264.690 ;
        RECT 2867.280 2621.750 2867.540 2622.070 ;
        RECT 2900.860 2621.750 2901.120 2622.070 ;
        RECT 2900.920 2619.885 2901.060 2621.750 ;
        RECT 2900.850 2619.515 2901.130 2619.885 ;
      LAYER via2 ;
        RECT 2900.850 2619.560 2901.130 2619.840 ;
      LAYER met3 ;
        RECT 2900.825 2619.850 2901.155 2619.865 ;
        RECT 2917.600 2619.850 2924.800 2620.300 ;
        RECT 2900.825 2619.550 2924.800 2619.850 ;
        RECT 2900.825 2619.535 2901.155 2619.550 ;
        RECT 2917.600 2619.100 2924.800 2619.550 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.510 248.100 2214.830 248.160 ;
        RECT 2901.290 248.100 2901.610 248.160 ;
        RECT 2214.510 247.960 2901.610 248.100 ;
        RECT 2214.510 247.900 2214.830 247.960 ;
        RECT 2901.290 247.900 2901.610 247.960 ;
      LAYER via ;
        RECT 2214.540 247.900 2214.800 248.160 ;
        RECT 2901.320 247.900 2901.580 248.160 ;
      LAYER met2 ;
        RECT 2901.310 2854.115 2901.590 2854.485 ;
        RECT 2214.490 260.000 2214.770 264.000 ;
        RECT 2214.600 248.190 2214.740 260.000 ;
        RECT 2901.380 248.190 2901.520 2854.115 ;
        RECT 2214.540 247.870 2214.800 248.190 ;
        RECT 2901.320 247.870 2901.580 248.190 ;
      LAYER via2 ;
        RECT 2901.310 2854.160 2901.590 2854.440 ;
      LAYER met3 ;
        RECT 2901.285 2854.450 2901.615 2854.465 ;
        RECT 2917.600 2854.450 2924.800 2854.900 ;
        RECT 2901.285 2854.150 2924.800 2854.450 ;
        RECT 2901.285 2854.135 2901.615 2854.150 ;
        RECT 2917.600 2853.700 2924.800 2854.150 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2704.410 3084.720 2704.730 3084.780 ;
        RECT 2745.810 3084.720 2746.130 3084.780 ;
        RECT 2704.410 3084.580 2746.130 3084.720 ;
        RECT 2704.410 3084.520 2704.730 3084.580 ;
        RECT 2745.810 3084.520 2746.130 3084.580 ;
      LAYER via ;
        RECT 2704.440 3084.520 2704.700 3084.780 ;
        RECT 2745.840 3084.520 2746.100 3084.780 ;
      LAYER met2 ;
        RECT 2767.450 3085.570 2767.730 3085.685 ;
        RECT 2766.600 3085.430 2767.730 3085.570 ;
        RECT 2766.600 3085.005 2766.740 3085.430 ;
        RECT 2767.450 3085.315 2767.730 3085.430 ;
        RECT 2801.490 3085.570 2801.770 3085.685 ;
        RECT 2801.490 3085.430 2802.160 3085.570 ;
        RECT 2801.490 3085.315 2801.770 3085.430 ;
        RECT 2802.020 3085.005 2802.160 3085.430 ;
        RECT 2863.130 3085.315 2863.410 3085.685 ;
        RECT 2704.440 3084.490 2704.700 3084.810 ;
        RECT 2745.830 3084.635 2746.110 3085.005 ;
        RECT 2766.530 3084.635 2766.810 3085.005 ;
        RECT 2801.950 3084.635 2802.230 3085.005 ;
        RECT 2863.200 3084.890 2863.340 3085.315 ;
        RECT 2863.590 3084.890 2863.870 3085.005 ;
        RECT 2863.200 3084.750 2863.870 3084.890 ;
        RECT 2863.590 3084.635 2863.870 3084.750 ;
        RECT 2745.840 3084.490 2746.100 3084.635 ;
        RECT 2704.500 3064.605 2704.640 3084.490 ;
        RECT 2704.430 3064.235 2704.710 3064.605 ;
      LAYER via2 ;
        RECT 2767.450 3085.360 2767.730 3085.640 ;
        RECT 2801.490 3085.360 2801.770 3085.640 ;
        RECT 2863.130 3085.360 2863.410 3085.640 ;
        RECT 2745.830 3084.680 2746.110 3084.960 ;
        RECT 2766.530 3084.680 2766.810 3084.960 ;
        RECT 2801.950 3084.680 2802.230 3084.960 ;
        RECT 2863.590 3084.680 2863.870 3084.960 ;
        RECT 2704.430 3064.280 2704.710 3064.560 ;
      LAYER met3 ;
        RECT 2917.600 3089.050 2924.800 3089.500 ;
        RECT 2916.710 3088.750 2924.800 3089.050 ;
        RECT 2767.425 3085.650 2767.755 3085.665 ;
        RECT 2801.465 3085.650 2801.795 3085.665 ;
        RECT 2863.105 3085.650 2863.435 3085.665 ;
        RECT 2767.425 3085.350 2801.795 3085.650 ;
        RECT 2767.425 3085.335 2767.755 3085.350 ;
        RECT 2801.465 3085.335 2801.795 3085.350 ;
        RECT 2849.550 3085.350 2863.435 3085.650 ;
        RECT 2745.805 3084.970 2746.135 3084.985 ;
        RECT 2766.505 3084.970 2766.835 3084.985 ;
        RECT 2745.805 3084.670 2766.835 3084.970 ;
        RECT 2745.805 3084.655 2746.135 3084.670 ;
        RECT 2766.505 3084.655 2766.835 3084.670 ;
        RECT 2801.925 3084.970 2802.255 3084.985 ;
        RECT 2849.550 3084.970 2849.850 3085.350 ;
        RECT 2863.105 3085.335 2863.435 3085.350 ;
        RECT 2801.925 3084.670 2849.850 3084.970 ;
        RECT 2863.565 3084.970 2863.895 3084.985 ;
        RECT 2916.710 3084.970 2917.010 3088.750 ;
        RECT 2917.600 3088.300 2924.800 3088.750 ;
        RECT 2863.565 3084.670 2917.010 3084.970 ;
        RECT 2801.925 3084.655 2802.255 3084.670 ;
        RECT 2863.565 3084.655 2863.895 3084.670 ;
        RECT 2660.910 3064.570 2661.290 3064.580 ;
        RECT 2704.405 3064.570 2704.735 3064.585 ;
        RECT 2660.910 3064.270 2704.735 3064.570 ;
        RECT 2660.910 3064.260 2661.290 3064.270 ;
        RECT 2704.405 3064.255 2704.735 3064.270 ;
        RECT 307.550 1701.850 307.930 1701.860 ;
        RECT 307.550 1701.550 310.650 1701.850 ;
        RECT 307.550 1701.540 307.930 1701.550 ;
        RECT 310.350 1700.880 310.650 1701.550 ;
        RECT 310.000 1700.280 314.000 1700.880 ;
      LAYER via3 ;
        RECT 2660.940 3064.260 2661.260 3064.580 ;
        RECT 307.580 1701.540 307.900 1701.860 ;
      LAYER met4 ;
        RECT 2660.935 3064.255 2661.265 3064.585 ;
        RECT 2660.950 1702.290 2661.250 3064.255 ;
        RECT 307.150 1701.110 308.330 1702.290 ;
        RECT 2660.510 1701.110 2661.690 1702.290 ;
      LAYER met5 ;
        RECT 627.100 1711.100 666.420 1712.700 ;
        RECT 336.380 1702.500 338.900 1709.300 ;
        RECT 627.100 1705.900 628.700 1711.100 ;
        RECT 413.660 1704.300 435.500 1705.900 ;
        RECT 306.940 1700.900 405.140 1702.500 ;
        RECT 403.540 1695.700 405.140 1700.900 ;
        RECT 413.660 1695.700 415.260 1704.300 ;
        RECT 433.900 1702.500 435.500 1704.300 ;
        RECT 471.620 1704.300 556.020 1705.900 ;
        RECT 471.620 1702.500 473.220 1704.300 ;
        RECT 433.900 1700.900 473.220 1702.500 ;
        RECT 554.420 1702.500 556.020 1704.300 ;
        RECT 568.220 1704.300 628.700 1705.900 ;
        RECT 664.820 1705.900 666.420 1711.100 ;
        RECT 690.580 1711.100 735.420 1712.700 ;
        RECT 690.580 1709.300 692.180 1711.100 ;
        RECT 675.860 1707.700 692.180 1709.300 ;
        RECT 675.860 1705.900 677.460 1707.700 ;
        RECT 664.820 1704.300 677.460 1705.900 ;
        RECT 568.220 1702.500 569.820 1704.300 ;
        RECT 554.420 1700.900 569.820 1702.500 ;
        RECT 403.540 1694.100 415.260 1695.700 ;
        RECT 733.820 1695.700 735.420 1711.100 ;
        RECT 812.940 1711.100 832.020 1712.700 ;
        RECT 812.940 1709.300 814.540 1711.100 ;
        RECT 766.020 1707.700 814.540 1709.300 ;
        RECT 766.020 1699.100 767.620 1707.700 ;
        RECT 765.100 1697.500 767.620 1699.100 ;
        RECT 765.100 1695.700 766.700 1697.500 ;
        RECT 733.820 1694.100 766.700 1695.700 ;
        RECT 830.420 1695.700 832.020 1711.100 ;
        RECT 909.540 1711.100 928.620 1712.700 ;
        RECT 909.540 1709.300 911.140 1711.100 ;
        RECT 862.620 1707.700 911.140 1709.300 ;
        RECT 862.620 1699.100 864.220 1707.700 ;
        RECT 861.700 1697.500 864.220 1699.100 ;
        RECT 861.700 1695.700 863.300 1697.500 ;
        RECT 830.420 1694.100 863.300 1695.700 ;
        RECT 927.020 1695.700 928.620 1711.100 ;
        RECT 1006.140 1711.100 1025.220 1712.700 ;
        RECT 1006.140 1709.300 1007.740 1711.100 ;
        RECT 959.220 1707.700 1007.740 1709.300 ;
        RECT 959.220 1699.100 960.820 1707.700 ;
        RECT 958.300 1697.500 960.820 1699.100 ;
        RECT 958.300 1695.700 959.900 1697.500 ;
        RECT 927.020 1694.100 959.900 1695.700 ;
        RECT 1023.620 1695.700 1025.220 1711.100 ;
        RECT 1102.740 1711.100 1121.820 1712.700 ;
        RECT 1102.740 1709.300 1104.340 1711.100 ;
        RECT 1055.820 1707.700 1104.340 1709.300 ;
        RECT 1055.820 1699.100 1057.420 1707.700 ;
        RECT 1054.900 1697.500 1057.420 1699.100 ;
        RECT 1054.900 1695.700 1056.500 1697.500 ;
        RECT 1023.620 1694.100 1056.500 1695.700 ;
        RECT 1120.220 1695.700 1121.820 1711.100 ;
        RECT 1199.340 1711.100 1218.420 1712.700 ;
        RECT 1199.340 1709.300 1200.940 1711.100 ;
        RECT 1152.420 1707.700 1200.940 1709.300 ;
        RECT 1152.420 1699.100 1154.020 1707.700 ;
        RECT 1151.500 1697.500 1154.020 1699.100 ;
        RECT 1151.500 1695.700 1153.100 1697.500 ;
        RECT 1120.220 1694.100 1153.100 1695.700 ;
        RECT 1216.820 1695.700 1218.420 1711.100 ;
        RECT 1295.940 1711.100 1315.020 1712.700 ;
        RECT 1295.940 1709.300 1297.540 1711.100 ;
        RECT 1249.020 1707.700 1297.540 1709.300 ;
        RECT 1249.020 1699.100 1250.620 1707.700 ;
        RECT 1248.100 1697.500 1250.620 1699.100 ;
        RECT 1248.100 1695.700 1249.700 1697.500 ;
        RECT 1216.820 1694.100 1249.700 1695.700 ;
        RECT 1313.420 1695.700 1315.020 1711.100 ;
        RECT 1392.540 1711.100 1411.620 1712.700 ;
        RECT 1392.540 1709.300 1394.140 1711.100 ;
        RECT 1345.620 1707.700 1394.140 1709.300 ;
        RECT 1345.620 1699.100 1347.220 1707.700 ;
        RECT 1344.700 1697.500 1347.220 1699.100 ;
        RECT 1344.700 1695.700 1346.300 1697.500 ;
        RECT 1313.420 1694.100 1346.300 1695.700 ;
        RECT 1410.020 1695.700 1411.620 1711.100 ;
        RECT 1489.140 1711.100 1508.220 1712.700 ;
        RECT 1489.140 1709.300 1490.740 1711.100 ;
        RECT 1442.220 1707.700 1490.740 1709.300 ;
        RECT 1442.220 1699.100 1443.820 1707.700 ;
        RECT 1441.300 1697.500 1443.820 1699.100 ;
        RECT 1441.300 1695.700 1442.900 1697.500 ;
        RECT 1410.020 1694.100 1442.900 1695.700 ;
        RECT 1506.620 1695.700 1508.220 1711.100 ;
        RECT 1585.740 1711.100 1604.820 1712.700 ;
        RECT 1585.740 1709.300 1587.340 1711.100 ;
        RECT 1538.820 1707.700 1587.340 1709.300 ;
        RECT 1538.820 1699.100 1540.420 1707.700 ;
        RECT 1537.900 1697.500 1540.420 1699.100 ;
        RECT 1537.900 1695.700 1539.500 1697.500 ;
        RECT 1506.620 1694.100 1539.500 1695.700 ;
        RECT 1603.220 1695.700 1604.820 1711.100 ;
        RECT 1682.340 1711.100 1701.420 1712.700 ;
        RECT 1682.340 1709.300 1683.940 1711.100 ;
        RECT 1635.420 1707.700 1683.940 1709.300 ;
        RECT 1635.420 1699.100 1637.020 1707.700 ;
        RECT 1634.500 1697.500 1637.020 1699.100 ;
        RECT 1634.500 1695.700 1636.100 1697.500 ;
        RECT 1603.220 1694.100 1636.100 1695.700 ;
        RECT 1699.820 1695.700 1701.420 1711.100 ;
        RECT 1778.940 1711.100 1798.020 1712.700 ;
        RECT 1778.940 1709.300 1780.540 1711.100 ;
        RECT 1732.020 1707.700 1780.540 1709.300 ;
        RECT 1732.020 1699.100 1733.620 1707.700 ;
        RECT 1731.100 1697.500 1733.620 1699.100 ;
        RECT 1731.100 1695.700 1732.700 1697.500 ;
        RECT 1699.820 1694.100 1732.700 1695.700 ;
        RECT 1796.420 1695.700 1798.020 1711.100 ;
        RECT 1875.540 1711.100 1894.620 1712.700 ;
        RECT 1875.540 1709.300 1877.140 1711.100 ;
        RECT 1828.620 1707.700 1877.140 1709.300 ;
        RECT 1828.620 1699.100 1830.220 1707.700 ;
        RECT 1827.700 1697.500 1830.220 1699.100 ;
        RECT 1827.700 1695.700 1829.300 1697.500 ;
        RECT 1796.420 1694.100 1829.300 1695.700 ;
        RECT 1893.020 1695.700 1894.620 1711.100 ;
        RECT 1972.140 1711.100 1991.220 1712.700 ;
        RECT 1972.140 1709.300 1973.740 1711.100 ;
        RECT 1925.220 1707.700 1973.740 1709.300 ;
        RECT 1925.220 1699.100 1926.820 1707.700 ;
        RECT 1924.300 1697.500 1926.820 1699.100 ;
        RECT 1924.300 1695.700 1925.900 1697.500 ;
        RECT 1893.020 1694.100 1925.900 1695.700 ;
        RECT 1989.620 1695.700 1991.220 1711.100 ;
        RECT 2068.740 1711.100 2087.820 1712.700 ;
        RECT 2068.740 1709.300 2070.340 1711.100 ;
        RECT 2021.820 1707.700 2070.340 1709.300 ;
        RECT 2021.820 1699.100 2023.420 1707.700 ;
        RECT 2020.900 1697.500 2023.420 1699.100 ;
        RECT 2020.900 1695.700 2022.500 1697.500 ;
        RECT 1989.620 1694.100 2022.500 1695.700 ;
        RECT 2086.220 1695.700 2087.820 1711.100 ;
        RECT 2165.340 1711.100 2184.420 1712.700 ;
        RECT 2165.340 1709.300 2166.940 1711.100 ;
        RECT 2118.420 1707.700 2166.940 1709.300 ;
        RECT 2118.420 1699.100 2120.020 1707.700 ;
        RECT 2117.500 1697.500 2120.020 1699.100 ;
        RECT 2117.500 1695.700 2119.100 1697.500 ;
        RECT 2086.220 1694.100 2119.100 1695.700 ;
        RECT 2182.820 1695.700 2184.420 1711.100 ;
        RECT 2261.940 1711.100 2281.020 1712.700 ;
        RECT 2261.940 1709.300 2263.540 1711.100 ;
        RECT 2215.020 1707.700 2263.540 1709.300 ;
        RECT 2215.020 1699.100 2216.620 1707.700 ;
        RECT 2214.100 1697.500 2216.620 1699.100 ;
        RECT 2214.100 1695.700 2215.700 1697.500 ;
        RECT 2182.820 1694.100 2215.700 1695.700 ;
        RECT 2279.420 1695.700 2281.020 1711.100 ;
        RECT 2358.540 1711.100 2377.620 1712.700 ;
        RECT 2358.540 1709.300 2360.140 1711.100 ;
        RECT 2311.620 1707.700 2360.140 1709.300 ;
        RECT 2311.620 1699.100 2313.220 1707.700 ;
        RECT 2310.700 1697.500 2313.220 1699.100 ;
        RECT 2310.700 1695.700 2312.300 1697.500 ;
        RECT 2279.420 1694.100 2312.300 1695.700 ;
        RECT 2376.020 1695.700 2377.620 1711.100 ;
        RECT 2455.140 1709.300 2457.660 1712.700 ;
        RECT 2408.220 1707.700 2475.140 1709.300 ;
        RECT 2408.220 1699.100 2409.820 1707.700 ;
        RECT 2407.300 1697.500 2409.820 1699.100 ;
        RECT 2407.300 1695.700 2408.900 1697.500 ;
        RECT 2376.020 1694.100 2408.900 1695.700 ;
        RECT 2473.540 1695.700 2475.140 1707.700 ;
        RECT 2569.220 1704.300 2575.420 1705.900 ;
        RECT 2569.220 1695.700 2570.820 1704.300 ;
        RECT 2573.820 1699.100 2575.420 1704.300 ;
        RECT 2617.980 1704.300 2628.780 1705.900 ;
        RECT 2617.980 1699.100 2619.580 1704.300 ;
        RECT 2627.180 1702.500 2628.780 1704.300 ;
        RECT 2627.180 1700.900 2661.900 1702.500 ;
        RECT 2573.820 1697.500 2619.580 1699.100 ;
        RECT 2473.540 1694.100 2570.820 1695.700 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.250 3318.980 268.570 3319.040 ;
        RECT 2900.830 3318.980 2901.150 3319.040 ;
        RECT 268.250 3318.840 2901.150 3318.980 ;
        RECT 268.250 3318.780 268.570 3318.840 ;
        RECT 2900.830 3318.780 2901.150 3318.840 ;
        RECT 268.250 687.720 268.570 687.780 ;
        RECT 296.770 687.720 297.090 687.780 ;
        RECT 268.250 687.580 297.090 687.720 ;
        RECT 268.250 687.520 268.570 687.580 ;
        RECT 296.770 687.520 297.090 687.580 ;
      LAYER via ;
        RECT 268.280 3318.780 268.540 3319.040 ;
        RECT 2900.860 3318.780 2901.120 3319.040 ;
        RECT 268.280 687.520 268.540 687.780 ;
        RECT 296.800 687.520 297.060 687.780 ;
      LAYER met2 ;
        RECT 2900.850 3323.315 2901.130 3323.685 ;
        RECT 2900.920 3319.070 2901.060 3323.315 ;
        RECT 268.280 3318.750 268.540 3319.070 ;
        RECT 2900.860 3318.750 2901.120 3319.070 ;
        RECT 268.340 687.810 268.480 3318.750 ;
        RECT 268.280 687.490 268.540 687.810 ;
        RECT 296.800 687.490 297.060 687.810 ;
        RECT 296.860 685.965 297.000 687.490 ;
        RECT 296.790 685.595 297.070 685.965 ;
      LAYER via2 ;
        RECT 2900.850 3323.360 2901.130 3323.640 ;
        RECT 296.790 685.640 297.070 685.920 ;
      LAYER met3 ;
        RECT 2900.825 3323.650 2901.155 3323.665 ;
        RECT 2917.600 3323.650 2924.800 3324.100 ;
        RECT 2900.825 3323.350 2924.800 3323.650 ;
        RECT 2900.825 3323.335 2901.155 3323.350 ;
        RECT 2917.600 3322.900 2924.800 3323.350 ;
        RECT 296.765 685.930 297.095 685.945 ;
        RECT 310.000 685.930 314.000 686.320 ;
        RECT 296.765 685.720 314.000 685.930 ;
        RECT 296.765 685.630 310.500 685.720 ;
        RECT 296.765 685.615 297.095 685.630 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 3501.560 393.230 3501.620 ;
        RECT 2865.410 3501.560 2865.730 3501.620 ;
        RECT 392.910 3501.420 2865.730 3501.560 ;
        RECT 392.910 3501.360 393.230 3501.420 ;
        RECT 2865.410 3501.360 2865.730 3501.420 ;
      LAYER via ;
        RECT 392.940 3501.360 393.200 3501.620 ;
        RECT 2865.440 3501.360 2865.700 3501.620 ;
      LAYER met2 ;
        RECT 2865.290 3517.600 2865.850 3524.800 ;
        RECT 2865.500 3501.650 2865.640 3517.600 ;
        RECT 392.940 3501.330 393.200 3501.650 ;
        RECT 2865.440 3501.330 2865.700 3501.650 ;
        RECT 393.000 3260.330 393.140 3501.330 ;
        RECT 391.620 3260.190 393.140 3260.330 ;
        RECT 390.130 3259.650 390.410 3260.000 ;
        RECT 391.620 3259.650 391.760 3260.190 ;
        RECT 390.130 3259.510 391.760 3259.650 ;
        RECT 390.130 3256.000 390.410 3259.510 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2541.110 3501.900 2541.430 3501.960 ;
        RECT 2654.270 3501.900 2654.590 3501.960 ;
        RECT 2541.110 3501.760 2654.590 3501.900 ;
        RECT 2541.110 3501.700 2541.430 3501.760 ;
        RECT 2654.270 3501.700 2654.590 3501.760 ;
      LAYER via ;
        RECT 2541.140 3501.700 2541.400 3501.960 ;
        RECT 2654.300 3501.700 2654.560 3501.960 ;
      LAYER met2 ;
        RECT 2540.990 3517.600 2541.550 3524.800 ;
        RECT 2541.200 3501.990 2541.340 3517.600 ;
        RECT 2541.140 3501.670 2541.400 3501.990 ;
        RECT 2654.300 3501.670 2654.560 3501.990 ;
        RECT 827.130 260.000 827.410 264.000 ;
        RECT 827.240 243.965 827.380 260.000 ;
        RECT 2654.360 243.965 2654.500 3501.670 ;
        RECT 827.170 243.595 827.450 243.965 ;
        RECT 2654.290 243.595 2654.570 243.965 ;
      LAYER via2 ;
        RECT 827.170 243.640 827.450 243.920 ;
        RECT 2654.290 243.640 2654.570 243.920 ;
      LAYER met3 ;
        RECT 827.145 243.930 827.475 243.945 ;
        RECT 2654.265 243.930 2654.595 243.945 ;
        RECT 827.145 243.630 2654.595 243.930 ;
        RECT 827.145 243.615 827.475 243.630 ;
        RECT 2654.265 243.615 2654.595 243.630 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1552.110 3503.260 1552.430 3503.320 ;
        RECT 2216.810 3503.260 2217.130 3503.320 ;
        RECT 1552.110 3503.120 2217.130 3503.260 ;
        RECT 1552.110 3503.060 1552.430 3503.120 ;
        RECT 2216.810 3503.060 2217.130 3503.120 ;
        RECT 1548.430 3277.500 1548.750 3277.560 ;
        RECT 1552.110 3277.500 1552.430 3277.560 ;
        RECT 1548.430 3277.360 1552.430 3277.500 ;
        RECT 1548.430 3277.300 1548.750 3277.360 ;
        RECT 1552.110 3277.300 1552.430 3277.360 ;
      LAYER via ;
        RECT 1552.140 3503.060 1552.400 3503.320 ;
        RECT 2216.840 3503.060 2217.100 3503.320 ;
        RECT 1548.460 3277.300 1548.720 3277.560 ;
        RECT 1552.140 3277.300 1552.400 3277.560 ;
      LAYER met2 ;
        RECT 2216.690 3517.600 2217.250 3524.800 ;
        RECT 2216.900 3503.350 2217.040 3517.600 ;
        RECT 1552.140 3503.030 1552.400 3503.350 ;
        RECT 2216.840 3503.030 2217.100 3503.350 ;
        RECT 1552.200 3277.590 1552.340 3503.030 ;
        RECT 1548.460 3277.270 1548.720 3277.590 ;
        RECT 1552.140 3277.270 1552.400 3277.590 ;
        RECT 1548.520 3260.000 1548.660 3277.270 ;
        RECT 1548.410 3256.000 1548.690 3260.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1892.050 3502.580 1892.370 3502.640 ;
        RECT 2651.510 3502.580 2651.830 3502.640 ;
        RECT 1892.050 3502.440 2651.830 3502.580 ;
        RECT 1892.050 3502.380 1892.370 3502.440 ;
        RECT 2651.510 3502.380 2651.830 3502.440 ;
      LAYER via ;
        RECT 1892.080 3502.380 1892.340 3502.640 ;
        RECT 2651.540 3502.380 2651.800 3502.640 ;
      LAYER met2 ;
        RECT 1891.930 3517.600 1892.490 3524.800 ;
        RECT 1892.140 3502.670 1892.280 3517.600 ;
        RECT 1892.080 3502.350 1892.340 3502.670 ;
        RECT 2651.540 3502.350 2651.800 3502.670 ;
        RECT 2586.170 260.000 2586.450 264.000 ;
        RECT 2586.280 248.045 2586.420 260.000 ;
        RECT 2651.600 248.045 2651.740 3502.350 ;
        RECT 2586.210 247.675 2586.490 248.045 ;
        RECT 2651.530 247.675 2651.810 248.045 ;
      LAYER via2 ;
        RECT 2586.210 247.720 2586.490 248.000 ;
        RECT 2651.530 247.720 2651.810 248.000 ;
      LAYER met3 ;
        RECT 2586.185 248.010 2586.515 248.025 ;
        RECT 2651.505 248.010 2651.835 248.025 ;
        RECT 2586.185 247.710 2651.835 248.010 ;
        RECT 2586.185 247.695 2586.515 247.710 ;
        RECT 2651.505 247.695 2651.835 247.710 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.910 3503.600 1152.230 3503.660 ;
        RECT 1567.750 3503.600 1568.070 3503.660 ;
        RECT 1151.910 3503.460 1568.070 3503.600 ;
        RECT 1151.910 3503.400 1152.230 3503.460 ;
        RECT 1567.750 3503.400 1568.070 3503.460 ;
        RECT 1148.230 3277.500 1148.550 3277.560 ;
        RECT 1151.910 3277.500 1152.230 3277.560 ;
        RECT 1148.230 3277.360 1152.230 3277.500 ;
        RECT 1148.230 3277.300 1148.550 3277.360 ;
        RECT 1151.910 3277.300 1152.230 3277.360 ;
      LAYER via ;
        RECT 1151.940 3503.400 1152.200 3503.660 ;
        RECT 1567.780 3503.400 1568.040 3503.660 ;
        RECT 1148.260 3277.300 1148.520 3277.560 ;
        RECT 1151.940 3277.300 1152.200 3277.560 ;
      LAYER met2 ;
        RECT 1567.630 3517.600 1568.190 3524.800 ;
        RECT 1567.840 3503.690 1567.980 3517.600 ;
        RECT 1151.940 3503.370 1152.200 3503.690 ;
        RECT 1567.780 3503.370 1568.040 3503.690 ;
        RECT 1152.000 3277.590 1152.140 3503.370 ;
        RECT 1148.260 3277.270 1148.520 3277.590 ;
        RECT 1151.940 3277.270 1152.200 3277.590 ;
        RECT 1148.320 3260.000 1148.460 3277.270 ;
        RECT 1148.210 3256.000 1148.490 3260.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1200.780 2614.570 1200.840 ;
        RECT 2701.650 1200.780 2701.970 1200.840 ;
        RECT 2614.250 1200.640 2701.970 1200.780 ;
        RECT 2614.250 1200.580 2614.570 1200.640 ;
        RECT 2701.650 1200.580 2701.970 1200.640 ;
        RECT 2701.650 275.980 2701.970 276.040 ;
        RECT 2898.990 275.980 2899.310 276.040 ;
        RECT 2701.650 275.840 2899.310 275.980 ;
        RECT 2701.650 275.780 2701.970 275.840 ;
        RECT 2898.990 275.780 2899.310 275.840 ;
      LAYER via ;
        RECT 2614.280 1200.580 2614.540 1200.840 ;
        RECT 2701.680 1200.580 2701.940 1200.840 ;
        RECT 2701.680 275.780 2701.940 276.040 ;
        RECT 2899.020 275.780 2899.280 276.040 ;
      LAYER met2 ;
        RECT 2614.270 1205.115 2614.550 1205.485 ;
        RECT 2614.340 1200.870 2614.480 1205.115 ;
        RECT 2614.280 1200.550 2614.540 1200.870 ;
        RECT 2701.680 1200.550 2701.940 1200.870 ;
        RECT 2701.740 276.070 2701.880 1200.550 ;
        RECT 2701.680 275.750 2701.940 276.070 ;
        RECT 2899.020 275.750 2899.280 276.070 ;
        RECT 2899.080 273.885 2899.220 275.750 ;
        RECT 2899.010 273.515 2899.290 273.885 ;
      LAYER via2 ;
        RECT 2614.270 1205.160 2614.550 1205.440 ;
        RECT 2899.010 273.560 2899.290 273.840 ;
      LAYER met3 ;
        RECT 2606.000 1205.450 2610.000 1205.840 ;
        RECT 2614.245 1205.450 2614.575 1205.465 ;
        RECT 2606.000 1205.240 2614.575 1205.450 ;
        RECT 2609.580 1205.150 2614.575 1205.240 ;
        RECT 2614.245 1205.135 2614.575 1205.150 ;
        RECT 2898.985 273.850 2899.315 273.865 ;
        RECT 2917.600 273.850 2924.800 274.300 ;
        RECT 2898.985 273.550 2924.800 273.850 ;
        RECT 2898.985 273.535 2899.315 273.550 ;
        RECT 2917.600 273.100 2924.800 273.550 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 275.610 3503.260 275.930 3503.320 ;
        RECT 1243.450 3503.260 1243.770 3503.320 ;
        RECT 275.610 3503.120 1243.770 3503.260 ;
        RECT 275.610 3503.060 275.930 3503.120 ;
        RECT 1243.450 3503.060 1243.770 3503.120 ;
      LAYER via ;
        RECT 275.640 3503.060 275.900 3503.320 ;
        RECT 1243.480 3503.060 1243.740 3503.320 ;
      LAYER met2 ;
        RECT 1243.330 3517.600 1243.890 3524.800 ;
        RECT 1243.540 3503.350 1243.680 3517.600 ;
        RECT 275.640 3503.030 275.900 3503.350 ;
        RECT 1243.480 3503.030 1243.740 3503.350 ;
        RECT 275.700 243.965 275.840 3503.030 ;
        RECT 483.970 260.000 484.250 264.000 ;
        RECT 484.080 243.965 484.220 260.000 ;
        RECT 275.630 243.595 275.910 243.965 ;
        RECT 484.010 243.595 484.290 243.965 ;
      LAYER via2 ;
        RECT 275.630 243.640 275.910 243.920 ;
        RECT 484.010 243.640 484.290 243.920 ;
      LAYER met3 ;
        RECT 275.605 243.930 275.935 243.945 ;
        RECT 483.985 243.930 484.315 243.945 ;
        RECT 275.605 243.630 484.315 243.930 ;
        RECT 275.605 243.615 275.935 243.630 ;
        RECT 483.985 243.615 484.315 243.630 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 304.590 3287.700 304.910 3287.760 ;
        RECT 918.230 3287.700 918.550 3287.760 ;
        RECT 304.590 3287.560 918.550 3287.700 ;
        RECT 304.590 3287.500 304.910 3287.560 ;
        RECT 918.230 3287.500 918.550 3287.560 ;
      LAYER via ;
        RECT 304.620 3287.500 304.880 3287.760 ;
        RECT 918.260 3287.500 918.520 3287.760 ;
      LAYER met2 ;
        RECT 918.570 3517.600 919.130 3524.800 ;
        RECT 918.780 3443.250 918.920 3517.600 ;
        RECT 918.780 3443.110 919.380 3443.250 ;
        RECT 919.240 3346.690 919.380 3443.110 ;
        RECT 918.320 3346.550 919.380 3346.690 ;
        RECT 918.320 3287.790 918.460 3346.550 ;
        RECT 304.620 3287.470 304.880 3287.790 ;
        RECT 918.260 3287.470 918.520 3287.790 ;
        RECT 304.680 1321.085 304.820 3287.470 ;
        RECT 304.610 1320.715 304.890 1321.085 ;
      LAYER via2 ;
        RECT 304.610 1320.760 304.890 1321.040 ;
      LAYER met3 ;
        RECT 304.585 1321.050 304.915 1321.065 ;
        RECT 310.000 1321.050 314.000 1321.440 ;
        RECT 304.585 1320.840 314.000 1321.050 ;
        RECT 304.585 1320.750 310.500 1320.840 ;
        RECT 304.585 1320.735 304.915 1320.750 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 3502.580 241.430 3502.640 ;
        RECT 594.390 3502.580 594.710 3502.640 ;
        RECT 241.110 3502.440 594.710 3502.580 ;
        RECT 241.110 3502.380 241.430 3502.440 ;
        RECT 594.390 3502.380 594.710 3502.440 ;
        RECT 241.110 247.420 241.430 247.480 ;
        RECT 783.910 247.420 784.230 247.480 ;
        RECT 241.110 247.280 784.230 247.420 ;
        RECT 241.110 247.220 241.430 247.280 ;
        RECT 783.910 247.220 784.230 247.280 ;
      LAYER via ;
        RECT 241.140 3502.380 241.400 3502.640 ;
        RECT 594.420 3502.380 594.680 3502.640 ;
        RECT 241.140 247.220 241.400 247.480 ;
        RECT 783.940 247.220 784.200 247.480 ;
      LAYER met2 ;
        RECT 594.270 3517.600 594.830 3524.800 ;
        RECT 594.480 3502.670 594.620 3517.600 ;
        RECT 241.140 3502.350 241.400 3502.670 ;
        RECT 594.420 3502.350 594.680 3502.670 ;
        RECT 241.200 247.510 241.340 3502.350 ;
        RECT 783.890 260.000 784.170 264.000 ;
        RECT 784.000 247.510 784.140 260.000 ;
        RECT 241.140 247.190 241.400 247.510 ;
        RECT 783.940 247.190 784.200 247.510 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 270.090 3502.240 270.410 3502.300 ;
        RECT 1959.670 3502.240 1959.990 3502.300 ;
        RECT 270.090 3502.100 1959.990 3502.240 ;
        RECT 270.090 3502.040 270.410 3502.100 ;
        RECT 1959.670 3502.040 1959.990 3502.100 ;
      LAYER via ;
        RECT 270.120 3502.040 270.380 3502.300 ;
        RECT 1959.700 3502.040 1959.960 3502.300 ;
      LAYER met2 ;
        RECT 269.970 3517.600 270.530 3524.800 ;
        RECT 270.180 3502.330 270.320 3517.600 ;
        RECT 270.120 3502.010 270.380 3502.330 ;
        RECT 1959.700 3502.010 1959.960 3502.330 ;
        RECT 1959.760 3259.650 1959.900 3502.010 ;
        RECT 1963.330 3259.650 1963.610 3260.000 ;
        RECT 1959.760 3259.510 1963.610 3259.650 ;
        RECT 1963.330 3256.000 1963.610 3259.510 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.790 3470.960 15.110 3471.020 ;
        RECT 2644.610 3470.960 2644.930 3471.020 ;
        RECT 14.790 3470.820 2644.930 3470.960 ;
        RECT 14.790 3470.760 15.110 3470.820 ;
        RECT 2644.610 3470.760 2644.930 3470.820 ;
        RECT 2615.170 528.260 2615.490 528.320 ;
        RECT 2644.610 528.260 2644.930 528.320 ;
        RECT 2615.170 528.120 2644.930 528.260 ;
        RECT 2615.170 528.060 2615.490 528.120 ;
        RECT 2644.610 528.060 2644.930 528.120 ;
      LAYER via ;
        RECT 14.820 3470.760 15.080 3471.020 ;
        RECT 2644.640 3470.760 2644.900 3471.020 ;
        RECT 2615.200 528.060 2615.460 528.320 ;
        RECT 2644.640 528.060 2644.900 528.320 ;
      LAYER met2 ;
        RECT 14.810 3476.995 15.090 3477.365 ;
        RECT 14.880 3471.050 15.020 3476.995 ;
        RECT 14.820 3470.730 15.080 3471.050 ;
        RECT 2644.640 3470.730 2644.900 3471.050 ;
        RECT 2644.700 528.350 2644.840 3470.730 ;
        RECT 2615.200 528.205 2615.460 528.350 ;
        RECT 2615.190 527.835 2615.470 528.205 ;
        RECT 2644.640 528.030 2644.900 528.350 ;
      LAYER via2 ;
        RECT 14.810 3477.040 15.090 3477.320 ;
        RECT 2615.190 527.880 2615.470 528.160 ;
      LAYER met3 ;
        RECT -4.800 3477.330 2.400 3477.780 ;
        RECT 14.785 3477.330 15.115 3477.345 ;
        RECT -4.800 3477.030 15.115 3477.330 ;
        RECT -4.800 3476.580 2.400 3477.030 ;
        RECT 14.785 3477.015 15.115 3477.030 ;
        RECT 2606.000 528.170 2610.000 528.560 ;
        RECT 2615.165 528.170 2615.495 528.185 ;
        RECT 2606.000 527.960 2615.495 528.170 ;
        RECT 2609.580 527.870 2615.495 527.960 ;
        RECT 2615.165 527.855 2615.495 527.870 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 3222.420 15.570 3222.480 ;
        RECT 72.750 3222.420 73.070 3222.480 ;
        RECT 15.250 3222.280 73.070 3222.420 ;
        RECT 15.250 3222.220 15.570 3222.280 ;
        RECT 72.750 3222.220 73.070 3222.280 ;
        RECT 72.750 1028.060 73.070 1028.120 ;
        RECT 296.770 1028.060 297.090 1028.120 ;
        RECT 72.750 1027.920 297.090 1028.060 ;
        RECT 72.750 1027.860 73.070 1027.920 ;
        RECT 296.770 1027.860 297.090 1027.920 ;
      LAYER via ;
        RECT 15.280 3222.220 15.540 3222.480 ;
        RECT 72.780 3222.220 73.040 3222.480 ;
        RECT 72.780 1027.860 73.040 1028.120 ;
        RECT 296.800 1027.860 297.060 1028.120 ;
      LAYER met2 ;
        RECT 15.270 3226.075 15.550 3226.445 ;
        RECT 15.340 3222.510 15.480 3226.075 ;
        RECT 15.280 3222.190 15.540 3222.510 ;
        RECT 72.780 3222.190 73.040 3222.510 ;
        RECT 72.840 1028.150 72.980 3222.190 ;
        RECT 72.780 1027.830 73.040 1028.150 ;
        RECT 296.800 1027.830 297.060 1028.150 ;
        RECT 296.860 1024.605 297.000 1027.830 ;
        RECT 296.790 1024.235 297.070 1024.605 ;
      LAYER via2 ;
        RECT 15.270 3226.120 15.550 3226.400 ;
        RECT 296.790 1024.280 297.070 1024.560 ;
      LAYER met3 ;
        RECT -4.800 3226.410 2.400 3226.860 ;
        RECT 15.245 3226.410 15.575 3226.425 ;
        RECT -4.800 3226.110 15.575 3226.410 ;
        RECT -4.800 3225.660 2.400 3226.110 ;
        RECT 15.245 3226.095 15.575 3226.110 ;
        RECT 296.765 1024.570 297.095 1024.585 ;
        RECT 310.000 1024.570 314.000 1024.960 ;
        RECT 296.765 1024.360 314.000 1024.570 ;
        RECT 296.765 1024.270 310.500 1024.360 ;
        RECT 296.765 1024.255 297.095 1024.270 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2974.220 17.870 2974.280 ;
        RECT 65.390 2974.220 65.710 2974.280 ;
        RECT 17.550 2974.080 65.710 2974.220 ;
        RECT 17.550 2974.020 17.870 2974.080 ;
        RECT 65.390 2974.020 65.710 2974.080 ;
        RECT 65.390 255.580 65.710 255.640 ;
        RECT 584.270 255.580 584.590 255.640 ;
        RECT 65.390 255.440 584.590 255.580 ;
        RECT 65.390 255.380 65.710 255.440 ;
        RECT 584.270 255.380 584.590 255.440 ;
      LAYER via ;
        RECT 17.580 2974.020 17.840 2974.280 ;
        RECT 65.420 2974.020 65.680 2974.280 ;
        RECT 65.420 255.380 65.680 255.640 ;
        RECT 584.300 255.380 584.560 255.640 ;
      LAYER met2 ;
        RECT 17.570 2974.475 17.850 2974.845 ;
        RECT 17.640 2974.310 17.780 2974.475 ;
        RECT 17.580 2973.990 17.840 2974.310 ;
        RECT 65.420 2973.990 65.680 2974.310 ;
        RECT 65.480 255.670 65.620 2973.990 ;
        RECT 584.250 260.000 584.530 264.000 ;
        RECT 584.360 255.670 584.500 260.000 ;
        RECT 65.420 255.350 65.680 255.670 ;
        RECT 584.300 255.350 584.560 255.670 ;
      LAYER via2 ;
        RECT 17.570 2974.520 17.850 2974.800 ;
      LAYER met3 ;
        RECT -4.800 2974.810 2.400 2975.260 ;
        RECT 17.545 2974.810 17.875 2974.825 ;
        RECT -4.800 2974.510 17.875 2974.810 ;
        RECT -4.800 2974.060 2.400 2974.510 ;
        RECT 17.545 2974.495 17.875 2974.510 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2718.880 20.630 2718.940 ;
        RECT 169.810 2718.880 170.130 2718.940 ;
        RECT 20.310 2718.740 170.130 2718.880 ;
        RECT 20.310 2718.680 20.630 2718.740 ;
        RECT 169.810 2718.680 170.130 2718.740 ;
        RECT 169.810 1366.020 170.130 1366.080 ;
        RECT 296.770 1366.020 297.090 1366.080 ;
        RECT 169.810 1365.880 297.090 1366.020 ;
        RECT 169.810 1365.820 170.130 1365.880 ;
        RECT 296.770 1365.820 297.090 1365.880 ;
      LAYER via ;
        RECT 20.340 2718.680 20.600 2718.940 ;
        RECT 169.840 2718.680 170.100 2718.940 ;
        RECT 169.840 1365.820 170.100 1366.080 ;
        RECT 296.800 1365.820 297.060 1366.080 ;
      LAYER met2 ;
        RECT 20.330 2722.875 20.610 2723.245 ;
        RECT 20.400 2718.970 20.540 2722.875 ;
        RECT 20.340 2718.650 20.600 2718.970 ;
        RECT 169.840 2718.650 170.100 2718.970 ;
        RECT 169.900 1366.110 170.040 2718.650 ;
        RECT 169.840 1365.790 170.100 1366.110 ;
        RECT 296.800 1365.790 297.060 1366.110 ;
        RECT 296.860 1363.245 297.000 1365.790 ;
        RECT 296.790 1362.875 297.070 1363.245 ;
      LAYER via2 ;
        RECT 20.330 2722.920 20.610 2723.200 ;
        RECT 296.790 1362.920 297.070 1363.200 ;
      LAYER met3 ;
        RECT -4.800 2723.210 2.400 2723.660 ;
        RECT 20.305 2723.210 20.635 2723.225 ;
        RECT -4.800 2722.910 20.635 2723.210 ;
        RECT -4.800 2722.460 2.400 2722.910 ;
        RECT 20.305 2722.895 20.635 2722.910 ;
        RECT 296.765 1363.210 297.095 1363.225 ;
        RECT 310.000 1363.210 314.000 1363.600 ;
        RECT 296.765 1363.000 314.000 1363.210 ;
        RECT 296.765 1362.910 310.500 1363.000 ;
        RECT 296.765 1362.895 297.095 1362.910 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2606.910 2704.515 2607.190 2704.885 ;
        RECT 2606.980 2698.085 2607.120 2704.515 ;
        RECT 2606.910 2697.715 2607.190 2698.085 ;
        RECT 20.330 2476.715 20.610 2477.085 ;
        RECT 20.400 2471.645 20.540 2476.715 ;
        RECT 20.330 2471.275 20.610 2471.645 ;
      LAYER via2 ;
        RECT 2606.910 2704.560 2607.190 2704.840 ;
        RECT 2606.910 2697.760 2607.190 2698.040 ;
        RECT 20.330 2476.760 20.610 2477.040 ;
        RECT 20.330 2471.320 20.610 2471.600 ;
      LAYER met3 ;
        RECT 156.670 2705.530 157.050 2705.540 ;
        RECT 209.110 2705.530 209.490 2705.540 ;
        RECT 156.670 2705.230 209.490 2705.530 ;
        RECT 2606.000 2705.320 2610.000 2705.920 ;
        RECT 156.670 2705.220 157.050 2705.230 ;
        RECT 209.110 2705.220 209.490 2705.230 ;
        RECT 2606.670 2704.865 2606.970 2705.320 ;
        RECT 2606.670 2704.550 2607.215 2704.865 ;
        RECT 2606.885 2704.535 2607.215 2704.550 ;
        RECT 2606.885 2698.060 2607.215 2698.065 ;
        RECT 2606.630 2698.050 2607.215 2698.060 ;
        RECT 2606.430 2697.750 2607.215 2698.050 ;
        RECT 2606.630 2697.740 2607.215 2697.750 ;
        RECT 2606.885 2697.735 2607.215 2697.740 ;
        RECT 20.305 2477.050 20.635 2477.065 ;
        RECT 156.670 2477.050 157.050 2477.060 ;
        RECT 20.305 2476.750 157.050 2477.050 ;
        RECT 20.305 2476.735 20.635 2476.750 ;
        RECT 156.670 2476.740 157.050 2476.750 ;
        RECT -4.800 2471.610 2.400 2472.060 ;
        RECT 20.305 2471.610 20.635 2471.625 ;
        RECT -4.800 2471.310 20.635 2471.610 ;
        RECT -4.800 2470.860 2.400 2471.310 ;
        RECT 20.305 2471.295 20.635 2471.310 ;
      LAYER via3 ;
        RECT 156.700 2705.220 157.020 2705.540 ;
        RECT 209.140 2705.220 209.460 2705.540 ;
        RECT 2606.660 2697.740 2606.980 2698.060 ;
        RECT 156.700 2476.740 157.020 2477.060 ;
      LAYER met4 ;
        RECT 156.695 2705.215 157.025 2705.545 ;
        RECT 209.135 2705.215 209.465 2705.545 ;
        RECT 156.710 2477.065 157.010 2705.215 ;
        RECT 209.150 2698.490 209.450 2705.215 ;
        RECT 208.710 2697.310 209.890 2698.490 ;
        RECT 2606.230 2697.310 2607.410 2698.490 ;
        RECT 156.695 2476.735 157.025 2477.065 ;
      LAYER met5 ;
        RECT 313.380 2703.900 338.900 2705.500 ;
        RECT 313.380 2702.100 314.980 2703.900 ;
        RECT 240.700 2700.500 256.100 2702.100 ;
        RECT 240.700 2698.700 242.300 2700.500 ;
        RECT 208.500 2697.100 242.300 2698.700 ;
        RECT 254.500 2698.700 256.100 2700.500 ;
        RECT 288.540 2700.500 314.980 2702.100 ;
        RECT 288.540 2698.700 290.140 2700.500 ;
        RECT 254.500 2697.100 290.140 2698.700 ;
        RECT 337.300 2695.300 338.900 2703.900 ;
        RECT 481.740 2703.900 498.060 2705.500 ;
        RECT 481.740 2698.700 483.340 2703.900 ;
        RECT 496.460 2702.100 498.060 2703.900 ;
        RECT 496.460 2700.500 544.980 2702.100 ;
        RECT 372.260 2697.100 406.980 2698.700 ;
        RECT 337.300 2693.700 366.500 2695.300 ;
        RECT 364.900 2691.900 366.500 2693.700 ;
        RECT 372.260 2691.900 373.860 2697.100 ;
        RECT 405.380 2695.300 406.980 2697.100 ;
        RECT 409.060 2697.100 483.340 2698.700 ;
        RECT 543.380 2698.700 544.980 2700.500 ;
        RECT 603.180 2700.500 641.580 2702.100 ;
        RECT 543.380 2697.100 590.060 2698.700 ;
        RECT 409.060 2695.300 410.660 2697.100 ;
        RECT 405.380 2693.700 410.660 2695.300 ;
        RECT 364.900 2690.300 373.860 2691.900 ;
        RECT 588.460 2691.900 590.060 2697.100 ;
        RECT 603.180 2691.900 604.780 2700.500 ;
        RECT 639.980 2698.700 641.580 2700.500 ;
        RECT 699.780 2700.500 738.180 2702.100 ;
        RECT 639.980 2697.100 686.660 2698.700 ;
        RECT 588.460 2690.300 604.780 2691.900 ;
        RECT 685.060 2691.900 686.660 2697.100 ;
        RECT 699.780 2691.900 701.380 2700.500 ;
        RECT 736.580 2698.700 738.180 2700.500 ;
        RECT 796.380 2700.500 834.780 2702.100 ;
        RECT 736.580 2697.100 783.260 2698.700 ;
        RECT 685.060 2690.300 701.380 2691.900 ;
        RECT 781.660 2691.900 783.260 2697.100 ;
        RECT 796.380 2691.900 797.980 2700.500 ;
        RECT 833.180 2698.700 834.780 2700.500 ;
        RECT 892.980 2700.500 931.380 2702.100 ;
        RECT 833.180 2697.100 879.860 2698.700 ;
        RECT 781.660 2690.300 797.980 2691.900 ;
        RECT 878.260 2691.900 879.860 2697.100 ;
        RECT 892.980 2691.900 894.580 2700.500 ;
        RECT 929.780 2698.700 931.380 2700.500 ;
        RECT 989.580 2700.500 2404.300 2702.100 ;
        RECT 929.780 2697.100 976.460 2698.700 ;
        RECT 878.260 2690.300 894.580 2691.900 ;
        RECT 974.860 2691.900 976.460 2697.100 ;
        RECT 989.580 2691.900 991.180 2700.500 ;
        RECT 1026.380 2698.700 1027.980 2700.500 ;
        RECT 1076.060 2698.700 1077.660 2700.500 ;
        RECT 1026.380 2697.100 1077.660 2698.700 ;
        RECT 2402.700 2695.300 2404.300 2700.500 ;
        RECT 2414.660 2700.500 2450.300 2702.100 ;
        RECT 2414.660 2695.300 2416.260 2700.500 ;
        RECT 2402.700 2693.700 2416.260 2695.300 ;
        RECT 2448.700 2695.300 2450.300 2700.500 ;
        RECT 2495.620 2700.500 2500.900 2702.100 ;
        RECT 2495.620 2695.300 2497.220 2700.500 ;
        RECT 2448.700 2693.700 2497.220 2695.300 ;
        RECT 2499.300 2695.300 2500.900 2700.500 ;
        RECT 2512.180 2700.500 2559.780 2702.100 ;
        RECT 2512.180 2695.300 2513.780 2700.500 ;
        RECT 2558.180 2698.700 2559.780 2700.500 ;
        RECT 2558.180 2697.100 2607.620 2698.700 ;
        RECT 2499.300 2693.700 2513.780 2695.300 ;
        RECT 974.860 2690.300 991.180 2691.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2215.000 16.950 2215.060 ;
        RECT 168.890 2215.000 169.210 2215.060 ;
        RECT 16.630 2214.860 169.210 2215.000 ;
        RECT 16.630 2214.800 16.950 2214.860 ;
        RECT 168.890 2214.800 169.210 2214.860 ;
        RECT 168.890 248.100 169.210 248.160 ;
        RECT 870.390 248.100 870.710 248.160 ;
        RECT 168.890 247.960 870.710 248.100 ;
        RECT 168.890 247.900 169.210 247.960 ;
        RECT 870.390 247.900 870.710 247.960 ;
      LAYER via ;
        RECT 16.660 2214.800 16.920 2215.060 ;
        RECT 168.920 2214.800 169.180 2215.060 ;
        RECT 168.920 247.900 169.180 248.160 ;
        RECT 870.420 247.900 870.680 248.160 ;
      LAYER met2 ;
        RECT 16.650 2220.355 16.930 2220.725 ;
        RECT 16.720 2215.090 16.860 2220.355 ;
        RECT 16.660 2214.770 16.920 2215.090 ;
        RECT 168.920 2214.770 169.180 2215.090 ;
        RECT 168.980 248.190 169.120 2214.770 ;
        RECT 870.370 260.000 870.650 264.000 ;
        RECT 870.480 248.190 870.620 260.000 ;
        RECT 168.920 247.870 169.180 248.190 ;
        RECT 870.420 247.870 870.680 248.190 ;
      LAYER via2 ;
        RECT 16.650 2220.400 16.930 2220.680 ;
      LAYER met3 ;
        RECT -4.800 2220.690 2.400 2221.140 ;
        RECT 16.625 2220.690 16.955 2220.705 ;
        RECT -4.800 2220.390 16.955 2220.690 ;
        RECT -4.800 2219.940 2.400 2220.390 ;
        RECT 16.625 2220.375 16.955 2220.390 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2659.790 510.580 2660.110 510.640 ;
        RECT 2900.830 510.580 2901.150 510.640 ;
        RECT 2659.790 510.440 2901.150 510.580 ;
        RECT 2659.790 510.380 2660.110 510.440 ;
        RECT 2900.830 510.380 2901.150 510.440 ;
      LAYER via ;
        RECT 2659.820 510.380 2660.080 510.640 ;
        RECT 2900.860 510.380 2901.120 510.640 ;
      LAYER met2 ;
        RECT 2659.810 2815.355 2660.090 2815.725 ;
        RECT 2659.880 510.670 2660.020 2815.355 ;
        RECT 2659.820 510.350 2660.080 510.670 ;
        RECT 2900.860 510.350 2901.120 510.670 ;
        RECT 2900.920 508.485 2901.060 510.350 ;
        RECT 2900.850 508.115 2901.130 508.485 ;
      LAYER via2 ;
        RECT 2659.810 2815.400 2660.090 2815.680 ;
        RECT 2900.850 508.160 2901.130 508.440 ;
      LAYER met3 ;
        RECT 310.000 2820.920 314.000 2821.520 ;
        RECT 312.190 2818.420 312.490 2820.920 ;
        RECT 312.150 2818.100 312.530 2818.420 ;
        RECT 2606.630 2815.690 2607.010 2815.700 ;
        RECT 2659.785 2815.690 2660.115 2815.705 ;
        RECT 2606.630 2815.390 2660.115 2815.690 ;
        RECT 2606.630 2815.380 2607.010 2815.390 ;
        RECT 2659.785 2815.375 2660.115 2815.390 ;
        RECT 2606.630 2810.250 2607.010 2810.260 ;
        RECT 2611.230 2810.250 2611.610 2810.260 ;
        RECT 2606.630 2809.950 2611.610 2810.250 ;
        RECT 2606.630 2809.940 2607.010 2809.950 ;
        RECT 2611.230 2809.940 2611.610 2809.950 ;
        RECT 2900.825 508.450 2901.155 508.465 ;
        RECT 2917.600 508.450 2924.800 508.900 ;
        RECT 2900.825 508.150 2924.800 508.450 ;
        RECT 2900.825 508.135 2901.155 508.150 ;
        RECT 2917.600 507.700 2924.800 508.150 ;
      LAYER via3 ;
        RECT 312.180 2818.100 312.500 2818.420 ;
        RECT 2606.660 2815.380 2606.980 2815.700 ;
        RECT 2606.660 2809.940 2606.980 2810.260 ;
        RECT 2611.260 2809.940 2611.580 2810.260 ;
      LAYER met4 ;
        RECT 312.175 2818.095 312.505 2818.425 ;
        RECT 312.190 2814.090 312.490 2818.095 ;
        RECT 2606.655 2815.375 2606.985 2815.705 ;
        RECT 311.750 2812.910 312.930 2814.090 ;
        RECT 2606.670 2810.265 2606.970 2815.375 ;
        RECT 2606.655 2809.935 2606.985 2810.265 ;
        RECT 2610.830 2809.510 2612.010 2810.690 ;
      LAYER met5 ;
        RECT 311.540 2812.700 352.700 2814.300 ;
        RECT 351.100 2810.900 352.700 2812.700 ;
        RECT 393.420 2812.700 408.820 2814.300 ;
        RECT 393.420 2810.900 395.020 2812.700 ;
        RECT 351.100 2809.300 395.020 2810.900 ;
        RECT 407.220 2810.900 408.820 2812.700 ;
        RECT 515.780 2812.700 567.060 2814.300 ;
        RECT 407.220 2809.300 497.140 2810.900 ;
        RECT 495.540 2807.500 497.140 2809.300 ;
        RECT 515.780 2807.500 517.380 2812.700 ;
        RECT 495.540 2805.900 517.380 2807.500 ;
        RECT 565.460 2807.500 567.060 2812.700 ;
        RECT 612.380 2812.700 663.660 2814.300 ;
        RECT 612.380 2807.500 613.980 2812.700 ;
        RECT 565.460 2805.900 613.980 2807.500 ;
        RECT 662.060 2807.500 663.660 2812.700 ;
        RECT 708.980 2812.700 760.260 2814.300 ;
        RECT 708.980 2807.500 710.580 2812.700 ;
        RECT 662.060 2805.900 710.580 2807.500 ;
        RECT 758.660 2807.500 760.260 2812.700 ;
        RECT 805.580 2812.700 856.860 2814.300 ;
        RECT 805.580 2807.500 807.180 2812.700 ;
        RECT 758.660 2805.900 807.180 2807.500 ;
        RECT 855.260 2807.500 856.860 2812.700 ;
        RECT 902.180 2812.700 953.460 2814.300 ;
        RECT 902.180 2807.500 903.780 2812.700 ;
        RECT 855.260 2805.900 903.780 2807.500 ;
        RECT 951.860 2807.500 953.460 2812.700 ;
        RECT 998.780 2812.700 1050.060 2814.300 ;
        RECT 998.780 2807.500 1000.380 2812.700 ;
        RECT 951.860 2805.900 1000.380 2807.500 ;
        RECT 1048.460 2807.500 1050.060 2812.700 ;
        RECT 1095.380 2812.700 1146.660 2814.300 ;
        RECT 1095.380 2807.500 1096.980 2812.700 ;
        RECT 1048.460 2805.900 1096.980 2807.500 ;
        RECT 1145.060 2807.500 1146.660 2812.700 ;
        RECT 1191.980 2812.700 1243.260 2814.300 ;
        RECT 1191.980 2807.500 1193.580 2812.700 ;
        RECT 1145.060 2805.900 1193.580 2807.500 ;
        RECT 1241.660 2807.500 1243.260 2812.700 ;
        RECT 1288.580 2812.700 1339.860 2814.300 ;
        RECT 1288.580 2807.500 1290.180 2812.700 ;
        RECT 1241.660 2805.900 1290.180 2807.500 ;
        RECT 1338.260 2807.500 1339.860 2812.700 ;
        RECT 1385.180 2812.700 1436.460 2814.300 ;
        RECT 1385.180 2807.500 1386.780 2812.700 ;
        RECT 1338.260 2805.900 1386.780 2807.500 ;
        RECT 1434.860 2807.500 1436.460 2812.700 ;
        RECT 1481.780 2812.700 1533.060 2814.300 ;
        RECT 1481.780 2807.500 1483.380 2812.700 ;
        RECT 1434.860 2805.900 1483.380 2807.500 ;
        RECT 1531.460 2807.500 1533.060 2812.700 ;
        RECT 1578.380 2812.700 1629.660 2814.300 ;
        RECT 1578.380 2807.500 1579.980 2812.700 ;
        RECT 1531.460 2805.900 1579.980 2807.500 ;
        RECT 1628.060 2807.500 1629.660 2812.700 ;
        RECT 1674.980 2812.700 1726.260 2814.300 ;
        RECT 1674.980 2807.500 1676.580 2812.700 ;
        RECT 1628.060 2805.900 1676.580 2807.500 ;
        RECT 1724.660 2807.500 1726.260 2812.700 ;
        RECT 1771.580 2812.700 1822.860 2814.300 ;
        RECT 1771.580 2807.500 1773.180 2812.700 ;
        RECT 1724.660 2805.900 1773.180 2807.500 ;
        RECT 1821.260 2807.500 1822.860 2812.700 ;
        RECT 1868.180 2812.700 1919.460 2814.300 ;
        RECT 1868.180 2807.500 1869.780 2812.700 ;
        RECT 1821.260 2805.900 1869.780 2807.500 ;
        RECT 1917.860 2807.500 1919.460 2812.700 ;
        RECT 1964.780 2812.700 2016.060 2814.300 ;
        RECT 1964.780 2807.500 1966.380 2812.700 ;
        RECT 1917.860 2805.900 1966.380 2807.500 ;
        RECT 2014.460 2807.500 2016.060 2812.700 ;
        RECT 2061.380 2812.700 2112.660 2814.300 ;
        RECT 2061.380 2807.500 2062.980 2812.700 ;
        RECT 2014.460 2805.900 2062.980 2807.500 ;
        RECT 2111.060 2807.500 2112.660 2812.700 ;
        RECT 2157.980 2812.700 2209.260 2814.300 ;
        RECT 2157.980 2807.500 2159.580 2812.700 ;
        RECT 2111.060 2805.900 2159.580 2807.500 ;
        RECT 2207.660 2807.500 2209.260 2812.700 ;
        RECT 2254.580 2812.700 2305.860 2814.300 ;
        RECT 2254.580 2807.500 2256.180 2812.700 ;
        RECT 2207.660 2805.900 2256.180 2807.500 ;
        RECT 2304.260 2807.500 2305.860 2812.700 ;
        RECT 2351.180 2812.700 2381.300 2814.300 ;
        RECT 2351.180 2807.500 2352.780 2812.700 ;
        RECT 2379.700 2810.900 2381.300 2812.700 ;
        RECT 2447.780 2812.700 2477.900 2814.300 ;
        RECT 2379.700 2809.300 2429.140 2810.900 ;
        RECT 2304.260 2805.900 2352.780 2807.500 ;
        RECT 2427.540 2807.500 2429.140 2809.300 ;
        RECT 2447.780 2807.500 2449.380 2812.700 ;
        RECT 2476.300 2810.900 2477.900 2812.700 ;
        RECT 2476.300 2809.300 2612.220 2810.900 ;
        RECT 2427.540 2805.900 2449.380 2807.500 ;
        RECT 2524.140 2805.900 2526.660 2809.300 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 1966.800 20.630 1966.860 ;
        RECT 265.950 1966.800 266.270 1966.860 ;
        RECT 20.310 1966.660 266.270 1966.800 ;
        RECT 20.310 1966.600 20.630 1966.660 ;
        RECT 265.950 1966.600 266.270 1966.660 ;
        RECT 265.950 241.300 266.270 241.360 ;
        RECT 2033.730 241.300 2034.050 241.360 ;
        RECT 265.950 241.160 2034.050 241.300 ;
        RECT 265.950 241.100 266.270 241.160 ;
        RECT 2033.730 241.100 2034.050 241.160 ;
        RECT 2037.410 241.300 2037.730 241.360 ;
        RECT 2100.890 241.300 2101.210 241.360 ;
        RECT 2037.410 241.160 2101.210 241.300 ;
        RECT 2037.410 241.100 2037.730 241.160 ;
        RECT 2100.890 241.100 2101.210 241.160 ;
        RECT 2120.210 241.300 2120.530 241.360 ;
        RECT 2542.950 241.300 2543.270 241.360 ;
        RECT 2120.210 241.160 2543.270 241.300 ;
        RECT 2120.210 241.100 2120.530 241.160 ;
        RECT 2542.950 241.100 2543.270 241.160 ;
      LAYER via ;
        RECT 20.340 1966.600 20.600 1966.860 ;
        RECT 265.980 1966.600 266.240 1966.860 ;
        RECT 265.980 241.100 266.240 241.360 ;
        RECT 2033.760 241.100 2034.020 241.360 ;
        RECT 2037.440 241.100 2037.700 241.360 ;
        RECT 2100.920 241.100 2101.180 241.360 ;
        RECT 2120.240 241.100 2120.500 241.360 ;
        RECT 2542.980 241.100 2543.240 241.360 ;
      LAYER met2 ;
        RECT 20.330 1968.755 20.610 1969.125 ;
        RECT 20.400 1966.890 20.540 1968.755 ;
        RECT 20.340 1966.570 20.600 1966.890 ;
        RECT 265.980 1966.570 266.240 1966.890 ;
        RECT 266.040 241.390 266.180 1966.570 ;
        RECT 2542.930 260.000 2543.210 264.000 ;
        RECT 2543.040 241.390 2543.180 260.000 ;
        RECT 265.980 241.070 266.240 241.390 ;
        RECT 2033.760 241.070 2034.020 241.390 ;
        RECT 2037.440 241.070 2037.700 241.390 ;
        RECT 2100.920 241.070 2101.180 241.390 ;
        RECT 2120.240 241.070 2120.500 241.390 ;
        RECT 2542.980 241.070 2543.240 241.390 ;
        RECT 2033.820 240.565 2033.960 241.070 ;
        RECT 2037.500 240.565 2037.640 241.070 ;
        RECT 2100.980 240.565 2101.120 241.070 ;
        RECT 2120.300 240.565 2120.440 241.070 ;
        RECT 2033.750 240.195 2034.030 240.565 ;
        RECT 2037.430 240.195 2037.710 240.565 ;
        RECT 2100.910 240.195 2101.190 240.565 ;
        RECT 2120.230 240.195 2120.510 240.565 ;
      LAYER via2 ;
        RECT 20.330 1968.800 20.610 1969.080 ;
        RECT 2033.750 240.240 2034.030 240.520 ;
        RECT 2037.430 240.240 2037.710 240.520 ;
        RECT 2100.910 240.240 2101.190 240.520 ;
        RECT 2120.230 240.240 2120.510 240.520 ;
      LAYER met3 ;
        RECT -4.800 1969.090 2.400 1969.540 ;
        RECT 20.305 1969.090 20.635 1969.105 ;
        RECT -4.800 1968.790 20.635 1969.090 ;
        RECT -4.800 1968.340 2.400 1968.790 ;
        RECT 20.305 1968.775 20.635 1968.790 ;
        RECT 2033.725 240.530 2034.055 240.545 ;
        RECT 2037.405 240.530 2037.735 240.545 ;
        RECT 2033.725 240.230 2037.735 240.530 ;
        RECT 2033.725 240.215 2034.055 240.230 ;
        RECT 2037.405 240.215 2037.735 240.230 ;
        RECT 2100.885 240.530 2101.215 240.545 ;
        RECT 2120.205 240.530 2120.535 240.545 ;
        RECT 2100.885 240.230 2120.535 240.530 ;
        RECT 2100.885 240.215 2101.215 240.230 ;
        RECT 2120.205 240.215 2120.535 240.230 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 3266.620 45.010 3266.680 ;
        RECT 1134.430 3266.620 1134.750 3266.680 ;
        RECT 44.690 3266.480 1134.750 3266.620 ;
        RECT 44.690 3266.420 45.010 3266.480 ;
        RECT 1134.430 3266.420 1134.750 3266.480 ;
        RECT 20.310 1717.580 20.630 1717.640 ;
        RECT 44.690 1717.580 45.010 1717.640 ;
        RECT 20.310 1717.440 45.010 1717.580 ;
        RECT 20.310 1717.380 20.630 1717.440 ;
        RECT 44.690 1717.380 45.010 1717.440 ;
      LAYER via ;
        RECT 44.720 3266.420 44.980 3266.680 ;
        RECT 1134.460 3266.420 1134.720 3266.680 ;
        RECT 20.340 1717.380 20.600 1717.640 ;
        RECT 44.720 1717.380 44.980 1717.640 ;
      LAYER met2 ;
        RECT 44.720 3266.390 44.980 3266.710 ;
        RECT 1134.460 3266.390 1134.720 3266.710 ;
        RECT 44.780 1717.670 44.920 3266.390 ;
        RECT 1134.520 3260.000 1134.660 3266.390 ;
        RECT 1134.410 3256.000 1134.690 3260.000 ;
        RECT 20.340 1717.525 20.600 1717.670 ;
        RECT 20.330 1717.155 20.610 1717.525 ;
        RECT 44.720 1717.350 44.980 1717.670 ;
      LAYER via2 ;
        RECT 20.330 1717.200 20.610 1717.480 ;
      LAYER met3 ;
        RECT -4.800 1717.490 2.400 1717.940 ;
        RECT 20.305 1717.490 20.635 1717.505 ;
        RECT -4.800 1717.190 20.635 1717.490 ;
        RECT -4.800 1716.740 2.400 1717.190 ;
        RECT 20.305 1717.175 20.635 1717.190 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 1462.920 20.630 1462.980 ;
        RECT 169.350 1462.920 169.670 1462.980 ;
        RECT 20.310 1462.780 169.670 1462.920 ;
        RECT 20.310 1462.720 20.630 1462.780 ;
        RECT 169.350 1462.720 169.670 1462.780 ;
        RECT 169.350 455.160 169.670 455.220 ;
        RECT 296.770 455.160 297.090 455.220 ;
        RECT 169.350 455.020 297.090 455.160 ;
        RECT 169.350 454.960 169.670 455.020 ;
        RECT 296.770 454.960 297.090 455.020 ;
      LAYER via ;
        RECT 20.340 1462.720 20.600 1462.980 ;
        RECT 169.380 1462.720 169.640 1462.980 ;
        RECT 169.380 454.960 169.640 455.220 ;
        RECT 296.800 454.960 297.060 455.220 ;
      LAYER met2 ;
        RECT 20.330 1466.235 20.610 1466.605 ;
        RECT 20.400 1463.010 20.540 1466.235 ;
        RECT 20.340 1462.690 20.600 1463.010 ;
        RECT 169.380 1462.690 169.640 1463.010 ;
        RECT 169.440 455.250 169.580 1462.690 ;
        RECT 169.380 454.930 169.640 455.250 ;
        RECT 296.800 454.930 297.060 455.250 ;
        RECT 296.860 453.405 297.000 454.930 ;
        RECT 296.790 453.035 297.070 453.405 ;
      LAYER via2 ;
        RECT 20.330 1466.280 20.610 1466.560 ;
        RECT 296.790 453.080 297.070 453.360 ;
      LAYER met3 ;
        RECT -4.800 1466.570 2.400 1467.020 ;
        RECT 20.305 1466.570 20.635 1466.585 ;
        RECT -4.800 1466.270 20.635 1466.570 ;
        RECT -4.800 1465.820 2.400 1466.270 ;
        RECT 20.305 1466.255 20.635 1466.270 ;
        RECT 296.765 453.370 297.095 453.385 ;
        RECT 310.000 453.370 314.000 453.760 ;
        RECT 296.765 453.160 314.000 453.370 ;
        RECT 296.765 453.070 310.500 453.160 ;
        RECT 296.765 453.055 297.095 453.070 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.290 3265.940 141.610 3266.000 ;
        RECT 1248.510 3265.940 1248.830 3266.000 ;
        RECT 141.290 3265.800 1248.830 3265.940 ;
        RECT 141.290 3265.740 141.610 3265.800 ;
        RECT 1248.510 3265.740 1248.830 3265.800 ;
        RECT 20.310 1221.180 20.630 1221.240 ;
        RECT 141.290 1221.180 141.610 1221.240 ;
        RECT 20.310 1221.040 141.610 1221.180 ;
        RECT 20.310 1220.980 20.630 1221.040 ;
        RECT 141.290 1220.980 141.610 1221.040 ;
      LAYER via ;
        RECT 141.320 3265.740 141.580 3266.000 ;
        RECT 1248.540 3265.740 1248.800 3266.000 ;
        RECT 20.340 1220.980 20.600 1221.240 ;
        RECT 141.320 1220.980 141.580 1221.240 ;
      LAYER met2 ;
        RECT 141.320 3265.710 141.580 3266.030 ;
        RECT 1248.540 3265.710 1248.800 3266.030 ;
        RECT 141.380 1221.270 141.520 3265.710 ;
        RECT 1248.600 3260.000 1248.740 3265.710 ;
        RECT 1248.490 3256.000 1248.770 3260.000 ;
        RECT 20.340 1220.950 20.600 1221.270 ;
        RECT 141.320 1220.950 141.580 1221.270 ;
        RECT 20.400 1215.005 20.540 1220.950 ;
        RECT 20.330 1214.635 20.610 1215.005 ;
      LAYER via2 ;
        RECT 20.330 1214.680 20.610 1214.960 ;
      LAYER met3 ;
        RECT -4.800 1214.970 2.400 1215.420 ;
        RECT 20.305 1214.970 20.635 1214.985 ;
        RECT -4.800 1214.670 20.635 1214.970 ;
        RECT -4.800 1214.220 2.400 1214.670 ;
        RECT 20.305 1214.655 20.635 1214.670 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 237.890 3267.300 238.210 3267.360 ;
        RECT 1076.470 3267.300 1076.790 3267.360 ;
        RECT 237.890 3267.160 1076.790 3267.300 ;
        RECT 237.890 3267.100 238.210 3267.160 ;
        RECT 1076.470 3267.100 1076.790 3267.160 ;
        RECT 18.930 965.840 19.250 965.900 ;
        RECT 237.890 965.840 238.210 965.900 ;
        RECT 18.930 965.700 238.210 965.840 ;
        RECT 18.930 965.640 19.250 965.700 ;
        RECT 237.890 965.640 238.210 965.700 ;
      LAYER via ;
        RECT 237.920 3267.100 238.180 3267.360 ;
        RECT 1076.500 3267.100 1076.760 3267.360 ;
        RECT 18.960 965.640 19.220 965.900 ;
        RECT 237.920 965.640 238.180 965.900 ;
      LAYER met2 ;
        RECT 237.920 3267.070 238.180 3267.390 ;
        RECT 1076.500 3267.070 1076.760 3267.390 ;
        RECT 237.980 965.930 238.120 3267.070 ;
        RECT 1076.560 3260.000 1076.700 3267.070 ;
        RECT 1076.450 3256.000 1076.730 3260.000 ;
        RECT 18.960 965.610 19.220 965.930 ;
        RECT 237.920 965.610 238.180 965.930 ;
        RECT 19.020 963.405 19.160 965.610 ;
        RECT 18.950 963.035 19.230 963.405 ;
      LAYER via2 ;
        RECT 18.950 963.080 19.230 963.360 ;
      LAYER met3 ;
        RECT -4.800 963.370 2.400 963.820 ;
        RECT 18.925 963.370 19.255 963.385 ;
        RECT -4.800 963.070 19.255 963.370 ;
        RECT -4.800 962.620 2.400 963.070 ;
        RECT 18.925 963.055 19.255 963.070 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 710.840 16.950 710.900 ;
        RECT 265.030 710.840 265.350 710.900 ;
        RECT 16.630 710.700 265.350 710.840 ;
        RECT 16.630 710.640 16.950 710.700 ;
        RECT 265.030 710.640 265.350 710.700 ;
        RECT 265.030 248.440 265.350 248.500 ;
        RECT 1484.950 248.440 1485.270 248.500 ;
        RECT 265.030 248.300 1485.270 248.440 ;
        RECT 265.030 248.240 265.350 248.300 ;
        RECT 1484.950 248.240 1485.270 248.300 ;
      LAYER via ;
        RECT 16.660 710.640 16.920 710.900 ;
        RECT 265.060 710.640 265.320 710.900 ;
        RECT 265.060 248.240 265.320 248.500 ;
        RECT 1484.980 248.240 1485.240 248.500 ;
      LAYER met2 ;
        RECT 16.650 711.435 16.930 711.805 ;
        RECT 16.720 710.930 16.860 711.435 ;
        RECT 16.660 710.610 16.920 710.930 ;
        RECT 265.060 710.610 265.320 710.930 ;
        RECT 265.120 248.530 265.260 710.610 ;
        RECT 1484.930 260.000 1485.210 264.000 ;
        RECT 1485.040 248.530 1485.180 260.000 ;
        RECT 265.060 248.210 265.320 248.530 ;
        RECT 1484.980 248.210 1485.240 248.530 ;
      LAYER via2 ;
        RECT 16.650 711.480 16.930 711.760 ;
      LAYER met3 ;
        RECT -4.800 711.770 2.400 712.220 ;
        RECT 16.625 711.770 16.955 711.785 ;
        RECT -4.800 711.470 16.955 711.770 ;
        RECT -4.800 711.020 2.400 711.470 ;
        RECT 16.625 711.455 16.955 711.470 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 193.470 2772.850 193.850 2772.860 ;
        RECT 207.270 2772.850 207.650 2772.860 ;
        RECT 193.470 2772.550 207.650 2772.850 ;
        RECT 193.470 2772.540 193.850 2772.550 ;
        RECT 207.270 2772.540 207.650 2772.550 ;
        RECT 154.830 2769.450 155.210 2769.460 ;
        RECT 178.750 2769.450 179.130 2769.460 ;
        RECT 154.830 2769.150 179.130 2769.450 ;
        RECT 2606.000 2769.450 2610.000 2769.840 ;
        RECT 2611.230 2769.450 2611.610 2769.460 ;
        RECT 2606.000 2769.240 2611.610 2769.450 ;
        RECT 2609.580 2769.150 2611.610 2769.240 ;
        RECT 154.830 2769.140 155.210 2769.150 ;
        RECT 178.750 2769.140 179.130 2769.150 ;
        RECT 2611.230 2769.140 2611.610 2769.150 ;
        RECT 154.830 462.210 155.210 462.220 ;
        RECT 3.070 461.910 155.210 462.210 ;
        RECT -4.800 460.850 2.400 461.300 ;
        RECT 3.070 460.850 3.370 461.910 ;
        RECT 154.830 461.900 155.210 461.910 ;
        RECT -4.800 460.550 3.370 460.850 ;
        RECT -4.800 460.100 2.400 460.550 ;
      LAYER via3 ;
        RECT 193.500 2772.540 193.820 2772.860 ;
        RECT 207.300 2772.540 207.620 2772.860 ;
        RECT 154.860 2769.140 155.180 2769.460 ;
        RECT 178.780 2769.140 179.100 2769.460 ;
        RECT 2611.260 2769.140 2611.580 2769.460 ;
        RECT 154.860 461.900 155.180 462.220 ;
      LAYER met4 ;
        RECT 193.070 2772.110 194.250 2773.290 ;
        RECT 206.870 2772.110 208.050 2773.290 ;
        RECT 154.855 2769.135 155.185 2769.465 ;
        RECT 154.870 462.225 155.170 2769.135 ;
        RECT 178.350 2768.710 179.530 2769.890 ;
        RECT 2610.830 2768.710 2612.010 2769.890 ;
        RECT 154.855 461.895 155.185 462.225 ;
      LAYER met5 ;
        RECT 239.780 2775.300 289.220 2776.900 ;
        RECT 239.780 2773.500 241.380 2775.300 ;
        RECT 179.060 2771.900 194.460 2773.500 ;
        RECT 206.660 2771.900 241.380 2773.500 ;
        RECT 179.060 2770.100 180.660 2771.900 ;
        RECT 177.360 2768.500 180.660 2770.100 ;
        RECT 287.620 2770.100 289.220 2775.300 ;
        RECT 337.300 2775.300 355.460 2776.900 ;
        RECT 337.300 2770.100 338.900 2775.300 ;
        RECT 287.620 2768.500 338.900 2770.100 ;
        RECT 353.860 2770.100 355.460 2775.300 ;
        RECT 444.940 2775.300 497.140 2776.900 ;
        RECT 444.940 2773.500 446.540 2775.300 ;
        RECT 416.420 2771.900 446.540 2773.500 ;
        RECT 416.420 2770.100 418.020 2771.900 ;
        RECT 353.860 2768.500 418.020 2770.100 ;
        RECT 495.540 2770.100 497.140 2775.300 ;
        RECT 516.700 2775.300 566.140 2776.900 ;
        RECT 516.700 2770.100 518.300 2775.300 ;
        RECT 495.540 2768.500 518.300 2770.100 ;
        RECT 564.540 2770.100 566.140 2775.300 ;
        RECT 613.300 2775.300 662.740 2776.900 ;
        RECT 613.300 2770.100 614.900 2775.300 ;
        RECT 564.540 2768.500 614.900 2770.100 ;
        RECT 661.140 2770.100 662.740 2775.300 ;
        RECT 709.900 2775.300 759.340 2776.900 ;
        RECT 709.900 2770.100 711.500 2775.300 ;
        RECT 661.140 2768.500 711.500 2770.100 ;
        RECT 757.740 2770.100 759.340 2775.300 ;
        RECT 806.500 2775.300 855.940 2776.900 ;
        RECT 806.500 2770.100 808.100 2775.300 ;
        RECT 757.740 2768.500 808.100 2770.100 ;
        RECT 854.340 2770.100 855.940 2775.300 ;
        RECT 903.100 2775.300 952.540 2776.900 ;
        RECT 903.100 2770.100 904.700 2775.300 ;
        RECT 854.340 2768.500 904.700 2770.100 ;
        RECT 950.940 2770.100 952.540 2775.300 ;
        RECT 999.700 2775.300 1049.140 2776.900 ;
        RECT 999.700 2770.100 1001.300 2775.300 ;
        RECT 950.940 2768.500 1001.300 2770.100 ;
        RECT 1047.540 2770.100 1049.140 2775.300 ;
        RECT 1096.300 2775.300 1145.740 2776.900 ;
        RECT 1096.300 2770.100 1097.900 2775.300 ;
        RECT 1047.540 2768.500 1097.900 2770.100 ;
        RECT 1144.140 2770.100 1145.740 2775.300 ;
        RECT 1192.900 2775.300 1242.340 2776.900 ;
        RECT 1192.900 2770.100 1194.500 2775.300 ;
        RECT 1144.140 2768.500 1194.500 2770.100 ;
        RECT 1240.740 2770.100 1242.340 2775.300 ;
        RECT 1289.500 2775.300 1338.940 2776.900 ;
        RECT 1289.500 2770.100 1291.100 2775.300 ;
        RECT 1240.740 2768.500 1291.100 2770.100 ;
        RECT 1337.340 2770.100 1338.940 2775.300 ;
        RECT 1386.100 2775.300 1435.540 2776.900 ;
        RECT 1386.100 2770.100 1387.700 2775.300 ;
        RECT 1337.340 2768.500 1387.700 2770.100 ;
        RECT 1433.940 2770.100 1435.540 2775.300 ;
        RECT 1482.700 2775.300 1532.140 2776.900 ;
        RECT 1482.700 2770.100 1484.300 2775.300 ;
        RECT 1433.940 2768.500 1484.300 2770.100 ;
        RECT 1530.540 2770.100 1532.140 2775.300 ;
        RECT 1579.300 2775.300 1628.740 2776.900 ;
        RECT 1579.300 2770.100 1580.900 2775.300 ;
        RECT 1530.540 2768.500 1580.900 2770.100 ;
        RECT 1627.140 2770.100 1628.740 2775.300 ;
        RECT 1675.900 2775.300 1725.340 2776.900 ;
        RECT 1675.900 2770.100 1677.500 2775.300 ;
        RECT 1627.140 2768.500 1677.500 2770.100 ;
        RECT 1723.740 2770.100 1725.340 2775.300 ;
        RECT 1772.500 2775.300 1821.940 2776.900 ;
        RECT 1772.500 2770.100 1774.100 2775.300 ;
        RECT 1723.740 2768.500 1774.100 2770.100 ;
        RECT 1820.340 2770.100 1821.940 2775.300 ;
        RECT 1869.100 2775.300 1918.540 2776.900 ;
        RECT 1869.100 2770.100 1870.700 2775.300 ;
        RECT 1820.340 2768.500 1870.700 2770.100 ;
        RECT 1916.940 2770.100 1918.540 2775.300 ;
        RECT 1965.700 2775.300 2015.140 2776.900 ;
        RECT 1965.700 2770.100 1967.300 2775.300 ;
        RECT 1916.940 2768.500 1967.300 2770.100 ;
        RECT 2013.540 2770.100 2015.140 2775.300 ;
        RECT 2062.300 2775.300 2111.740 2776.900 ;
        RECT 2062.300 2770.100 2063.900 2775.300 ;
        RECT 2013.540 2768.500 2063.900 2770.100 ;
        RECT 2110.140 2770.100 2111.740 2775.300 ;
        RECT 2158.900 2775.300 2208.340 2776.900 ;
        RECT 2158.900 2770.100 2160.500 2775.300 ;
        RECT 2110.140 2768.500 2160.500 2770.100 ;
        RECT 2206.740 2770.100 2208.340 2775.300 ;
        RECT 2255.500 2775.300 2304.940 2776.900 ;
        RECT 2255.500 2770.100 2257.100 2775.300 ;
        RECT 2206.740 2768.500 2257.100 2770.100 ;
        RECT 2303.340 2770.100 2304.940 2775.300 ;
        RECT 2352.100 2775.300 2429.140 2776.900 ;
        RECT 2352.100 2770.100 2353.700 2775.300 ;
        RECT 2303.340 2768.500 2353.700 2770.100 ;
        RECT 2427.540 2770.100 2429.140 2775.300 ;
        RECT 2448.700 2775.300 2525.740 2776.900 ;
        RECT 2448.700 2770.100 2450.300 2775.300 ;
        RECT 2427.540 2768.500 2450.300 2770.100 ;
        RECT 2524.140 2773.500 2525.740 2775.300 ;
        RECT 2571.980 2775.300 2594.740 2776.900 ;
        RECT 2571.980 2773.500 2573.580 2775.300 ;
        RECT 2524.140 2771.900 2573.580 2773.500 ;
        RECT 2524.140 2768.500 2526.660 2771.900 ;
        RECT 2593.140 2770.100 2594.740 2775.300 ;
        RECT 2593.140 2768.500 2612.220 2770.100 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1991.890 3272.315 1992.170 3272.685 ;
        RECT 2478.570 3272.315 2478.850 3272.685 ;
        RECT 1991.960 3267.245 1992.100 3272.315 ;
        RECT 17.110 3266.875 17.390 3267.245 ;
        RECT 1991.890 3266.875 1992.170 3267.245 ;
        RECT 17.180 209.285 17.320 3266.875 ;
        RECT 2478.640 3260.000 2478.780 3272.315 ;
        RECT 2478.530 3256.000 2478.810 3260.000 ;
        RECT 17.110 208.915 17.390 209.285 ;
      LAYER via2 ;
        RECT 1991.890 3272.360 1992.170 3272.640 ;
        RECT 2478.570 3272.360 2478.850 3272.640 ;
        RECT 17.110 3266.920 17.390 3267.200 ;
        RECT 1991.890 3266.920 1992.170 3267.200 ;
        RECT 17.110 208.960 17.390 209.240 ;
      LAYER met3 ;
        RECT 1991.865 3272.650 1992.195 3272.665 ;
        RECT 2478.545 3272.650 2478.875 3272.665 ;
        RECT 1991.865 3272.350 2478.875 3272.650 ;
        RECT 1991.865 3272.335 1992.195 3272.350 ;
        RECT 2478.545 3272.335 2478.875 3272.350 ;
        RECT 17.085 3267.210 17.415 3267.225 ;
        RECT 1991.865 3267.210 1992.195 3267.225 ;
        RECT 17.085 3266.910 1992.195 3267.210 ;
        RECT 17.085 3266.895 17.415 3266.910 ;
        RECT 1991.865 3266.895 1992.195 3266.910 ;
        RECT -4.800 209.250 2.400 209.700 ;
        RECT 17.085 209.250 17.415 209.265 ;
        RECT -4.800 208.950 17.415 209.250 ;
        RECT -4.800 208.500 2.400 208.950 ;
        RECT 17.085 208.935 17.415 208.950 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2111.640 2615.490 2111.700 ;
        RECT 2694.750 2111.640 2695.070 2111.700 ;
        RECT 2615.170 2111.500 2695.070 2111.640 ;
        RECT 2615.170 2111.440 2615.490 2111.500 ;
        RECT 2694.750 2111.440 2695.070 2111.500 ;
        RECT 2694.750 745.180 2695.070 745.240 ;
        RECT 2900.830 745.180 2901.150 745.240 ;
        RECT 2694.750 745.040 2901.150 745.180 ;
        RECT 2694.750 744.980 2695.070 745.040 ;
        RECT 2900.830 744.980 2901.150 745.040 ;
      LAYER via ;
        RECT 2615.200 2111.440 2615.460 2111.700 ;
        RECT 2694.780 2111.440 2695.040 2111.700 ;
        RECT 2694.780 744.980 2695.040 745.240 ;
        RECT 2900.860 744.980 2901.120 745.240 ;
      LAYER met2 ;
        RECT 2615.190 2113.595 2615.470 2113.965 ;
        RECT 2615.260 2111.730 2615.400 2113.595 ;
        RECT 2615.200 2111.410 2615.460 2111.730 ;
        RECT 2694.780 2111.410 2695.040 2111.730 ;
        RECT 2694.840 745.270 2694.980 2111.410 ;
        RECT 2694.780 744.950 2695.040 745.270 ;
        RECT 2900.860 744.950 2901.120 745.270 ;
        RECT 2900.920 743.085 2901.060 744.950 ;
        RECT 2900.850 742.715 2901.130 743.085 ;
      LAYER via2 ;
        RECT 2615.190 2113.640 2615.470 2113.920 ;
        RECT 2900.850 742.760 2901.130 743.040 ;
      LAYER met3 ;
        RECT 2606.000 2113.930 2610.000 2114.320 ;
        RECT 2615.165 2113.930 2615.495 2113.945 ;
        RECT 2606.000 2113.720 2615.495 2113.930 ;
        RECT 2609.580 2113.630 2615.495 2113.720 ;
        RECT 2615.165 2113.615 2615.495 2113.630 ;
        RECT 2900.825 743.050 2901.155 743.065 ;
        RECT 2917.600 743.050 2924.800 743.500 ;
        RECT 2900.825 742.750 2924.800 743.050 ;
        RECT 2900.825 742.735 2901.155 742.750 ;
        RECT 2917.600 742.300 2924.800 742.750 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2674.510 972.980 2674.830 973.040 ;
        RECT 2900.830 972.980 2901.150 973.040 ;
        RECT 2674.510 972.840 2901.150 972.980 ;
        RECT 2674.510 972.780 2674.830 972.840 ;
        RECT 2900.830 972.780 2901.150 972.840 ;
        RECT 1255.870 253.540 1256.190 253.600 ;
        RECT 2674.510 253.540 2674.830 253.600 ;
        RECT 1255.870 253.400 2674.830 253.540 ;
        RECT 1255.870 253.340 1256.190 253.400 ;
        RECT 2674.510 253.340 2674.830 253.400 ;
      LAYER via ;
        RECT 2674.540 972.780 2674.800 973.040 ;
        RECT 2900.860 972.780 2901.120 973.040 ;
        RECT 1255.900 253.340 1256.160 253.600 ;
        RECT 2674.540 253.340 2674.800 253.600 ;
      LAYER met2 ;
        RECT 2900.850 977.315 2901.130 977.685 ;
        RECT 2900.920 973.070 2901.060 977.315 ;
        RECT 2674.540 972.750 2674.800 973.070 ;
        RECT 2900.860 972.750 2901.120 973.070 ;
        RECT 1255.850 260.000 1256.130 264.000 ;
        RECT 1255.960 253.630 1256.100 260.000 ;
        RECT 2674.600 253.630 2674.740 972.750 ;
        RECT 1255.900 253.310 1256.160 253.630 ;
        RECT 2674.540 253.310 2674.800 253.630 ;
      LAYER via2 ;
        RECT 2900.850 977.360 2901.130 977.640 ;
      LAYER met3 ;
        RECT 2900.825 977.650 2901.155 977.665 ;
        RECT 2917.600 977.650 2924.800 978.100 ;
        RECT 2900.825 977.350 2924.800 977.650 ;
        RECT 2900.825 977.335 2901.155 977.350 ;
        RECT 2917.600 976.900 2924.800 977.350 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2680.950 1207.580 2681.270 1207.640 ;
        RECT 2900.830 1207.580 2901.150 1207.640 ;
        RECT 2680.950 1207.440 2901.150 1207.580 ;
        RECT 2680.950 1207.380 2681.270 1207.440 ;
        RECT 2900.830 1207.380 2901.150 1207.440 ;
        RECT 684.550 240.960 684.870 241.020 ;
        RECT 2680.950 240.960 2681.270 241.020 ;
        RECT 684.550 240.820 2681.270 240.960 ;
        RECT 684.550 240.760 684.870 240.820 ;
        RECT 2680.950 240.760 2681.270 240.820 ;
      LAYER via ;
        RECT 2680.980 1207.380 2681.240 1207.640 ;
        RECT 2900.860 1207.380 2901.120 1207.640 ;
        RECT 684.580 240.760 684.840 241.020 ;
        RECT 2680.980 240.760 2681.240 241.020 ;
      LAYER met2 ;
        RECT 2900.850 1211.915 2901.130 1212.285 ;
        RECT 2900.920 1207.670 2901.060 1211.915 ;
        RECT 2680.980 1207.350 2681.240 1207.670 ;
        RECT 2900.860 1207.350 2901.120 1207.670 ;
        RECT 684.530 260.000 684.810 264.000 ;
        RECT 684.640 241.050 684.780 260.000 ;
        RECT 2681.040 241.050 2681.180 1207.350 ;
        RECT 684.580 240.730 684.840 241.050 ;
        RECT 2680.980 240.730 2681.240 241.050 ;
      LAYER via2 ;
        RECT 2900.850 1211.960 2901.130 1212.240 ;
      LAYER met3 ;
        RECT 2900.825 1212.250 2901.155 1212.265 ;
        RECT 2917.600 1212.250 2924.800 1212.700 ;
        RECT 2900.825 1211.950 2924.800 1212.250 ;
        RECT 2900.825 1211.935 2901.155 1211.950 ;
        RECT 2917.600 1211.500 2924.800 1211.950 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2606.430 3271.720 2606.750 3271.780 ;
        RECT 2860.350 3271.720 2860.670 3271.780 ;
        RECT 2606.430 3271.580 2860.670 3271.720 ;
        RECT 2606.430 3271.520 2606.750 3271.580 ;
        RECT 2860.350 3271.520 2860.670 3271.580 ;
        RECT 2860.350 1448.980 2860.670 1449.040 ;
        RECT 2900.830 1448.980 2901.150 1449.040 ;
        RECT 2860.350 1448.840 2901.150 1448.980 ;
        RECT 2860.350 1448.780 2860.670 1448.840 ;
        RECT 2900.830 1448.780 2901.150 1448.840 ;
      LAYER via ;
        RECT 2606.460 3271.520 2606.720 3271.780 ;
        RECT 2860.380 3271.520 2860.640 3271.780 ;
        RECT 2860.380 1448.780 2860.640 1449.040 ;
        RECT 2900.860 1448.780 2901.120 1449.040 ;
      LAYER met2 ;
        RECT 2606.460 3271.490 2606.720 3271.810 ;
        RECT 2860.380 3271.490 2860.640 3271.810 ;
        RECT 2606.520 3260.000 2606.660 3271.490 ;
        RECT 2606.410 3256.000 2606.690 3260.000 ;
        RECT 2860.440 1449.070 2860.580 3271.490 ;
        RECT 2860.380 1448.750 2860.640 1449.070 ;
        RECT 2900.860 1448.750 2901.120 1449.070 ;
        RECT 2900.920 1446.885 2901.060 1448.750 ;
        RECT 2900.850 1446.515 2901.130 1446.885 ;
      LAYER via2 ;
        RECT 2900.850 1446.560 2901.130 1446.840 ;
      LAYER met3 ;
        RECT 2900.825 1446.850 2901.155 1446.865 ;
        RECT 2917.600 1446.850 2924.800 1447.300 ;
        RECT 2900.825 1446.550 2924.800 1446.850 ;
        RECT 2900.825 1446.535 2901.155 1446.550 ;
        RECT 2917.600 1446.100 2924.800 1446.550 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1506.110 3265.600 1506.430 3265.660 ;
        RECT 2749.950 3265.600 2750.270 3265.660 ;
        RECT 1506.110 3265.460 2750.270 3265.600 ;
        RECT 1506.110 3265.400 1506.430 3265.460 ;
        RECT 2749.950 3265.400 2750.270 3265.460 ;
        RECT 2749.950 1683.580 2750.270 1683.640 ;
        RECT 2900.830 1683.580 2901.150 1683.640 ;
        RECT 2749.950 1683.440 2901.150 1683.580 ;
        RECT 2749.950 1683.380 2750.270 1683.440 ;
        RECT 2900.830 1683.380 2901.150 1683.440 ;
      LAYER via ;
        RECT 1506.140 3265.400 1506.400 3265.660 ;
        RECT 2749.980 3265.400 2750.240 3265.660 ;
        RECT 2749.980 1683.380 2750.240 1683.640 ;
        RECT 2900.860 1683.380 2901.120 1683.640 ;
      LAYER met2 ;
        RECT 1506.140 3265.370 1506.400 3265.690 ;
        RECT 2749.980 3265.370 2750.240 3265.690 ;
        RECT 1506.200 3260.000 1506.340 3265.370 ;
        RECT 1506.090 3256.000 1506.370 3260.000 ;
        RECT 2750.040 1683.670 2750.180 3265.370 ;
        RECT 2749.980 1683.350 2750.240 1683.670 ;
        RECT 2900.860 1683.350 2901.120 1683.670 ;
        RECT 2900.920 1681.485 2901.060 1683.350 ;
        RECT 2900.850 1681.115 2901.130 1681.485 ;
      LAYER via2 ;
        RECT 2900.850 1681.160 2901.130 1681.440 ;
      LAYER met3 ;
        RECT 2900.825 1681.450 2901.155 1681.465 ;
        RECT 2917.600 1681.450 2924.800 1681.900 ;
        RECT 2900.825 1681.150 2924.800 1681.450 ;
        RECT 2900.825 1681.135 2901.155 1681.150 ;
        RECT 2917.600 1680.700 2924.800 1681.150 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 333.110 3263.900 333.430 3263.960 ;
        RECT 2846.550 3263.900 2846.870 3263.960 ;
        RECT 333.110 3263.760 2846.870 3263.900 ;
        RECT 333.110 3263.700 333.430 3263.760 ;
        RECT 2846.550 3263.700 2846.870 3263.760 ;
        RECT 2846.550 1918.180 2846.870 1918.240 ;
        RECT 2900.830 1918.180 2901.150 1918.240 ;
        RECT 2846.550 1918.040 2901.150 1918.180 ;
        RECT 2846.550 1917.980 2846.870 1918.040 ;
        RECT 2900.830 1917.980 2901.150 1918.040 ;
      LAYER via ;
        RECT 333.140 3263.700 333.400 3263.960 ;
        RECT 2846.580 3263.700 2846.840 3263.960 ;
        RECT 2846.580 1917.980 2846.840 1918.240 ;
        RECT 2900.860 1917.980 2901.120 1918.240 ;
      LAYER met2 ;
        RECT 333.140 3263.670 333.400 3263.990 ;
        RECT 2846.580 3263.670 2846.840 3263.990 ;
        RECT 333.200 3260.000 333.340 3263.670 ;
        RECT 333.090 3256.000 333.370 3260.000 ;
        RECT 2846.640 1918.270 2846.780 3263.670 ;
        RECT 2846.580 1917.950 2846.840 1918.270 ;
        RECT 2900.860 1917.950 2901.120 1918.270 ;
        RECT 2900.920 1916.085 2901.060 1917.950 ;
        RECT 2900.850 1915.715 2901.130 1916.085 ;
      LAYER via2 ;
        RECT 2900.850 1915.760 2901.130 1916.040 ;
      LAYER met3 ;
        RECT 2900.825 1916.050 2901.155 1916.065 ;
        RECT 2917.600 1916.050 2924.800 1916.500 ;
        RECT 2900.825 1915.750 2924.800 1916.050 ;
        RECT 2900.825 1915.735 2901.155 1915.750 ;
        RECT 2917.600 1915.300 2924.800 1915.750 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 647.750 3270.700 648.070 3270.760 ;
        RECT 2660.710 3270.700 2661.030 3270.760 ;
        RECT 647.750 3270.560 2661.030 3270.700 ;
        RECT 647.750 3270.500 648.070 3270.560 ;
        RECT 2660.710 3270.500 2661.030 3270.560 ;
        RECT 2660.710 2152.780 2661.030 2152.840 ;
        RECT 2900.830 2152.780 2901.150 2152.840 ;
        RECT 2660.710 2152.640 2901.150 2152.780 ;
        RECT 2660.710 2152.580 2661.030 2152.640 ;
        RECT 2900.830 2152.580 2901.150 2152.640 ;
      LAYER via ;
        RECT 647.780 3270.500 648.040 3270.760 ;
        RECT 2660.740 3270.500 2661.000 3270.760 ;
        RECT 2660.740 2152.580 2661.000 2152.840 ;
        RECT 2900.860 2152.580 2901.120 2152.840 ;
      LAYER met2 ;
        RECT 647.780 3270.470 648.040 3270.790 ;
        RECT 2660.740 3270.470 2661.000 3270.790 ;
        RECT 647.840 3260.000 647.980 3270.470 ;
        RECT 647.730 3256.000 648.010 3260.000 ;
        RECT 2660.800 2152.870 2660.940 3270.470 ;
        RECT 2660.740 2152.550 2661.000 2152.870 ;
        RECT 2900.860 2152.550 2901.120 2152.870 ;
        RECT 2900.920 2150.685 2901.060 2152.550 ;
        RECT 2900.850 2150.315 2901.130 2150.685 ;
      LAYER via2 ;
        RECT 2900.850 2150.360 2901.130 2150.640 ;
      LAYER met3 ;
        RECT 2900.825 2150.650 2901.155 2150.665 ;
        RECT 2917.600 2150.650 2924.800 2151.100 ;
        RECT 2900.825 2150.350 2924.800 2150.650 ;
        RECT 2900.825 2150.335 2901.155 2150.350 ;
        RECT 2917.600 2149.900 2924.800 2150.350 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2090.900 2615.490 2090.960 ;
        RECT 2846.090 2090.900 2846.410 2090.960 ;
        RECT 2615.170 2090.760 2846.410 2090.900 ;
        RECT 2615.170 2090.700 2615.490 2090.760 ;
        RECT 2846.090 2090.700 2846.410 2090.760 ;
        RECT 2846.090 200.160 2846.410 200.220 ;
        RECT 2900.830 200.160 2901.150 200.220 ;
        RECT 2846.090 200.020 2901.150 200.160 ;
        RECT 2846.090 199.960 2846.410 200.020 ;
        RECT 2900.830 199.960 2901.150 200.020 ;
      LAYER via ;
        RECT 2615.200 2090.700 2615.460 2090.960 ;
        RECT 2846.120 2090.700 2846.380 2090.960 ;
        RECT 2846.120 199.960 2846.380 200.220 ;
        RECT 2900.860 199.960 2901.120 200.220 ;
      LAYER met2 ;
        RECT 2615.190 2093.195 2615.470 2093.565 ;
        RECT 2615.260 2090.990 2615.400 2093.195 ;
        RECT 2615.200 2090.670 2615.460 2090.990 ;
        RECT 2846.120 2090.670 2846.380 2090.990 ;
        RECT 2846.180 200.250 2846.320 2090.670 ;
        RECT 2846.120 199.930 2846.380 200.250 ;
        RECT 2900.860 199.930 2901.120 200.250 ;
        RECT 2900.920 195.685 2901.060 199.930 ;
        RECT 2900.850 195.315 2901.130 195.685 ;
      LAYER via2 ;
        RECT 2615.190 2093.240 2615.470 2093.520 ;
        RECT 2900.850 195.360 2901.130 195.640 ;
      LAYER met3 ;
        RECT 2606.000 2093.530 2610.000 2093.920 ;
        RECT 2615.165 2093.530 2615.495 2093.545 ;
        RECT 2606.000 2093.320 2615.495 2093.530 ;
        RECT 2609.580 2093.230 2615.495 2093.320 ;
        RECT 2615.165 2093.215 2615.495 2093.230 ;
        RECT 2900.825 195.650 2901.155 195.665 ;
        RECT 2917.600 195.650 2924.800 196.100 ;
        RECT 2900.825 195.350 2924.800 195.650 ;
        RECT 2900.825 195.335 2901.155 195.350 ;
        RECT 2917.600 194.900 2924.800 195.350 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 3001.760 2615.490 3001.820 ;
        RECT 2639.090 3001.760 2639.410 3001.820 ;
        RECT 2615.170 3001.620 2639.410 3001.760 ;
        RECT 2615.170 3001.560 2615.490 3001.620 ;
        RECT 2639.090 3001.560 2639.410 3001.620 ;
        RECT 2639.090 2546.160 2639.410 2546.220 ;
        RECT 2900.830 2546.160 2901.150 2546.220 ;
        RECT 2639.090 2546.020 2901.150 2546.160 ;
        RECT 2639.090 2545.960 2639.410 2546.020 ;
        RECT 2900.830 2545.960 2901.150 2546.020 ;
      LAYER via ;
        RECT 2615.200 3001.560 2615.460 3001.820 ;
        RECT 2639.120 3001.560 2639.380 3001.820 ;
        RECT 2639.120 2545.960 2639.380 2546.220 ;
        RECT 2900.860 2545.960 2901.120 2546.220 ;
      LAYER met2 ;
        RECT 2615.190 3001.675 2615.470 3002.045 ;
        RECT 2615.200 3001.530 2615.460 3001.675 ;
        RECT 2639.120 3001.530 2639.380 3001.850 ;
        RECT 2639.180 2546.250 2639.320 3001.530 ;
        RECT 2639.120 2545.930 2639.380 2546.250 ;
        RECT 2900.860 2545.930 2901.120 2546.250 ;
        RECT 2900.920 2541.685 2901.060 2545.930 ;
        RECT 2900.850 2541.315 2901.130 2541.685 ;
      LAYER via2 ;
        RECT 2615.190 3001.720 2615.470 3002.000 ;
        RECT 2900.850 2541.360 2901.130 2541.640 ;
      LAYER met3 ;
        RECT 2606.000 3002.010 2610.000 3002.400 ;
        RECT 2615.165 3002.010 2615.495 3002.025 ;
        RECT 2606.000 3001.800 2615.495 3002.010 ;
        RECT 2609.580 3001.710 2615.495 3001.800 ;
        RECT 2615.165 3001.695 2615.495 3001.710 ;
        RECT 2900.825 2541.650 2901.155 2541.665 ;
        RECT 2917.600 2541.650 2924.800 2542.100 ;
        RECT 2900.825 2541.350 2924.800 2541.650 ;
        RECT 2900.825 2541.335 2901.155 2541.350 ;
        RECT 2917.600 2540.900 2924.800 2541.350 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2701.650 2773.960 2701.970 2774.020 ;
        RECT 2900.830 2773.960 2901.150 2774.020 ;
        RECT 2701.650 2773.820 2901.150 2773.960 ;
        RECT 2701.650 2773.760 2701.970 2773.820 ;
        RECT 2900.830 2773.760 2901.150 2773.820 ;
        RECT 2615.170 1800.880 2615.490 1800.940 ;
        RECT 2701.650 1800.880 2701.970 1800.940 ;
        RECT 2615.170 1800.740 2701.970 1800.880 ;
        RECT 2615.170 1800.680 2615.490 1800.740 ;
        RECT 2701.650 1800.680 2701.970 1800.740 ;
      LAYER via ;
        RECT 2701.680 2773.760 2701.940 2774.020 ;
        RECT 2900.860 2773.760 2901.120 2774.020 ;
        RECT 2615.200 1800.680 2615.460 1800.940 ;
        RECT 2701.680 1800.680 2701.940 1800.940 ;
      LAYER met2 ;
        RECT 2900.850 2775.915 2901.130 2776.285 ;
        RECT 2900.920 2774.050 2901.060 2775.915 ;
        RECT 2701.680 2773.730 2701.940 2774.050 ;
        RECT 2900.860 2773.730 2901.120 2774.050 ;
        RECT 2701.740 1800.970 2701.880 2773.730 ;
        RECT 2615.200 1800.650 2615.460 1800.970 ;
        RECT 2701.680 1800.650 2701.940 1800.970 ;
        RECT 2615.260 1797.085 2615.400 1800.650 ;
        RECT 2615.190 1796.715 2615.470 1797.085 ;
      LAYER via2 ;
        RECT 2900.850 2775.960 2901.130 2776.240 ;
        RECT 2615.190 1796.760 2615.470 1797.040 ;
      LAYER met3 ;
        RECT 2900.825 2776.250 2901.155 2776.265 ;
        RECT 2917.600 2776.250 2924.800 2776.700 ;
        RECT 2900.825 2775.950 2924.800 2776.250 ;
        RECT 2900.825 2775.935 2901.155 2775.950 ;
        RECT 2917.600 2775.500 2924.800 2775.950 ;
        RECT 2606.000 1797.050 2610.000 1797.440 ;
        RECT 2615.165 1797.050 2615.495 1797.065 ;
        RECT 2606.000 1796.840 2615.495 1797.050 ;
        RECT 2609.580 1796.750 2615.495 1796.840 ;
        RECT 2615.165 1796.735 2615.495 1796.750 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2801.030 3011.195 2801.310 3011.565 ;
        RECT 2801.100 3009.525 2801.240 3011.195 ;
        RECT 2825.410 3010.515 2825.690 3010.885 ;
        RECT 2801.030 3009.155 2801.310 3009.525 ;
        RECT 2825.480 3008.845 2825.620 3010.515 ;
        RECT 2863.130 3009.155 2863.410 3009.525 ;
        RECT 2825.410 3008.475 2825.690 3008.845 ;
        RECT 2863.200 3008.730 2863.340 3009.155 ;
        RECT 2863.590 3008.730 2863.870 3008.845 ;
        RECT 2863.200 3008.590 2863.870 3008.730 ;
        RECT 2863.590 3008.475 2863.870 3008.590 ;
        RECT 2659.350 2352.275 2659.630 2352.645 ;
        RECT 2659.420 2305.725 2659.560 2352.275 ;
        RECT 2659.350 2305.355 2659.630 2305.725 ;
        RECT 2658.430 2213.555 2658.710 2213.925 ;
        RECT 2658.500 2167.005 2658.640 2213.555 ;
        RECT 2658.430 2166.635 2658.710 2167.005 ;
        RECT 2658.430 2165.955 2658.710 2166.325 ;
        RECT 2658.500 2118.725 2658.640 2165.955 ;
        RECT 2658.430 2118.355 2658.710 2118.725 ;
        RECT 2659.350 2027.235 2659.630 2027.605 ;
        RECT 2659.420 1980.685 2659.560 2027.235 ;
        RECT 2659.350 1980.315 2659.630 1980.685 ;
        RECT 2660.730 1979.635 2661.010 1980.005 ;
        RECT 2660.800 1932.405 2660.940 1979.635 ;
        RECT 2660.730 1932.035 2661.010 1932.405 ;
        RECT 2658.890 1827.315 2659.170 1827.685 ;
        RECT 2658.960 1780.765 2659.100 1827.315 ;
        RECT 2658.890 1780.395 2659.170 1780.765 ;
        RECT 2659.350 1669.555 2659.630 1669.925 ;
        RECT 2659.420 1594.445 2659.560 1669.555 ;
        RECT 2659.350 1594.075 2659.630 1594.445 ;
        RECT 2660.270 1586.595 2660.550 1586.965 ;
        RECT 2660.340 1538.685 2660.480 1586.595 ;
        RECT 2660.270 1538.315 2660.550 1538.685 ;
        RECT 2659.350 1531.515 2659.630 1531.885 ;
        RECT 2659.420 1484.965 2659.560 1531.515 ;
        RECT 2659.350 1484.595 2659.630 1484.965 ;
        RECT 2659.350 1434.955 2659.630 1435.325 ;
        RECT 2659.420 1388.405 2659.560 1434.955 ;
        RECT 2659.350 1388.035 2659.630 1388.405 ;
        RECT 2660.730 1120.795 2661.010 1121.165 ;
        RECT 2660.800 1064.045 2660.940 1120.795 ;
        RECT 2660.730 1063.675 2661.010 1064.045 ;
        RECT 2660.730 1014.035 2661.010 1014.405 ;
        RECT 2660.800 966.805 2660.940 1014.035 ;
        RECT 2660.730 966.435 2661.010 966.805 ;
      LAYER via2 ;
        RECT 2801.030 3011.240 2801.310 3011.520 ;
        RECT 2825.410 3010.560 2825.690 3010.840 ;
        RECT 2801.030 3009.200 2801.310 3009.480 ;
        RECT 2863.130 3009.200 2863.410 3009.480 ;
        RECT 2825.410 3008.520 2825.690 3008.800 ;
        RECT 2863.590 3008.520 2863.870 3008.800 ;
        RECT 2659.350 2352.320 2659.630 2352.600 ;
        RECT 2659.350 2305.400 2659.630 2305.680 ;
        RECT 2658.430 2213.600 2658.710 2213.880 ;
        RECT 2658.430 2166.680 2658.710 2166.960 ;
        RECT 2658.430 2166.000 2658.710 2166.280 ;
        RECT 2658.430 2118.400 2658.710 2118.680 ;
        RECT 2659.350 2027.280 2659.630 2027.560 ;
        RECT 2659.350 1980.360 2659.630 1980.640 ;
        RECT 2660.730 1979.680 2661.010 1979.960 ;
        RECT 2660.730 1932.080 2661.010 1932.360 ;
        RECT 2658.890 1827.360 2659.170 1827.640 ;
        RECT 2658.890 1780.440 2659.170 1780.720 ;
        RECT 2659.350 1669.600 2659.630 1669.880 ;
        RECT 2659.350 1594.120 2659.630 1594.400 ;
        RECT 2660.270 1586.640 2660.550 1586.920 ;
        RECT 2660.270 1538.360 2660.550 1538.640 ;
        RECT 2659.350 1531.560 2659.630 1531.840 ;
        RECT 2659.350 1484.640 2659.630 1484.920 ;
        RECT 2659.350 1435.000 2659.630 1435.280 ;
        RECT 2659.350 1388.080 2659.630 1388.360 ;
        RECT 2660.730 1120.840 2661.010 1121.120 ;
        RECT 2660.730 1063.720 2661.010 1064.000 ;
        RECT 2660.730 1014.080 2661.010 1014.360 ;
        RECT 2660.730 966.480 2661.010 966.760 ;
      LAYER met3 ;
        RECT 2752.910 3011.530 2753.290 3011.540 ;
        RECT 2801.005 3011.530 2801.335 3011.545 ;
        RECT 2752.910 3011.230 2801.335 3011.530 ;
        RECT 2752.910 3011.220 2753.290 3011.230 ;
        RECT 2801.005 3011.215 2801.335 3011.230 ;
        RECT 2825.385 3010.850 2825.715 3010.865 ;
        RECT 2917.600 3010.850 2924.800 3011.300 ;
        RECT 2801.710 3010.550 2825.715 3010.850 ;
        RECT 2659.070 3010.170 2659.450 3010.180 ;
        RECT 2752.910 3010.170 2753.290 3010.180 ;
        RECT 2659.070 3009.870 2670.450 3010.170 ;
        RECT 2659.070 3009.860 2659.450 3009.870 ;
        RECT 2670.150 3008.810 2670.450 3009.870 ;
        RECT 2718.910 3009.870 2753.290 3010.170 ;
        RECT 2718.910 3008.810 2719.210 3009.870 ;
        RECT 2752.910 3009.860 2753.290 3009.870 ;
        RECT 2801.005 3009.490 2801.335 3009.505 ;
        RECT 2801.710 3009.490 2802.010 3010.550 ;
        RECT 2825.385 3010.535 2825.715 3010.550 ;
        RECT 2916.710 3010.550 2924.800 3010.850 ;
        RECT 2863.105 3009.490 2863.435 3009.505 ;
        RECT 2801.005 3009.190 2802.010 3009.490 ;
        RECT 2849.550 3009.190 2863.435 3009.490 ;
        RECT 2801.005 3009.175 2801.335 3009.190 ;
        RECT 2670.150 3008.510 2719.210 3008.810 ;
        RECT 2825.385 3008.810 2825.715 3008.825 ;
        RECT 2849.550 3008.810 2849.850 3009.190 ;
        RECT 2863.105 3009.175 2863.435 3009.190 ;
        RECT 2825.385 3008.510 2849.850 3008.810 ;
        RECT 2863.565 3008.810 2863.895 3008.825 ;
        RECT 2916.710 3008.810 2917.010 3010.550 ;
        RECT 2917.600 3010.100 2924.800 3010.550 ;
        RECT 2863.565 3008.510 2917.010 3008.810 ;
        RECT 2825.385 3008.495 2825.715 3008.510 ;
        RECT 2863.565 3008.495 2863.895 3008.510 ;
        RECT 2659.325 2352.610 2659.655 2352.625 ;
        RECT 2659.990 2352.610 2660.370 2352.620 ;
        RECT 2659.325 2352.310 2660.370 2352.610 ;
        RECT 2659.325 2352.295 2659.655 2352.310 ;
        RECT 2659.990 2352.300 2660.370 2352.310 ;
        RECT 2659.325 2305.690 2659.655 2305.705 ;
        RECT 2658.190 2305.390 2659.655 2305.690 ;
        RECT 2658.190 2305.020 2658.490 2305.390 ;
        RECT 2659.325 2305.375 2659.655 2305.390 ;
        RECT 2658.150 2304.700 2658.530 2305.020 ;
        RECT 2658.150 2284.300 2658.530 2284.620 ;
        RECT 2658.190 2283.250 2658.490 2284.300 ;
        RECT 2659.070 2283.250 2659.450 2283.260 ;
        RECT 2658.190 2282.950 2659.450 2283.250 ;
        RECT 2659.070 2282.940 2659.450 2282.950 ;
        RECT 2658.150 2215.250 2658.530 2215.260 ;
        RECT 2659.070 2215.250 2659.450 2215.260 ;
        RECT 2658.150 2214.950 2659.450 2215.250 ;
        RECT 2658.150 2214.940 2658.530 2214.950 ;
        RECT 2659.070 2214.940 2659.450 2214.950 ;
        RECT 2658.405 2213.900 2658.735 2213.905 ;
        RECT 2658.150 2213.890 2658.735 2213.900 ;
        RECT 2657.950 2213.590 2658.735 2213.890 ;
        RECT 2658.150 2213.580 2658.735 2213.590 ;
        RECT 2658.405 2213.575 2658.735 2213.580 ;
        RECT 2658.405 2166.970 2658.735 2166.985 ;
        RECT 2659.070 2166.970 2659.450 2166.980 ;
        RECT 2658.405 2166.670 2659.450 2166.970 ;
        RECT 2658.405 2166.655 2658.735 2166.670 ;
        RECT 2659.070 2166.660 2659.450 2166.670 ;
        RECT 2658.405 2166.290 2658.735 2166.305 ;
        RECT 2659.070 2166.290 2659.450 2166.300 ;
        RECT 2658.405 2165.990 2659.450 2166.290 ;
        RECT 2658.405 2165.975 2658.735 2165.990 ;
        RECT 2659.070 2165.980 2659.450 2165.990 ;
        RECT 2658.405 2118.700 2658.735 2118.705 ;
        RECT 2658.150 2118.690 2658.735 2118.700 ;
        RECT 2657.950 2118.390 2658.735 2118.690 ;
        RECT 2658.150 2118.380 2658.735 2118.390 ;
        RECT 2658.405 2118.375 2658.735 2118.380 ;
        RECT 2659.070 2043.210 2659.450 2043.220 ;
        RECT 2658.190 2042.910 2659.450 2043.210 ;
        RECT 2658.190 2041.860 2658.490 2042.910 ;
        RECT 2659.070 2042.900 2659.450 2042.910 ;
        RECT 2658.150 2041.540 2658.530 2041.860 ;
        RECT 2658.150 2027.940 2658.530 2028.260 ;
        RECT 2658.190 2027.570 2658.490 2027.940 ;
        RECT 2659.325 2027.570 2659.655 2027.585 ;
        RECT 2658.190 2027.270 2659.655 2027.570 ;
        RECT 2659.325 2027.255 2659.655 2027.270 ;
        RECT 2659.325 1980.650 2659.655 1980.665 ;
        RECT 2659.990 1980.650 2660.370 1980.660 ;
        RECT 2659.325 1980.350 2660.370 1980.650 ;
        RECT 2659.325 1980.335 2659.655 1980.350 ;
        RECT 2659.990 1980.340 2660.370 1980.350 ;
        RECT 2659.990 1979.970 2660.370 1979.980 ;
        RECT 2660.705 1979.970 2661.035 1979.985 ;
        RECT 2659.990 1979.670 2661.035 1979.970 ;
        RECT 2659.990 1979.660 2660.370 1979.670 ;
        RECT 2660.705 1979.655 2661.035 1979.670 ;
        RECT 2659.990 1932.370 2660.370 1932.380 ;
        RECT 2660.705 1932.370 2661.035 1932.385 ;
        RECT 2659.990 1932.070 2661.035 1932.370 ;
        RECT 2659.990 1932.060 2660.370 1932.070 ;
        RECT 2660.705 1932.055 2661.035 1932.070 ;
        RECT 2659.990 1829.690 2660.370 1829.700 ;
        RECT 2658.190 1829.390 2660.370 1829.690 ;
        RECT 2658.190 1829.020 2658.490 1829.390 ;
        RECT 2659.990 1829.380 2660.370 1829.390 ;
        RECT 2658.150 1828.700 2658.530 1829.020 ;
        RECT 2658.150 1827.650 2658.530 1827.660 ;
        RECT 2658.865 1827.650 2659.195 1827.665 ;
        RECT 2658.150 1827.350 2659.195 1827.650 ;
        RECT 2658.150 1827.340 2658.530 1827.350 ;
        RECT 2658.865 1827.335 2659.195 1827.350 ;
        RECT 2658.865 1780.740 2659.195 1780.745 ;
        RECT 2658.865 1780.730 2659.450 1780.740 ;
        RECT 2658.640 1780.430 2659.450 1780.730 ;
        RECT 2658.865 1780.420 2659.450 1780.430 ;
        RECT 2658.865 1780.415 2659.195 1780.420 ;
        RECT 2659.070 1753.220 2659.450 1753.540 ;
        RECT 2659.110 1752.180 2659.410 1753.220 ;
        RECT 2659.070 1751.860 2659.450 1752.180 ;
        RECT 2658.150 1704.940 2658.530 1705.260 ;
        RECT 2658.190 1703.890 2658.490 1704.940 ;
        RECT 2659.070 1703.890 2659.450 1703.900 ;
        RECT 2658.190 1703.590 2659.450 1703.890 ;
        RECT 2659.070 1703.580 2659.450 1703.590 ;
        RECT 2659.325 1669.900 2659.655 1669.905 ;
        RECT 2659.070 1669.890 2659.655 1669.900 ;
        RECT 2658.870 1669.590 2659.655 1669.890 ;
        RECT 2659.070 1669.580 2659.655 1669.590 ;
        RECT 2659.325 1669.575 2659.655 1669.580 ;
        RECT 2659.325 1594.410 2659.655 1594.425 ;
        RECT 2659.990 1594.410 2660.370 1594.420 ;
        RECT 2659.325 1594.110 2660.370 1594.410 ;
        RECT 2659.325 1594.095 2659.655 1594.110 ;
        RECT 2659.990 1594.100 2660.370 1594.110 ;
        RECT 2660.245 1586.940 2660.575 1586.945 ;
        RECT 2659.990 1586.930 2660.575 1586.940 ;
        RECT 2659.990 1586.630 2660.800 1586.930 ;
        RECT 2659.990 1586.620 2660.575 1586.630 ;
        RECT 2660.245 1586.615 2660.575 1586.620 ;
        RECT 2659.070 1538.650 2659.450 1538.660 ;
        RECT 2660.245 1538.650 2660.575 1538.665 ;
        RECT 2659.070 1538.350 2660.575 1538.650 ;
        RECT 2659.070 1538.340 2659.450 1538.350 ;
        RECT 2660.245 1538.335 2660.575 1538.350 ;
        RECT 2659.325 1531.860 2659.655 1531.865 ;
        RECT 2659.070 1531.850 2659.655 1531.860 ;
        RECT 2659.070 1531.550 2659.880 1531.850 ;
        RECT 2659.070 1531.540 2659.655 1531.550 ;
        RECT 2659.325 1531.535 2659.655 1531.540 ;
        RECT 2659.325 1484.930 2659.655 1484.945 ;
        RECT 2659.110 1484.615 2659.655 1484.930 ;
        RECT 2659.110 1484.260 2659.410 1484.615 ;
        RECT 2659.070 1483.940 2659.450 1484.260 ;
        RECT 2658.150 1436.650 2658.530 1436.660 ;
        RECT 2659.990 1436.650 2660.370 1436.660 ;
        RECT 2658.150 1436.350 2660.370 1436.650 ;
        RECT 2658.150 1436.340 2658.530 1436.350 ;
        RECT 2659.990 1436.340 2660.370 1436.350 ;
        RECT 2659.325 1435.290 2659.655 1435.305 ;
        RECT 2659.990 1435.290 2660.370 1435.300 ;
        RECT 2659.325 1434.990 2660.370 1435.290 ;
        RECT 2659.325 1434.975 2659.655 1434.990 ;
        RECT 2659.990 1434.980 2660.370 1434.990 ;
        RECT 2659.325 1388.370 2659.655 1388.385 ;
        RECT 2658.190 1388.070 2659.655 1388.370 ;
        RECT 2658.190 1387.700 2658.490 1388.070 ;
        RECT 2659.325 1388.055 2659.655 1388.070 ;
        RECT 2658.150 1387.380 2658.530 1387.700 ;
        RECT 2658.150 1221.460 2658.530 1221.780 ;
        RECT 2658.190 1220.410 2658.490 1221.460 ;
        RECT 2659.070 1220.410 2659.450 1220.420 ;
        RECT 2658.190 1220.110 2659.450 1220.410 ;
        RECT 2659.070 1220.100 2659.450 1220.110 ;
        RECT 2659.990 1121.130 2660.370 1121.140 ;
        RECT 2660.705 1121.130 2661.035 1121.145 ;
        RECT 2659.990 1120.830 2661.035 1121.130 ;
        RECT 2659.990 1120.820 2660.370 1120.830 ;
        RECT 2660.705 1120.815 2661.035 1120.830 ;
        RECT 2660.705 1064.010 2661.035 1064.025 ;
        RECT 2660.030 1063.710 2661.035 1064.010 ;
        RECT 2660.030 1063.340 2660.330 1063.710 ;
        RECT 2660.705 1063.695 2661.035 1063.710 ;
        RECT 2659.990 1063.020 2660.370 1063.340 ;
        RECT 2659.990 1014.370 2660.370 1014.380 ;
        RECT 2660.705 1014.370 2661.035 1014.385 ;
        RECT 2659.990 1014.070 2661.035 1014.370 ;
        RECT 2659.990 1014.060 2660.370 1014.070 ;
        RECT 2660.705 1014.055 2661.035 1014.070 ;
        RECT 2660.705 966.770 2661.035 966.785 ;
        RECT 2660.030 966.470 2661.035 966.770 ;
        RECT 2659.070 966.260 2659.450 966.270 ;
        RECT 2660.030 966.260 2660.330 966.470 ;
        RECT 2660.705 966.455 2661.035 966.470 ;
        RECT 2659.070 965.960 2660.330 966.260 ;
        RECT 2659.070 965.950 2659.450 965.960 ;
        RECT 310.000 940.040 314.000 940.640 ;
        RECT 309.390 939.570 309.770 939.580 ;
        RECT 310.350 939.570 310.650 940.040 ;
        RECT 309.390 939.270 310.650 939.570 ;
        RECT 309.390 939.260 309.770 939.270 ;
      LAYER via3 ;
        RECT 2752.940 3011.220 2753.260 3011.540 ;
        RECT 2659.100 3009.860 2659.420 3010.180 ;
        RECT 2752.940 3009.860 2753.260 3010.180 ;
        RECT 2660.020 2352.300 2660.340 2352.620 ;
        RECT 2658.180 2304.700 2658.500 2305.020 ;
        RECT 2658.180 2284.300 2658.500 2284.620 ;
        RECT 2659.100 2282.940 2659.420 2283.260 ;
        RECT 2658.180 2214.940 2658.500 2215.260 ;
        RECT 2659.100 2214.940 2659.420 2215.260 ;
        RECT 2658.180 2213.580 2658.500 2213.900 ;
        RECT 2659.100 2166.660 2659.420 2166.980 ;
        RECT 2659.100 2165.980 2659.420 2166.300 ;
        RECT 2658.180 2118.380 2658.500 2118.700 ;
        RECT 2659.100 2042.900 2659.420 2043.220 ;
        RECT 2658.180 2041.540 2658.500 2041.860 ;
        RECT 2658.180 2027.940 2658.500 2028.260 ;
        RECT 2660.020 1980.340 2660.340 1980.660 ;
        RECT 2660.020 1979.660 2660.340 1979.980 ;
        RECT 2660.020 1932.060 2660.340 1932.380 ;
        RECT 2660.020 1829.380 2660.340 1829.700 ;
        RECT 2658.180 1828.700 2658.500 1829.020 ;
        RECT 2658.180 1827.340 2658.500 1827.660 ;
        RECT 2659.100 1780.420 2659.420 1780.740 ;
        RECT 2659.100 1753.220 2659.420 1753.540 ;
        RECT 2659.100 1751.860 2659.420 1752.180 ;
        RECT 2658.180 1704.940 2658.500 1705.260 ;
        RECT 2659.100 1703.580 2659.420 1703.900 ;
        RECT 2659.100 1669.580 2659.420 1669.900 ;
        RECT 2660.020 1594.100 2660.340 1594.420 ;
        RECT 2660.020 1586.620 2660.340 1586.940 ;
        RECT 2659.100 1538.340 2659.420 1538.660 ;
        RECT 2659.100 1531.540 2659.420 1531.860 ;
        RECT 2659.100 1483.940 2659.420 1484.260 ;
        RECT 2658.180 1436.340 2658.500 1436.660 ;
        RECT 2660.020 1436.340 2660.340 1436.660 ;
        RECT 2660.020 1434.980 2660.340 1435.300 ;
        RECT 2658.180 1387.380 2658.500 1387.700 ;
        RECT 2658.180 1221.460 2658.500 1221.780 ;
        RECT 2659.100 1220.100 2659.420 1220.420 ;
        RECT 2660.020 1120.820 2660.340 1121.140 ;
        RECT 2660.020 1063.020 2660.340 1063.340 ;
        RECT 2660.020 1014.060 2660.340 1014.380 ;
        RECT 2659.100 965.950 2659.420 966.270 ;
        RECT 309.420 939.260 309.740 939.580 ;
      LAYER met4 ;
        RECT 2752.935 3011.215 2753.265 3011.545 ;
        RECT 2752.950 3010.185 2753.250 3011.215 ;
        RECT 2659.095 3009.855 2659.425 3010.185 ;
        RECT 2752.935 3009.855 2753.265 3010.185 ;
        RECT 2659.110 2963.250 2659.410 3009.855 ;
        RECT 2657.270 2962.950 2659.410 2963.250 ;
        RECT 2657.270 2959.850 2657.570 2962.950 ;
        RECT 2657.270 2959.550 2658.490 2959.850 ;
        RECT 2658.190 2956.450 2658.490 2959.550 ;
        RECT 2658.190 2956.150 2659.410 2956.450 ;
        RECT 2659.110 2524.650 2659.410 2956.150 ;
        RECT 2659.110 2524.350 2660.330 2524.650 ;
        RECT 2660.030 2352.625 2660.330 2524.350 ;
        RECT 2660.015 2352.295 2660.345 2352.625 ;
        RECT 2658.175 2304.695 2658.505 2305.025 ;
        RECT 2658.190 2284.625 2658.490 2304.695 ;
        RECT 2658.175 2284.295 2658.505 2284.625 ;
        RECT 2659.095 2282.935 2659.425 2283.265 ;
        RECT 2659.110 2215.265 2659.410 2282.935 ;
        RECT 2658.175 2214.935 2658.505 2215.265 ;
        RECT 2659.095 2214.935 2659.425 2215.265 ;
        RECT 2658.190 2213.905 2658.490 2214.935 ;
        RECT 2658.175 2213.575 2658.505 2213.905 ;
        RECT 2659.095 2166.655 2659.425 2166.985 ;
        RECT 2659.110 2166.305 2659.410 2166.655 ;
        RECT 2659.095 2165.975 2659.425 2166.305 ;
        RECT 2658.175 2118.375 2658.505 2118.705 ;
        RECT 2658.190 2089.450 2658.490 2118.375 ;
        RECT 2658.190 2089.150 2659.410 2089.450 ;
        RECT 2659.110 2043.225 2659.410 2089.150 ;
        RECT 2659.095 2042.895 2659.425 2043.225 ;
        RECT 2658.175 2041.535 2658.505 2041.865 ;
        RECT 2658.190 2028.265 2658.490 2041.535 ;
        RECT 2658.175 2027.935 2658.505 2028.265 ;
        RECT 2660.015 1980.335 2660.345 1980.665 ;
        RECT 2660.030 1979.985 2660.330 1980.335 ;
        RECT 2660.015 1979.655 2660.345 1979.985 ;
        RECT 2660.015 1932.055 2660.345 1932.385 ;
        RECT 2660.030 1829.705 2660.330 1932.055 ;
        RECT 2660.015 1829.375 2660.345 1829.705 ;
        RECT 2658.175 1828.695 2658.505 1829.025 ;
        RECT 2658.190 1827.665 2658.490 1828.695 ;
        RECT 2658.175 1827.335 2658.505 1827.665 ;
        RECT 2659.095 1780.415 2659.425 1780.745 ;
        RECT 2659.110 1753.545 2659.410 1780.415 ;
        RECT 2659.095 1753.215 2659.425 1753.545 ;
        RECT 2659.095 1751.855 2659.425 1752.185 ;
        RECT 2659.110 1739.250 2659.410 1751.855 ;
        RECT 2658.190 1738.950 2659.410 1739.250 ;
        RECT 2658.190 1705.265 2658.490 1738.950 ;
        RECT 2658.175 1704.935 2658.505 1705.265 ;
        RECT 2659.095 1703.575 2659.425 1703.905 ;
        RECT 2659.110 1669.905 2659.410 1703.575 ;
        RECT 2659.095 1669.575 2659.425 1669.905 ;
        RECT 2660.015 1594.095 2660.345 1594.425 ;
        RECT 2660.030 1586.945 2660.330 1594.095 ;
        RECT 2660.015 1586.615 2660.345 1586.945 ;
        RECT 2659.095 1538.335 2659.425 1538.665 ;
        RECT 2659.110 1531.865 2659.410 1538.335 ;
        RECT 2659.095 1531.535 2659.425 1531.865 ;
        RECT 2659.095 1483.935 2659.425 1484.265 ;
        RECT 2659.110 1463.850 2659.410 1483.935 ;
        RECT 2658.190 1463.550 2659.410 1463.850 ;
        RECT 2658.190 1436.665 2658.490 1463.550 ;
        RECT 2658.175 1436.335 2658.505 1436.665 ;
        RECT 2660.015 1436.335 2660.345 1436.665 ;
        RECT 2660.030 1435.305 2660.330 1436.335 ;
        RECT 2660.015 1434.975 2660.345 1435.305 ;
        RECT 2658.175 1387.375 2658.505 1387.705 ;
        RECT 2658.190 1361.850 2658.490 1387.375 ;
        RECT 2658.190 1361.550 2660.330 1361.850 ;
        RECT 2660.030 1273.450 2660.330 1361.550 ;
        RECT 2659.110 1273.150 2660.330 1273.450 ;
        RECT 2659.110 1270.050 2659.410 1273.150 ;
        RECT 2658.190 1269.750 2659.410 1270.050 ;
        RECT 2658.190 1221.785 2658.490 1269.750 ;
        RECT 2658.175 1221.455 2658.505 1221.785 ;
        RECT 2659.095 1220.095 2659.425 1220.425 ;
        RECT 2659.110 1174.850 2659.410 1220.095 ;
        RECT 2659.110 1174.550 2660.330 1174.850 ;
        RECT 2660.030 1121.145 2660.330 1174.550 ;
        RECT 2660.015 1120.815 2660.345 1121.145 ;
        RECT 2660.015 1063.015 2660.345 1063.345 ;
        RECT 2660.030 1014.385 2660.330 1063.015 ;
        RECT 2660.015 1014.055 2660.345 1014.385 ;
        RECT 2659.095 965.945 2659.425 966.275 ;
        RECT 2659.110 940.690 2659.410 965.945 ;
        RECT 309.415 939.255 309.745 939.585 ;
        RECT 2658.670 939.510 2659.850 940.690 ;
        RECT 309.430 937.290 309.730 939.255 ;
        RECT 308.990 936.110 310.170 937.290 ;
      LAYER met5 ;
        RECT 515.780 937.500 518.300 940.900 ;
        RECT 612.380 937.500 614.900 940.900 ;
        RECT 308.780 935.900 351.780 937.500 ;
        RECT 350.180 934.100 351.780 935.900 ;
        RECT 402.620 935.900 451.140 937.500 ;
        RECT 402.620 934.100 404.220 935.900 ;
        RECT 350.180 932.500 404.220 934.100 ;
        RECT 449.540 934.100 451.140 935.900 ;
        RECT 515.780 935.900 547.740 937.500 ;
        RECT 515.780 934.100 517.380 935.900 ;
        RECT 449.540 932.500 517.380 934.100 ;
        RECT 546.140 934.100 547.740 935.900 ;
        RECT 612.380 935.900 644.340 937.500 ;
        RECT 612.380 934.100 613.980 935.900 ;
        RECT 546.140 932.500 613.980 934.100 ;
        RECT 642.740 934.100 644.340 935.900 ;
        RECT 708.980 934.100 711.500 940.900 ;
        RECT 785.340 939.300 808.100 940.900 ;
        RECT 785.340 937.500 786.940 939.300 ;
        RECT 737.500 935.900 786.940 937.500 ;
        RECT 737.500 934.100 739.100 935.900 ;
        RECT 642.740 932.500 739.100 934.100 ;
        RECT 806.500 934.100 808.100 939.300 ;
        RECT 854.340 939.300 904.700 940.900 ;
        RECT 854.340 934.100 855.940 939.300 ;
        RECT 806.500 932.500 855.940 934.100 ;
        RECT 903.100 934.100 904.700 939.300 ;
        RECT 950.940 939.300 1001.300 940.900 ;
        RECT 950.940 934.100 952.540 939.300 ;
        RECT 903.100 932.500 952.540 934.100 ;
        RECT 999.700 934.100 1001.300 939.300 ;
        RECT 1047.540 939.300 1097.900 940.900 ;
        RECT 1047.540 934.100 1049.140 939.300 ;
        RECT 999.700 932.500 1049.140 934.100 ;
        RECT 1096.300 934.100 1097.900 939.300 ;
        RECT 1144.140 939.300 1194.500 940.900 ;
        RECT 1144.140 934.100 1145.740 939.300 ;
        RECT 1096.300 932.500 1145.740 934.100 ;
        RECT 1192.900 934.100 1194.500 939.300 ;
        RECT 1240.740 939.300 1291.100 940.900 ;
        RECT 1240.740 934.100 1242.340 939.300 ;
        RECT 1192.900 932.500 1242.340 934.100 ;
        RECT 1289.500 934.100 1291.100 939.300 ;
        RECT 1337.340 939.300 1387.700 940.900 ;
        RECT 1337.340 934.100 1338.940 939.300 ;
        RECT 1289.500 932.500 1338.940 934.100 ;
        RECT 1386.100 934.100 1387.700 939.300 ;
        RECT 1433.940 939.300 1484.300 940.900 ;
        RECT 1433.940 934.100 1435.540 939.300 ;
        RECT 1386.100 932.500 1435.540 934.100 ;
        RECT 1482.700 934.100 1484.300 939.300 ;
        RECT 1530.540 939.300 1580.900 940.900 ;
        RECT 1530.540 934.100 1532.140 939.300 ;
        RECT 1482.700 932.500 1532.140 934.100 ;
        RECT 1579.300 934.100 1580.900 939.300 ;
        RECT 1627.140 939.300 1677.500 940.900 ;
        RECT 1627.140 934.100 1628.740 939.300 ;
        RECT 1579.300 932.500 1628.740 934.100 ;
        RECT 1675.900 934.100 1677.500 939.300 ;
        RECT 1723.740 939.300 1774.100 940.900 ;
        RECT 1723.740 934.100 1725.340 939.300 ;
        RECT 1675.900 932.500 1725.340 934.100 ;
        RECT 1772.500 934.100 1774.100 939.300 ;
        RECT 1820.340 939.300 1870.700 940.900 ;
        RECT 1820.340 934.100 1821.940 939.300 ;
        RECT 1772.500 932.500 1821.940 934.100 ;
        RECT 1869.100 934.100 1870.700 939.300 ;
        RECT 1916.940 939.300 1967.300 940.900 ;
        RECT 1916.940 934.100 1918.540 939.300 ;
        RECT 1869.100 932.500 1918.540 934.100 ;
        RECT 1965.700 934.100 1967.300 939.300 ;
        RECT 2013.540 939.300 2063.900 940.900 ;
        RECT 2013.540 934.100 2015.140 939.300 ;
        RECT 1965.700 932.500 2015.140 934.100 ;
        RECT 2062.300 934.100 2063.900 939.300 ;
        RECT 2110.140 939.300 2160.500 940.900 ;
        RECT 2110.140 934.100 2111.740 939.300 ;
        RECT 2062.300 932.500 2111.740 934.100 ;
        RECT 2158.900 934.100 2160.500 939.300 ;
        RECT 2206.740 939.300 2257.100 940.900 ;
        RECT 2206.740 934.100 2208.340 939.300 ;
        RECT 2158.900 932.500 2208.340 934.100 ;
        RECT 2255.500 934.100 2257.100 939.300 ;
        RECT 2303.340 939.300 2353.700 940.900 ;
        RECT 2303.340 934.100 2304.940 939.300 ;
        RECT 2255.500 932.500 2304.940 934.100 ;
        RECT 2352.100 934.100 2353.700 939.300 ;
        RECT 2399.940 939.300 2450.300 940.900 ;
        RECT 2399.940 934.100 2401.540 939.300 ;
        RECT 2352.100 932.500 2401.540 934.100 ;
        RECT 2448.700 934.100 2450.300 939.300 ;
        RECT 2524.140 939.300 2546.900 940.900 ;
        RECT 2524.140 937.500 2525.740 939.300 ;
        RECT 2476.300 935.900 2525.740 937.500 ;
        RECT 2476.300 934.100 2477.900 935.900 ;
        RECT 2448.700 932.500 2477.900 934.100 ;
        RECT 2545.300 934.100 2546.900 939.300 ;
        RECT 2575.660 939.300 2660.060 940.900 ;
        RECT 2575.660 934.100 2577.260 939.300 ;
        RECT 2545.300 932.500 2577.260 934.100 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 676.270 3264.580 676.590 3264.640 ;
        RECT 2614.710 3264.580 2615.030 3264.640 ;
        RECT 676.270 3264.440 2615.030 3264.580 ;
        RECT 676.270 3264.380 676.590 3264.440 ;
        RECT 2614.710 3264.380 2615.030 3264.440 ;
        RECT 2614.710 3249.960 2615.030 3250.020 ;
        RECT 2900.830 3249.960 2901.150 3250.020 ;
        RECT 2614.710 3249.820 2901.150 3249.960 ;
        RECT 2614.710 3249.760 2615.030 3249.820 ;
        RECT 2900.830 3249.760 2901.150 3249.820 ;
      LAYER via ;
        RECT 676.300 3264.380 676.560 3264.640 ;
        RECT 2614.740 3264.380 2615.000 3264.640 ;
        RECT 2614.740 3249.760 2615.000 3250.020 ;
        RECT 2900.860 3249.760 2901.120 3250.020 ;
      LAYER met2 ;
        RECT 676.300 3264.350 676.560 3264.670 ;
        RECT 2614.740 3264.350 2615.000 3264.670 ;
        RECT 676.360 3260.000 676.500 3264.350 ;
        RECT 676.250 3256.000 676.530 3260.000 ;
        RECT 2614.800 3250.050 2614.940 3264.350 ;
        RECT 2614.740 3249.730 2615.000 3250.050 ;
        RECT 2900.860 3249.730 2901.120 3250.050 ;
        RECT 2900.920 3245.485 2901.060 3249.730 ;
        RECT 2900.850 3245.115 2901.130 3245.485 ;
      LAYER via2 ;
        RECT 2900.850 3245.160 2901.130 3245.440 ;
      LAYER met3 ;
        RECT 2900.825 3245.450 2901.155 3245.465 ;
        RECT 2917.600 3245.450 2924.800 3245.900 ;
        RECT 2900.825 3245.150 2924.800 3245.450 ;
        RECT 2900.825 3245.135 2901.155 3245.150 ;
        RECT 2917.600 3244.700 2924.800 3245.150 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2866.790 3477.760 2867.110 3477.820 ;
        RECT 2900.830 3477.760 2901.150 3477.820 ;
        RECT 2866.790 3477.620 2901.150 3477.760 ;
        RECT 2866.790 3477.560 2867.110 3477.620 ;
        RECT 2900.830 3477.560 2901.150 3477.620 ;
        RECT 770.110 255.240 770.430 255.300 ;
        RECT 2866.790 255.240 2867.110 255.300 ;
        RECT 770.110 255.100 2867.110 255.240 ;
        RECT 770.110 255.040 770.430 255.100 ;
        RECT 2866.790 255.040 2867.110 255.100 ;
      LAYER via ;
        RECT 2866.820 3477.560 2867.080 3477.820 ;
        RECT 2900.860 3477.560 2901.120 3477.820 ;
        RECT 770.140 255.040 770.400 255.300 ;
        RECT 2866.820 255.040 2867.080 255.300 ;
      LAYER met2 ;
        RECT 2900.850 3479.715 2901.130 3480.085 ;
        RECT 2900.920 3477.850 2901.060 3479.715 ;
        RECT 2866.820 3477.530 2867.080 3477.850 ;
        RECT 2900.860 3477.530 2901.120 3477.850 ;
        RECT 770.090 260.000 770.370 264.000 ;
        RECT 770.200 255.330 770.340 260.000 ;
        RECT 2866.880 255.330 2867.020 3477.530 ;
        RECT 770.140 255.010 770.400 255.330 ;
        RECT 2866.820 255.010 2867.080 255.330 ;
      LAYER via2 ;
        RECT 2900.850 3479.760 2901.130 3480.040 ;
      LAYER met3 ;
        RECT 2900.825 3480.050 2901.155 3480.065 ;
        RECT 2917.600 3480.050 2924.800 3480.500 ;
        RECT 2900.825 3479.750 2924.800 3480.050 ;
        RECT 2900.825 3479.735 2901.155 3479.750 ;
        RECT 2917.600 3479.300 2924.800 3479.750 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2642.770 3487.960 2643.090 3488.020 ;
        RECT 2649.210 3487.960 2649.530 3488.020 ;
        RECT 2642.770 3487.820 2649.530 3487.960 ;
        RECT 2642.770 3487.760 2643.090 3487.820 ;
        RECT 2649.210 3487.760 2649.530 3487.820 ;
        RECT 2615.170 847.180 2615.490 847.240 ;
        RECT 2642.770 847.180 2643.090 847.240 ;
        RECT 2615.170 847.040 2643.090 847.180 ;
        RECT 2615.170 846.980 2615.490 847.040 ;
        RECT 2642.770 846.980 2643.090 847.040 ;
      LAYER via ;
        RECT 2642.800 3487.760 2643.060 3488.020 ;
        RECT 2649.240 3487.760 2649.500 3488.020 ;
        RECT 2615.200 846.980 2615.460 847.240 ;
        RECT 2642.800 846.980 2643.060 847.240 ;
      LAYER met2 ;
        RECT 2649.090 3517.600 2649.650 3524.800 ;
        RECT 2649.300 3488.050 2649.440 3517.600 ;
        RECT 2642.800 3487.730 2643.060 3488.050 ;
        RECT 2649.240 3487.730 2649.500 3488.050 ;
        RECT 2642.860 847.270 2643.000 3487.730 ;
        RECT 2615.200 846.950 2615.460 847.270 ;
        RECT 2642.800 846.950 2643.060 847.270 ;
        RECT 2615.260 846.445 2615.400 846.950 ;
        RECT 2615.190 846.075 2615.470 846.445 ;
      LAYER via2 ;
        RECT 2615.190 846.120 2615.470 846.400 ;
      LAYER met3 ;
        RECT 2606.000 846.410 2610.000 846.800 ;
        RECT 2615.165 846.410 2615.495 846.425 ;
        RECT 2606.000 846.200 2615.495 846.410 ;
        RECT 2609.580 846.110 2615.495 846.200 ;
        RECT 2615.165 846.095 2615.495 846.110 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 260.890 3501.900 261.210 3501.960 ;
        RECT 2324.910 3501.900 2325.230 3501.960 ;
        RECT 260.890 3501.760 2325.230 3501.900 ;
        RECT 260.890 3501.700 261.210 3501.760 ;
        RECT 2324.910 3501.700 2325.230 3501.760 ;
        RECT 260.890 793.460 261.210 793.520 ;
        RECT 296.770 793.460 297.090 793.520 ;
        RECT 260.890 793.320 297.090 793.460 ;
        RECT 260.890 793.260 261.210 793.320 ;
        RECT 296.770 793.260 297.090 793.320 ;
      LAYER via ;
        RECT 260.920 3501.700 261.180 3501.960 ;
        RECT 2324.940 3501.700 2325.200 3501.960 ;
        RECT 260.920 793.260 261.180 793.520 ;
        RECT 296.800 793.260 297.060 793.520 ;
      LAYER met2 ;
        RECT 2324.790 3517.600 2325.350 3524.800 ;
        RECT 2325.000 3501.990 2325.140 3517.600 ;
        RECT 260.920 3501.670 261.180 3501.990 ;
        RECT 2324.940 3501.670 2325.200 3501.990 ;
        RECT 260.980 793.550 261.120 3501.670 ;
        RECT 260.920 793.230 261.180 793.550 ;
        RECT 296.800 793.230 297.060 793.550 ;
        RECT 296.860 792.045 297.000 793.230 ;
        RECT 296.790 791.675 297.070 792.045 ;
      LAYER via2 ;
        RECT 296.790 791.720 297.070 792.000 ;
      LAYER met3 ;
        RECT 296.765 792.010 297.095 792.025 ;
        RECT 310.000 792.010 314.000 792.400 ;
        RECT 296.765 791.800 314.000 792.010 ;
        RECT 296.765 791.710 310.500 791.800 ;
        RECT 296.765 791.695 297.095 791.710 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2000.610 3329.180 2000.930 3329.240 ;
        RECT 2609.650 3329.180 2609.970 3329.240 ;
        RECT 2000.610 3329.040 2609.970 3329.180 ;
        RECT 2000.610 3328.980 2000.930 3329.040 ;
        RECT 2609.650 3328.980 2609.970 3329.040 ;
      LAYER via ;
        RECT 2000.640 3328.980 2000.900 3329.240 ;
        RECT 2609.680 3328.980 2609.940 3329.240 ;
      LAYER met2 ;
        RECT 2000.490 3517.600 2001.050 3524.800 ;
        RECT 2000.700 3329.270 2000.840 3517.600 ;
        RECT 2000.640 3328.950 2000.900 3329.270 ;
        RECT 2609.680 3328.950 2609.940 3329.270 ;
        RECT 2609.740 1757.645 2609.880 3328.950 ;
        RECT 2609.670 1757.275 2609.950 1757.645 ;
      LAYER via2 ;
        RECT 2609.670 1757.320 2609.950 1757.600 ;
      LAYER met3 ;
        RECT 2609.645 1757.610 2609.975 1757.625 ;
        RECT 2609.430 1757.295 2609.975 1757.610 ;
        RECT 2609.430 1755.280 2609.730 1757.295 ;
        RECT 2606.000 1754.680 2610.000 1755.280 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1675.850 3502.920 1676.170 3502.980 ;
        RECT 2671.290 3502.920 2671.610 3502.980 ;
        RECT 1675.850 3502.780 2671.610 3502.920 ;
        RECT 1675.850 3502.720 1676.170 3502.780 ;
        RECT 2671.290 3502.720 2671.610 3502.780 ;
      LAYER via ;
        RECT 1675.880 3502.720 1676.140 3502.980 ;
        RECT 2671.320 3502.720 2671.580 3502.980 ;
      LAYER met2 ;
        RECT 1675.730 3517.600 1676.290 3524.800 ;
        RECT 1675.940 3503.010 1676.080 3517.600 ;
        RECT 1675.880 3502.690 1676.140 3503.010 ;
        RECT 2671.320 3502.690 2671.580 3503.010 ;
        RECT 2157.450 260.000 2157.730 264.000 ;
        RECT 2157.560 247.365 2157.700 260.000 ;
        RECT 2671.380 247.365 2671.520 3502.690 ;
        RECT 2157.490 246.995 2157.770 247.365 ;
        RECT 2671.310 246.995 2671.590 247.365 ;
      LAYER via2 ;
        RECT 2157.490 247.040 2157.770 247.320 ;
        RECT 2671.310 247.040 2671.590 247.320 ;
      LAYER met3 ;
        RECT 2157.465 247.330 2157.795 247.345 ;
        RECT 2671.285 247.330 2671.615 247.345 ;
        RECT 2157.465 247.030 2671.615 247.330 ;
        RECT 2157.465 247.015 2157.795 247.030 ;
        RECT 2671.285 247.015 2671.615 247.030 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 230.070 3502.920 230.390 3502.980 ;
        RECT 1351.550 3502.920 1351.870 3502.980 ;
        RECT 230.070 3502.780 1351.870 3502.920 ;
        RECT 230.070 3502.720 230.390 3502.780 ;
        RECT 1351.550 3502.720 1351.870 3502.780 ;
      LAYER via ;
        RECT 230.100 3502.720 230.360 3502.980 ;
        RECT 1351.580 3502.720 1351.840 3502.980 ;
      LAYER met2 ;
        RECT 1351.430 3517.600 1351.990 3524.800 ;
        RECT 1351.640 3503.010 1351.780 3517.600 ;
        RECT 230.100 3502.690 230.360 3503.010 ;
        RECT 1351.580 3502.690 1351.840 3503.010 ;
        RECT 230.160 248.045 230.300 3502.690 ;
        RECT 656.010 260.000 656.290 264.000 ;
        RECT 656.120 248.045 656.260 260.000 ;
        RECT 230.090 247.675 230.370 248.045 ;
        RECT 656.050 247.675 656.330 248.045 ;
      LAYER via2 ;
        RECT 230.090 247.720 230.370 248.000 ;
        RECT 656.050 247.720 656.330 248.000 ;
      LAYER met3 ;
        RECT 230.065 248.010 230.395 248.025 ;
        RECT 656.025 248.010 656.355 248.025 ;
        RECT 230.065 247.710 656.355 248.010 ;
        RECT 230.065 247.695 230.395 247.710 ;
        RECT 656.025 247.695 656.355 247.710 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 776.550 3278.520 776.870 3278.580 ;
        RECT 2770.190 3278.520 2770.510 3278.580 ;
        RECT 776.550 3278.380 2770.510 3278.520 ;
        RECT 776.550 3278.320 776.870 3278.380 ;
        RECT 2770.190 3278.320 2770.510 3278.380 ;
        RECT 2770.190 434.760 2770.510 434.820 ;
        RECT 2900.830 434.760 2901.150 434.820 ;
        RECT 2770.190 434.620 2901.150 434.760 ;
        RECT 2770.190 434.560 2770.510 434.620 ;
        RECT 2900.830 434.560 2901.150 434.620 ;
      LAYER via ;
        RECT 776.580 3278.320 776.840 3278.580 ;
        RECT 2770.220 3278.320 2770.480 3278.580 ;
        RECT 2770.220 434.560 2770.480 434.820 ;
        RECT 2900.860 434.560 2901.120 434.820 ;
      LAYER met2 ;
        RECT 776.580 3278.290 776.840 3278.610 ;
        RECT 2770.220 3278.290 2770.480 3278.610 ;
        RECT 776.640 3260.000 776.780 3278.290 ;
        RECT 776.530 3256.000 776.810 3260.000 ;
        RECT 2770.280 434.850 2770.420 3278.290 ;
        RECT 2770.220 434.530 2770.480 434.850 ;
        RECT 2900.860 434.530 2901.120 434.850 ;
        RECT 2900.920 430.285 2901.060 434.530 ;
        RECT 2900.850 429.915 2901.130 430.285 ;
      LAYER via2 ;
        RECT 2900.850 429.960 2901.130 430.240 ;
      LAYER met3 ;
        RECT 2900.825 430.250 2901.155 430.265 ;
        RECT 2917.600 430.250 2924.800 430.700 ;
        RECT 2900.825 429.950 2924.800 430.250 ;
        RECT 2900.825 429.935 2901.155 429.950 ;
        RECT 2917.600 429.500 2924.800 429.950 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1025.945 3429.325 1026.115 3477.435 ;
        RECT 1027.785 3332.765 1027.955 3380.875 ;
      LAYER mcon ;
        RECT 1025.945 3477.265 1026.115 3477.435 ;
        RECT 1027.785 3380.705 1027.955 3380.875 ;
      LAYER met1 ;
        RECT 1025.870 3477.420 1026.190 3477.480 ;
        RECT 1025.675 3477.280 1026.190 3477.420 ;
        RECT 1025.870 3477.220 1026.190 3477.280 ;
        RECT 1025.885 3429.480 1026.175 3429.525 ;
        RECT 1026.330 3429.480 1026.650 3429.540 ;
        RECT 1025.885 3429.340 1026.650 3429.480 ;
        RECT 1025.885 3429.295 1026.175 3429.340 ;
        RECT 1026.330 3429.280 1026.650 3429.340 ;
        RECT 1026.790 3394.800 1027.110 3394.860 ;
        RECT 1027.710 3394.800 1028.030 3394.860 ;
        RECT 1026.790 3394.660 1028.030 3394.800 ;
        RECT 1026.790 3394.600 1027.110 3394.660 ;
        RECT 1027.710 3394.600 1028.030 3394.660 ;
        RECT 1027.710 3380.860 1028.030 3380.920 ;
        RECT 1027.515 3380.720 1028.030 3380.860 ;
        RECT 1027.710 3380.660 1028.030 3380.720 ;
        RECT 1027.710 3332.920 1028.030 3332.980 ;
        RECT 1027.515 3332.780 1028.030 3332.920 ;
        RECT 1027.710 3332.720 1028.030 3332.780 ;
        RECT 1027.710 3287.700 1028.030 3287.760 ;
        RECT 2617.010 3287.700 2617.330 3287.760 ;
        RECT 1027.710 3287.560 2617.330 3287.700 ;
        RECT 1027.710 3287.500 1028.030 3287.560 ;
        RECT 2617.010 3287.500 2617.330 3287.560 ;
      LAYER via ;
        RECT 1025.900 3477.220 1026.160 3477.480 ;
        RECT 1026.360 3429.280 1026.620 3429.540 ;
        RECT 1026.820 3394.600 1027.080 3394.860 ;
        RECT 1027.740 3394.600 1028.000 3394.860 ;
        RECT 1027.740 3380.660 1028.000 3380.920 ;
        RECT 1027.740 3332.720 1028.000 3332.980 ;
        RECT 1027.740 3287.500 1028.000 3287.760 ;
        RECT 2617.040 3287.500 2617.300 3287.760 ;
      LAYER met2 ;
        RECT 1027.130 3517.600 1027.690 3524.800 ;
        RECT 1027.340 3517.370 1027.480 3517.600 ;
        RECT 1026.420 3517.230 1027.480 3517.370 ;
        RECT 1026.420 3491.530 1026.560 3517.230 ;
        RECT 1025.960 3491.390 1026.560 3491.530 ;
        RECT 1025.960 3477.510 1026.100 3491.390 ;
        RECT 1025.900 3477.190 1026.160 3477.510 ;
        RECT 1026.360 3429.250 1026.620 3429.570 ;
        RECT 1026.420 3394.970 1026.560 3429.250 ;
        RECT 1026.420 3394.890 1027.020 3394.970 ;
        RECT 1026.420 3394.830 1027.080 3394.890 ;
        RECT 1026.820 3394.570 1027.080 3394.830 ;
        RECT 1027.740 3394.570 1028.000 3394.890 ;
        RECT 1027.800 3380.950 1027.940 3394.570 ;
        RECT 1027.740 3380.630 1028.000 3380.950 ;
        RECT 1027.740 3332.690 1028.000 3333.010 ;
        RECT 1027.800 3287.790 1027.940 3332.690 ;
        RECT 1027.740 3287.470 1028.000 3287.790 ;
        RECT 2617.040 3287.470 2617.300 3287.790 ;
        RECT 2617.100 2959.885 2617.240 3287.470 ;
        RECT 2617.030 2959.515 2617.310 2959.885 ;
      LAYER via2 ;
        RECT 2617.030 2959.560 2617.310 2959.840 ;
      LAYER met3 ;
        RECT 2606.000 2959.850 2610.000 2960.240 ;
        RECT 2617.005 2959.850 2617.335 2959.865 ;
        RECT 2606.000 2959.640 2617.335 2959.850 ;
        RECT 2609.580 2959.550 2617.335 2959.640 ;
        RECT 2617.005 2959.535 2617.335 2959.550 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 702.490 3502.580 702.810 3502.640 ;
        RECT 1863.070 3502.580 1863.390 3502.640 ;
        RECT 702.490 3502.440 1863.390 3502.580 ;
        RECT 702.490 3502.380 702.810 3502.440 ;
        RECT 1863.070 3502.380 1863.390 3502.440 ;
      LAYER via ;
        RECT 702.520 3502.380 702.780 3502.640 ;
        RECT 1863.100 3502.380 1863.360 3502.640 ;
      LAYER met2 ;
        RECT 702.370 3517.600 702.930 3524.800 ;
        RECT 702.580 3502.670 702.720 3517.600 ;
        RECT 702.520 3502.350 702.780 3502.670 ;
        RECT 1863.100 3502.350 1863.360 3502.670 ;
        RECT 1863.160 3260.000 1863.300 3502.350 ;
        RECT 1863.050 3256.000 1863.330 3260.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 378.265 3429.325 378.435 3477.435 ;
      LAYER mcon ;
        RECT 378.265 3477.265 378.435 3477.435 ;
      LAYER met1 ;
        RECT 378.190 3477.420 378.510 3477.480 ;
        RECT 377.995 3477.280 378.510 3477.420 ;
        RECT 378.190 3477.220 378.510 3477.280 ;
        RECT 378.205 3429.480 378.495 3429.525 ;
        RECT 379.110 3429.480 379.430 3429.540 ;
        RECT 378.205 3429.340 379.430 3429.480 ;
        RECT 378.205 3429.295 378.495 3429.340 ;
        RECT 379.110 3429.280 379.430 3429.340 ;
        RECT 379.110 3301.640 379.430 3301.700 ;
        RECT 2610.110 3301.640 2610.430 3301.700 ;
        RECT 379.110 3301.500 2610.430 3301.640 ;
        RECT 379.110 3301.440 379.430 3301.500 ;
        RECT 2610.110 3301.440 2610.430 3301.500 ;
      LAYER via ;
        RECT 378.220 3477.220 378.480 3477.480 ;
        RECT 379.140 3429.280 379.400 3429.540 ;
        RECT 379.140 3301.440 379.400 3301.700 ;
        RECT 2610.140 3301.440 2610.400 3301.700 ;
      LAYER met2 ;
        RECT 378.070 3517.600 378.630 3524.800 ;
        RECT 378.280 3477.510 378.420 3517.600 ;
        RECT 378.220 3477.190 378.480 3477.510 ;
        RECT 379.140 3429.250 379.400 3429.570 ;
        RECT 379.200 3301.730 379.340 3429.250 ;
        RECT 379.140 3301.410 379.400 3301.730 ;
        RECT 2610.140 3301.410 2610.400 3301.730 ;
        RECT 2610.200 1735.885 2610.340 3301.410 ;
        RECT 2610.130 1735.515 2610.410 1735.885 ;
      LAYER via2 ;
        RECT 2610.130 1735.560 2610.410 1735.840 ;
      LAYER met3 ;
        RECT 2610.105 1735.850 2610.435 1735.865 ;
        RECT 2609.430 1735.550 2610.435 1735.850 ;
        RECT 2609.430 1733.520 2609.730 1735.550 ;
        RECT 2610.105 1735.535 2610.435 1735.550 ;
        RECT 2606.000 1732.920 2610.000 1733.520 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 53.965 3381.045 54.135 3429.155 ;
        RECT 53.505 2898.245 53.675 2946.355 ;
        RECT 53.965 2704.785 54.135 2719.235 ;
        RECT 53.965 2283.525 54.135 2318.375 ;
        RECT 53.965 2041.785 54.135 2063.035 ;
        RECT 54.425 1980.585 54.595 1994.695 ;
        RECT 53.965 1876.885 54.135 1924.995 ;
        RECT 54.425 1780.325 54.595 1801.575 ;
        RECT 53.965 1732.045 54.135 1779.815 ;
        RECT 53.505 1594.005 53.675 1642.115 ;
        RECT 54.425 1497.445 54.595 1545.555 ;
        RECT 54.425 1449.505 54.595 1463.275 ;
        RECT 54.425 1400.885 54.595 1448.995 ;
        RECT 54.425 1268.965 54.595 1303.815 ;
        RECT 54.425 882.725 54.595 883.915 ;
      LAYER mcon ;
        RECT 53.965 3428.985 54.135 3429.155 ;
        RECT 53.505 2946.185 53.675 2946.355 ;
        RECT 53.965 2719.065 54.135 2719.235 ;
        RECT 53.965 2318.205 54.135 2318.375 ;
        RECT 53.965 2062.865 54.135 2063.035 ;
        RECT 54.425 1994.525 54.595 1994.695 ;
        RECT 53.965 1924.825 54.135 1924.995 ;
        RECT 54.425 1801.405 54.595 1801.575 ;
        RECT 53.965 1779.645 54.135 1779.815 ;
        RECT 53.505 1641.945 53.675 1642.115 ;
        RECT 54.425 1545.385 54.595 1545.555 ;
        RECT 54.425 1463.105 54.595 1463.275 ;
        RECT 54.425 1448.825 54.595 1448.995 ;
        RECT 54.425 1303.645 54.595 1303.815 ;
        RECT 54.425 883.745 54.595 883.915 ;
      LAYER met1 ;
        RECT 53.430 3477.760 53.750 3477.820 ;
        RECT 53.890 3477.760 54.210 3477.820 ;
        RECT 53.430 3477.620 54.210 3477.760 ;
        RECT 53.430 3477.560 53.750 3477.620 ;
        RECT 53.890 3477.560 54.210 3477.620 ;
        RECT 53.430 3443.080 53.750 3443.140 ;
        RECT 54.350 3443.080 54.670 3443.140 ;
        RECT 53.430 3442.940 54.670 3443.080 ;
        RECT 53.430 3442.880 53.750 3442.940 ;
        RECT 54.350 3442.880 54.670 3442.940 ;
        RECT 53.905 3429.140 54.195 3429.185 ;
        RECT 54.350 3429.140 54.670 3429.200 ;
        RECT 53.905 3429.000 54.670 3429.140 ;
        RECT 53.905 3428.955 54.195 3429.000 ;
        RECT 54.350 3428.940 54.670 3429.000 ;
        RECT 53.890 3381.200 54.210 3381.260 ;
        RECT 53.695 3381.060 54.210 3381.200 ;
        RECT 53.890 3381.000 54.210 3381.060 ;
        RECT 53.890 3367.600 54.210 3367.660 ;
        RECT 54.810 3367.600 55.130 3367.660 ;
        RECT 53.890 3367.460 55.130 3367.600 ;
        RECT 53.890 3367.400 54.210 3367.460 ;
        RECT 54.810 3367.400 55.130 3367.460 ;
        RECT 53.890 3270.700 54.210 3270.760 ;
        RECT 54.810 3270.700 55.130 3270.760 ;
        RECT 53.890 3270.560 55.130 3270.700 ;
        RECT 53.890 3270.500 54.210 3270.560 ;
        RECT 54.810 3270.500 55.130 3270.560 ;
        RECT 53.890 3174.140 54.210 3174.200 ;
        RECT 54.810 3174.140 55.130 3174.200 ;
        RECT 53.890 3174.000 55.130 3174.140 ;
        RECT 53.890 3173.940 54.210 3174.000 ;
        RECT 54.810 3173.940 55.130 3174.000 ;
        RECT 53.890 3077.580 54.210 3077.640 ;
        RECT 54.810 3077.580 55.130 3077.640 ;
        RECT 53.890 3077.440 55.130 3077.580 ;
        RECT 53.890 3077.380 54.210 3077.440 ;
        RECT 54.810 3077.380 55.130 3077.440 ;
        RECT 53.890 2981.020 54.210 2981.080 ;
        RECT 54.810 2981.020 55.130 2981.080 ;
        RECT 53.890 2980.880 55.130 2981.020 ;
        RECT 53.890 2980.820 54.210 2980.880 ;
        RECT 54.810 2980.820 55.130 2980.880 ;
        RECT 53.445 2946.340 53.735 2946.385 ;
        RECT 53.890 2946.340 54.210 2946.400 ;
        RECT 53.445 2946.200 54.210 2946.340 ;
        RECT 53.445 2946.155 53.735 2946.200 ;
        RECT 53.890 2946.140 54.210 2946.200 ;
        RECT 53.430 2898.400 53.750 2898.460 ;
        RECT 53.235 2898.260 53.750 2898.400 ;
        RECT 53.430 2898.200 53.750 2898.260 ;
        RECT 53.890 2719.220 54.210 2719.280 ;
        RECT 53.695 2719.080 54.210 2719.220 ;
        RECT 53.890 2719.020 54.210 2719.080 ;
        RECT 53.890 2704.940 54.210 2705.000 ;
        RECT 53.695 2704.800 54.210 2704.940 ;
        RECT 53.890 2704.740 54.210 2704.800 ;
        RECT 53.890 2670.600 54.210 2670.660 ;
        RECT 54.810 2670.600 55.130 2670.660 ;
        RECT 53.890 2670.460 55.130 2670.600 ;
        RECT 53.890 2670.400 54.210 2670.460 ;
        RECT 54.810 2670.400 55.130 2670.460 ;
        RECT 54.350 2622.660 54.670 2622.720 ;
        RECT 53.980 2622.520 54.670 2622.660 ;
        RECT 53.980 2622.040 54.120 2622.520 ;
        RECT 54.350 2622.460 54.670 2622.520 ;
        RECT 53.890 2621.780 54.210 2622.040 ;
        RECT 52.970 2560.100 53.290 2560.160 ;
        RECT 54.350 2560.100 54.670 2560.160 ;
        RECT 52.970 2559.960 54.670 2560.100 ;
        RECT 52.970 2559.900 53.290 2559.960 ;
        RECT 54.350 2559.900 54.670 2559.960 ;
        RECT 54.350 2525.560 54.670 2525.820 ;
        RECT 54.440 2525.420 54.580 2525.560 ;
        RECT 54.810 2525.420 55.130 2525.480 ;
        RECT 54.440 2525.280 55.130 2525.420 ;
        RECT 54.810 2525.220 55.130 2525.280 ;
        RECT 53.890 2429.000 54.210 2429.260 ;
        RECT 53.980 2428.520 54.120 2429.000 ;
        RECT 54.350 2428.520 54.670 2428.580 ;
        RECT 53.980 2428.380 54.670 2428.520 ;
        RECT 54.350 2428.320 54.670 2428.380 ;
        RECT 52.970 2414.920 53.290 2414.980 ;
        RECT 54.350 2414.920 54.670 2414.980 ;
        RECT 52.970 2414.780 54.670 2414.920 ;
        RECT 52.970 2414.720 53.290 2414.780 ;
        RECT 54.350 2414.720 54.670 2414.780 ;
        RECT 53.890 2332.440 54.210 2332.700 ;
        RECT 53.980 2332.020 54.120 2332.440 ;
        RECT 53.890 2331.760 54.210 2332.020 ;
        RECT 53.890 2318.360 54.210 2318.420 ;
        RECT 53.695 2318.220 54.210 2318.360 ;
        RECT 53.890 2318.160 54.210 2318.220 ;
        RECT 53.890 2283.680 54.210 2283.740 ;
        RECT 53.695 2283.540 54.210 2283.680 ;
        RECT 53.890 2283.480 54.210 2283.540 ;
        RECT 53.430 2236.760 53.750 2236.820 ;
        RECT 54.350 2236.760 54.670 2236.820 ;
        RECT 53.430 2236.620 54.670 2236.760 ;
        RECT 53.430 2236.560 53.750 2236.620 ;
        RECT 54.350 2236.560 54.670 2236.620 ;
        RECT 53.890 2138.980 54.210 2139.240 ;
        RECT 53.980 2138.840 54.120 2138.980 ;
        RECT 54.350 2138.840 54.670 2138.900 ;
        RECT 53.980 2138.700 54.670 2138.840 ;
        RECT 54.350 2138.640 54.670 2138.700 ;
        RECT 53.890 2063.020 54.210 2063.080 ;
        RECT 53.695 2062.880 54.210 2063.020 ;
        RECT 53.890 2062.820 54.210 2062.880 ;
        RECT 53.905 2041.940 54.195 2041.985 ;
        RECT 54.350 2041.940 54.670 2042.000 ;
        RECT 53.905 2041.800 54.670 2041.940 ;
        RECT 53.905 2041.755 54.195 2041.800 ;
        RECT 54.350 2041.740 54.670 2041.800 ;
        RECT 54.350 1994.680 54.670 1994.740 ;
        RECT 54.155 1994.540 54.670 1994.680 ;
        RECT 54.350 1994.480 54.670 1994.540 ;
        RECT 53.890 1980.740 54.210 1980.800 ;
        RECT 54.365 1980.740 54.655 1980.785 ;
        RECT 53.890 1980.600 54.655 1980.740 ;
        RECT 53.890 1980.540 54.210 1980.600 ;
        RECT 54.365 1980.555 54.655 1980.600 ;
        RECT 53.430 1945.860 53.750 1946.120 ;
        RECT 53.520 1945.380 53.660 1945.860 ;
        RECT 53.890 1945.380 54.210 1945.440 ;
        RECT 53.520 1945.240 54.210 1945.380 ;
        RECT 53.890 1945.180 54.210 1945.240 ;
        RECT 53.890 1924.980 54.210 1925.040 ;
        RECT 53.695 1924.840 54.210 1924.980 ;
        RECT 53.890 1924.780 54.210 1924.840 ;
        RECT 53.905 1877.040 54.195 1877.085 ;
        RECT 54.810 1877.040 55.130 1877.100 ;
        RECT 53.905 1876.900 55.130 1877.040 ;
        RECT 53.905 1876.855 54.195 1876.900 ;
        RECT 54.810 1876.840 55.130 1876.900 ;
        RECT 54.350 1828.760 54.670 1828.820 ;
        RECT 54.810 1828.760 55.130 1828.820 ;
        RECT 54.350 1828.620 55.130 1828.760 ;
        RECT 54.350 1828.560 54.670 1828.620 ;
        RECT 54.810 1828.560 55.130 1828.620 ;
        RECT 54.350 1801.560 54.670 1801.620 ;
        RECT 54.155 1801.420 54.670 1801.560 ;
        RECT 54.350 1801.360 54.670 1801.420 ;
        RECT 54.350 1780.480 54.670 1780.540 ;
        RECT 54.155 1780.340 54.670 1780.480 ;
        RECT 54.350 1780.280 54.670 1780.340 ;
        RECT 53.905 1779.800 54.195 1779.845 ;
        RECT 54.350 1779.800 54.670 1779.860 ;
        RECT 53.905 1779.660 54.670 1779.800 ;
        RECT 53.905 1779.615 54.195 1779.660 ;
        RECT 54.350 1779.600 54.670 1779.660 ;
        RECT 53.890 1732.200 54.210 1732.260 ;
        RECT 53.695 1732.060 54.210 1732.200 ;
        RECT 53.890 1732.000 54.210 1732.060 ;
        RECT 53.890 1704.320 54.210 1704.380 ;
        RECT 54.810 1704.320 55.130 1704.380 ;
        RECT 53.890 1704.180 55.130 1704.320 ;
        RECT 53.890 1704.120 54.210 1704.180 ;
        RECT 54.810 1704.120 55.130 1704.180 ;
        RECT 53.430 1666.580 53.750 1666.640 ;
        RECT 54.810 1666.580 55.130 1666.640 ;
        RECT 53.430 1666.440 55.130 1666.580 ;
        RECT 53.430 1666.380 53.750 1666.440 ;
        RECT 54.810 1666.380 55.130 1666.440 ;
        RECT 53.430 1642.100 53.750 1642.160 ;
        RECT 53.235 1641.960 53.750 1642.100 ;
        RECT 53.430 1641.900 53.750 1641.960 ;
        RECT 53.445 1594.160 53.735 1594.205 ;
        RECT 53.890 1594.160 54.210 1594.220 ;
        RECT 53.445 1594.020 54.210 1594.160 ;
        RECT 53.445 1593.975 53.735 1594.020 ;
        RECT 53.890 1593.960 54.210 1594.020 ;
        RECT 54.365 1545.540 54.655 1545.585 ;
        RECT 54.810 1545.540 55.130 1545.600 ;
        RECT 54.365 1545.400 55.130 1545.540 ;
        RECT 54.365 1545.355 54.655 1545.400 ;
        RECT 54.810 1545.340 55.130 1545.400 ;
        RECT 54.350 1497.600 54.670 1497.660 ;
        RECT 54.155 1497.460 54.670 1497.600 ;
        RECT 54.350 1497.400 54.670 1497.460 ;
        RECT 54.350 1463.260 54.670 1463.320 ;
        RECT 54.155 1463.120 54.670 1463.260 ;
        RECT 54.350 1463.060 54.670 1463.120 ;
        RECT 54.365 1449.660 54.655 1449.705 ;
        RECT 54.810 1449.660 55.130 1449.720 ;
        RECT 54.365 1449.520 55.130 1449.660 ;
        RECT 54.365 1449.475 54.655 1449.520 ;
        RECT 54.810 1449.460 55.130 1449.520 ;
        RECT 54.350 1448.980 54.670 1449.040 ;
        RECT 54.155 1448.840 54.670 1448.980 ;
        RECT 54.350 1448.780 54.670 1448.840 ;
        RECT 54.365 1401.040 54.655 1401.085 ;
        RECT 54.810 1401.040 55.130 1401.100 ;
        RECT 54.365 1400.900 55.130 1401.040 ;
        RECT 54.365 1400.855 54.655 1400.900 ;
        RECT 54.810 1400.840 55.130 1400.900 ;
        RECT 53.890 1318.420 54.210 1318.480 ;
        RECT 53.520 1318.280 54.210 1318.420 ;
        RECT 53.520 1317.800 53.660 1318.280 ;
        RECT 53.890 1318.220 54.210 1318.280 ;
        RECT 53.430 1317.540 53.750 1317.800 ;
        RECT 53.430 1303.940 53.750 1304.200 ;
        RECT 53.520 1303.800 53.660 1303.940 ;
        RECT 54.365 1303.800 54.655 1303.845 ;
        RECT 53.520 1303.660 54.655 1303.800 ;
        RECT 54.365 1303.615 54.655 1303.660 ;
        RECT 54.350 1269.120 54.670 1269.180 ;
        RECT 54.155 1268.980 54.670 1269.120 ;
        RECT 54.350 1268.920 54.670 1268.980 ;
        RECT 54.350 1255.860 54.670 1255.920 ;
        RECT 54.810 1255.860 55.130 1255.920 ;
        RECT 54.350 1255.720 55.130 1255.860 ;
        RECT 54.350 1255.660 54.670 1255.720 ;
        RECT 54.810 1255.660 55.130 1255.720 ;
        RECT 54.810 1173.240 55.130 1173.300 ;
        RECT 54.440 1173.100 55.130 1173.240 ;
        RECT 54.440 1172.620 54.580 1173.100 ;
        RECT 54.810 1173.040 55.130 1173.100 ;
        RECT 54.350 1172.360 54.670 1172.620 ;
        RECT 53.430 1062.740 53.750 1062.800 ;
        RECT 53.890 1062.740 54.210 1062.800 ;
        RECT 53.430 1062.600 54.210 1062.740 ;
        RECT 53.430 1062.540 53.750 1062.600 ;
        RECT 53.890 1062.540 54.210 1062.600 ;
        RECT 53.430 1028.060 53.750 1028.120 ;
        RECT 54.350 1028.060 54.670 1028.120 ;
        RECT 53.430 1027.920 54.670 1028.060 ;
        RECT 53.430 1027.860 53.750 1027.920 ;
        RECT 54.350 1027.860 54.670 1027.920 ;
        RECT 54.350 980.460 54.670 980.520 ;
        RECT 53.980 980.320 54.670 980.460 ;
        RECT 53.980 979.840 54.120 980.320 ;
        RECT 54.350 980.260 54.670 980.320 ;
        RECT 53.890 979.580 54.210 979.840 ;
        RECT 52.970 917.900 53.290 917.960 ;
        RECT 54.350 917.900 54.670 917.960 ;
        RECT 52.970 917.760 54.670 917.900 ;
        RECT 52.970 917.700 53.290 917.760 ;
        RECT 54.350 917.700 54.670 917.760 ;
        RECT 54.350 883.900 54.670 883.960 ;
        RECT 54.155 883.760 54.670 883.900 ;
        RECT 54.350 883.700 54.670 883.760 ;
        RECT 54.350 882.880 54.670 882.940 ;
        RECT 54.155 882.740 54.670 882.880 ;
        RECT 54.350 882.680 54.670 882.740 ;
        RECT 52.970 845.480 53.290 845.540 ;
        RECT 53.890 845.480 54.210 845.540 ;
        RECT 52.970 845.340 54.210 845.480 ;
        RECT 52.970 845.280 53.290 845.340 ;
        RECT 53.890 845.280 54.210 845.340 ;
        RECT 53.890 786.800 54.210 787.060 ;
        RECT 53.980 786.320 54.120 786.800 ;
        RECT 54.810 786.320 55.130 786.380 ;
        RECT 53.980 786.180 55.130 786.320 ;
        RECT 54.810 786.120 55.130 786.180 ;
        RECT 54.810 772.720 55.130 772.780 ;
        RECT 55.730 772.720 56.050 772.780 ;
        RECT 54.810 772.580 56.050 772.720 ;
        RECT 54.810 772.520 55.130 772.580 ;
        RECT 55.730 772.520 56.050 772.580 ;
        RECT 54.350 690.440 54.670 690.500 ;
        RECT 53.980 690.300 54.670 690.440 ;
        RECT 53.980 689.820 54.120 690.300 ;
        RECT 54.350 690.240 54.670 690.300 ;
        RECT 53.890 689.560 54.210 689.820 ;
        RECT 52.510 676.160 52.830 676.220 ;
        RECT 53.890 676.160 54.210 676.220 ;
        RECT 52.510 676.020 54.210 676.160 ;
        RECT 52.510 675.960 52.830 676.020 ;
        RECT 53.890 675.960 54.210 676.020 ;
        RECT 53.430 593.340 53.750 593.600 ;
        RECT 53.520 593.200 53.660 593.340 ;
        RECT 54.350 593.200 54.670 593.260 ;
        RECT 53.520 593.060 54.670 593.200 ;
        RECT 54.350 593.000 54.670 593.060 ;
        RECT 52.970 579.600 53.290 579.660 ;
        RECT 54.350 579.600 54.670 579.660 ;
        RECT 52.970 579.460 54.670 579.600 ;
        RECT 52.970 579.400 53.290 579.460 ;
        RECT 54.350 579.400 54.670 579.460 ;
        RECT 53.890 496.780 54.210 497.040 ;
        RECT 53.980 496.640 54.120 496.780 ;
        RECT 54.810 496.640 55.130 496.700 ;
        RECT 53.980 496.500 55.130 496.640 ;
        RECT 54.810 496.440 55.130 496.500 ;
        RECT 53.890 414.020 54.210 414.080 ;
        RECT 296.770 414.020 297.090 414.080 ;
        RECT 53.890 413.880 297.090 414.020 ;
        RECT 53.890 413.820 54.210 413.880 ;
        RECT 296.770 413.820 297.090 413.880 ;
      LAYER via ;
        RECT 53.460 3477.560 53.720 3477.820 ;
        RECT 53.920 3477.560 54.180 3477.820 ;
        RECT 53.460 3442.880 53.720 3443.140 ;
        RECT 54.380 3442.880 54.640 3443.140 ;
        RECT 54.380 3428.940 54.640 3429.200 ;
        RECT 53.920 3381.000 54.180 3381.260 ;
        RECT 53.920 3367.400 54.180 3367.660 ;
        RECT 54.840 3367.400 55.100 3367.660 ;
        RECT 53.920 3270.500 54.180 3270.760 ;
        RECT 54.840 3270.500 55.100 3270.760 ;
        RECT 53.920 3173.940 54.180 3174.200 ;
        RECT 54.840 3173.940 55.100 3174.200 ;
        RECT 53.920 3077.380 54.180 3077.640 ;
        RECT 54.840 3077.380 55.100 3077.640 ;
        RECT 53.920 2980.820 54.180 2981.080 ;
        RECT 54.840 2980.820 55.100 2981.080 ;
        RECT 53.920 2946.140 54.180 2946.400 ;
        RECT 53.460 2898.200 53.720 2898.460 ;
        RECT 53.920 2719.020 54.180 2719.280 ;
        RECT 53.920 2704.740 54.180 2705.000 ;
        RECT 53.920 2670.400 54.180 2670.660 ;
        RECT 54.840 2670.400 55.100 2670.660 ;
        RECT 54.380 2622.460 54.640 2622.720 ;
        RECT 53.920 2621.780 54.180 2622.040 ;
        RECT 53.000 2559.900 53.260 2560.160 ;
        RECT 54.380 2559.900 54.640 2560.160 ;
        RECT 54.380 2525.560 54.640 2525.820 ;
        RECT 54.840 2525.220 55.100 2525.480 ;
        RECT 53.920 2429.000 54.180 2429.260 ;
        RECT 54.380 2428.320 54.640 2428.580 ;
        RECT 53.000 2414.720 53.260 2414.980 ;
        RECT 54.380 2414.720 54.640 2414.980 ;
        RECT 53.920 2332.440 54.180 2332.700 ;
        RECT 53.920 2331.760 54.180 2332.020 ;
        RECT 53.920 2318.160 54.180 2318.420 ;
        RECT 53.920 2283.480 54.180 2283.740 ;
        RECT 53.460 2236.560 53.720 2236.820 ;
        RECT 54.380 2236.560 54.640 2236.820 ;
        RECT 53.920 2138.980 54.180 2139.240 ;
        RECT 54.380 2138.640 54.640 2138.900 ;
        RECT 53.920 2062.820 54.180 2063.080 ;
        RECT 54.380 2041.740 54.640 2042.000 ;
        RECT 54.380 1994.480 54.640 1994.740 ;
        RECT 53.920 1980.540 54.180 1980.800 ;
        RECT 53.460 1945.860 53.720 1946.120 ;
        RECT 53.920 1945.180 54.180 1945.440 ;
        RECT 53.920 1924.780 54.180 1925.040 ;
        RECT 54.840 1876.840 55.100 1877.100 ;
        RECT 54.380 1828.560 54.640 1828.820 ;
        RECT 54.840 1828.560 55.100 1828.820 ;
        RECT 54.380 1801.360 54.640 1801.620 ;
        RECT 54.380 1780.280 54.640 1780.540 ;
        RECT 54.380 1779.600 54.640 1779.860 ;
        RECT 53.920 1732.000 54.180 1732.260 ;
        RECT 53.920 1704.120 54.180 1704.380 ;
        RECT 54.840 1704.120 55.100 1704.380 ;
        RECT 53.460 1666.380 53.720 1666.640 ;
        RECT 54.840 1666.380 55.100 1666.640 ;
        RECT 53.460 1641.900 53.720 1642.160 ;
        RECT 53.920 1593.960 54.180 1594.220 ;
        RECT 54.840 1545.340 55.100 1545.600 ;
        RECT 54.380 1497.400 54.640 1497.660 ;
        RECT 54.380 1463.060 54.640 1463.320 ;
        RECT 54.840 1449.460 55.100 1449.720 ;
        RECT 54.380 1448.780 54.640 1449.040 ;
        RECT 54.840 1400.840 55.100 1401.100 ;
        RECT 53.920 1318.220 54.180 1318.480 ;
        RECT 53.460 1317.540 53.720 1317.800 ;
        RECT 53.460 1303.940 53.720 1304.200 ;
        RECT 54.380 1268.920 54.640 1269.180 ;
        RECT 54.380 1255.660 54.640 1255.920 ;
        RECT 54.840 1255.660 55.100 1255.920 ;
        RECT 54.840 1173.040 55.100 1173.300 ;
        RECT 54.380 1172.360 54.640 1172.620 ;
        RECT 53.460 1062.540 53.720 1062.800 ;
        RECT 53.920 1062.540 54.180 1062.800 ;
        RECT 53.460 1027.860 53.720 1028.120 ;
        RECT 54.380 1027.860 54.640 1028.120 ;
        RECT 54.380 980.260 54.640 980.520 ;
        RECT 53.920 979.580 54.180 979.840 ;
        RECT 53.000 917.700 53.260 917.960 ;
        RECT 54.380 917.700 54.640 917.960 ;
        RECT 54.380 883.700 54.640 883.960 ;
        RECT 54.380 882.680 54.640 882.940 ;
        RECT 53.000 845.280 53.260 845.540 ;
        RECT 53.920 845.280 54.180 845.540 ;
        RECT 53.920 786.800 54.180 787.060 ;
        RECT 54.840 786.120 55.100 786.380 ;
        RECT 54.840 772.520 55.100 772.780 ;
        RECT 55.760 772.520 56.020 772.780 ;
        RECT 54.380 690.240 54.640 690.500 ;
        RECT 53.920 689.560 54.180 689.820 ;
        RECT 52.540 675.960 52.800 676.220 ;
        RECT 53.920 675.960 54.180 676.220 ;
        RECT 53.460 593.340 53.720 593.600 ;
        RECT 54.380 593.000 54.640 593.260 ;
        RECT 53.000 579.400 53.260 579.660 ;
        RECT 54.380 579.400 54.640 579.660 ;
        RECT 53.920 496.780 54.180 497.040 ;
        RECT 54.840 496.440 55.100 496.700 ;
        RECT 53.920 413.820 54.180 414.080 ;
        RECT 296.800 413.820 297.060 414.080 ;
      LAYER met2 ;
        RECT 53.770 3517.600 54.330 3524.800 ;
        RECT 53.980 3477.850 54.120 3517.600 ;
        RECT 53.460 3477.530 53.720 3477.850 ;
        RECT 53.920 3477.530 54.180 3477.850 ;
        RECT 53.520 3443.170 53.660 3477.530 ;
        RECT 53.460 3442.850 53.720 3443.170 ;
        RECT 54.380 3442.850 54.640 3443.170 ;
        RECT 54.440 3429.230 54.580 3442.850 ;
        RECT 54.380 3428.910 54.640 3429.230 ;
        RECT 53.920 3380.970 54.180 3381.290 ;
        RECT 53.980 3367.690 54.120 3380.970 ;
        RECT 53.920 3367.370 54.180 3367.690 ;
        RECT 54.840 3367.370 55.100 3367.690 ;
        RECT 54.900 3318.810 55.040 3367.370 ;
        RECT 53.980 3318.670 55.040 3318.810 ;
        RECT 53.980 3270.790 54.120 3318.670 ;
        RECT 53.920 3270.470 54.180 3270.790 ;
        RECT 54.840 3270.470 55.100 3270.790 ;
        RECT 54.900 3222.250 55.040 3270.470 ;
        RECT 53.980 3222.110 55.040 3222.250 ;
        RECT 53.980 3174.230 54.120 3222.110 ;
        RECT 53.920 3173.910 54.180 3174.230 ;
        RECT 54.840 3173.910 55.100 3174.230 ;
        RECT 54.900 3125.690 55.040 3173.910 ;
        RECT 53.980 3125.550 55.040 3125.690 ;
        RECT 53.980 3077.670 54.120 3125.550 ;
        RECT 53.920 3077.350 54.180 3077.670 ;
        RECT 54.840 3077.350 55.100 3077.670 ;
        RECT 54.900 3029.130 55.040 3077.350 ;
        RECT 53.980 3028.990 55.040 3029.130 ;
        RECT 53.980 2981.110 54.120 3028.990 ;
        RECT 53.920 2980.790 54.180 2981.110 ;
        RECT 54.840 2980.850 55.100 2981.110 ;
        RECT 54.440 2980.790 55.100 2980.850 ;
        RECT 54.440 2980.710 55.040 2980.790 ;
        RECT 54.440 2959.770 54.580 2980.710 ;
        RECT 53.980 2959.630 54.580 2959.770 ;
        RECT 53.980 2946.430 54.120 2959.630 ;
        RECT 53.920 2946.110 54.180 2946.430 ;
        RECT 53.460 2898.170 53.720 2898.490 ;
        RECT 53.520 2863.210 53.660 2898.170 ;
        RECT 53.520 2863.070 54.120 2863.210 ;
        RECT 53.980 2815.610 54.120 2863.070 ;
        RECT 53.980 2815.470 54.580 2815.610 ;
        RECT 54.440 2767.330 54.580 2815.470 ;
        RECT 54.440 2767.190 55.040 2767.330 ;
        RECT 54.900 2766.650 55.040 2767.190 ;
        RECT 54.440 2766.510 55.040 2766.650 ;
        RECT 54.440 2753.050 54.580 2766.510 ;
        RECT 53.980 2752.910 54.580 2753.050 ;
        RECT 53.980 2719.310 54.120 2752.910 ;
        RECT 53.920 2718.990 54.180 2719.310 ;
        RECT 53.920 2704.710 54.180 2705.030 ;
        RECT 53.980 2670.690 54.120 2704.710 ;
        RECT 53.920 2670.370 54.180 2670.690 ;
        RECT 54.840 2670.370 55.100 2670.690 ;
        RECT 54.900 2670.090 55.040 2670.370 ;
        RECT 54.440 2669.950 55.040 2670.090 ;
        RECT 54.440 2622.750 54.580 2669.950 ;
        RECT 54.380 2622.430 54.640 2622.750 ;
        RECT 53.920 2621.750 54.180 2622.070 ;
        RECT 53.980 2608.325 54.120 2621.750 ;
        RECT 52.990 2607.955 53.270 2608.325 ;
        RECT 53.910 2607.955 54.190 2608.325 ;
        RECT 53.060 2560.190 53.200 2607.955 ;
        RECT 53.000 2559.870 53.260 2560.190 ;
        RECT 54.380 2559.870 54.640 2560.190 ;
        RECT 54.440 2525.850 54.580 2559.870 ;
        RECT 54.380 2525.530 54.640 2525.850 ;
        RECT 54.840 2525.190 55.100 2525.510 ;
        RECT 54.900 2476.970 55.040 2525.190 ;
        RECT 53.980 2476.830 55.040 2476.970 ;
        RECT 53.980 2429.290 54.120 2476.830 ;
        RECT 53.920 2428.970 54.180 2429.290 ;
        RECT 54.380 2428.290 54.640 2428.610 ;
        RECT 54.440 2415.010 54.580 2428.290 ;
        RECT 53.000 2414.690 53.260 2415.010 ;
        RECT 54.380 2414.690 54.640 2415.010 ;
        RECT 53.060 2366.925 53.200 2414.690 ;
        RECT 52.990 2366.555 53.270 2366.925 ;
        RECT 53.910 2366.555 54.190 2366.925 ;
        RECT 53.980 2332.730 54.120 2366.555 ;
        RECT 53.920 2332.410 54.180 2332.730 ;
        RECT 53.920 2331.730 54.180 2332.050 ;
        RECT 53.980 2318.450 54.120 2331.730 ;
        RECT 53.920 2318.130 54.180 2318.450 ;
        RECT 53.920 2283.450 54.180 2283.770 ;
        RECT 53.980 2270.250 54.120 2283.450 ;
        RECT 53.980 2270.110 54.580 2270.250 ;
        RECT 54.440 2236.850 54.580 2270.110 ;
        RECT 53.460 2236.530 53.720 2236.850 ;
        RECT 54.380 2236.530 54.640 2236.850 ;
        RECT 53.520 2187.290 53.660 2236.530 ;
        RECT 53.520 2187.150 54.120 2187.290 ;
        RECT 53.980 2139.270 54.120 2187.150 ;
        RECT 53.920 2138.950 54.180 2139.270 ;
        RECT 54.380 2138.610 54.640 2138.930 ;
        RECT 54.440 2077.245 54.580 2138.610 ;
        RECT 54.370 2076.875 54.650 2077.245 ;
        RECT 53.910 2070.075 54.190 2070.445 ;
        RECT 53.980 2063.110 54.120 2070.075 ;
        RECT 53.920 2062.790 54.180 2063.110 ;
        RECT 54.380 2041.710 54.640 2042.030 ;
        RECT 54.440 1994.770 54.580 2041.710 ;
        RECT 54.380 1994.450 54.640 1994.770 ;
        RECT 53.920 1980.570 54.180 1980.830 ;
        RECT 53.520 1980.510 54.180 1980.570 ;
        RECT 53.520 1980.430 54.120 1980.510 ;
        RECT 53.520 1946.150 53.660 1980.430 ;
        RECT 53.460 1945.830 53.720 1946.150 ;
        RECT 53.920 1945.150 54.180 1945.470 ;
        RECT 53.980 1925.070 54.120 1945.150 ;
        RECT 53.920 1924.750 54.180 1925.070 ;
        RECT 54.840 1876.810 55.100 1877.130 ;
        RECT 54.900 1828.850 55.040 1876.810 ;
        RECT 54.380 1828.530 54.640 1828.850 ;
        RECT 54.840 1828.530 55.100 1828.850 ;
        RECT 54.440 1801.650 54.580 1828.530 ;
        RECT 54.380 1801.330 54.640 1801.650 ;
        RECT 54.380 1780.250 54.640 1780.570 ;
        RECT 54.440 1779.890 54.580 1780.250 ;
        RECT 54.380 1779.570 54.640 1779.890 ;
        RECT 53.920 1731.970 54.180 1732.290 ;
        RECT 53.980 1704.410 54.120 1731.970 ;
        RECT 53.920 1704.090 54.180 1704.410 ;
        RECT 54.840 1704.090 55.100 1704.410 ;
        RECT 54.900 1666.670 55.040 1704.090 ;
        RECT 53.460 1666.350 53.720 1666.670 ;
        RECT 54.840 1666.350 55.100 1666.670 ;
        RECT 53.520 1642.190 53.660 1666.350 ;
        RECT 53.460 1641.870 53.720 1642.190 ;
        RECT 53.920 1593.930 54.180 1594.250 ;
        RECT 53.980 1559.650 54.120 1593.930 ;
        RECT 53.980 1559.510 55.040 1559.650 ;
        RECT 54.900 1545.630 55.040 1559.510 ;
        RECT 54.840 1545.310 55.100 1545.630 ;
        RECT 54.380 1497.370 54.640 1497.690 ;
        RECT 54.440 1463.350 54.580 1497.370 ;
        RECT 54.380 1463.030 54.640 1463.350 ;
        RECT 54.840 1449.490 55.100 1449.750 ;
        RECT 54.440 1449.430 55.100 1449.490 ;
        RECT 54.440 1449.350 55.040 1449.430 ;
        RECT 54.440 1449.070 54.580 1449.350 ;
        RECT 54.380 1448.750 54.640 1449.070 ;
        RECT 54.840 1400.810 55.100 1401.130 ;
        RECT 54.900 1353.725 55.040 1400.810 ;
        RECT 54.830 1353.355 55.110 1353.725 ;
        RECT 53.450 1352.930 53.730 1353.045 ;
        RECT 53.450 1352.790 54.120 1352.930 ;
        RECT 53.450 1352.675 53.730 1352.790 ;
        RECT 53.980 1318.510 54.120 1352.790 ;
        RECT 53.920 1318.190 54.180 1318.510 ;
        RECT 53.460 1317.510 53.720 1317.830 ;
        RECT 53.520 1304.230 53.660 1317.510 ;
        RECT 53.460 1303.910 53.720 1304.230 ;
        RECT 54.380 1268.890 54.640 1269.210 ;
        RECT 54.440 1255.950 54.580 1268.890 ;
        RECT 54.380 1255.630 54.640 1255.950 ;
        RECT 54.840 1255.630 55.100 1255.950 ;
        RECT 54.900 1173.330 55.040 1255.630 ;
        RECT 54.840 1173.010 55.100 1173.330 ;
        RECT 54.380 1172.330 54.640 1172.650 ;
        RECT 54.440 1124.450 54.580 1172.330 ;
        RECT 53.980 1124.310 54.580 1124.450 ;
        RECT 53.980 1062.830 54.120 1124.310 ;
        RECT 53.460 1062.510 53.720 1062.830 ;
        RECT 53.920 1062.510 54.180 1062.830 ;
        RECT 53.520 1028.150 53.660 1062.510 ;
        RECT 53.460 1027.830 53.720 1028.150 ;
        RECT 54.380 1027.830 54.640 1028.150 ;
        RECT 54.440 980.550 54.580 1027.830 ;
        RECT 54.380 980.230 54.640 980.550 ;
        RECT 53.920 979.550 54.180 979.870 ;
        RECT 53.980 966.125 54.120 979.550 ;
        RECT 52.990 965.755 53.270 966.125 ;
        RECT 53.910 965.755 54.190 966.125 ;
        RECT 53.060 917.990 53.200 965.755 ;
        RECT 53.000 917.670 53.260 917.990 ;
        RECT 54.380 917.670 54.640 917.990 ;
        RECT 54.440 883.990 54.580 917.670 ;
        RECT 54.380 883.670 54.640 883.990 ;
        RECT 54.380 882.650 54.640 882.970 ;
        RECT 54.440 869.450 54.580 882.650 ;
        RECT 53.980 869.310 54.580 869.450 ;
        RECT 53.980 845.570 54.120 869.310 ;
        RECT 53.000 845.250 53.260 845.570 ;
        RECT 53.920 845.250 54.180 845.570 ;
        RECT 53.060 821.285 53.200 845.250 ;
        RECT 52.990 820.915 53.270 821.285 ;
        RECT 53.910 820.915 54.190 821.285 ;
        RECT 53.980 787.090 54.120 820.915 ;
        RECT 53.920 786.770 54.180 787.090 ;
        RECT 54.840 786.090 55.100 786.410 ;
        RECT 54.900 772.810 55.040 786.090 ;
        RECT 54.840 772.490 55.100 772.810 ;
        RECT 55.760 772.490 56.020 772.810 ;
        RECT 55.820 724.725 55.960 772.490 ;
        RECT 54.370 724.355 54.650 724.725 ;
        RECT 55.750 724.355 56.030 724.725 ;
        RECT 54.440 690.530 54.580 724.355 ;
        RECT 54.380 690.210 54.640 690.530 ;
        RECT 53.920 689.530 54.180 689.850 ;
        RECT 53.980 676.250 54.120 689.530 ;
        RECT 52.540 675.930 52.800 676.250 ;
        RECT 53.920 675.930 54.180 676.250 ;
        RECT 52.600 628.165 52.740 675.930 ;
        RECT 52.530 627.795 52.810 628.165 ;
        RECT 53.450 627.795 53.730 628.165 ;
        RECT 53.520 593.630 53.660 627.795 ;
        RECT 53.460 593.310 53.720 593.630 ;
        RECT 54.380 592.970 54.640 593.290 ;
        RECT 54.440 579.690 54.580 592.970 ;
        RECT 53.000 579.370 53.260 579.690 ;
        RECT 54.380 579.370 54.640 579.690 ;
        RECT 53.060 531.605 53.200 579.370 ;
        RECT 52.990 531.235 53.270 531.605 ;
        RECT 53.910 531.235 54.190 531.605 ;
        RECT 53.980 497.070 54.120 531.235 ;
        RECT 53.920 496.750 54.180 497.070 ;
        RECT 54.840 496.410 55.100 496.730 ;
        RECT 54.900 448.530 55.040 496.410 ;
        RECT 53.980 448.390 55.040 448.530 ;
        RECT 53.980 414.110 54.120 448.390 ;
        RECT 53.920 413.790 54.180 414.110 ;
        RECT 296.800 413.790 297.060 414.110 ;
        RECT 296.860 411.245 297.000 413.790 ;
        RECT 296.790 410.875 297.070 411.245 ;
      LAYER via2 ;
        RECT 52.990 2608.000 53.270 2608.280 ;
        RECT 53.910 2608.000 54.190 2608.280 ;
        RECT 52.990 2366.600 53.270 2366.880 ;
        RECT 53.910 2366.600 54.190 2366.880 ;
        RECT 54.370 2076.920 54.650 2077.200 ;
        RECT 53.910 2070.120 54.190 2070.400 ;
        RECT 54.830 1353.400 55.110 1353.680 ;
        RECT 53.450 1352.720 53.730 1353.000 ;
        RECT 52.990 965.800 53.270 966.080 ;
        RECT 53.910 965.800 54.190 966.080 ;
        RECT 52.990 820.960 53.270 821.240 ;
        RECT 53.910 820.960 54.190 821.240 ;
        RECT 54.370 724.400 54.650 724.680 ;
        RECT 55.750 724.400 56.030 724.680 ;
        RECT 52.530 627.840 52.810 628.120 ;
        RECT 53.450 627.840 53.730 628.120 ;
        RECT 52.990 531.280 53.270 531.560 ;
        RECT 53.910 531.280 54.190 531.560 ;
        RECT 296.790 410.920 297.070 411.200 ;
      LAYER met3 ;
        RECT 52.965 2608.290 53.295 2608.305 ;
        RECT 53.885 2608.290 54.215 2608.305 ;
        RECT 52.965 2607.990 54.215 2608.290 ;
        RECT 52.965 2607.975 53.295 2607.990 ;
        RECT 53.885 2607.975 54.215 2607.990 ;
        RECT 52.965 2366.890 53.295 2366.905 ;
        RECT 53.885 2366.890 54.215 2366.905 ;
        RECT 52.965 2366.590 54.215 2366.890 ;
        RECT 52.965 2366.575 53.295 2366.590 ;
        RECT 53.885 2366.575 54.215 2366.590 ;
        RECT 53.630 2077.210 54.010 2077.220 ;
        RECT 54.345 2077.210 54.675 2077.225 ;
        RECT 53.630 2076.910 54.675 2077.210 ;
        RECT 53.630 2076.900 54.010 2076.910 ;
        RECT 54.345 2076.895 54.675 2076.910 ;
        RECT 53.885 2070.420 54.215 2070.425 ;
        RECT 53.630 2070.410 54.215 2070.420 ;
        RECT 53.630 2070.110 54.440 2070.410 ;
        RECT 53.630 2070.100 54.215 2070.110 ;
        RECT 53.885 2070.095 54.215 2070.100 ;
        RECT 54.805 1353.690 55.135 1353.705 ;
        RECT 52.750 1353.390 55.135 1353.690 ;
        RECT 52.750 1353.010 53.050 1353.390 ;
        RECT 54.805 1353.375 55.135 1353.390 ;
        RECT 53.425 1353.010 53.755 1353.025 ;
        RECT 52.750 1352.710 53.755 1353.010 ;
        RECT 53.425 1352.695 53.755 1352.710 ;
        RECT 52.965 966.090 53.295 966.105 ;
        RECT 53.885 966.090 54.215 966.105 ;
        RECT 52.965 965.790 54.215 966.090 ;
        RECT 52.965 965.775 53.295 965.790 ;
        RECT 53.885 965.775 54.215 965.790 ;
        RECT 52.965 821.250 53.295 821.265 ;
        RECT 53.885 821.250 54.215 821.265 ;
        RECT 52.965 820.950 54.215 821.250 ;
        RECT 52.965 820.935 53.295 820.950 ;
        RECT 53.885 820.935 54.215 820.950 ;
        RECT 54.345 724.690 54.675 724.705 ;
        RECT 55.725 724.690 56.055 724.705 ;
        RECT 54.345 724.390 56.055 724.690 ;
        RECT 54.345 724.375 54.675 724.390 ;
        RECT 55.725 724.375 56.055 724.390 ;
        RECT 52.505 628.130 52.835 628.145 ;
        RECT 53.425 628.130 53.755 628.145 ;
        RECT 52.505 627.830 53.755 628.130 ;
        RECT 52.505 627.815 52.835 627.830 ;
        RECT 53.425 627.815 53.755 627.830 ;
        RECT 52.965 531.570 53.295 531.585 ;
        RECT 53.885 531.570 54.215 531.585 ;
        RECT 52.965 531.270 54.215 531.570 ;
        RECT 52.965 531.255 53.295 531.270 ;
        RECT 53.885 531.255 54.215 531.270 ;
        RECT 296.765 411.210 297.095 411.225 ;
        RECT 310.000 411.210 314.000 411.600 ;
        RECT 296.765 411.000 314.000 411.210 ;
        RECT 296.765 410.910 310.500 411.000 ;
        RECT 296.765 410.895 297.095 410.910 ;
      LAYER via3 ;
        RECT 53.660 2076.900 53.980 2077.220 ;
        RECT 53.660 2070.100 53.980 2070.420 ;
      LAYER met4 ;
        RECT 53.655 2076.895 53.985 2077.225 ;
        RECT 53.670 2070.425 53.970 2076.895 ;
        RECT 53.655 2070.095 53.985 2070.425 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3305.380 17.410 3305.440 ;
        RECT 175.790 3305.380 176.110 3305.440 ;
        RECT 17.090 3305.240 176.110 3305.380 ;
        RECT 17.090 3305.180 17.410 3305.240 ;
        RECT 175.790 3305.180 176.110 3305.240 ;
        RECT 175.790 1407.500 176.110 1407.560 ;
        RECT 296.770 1407.500 297.090 1407.560 ;
        RECT 175.790 1407.360 297.090 1407.500 ;
        RECT 175.790 1407.300 176.110 1407.360 ;
        RECT 296.770 1407.300 297.090 1407.360 ;
      LAYER via ;
        RECT 17.120 3305.180 17.380 3305.440 ;
        RECT 175.820 3305.180 176.080 3305.440 ;
        RECT 175.820 1407.300 176.080 1407.560 ;
        RECT 296.800 1407.300 297.060 1407.560 ;
      LAYER met2 ;
        RECT 17.110 3309.715 17.390 3310.085 ;
        RECT 17.180 3305.470 17.320 3309.715 ;
        RECT 17.120 3305.150 17.380 3305.470 ;
        RECT 175.820 3305.150 176.080 3305.470 ;
        RECT 175.880 1407.590 176.020 3305.150 ;
        RECT 175.820 1407.270 176.080 1407.590 ;
        RECT 296.800 1407.270 297.060 1407.590 ;
        RECT 296.860 1405.405 297.000 1407.270 ;
        RECT 296.790 1405.035 297.070 1405.405 ;
      LAYER via2 ;
        RECT 17.110 3309.760 17.390 3310.040 ;
        RECT 296.790 1405.080 297.070 1405.360 ;
      LAYER met3 ;
        RECT -4.800 3310.050 2.400 3310.500 ;
        RECT 17.085 3310.050 17.415 3310.065 ;
        RECT -4.800 3309.750 17.415 3310.050 ;
        RECT -4.800 3309.300 2.400 3309.750 ;
        RECT 17.085 3309.735 17.415 3309.750 ;
        RECT 296.765 1405.370 297.095 1405.385 ;
        RECT 310.000 1405.370 314.000 1405.760 ;
        RECT 296.765 1405.160 314.000 1405.370 ;
        RECT 296.765 1405.070 310.500 1405.160 ;
        RECT 296.765 1405.055 297.095 1405.070 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 3056.840 16.950 3056.900 ;
        RECT 258.590 3056.840 258.910 3056.900 ;
        RECT 16.630 3056.700 258.910 3056.840 ;
        RECT 16.630 3056.640 16.950 3056.700 ;
        RECT 258.590 3056.640 258.910 3056.700 ;
        RECT 258.590 1013.920 258.910 1014.180 ;
        RECT 258.680 1013.500 258.820 1013.920 ;
        RECT 258.590 1013.240 258.910 1013.500 ;
        RECT 258.590 250.820 258.910 250.880 ;
        RECT 2228.310 250.820 2228.630 250.880 ;
        RECT 258.590 250.680 2228.630 250.820 ;
        RECT 258.590 250.620 258.910 250.680 ;
        RECT 2228.310 250.620 2228.630 250.680 ;
      LAYER via ;
        RECT 16.660 3056.640 16.920 3056.900 ;
        RECT 258.620 3056.640 258.880 3056.900 ;
        RECT 258.620 1013.920 258.880 1014.180 ;
        RECT 258.620 1013.240 258.880 1013.500 ;
        RECT 258.620 250.620 258.880 250.880 ;
        RECT 2228.340 250.620 2228.600 250.880 ;
      LAYER met2 ;
        RECT 16.650 3058.115 16.930 3058.485 ;
        RECT 16.720 3056.930 16.860 3058.115 ;
        RECT 16.660 3056.610 16.920 3056.930 ;
        RECT 258.620 3056.610 258.880 3056.930 ;
        RECT 258.680 1014.210 258.820 3056.610 ;
        RECT 258.620 1013.890 258.880 1014.210 ;
        RECT 258.620 1013.210 258.880 1013.530 ;
        RECT 258.680 250.910 258.820 1013.210 ;
        RECT 2228.290 260.000 2228.570 264.000 ;
        RECT 2228.400 250.910 2228.540 260.000 ;
        RECT 258.620 250.590 258.880 250.910 ;
        RECT 2228.340 250.590 2228.600 250.910 ;
      LAYER via2 ;
        RECT 16.650 3058.160 16.930 3058.440 ;
      LAYER met3 ;
        RECT -4.800 3058.450 2.400 3058.900 ;
        RECT 16.625 3058.450 16.955 3058.465 ;
        RECT -4.800 3058.150 16.955 3058.450 ;
        RECT -4.800 3057.700 2.400 3058.150 ;
        RECT 16.625 3058.135 16.955 3058.150 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2801.500 16.950 2801.560 ;
        RECT 51.590 2801.500 51.910 2801.560 ;
        RECT 16.630 2801.360 51.910 2801.500 ;
        RECT 16.630 2801.300 16.950 2801.360 ;
        RECT 51.590 2801.300 51.910 2801.360 ;
        RECT 51.590 239.940 51.910 240.000 ;
        RECT 1842.830 239.940 1843.150 240.000 ;
        RECT 51.590 239.800 1843.150 239.940 ;
        RECT 51.590 239.740 51.910 239.800 ;
        RECT 1842.830 239.740 1843.150 239.800 ;
      LAYER via ;
        RECT 16.660 2801.300 16.920 2801.560 ;
        RECT 51.620 2801.300 51.880 2801.560 ;
        RECT 51.620 239.740 51.880 240.000 ;
        RECT 1842.860 239.740 1843.120 240.000 ;
      LAYER met2 ;
        RECT 16.650 2806.515 16.930 2806.885 ;
        RECT 16.720 2801.590 16.860 2806.515 ;
        RECT 16.660 2801.270 16.920 2801.590 ;
        RECT 51.620 2801.270 51.880 2801.590 ;
        RECT 51.680 240.030 51.820 2801.270 ;
        RECT 1842.810 260.000 1843.090 264.000 ;
        RECT 1842.920 240.030 1843.060 260.000 ;
        RECT 51.620 239.710 51.880 240.030 ;
        RECT 1842.860 239.710 1843.120 240.030 ;
      LAYER via2 ;
        RECT 16.650 2806.560 16.930 2806.840 ;
      LAYER met3 ;
        RECT -4.800 2806.850 2.400 2807.300 ;
        RECT 16.625 2806.850 16.955 2806.865 ;
        RECT -4.800 2806.550 16.955 2806.850 ;
        RECT -4.800 2806.100 2.400 2806.550 ;
        RECT 16.625 2806.535 16.955 2806.550 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 230.990 3277.840 231.310 3277.900 ;
        RECT 2577.910 3277.840 2578.230 3277.900 ;
        RECT 230.990 3277.700 2578.230 3277.840 ;
        RECT 230.990 3277.640 231.310 3277.700 ;
        RECT 2577.910 3277.640 2578.230 3277.700 ;
        RECT 19.850 2559.760 20.170 2559.820 ;
        RECT 230.990 2559.760 231.310 2559.820 ;
        RECT 19.850 2559.620 231.310 2559.760 ;
        RECT 19.850 2559.560 20.170 2559.620 ;
        RECT 230.990 2559.560 231.310 2559.620 ;
      LAYER via ;
        RECT 231.020 3277.640 231.280 3277.900 ;
        RECT 2577.940 3277.640 2578.200 3277.900 ;
        RECT 19.880 2559.560 20.140 2559.820 ;
        RECT 231.020 2559.560 231.280 2559.820 ;
      LAYER met2 ;
        RECT 231.020 3277.610 231.280 3277.930 ;
        RECT 2577.940 3277.610 2578.200 3277.930 ;
        RECT 231.080 2559.850 231.220 3277.610 ;
        RECT 2578.000 3260.000 2578.140 3277.610 ;
        RECT 2577.890 3256.000 2578.170 3260.000 ;
        RECT 19.880 2559.530 20.140 2559.850 ;
        RECT 231.020 2559.530 231.280 2559.850 ;
        RECT 19.940 2555.965 20.080 2559.530 ;
        RECT 19.870 2555.595 20.150 2555.965 ;
      LAYER via2 ;
        RECT 19.870 2555.640 20.150 2555.920 ;
      LAYER met3 ;
        RECT -4.800 2555.930 2.400 2556.380 ;
        RECT 19.845 2555.930 20.175 2555.945 ;
        RECT -4.800 2555.630 20.175 2555.930 ;
        RECT -4.800 2555.180 2.400 2555.630 ;
        RECT 19.845 2555.615 20.175 2555.630 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2319.465 3252.865 2319.635 3256.435 ;
      LAYER mcon ;
        RECT 2319.465 3256.265 2319.635 3256.435 ;
      LAYER met1 ;
        RECT 2319.390 3256.420 2319.710 3256.480 ;
        RECT 2319.195 3256.280 2319.710 3256.420 ;
        RECT 2319.390 3256.220 2319.710 3256.280 ;
        RECT 265.950 3253.020 266.270 3253.080 ;
        RECT 2319.405 3253.020 2319.695 3253.065 ;
        RECT 265.950 3252.880 2319.695 3253.020 ;
        RECT 265.950 3252.820 266.270 3252.880 ;
        RECT 2319.405 3252.835 2319.695 3252.880 ;
        RECT 20.310 2304.420 20.630 2304.480 ;
        RECT 265.950 2304.420 266.270 2304.480 ;
        RECT 20.310 2304.280 266.270 2304.420 ;
        RECT 20.310 2304.220 20.630 2304.280 ;
        RECT 265.950 2304.220 266.270 2304.280 ;
      LAYER via ;
        RECT 2319.420 3256.220 2319.680 3256.480 ;
        RECT 265.980 3252.820 266.240 3253.080 ;
        RECT 20.340 2304.220 20.600 2304.480 ;
        RECT 265.980 2304.220 266.240 2304.480 ;
      LAYER met2 ;
        RECT 2321.210 3256.930 2321.490 3260.000 ;
        RECT 2319.480 3256.790 2321.490 3256.930 ;
        RECT 2319.480 3256.510 2319.620 3256.790 ;
        RECT 2319.420 3256.190 2319.680 3256.510 ;
        RECT 2321.210 3256.000 2321.490 3256.790 ;
        RECT 265.980 3252.790 266.240 3253.110 ;
        RECT 266.040 2304.510 266.180 3252.790 ;
        RECT 20.340 2304.365 20.600 2304.510 ;
        RECT 20.330 2303.995 20.610 2304.365 ;
        RECT 265.980 2304.190 266.240 2304.510 ;
      LAYER via2 ;
        RECT 20.330 2304.040 20.610 2304.320 ;
      LAYER met3 ;
        RECT -4.800 2304.330 2.400 2304.780 ;
        RECT 20.305 2304.330 20.635 2304.345 ;
        RECT -4.800 2304.030 20.635 2304.330 ;
        RECT -4.800 2303.580 2.400 2304.030 ;
        RECT 20.305 2304.015 20.635 2304.030 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 2049.420 19.710 2049.480 ;
        RECT 259.510 2049.420 259.830 2049.480 ;
        RECT 19.390 2049.280 259.830 2049.420 ;
        RECT 19.390 2049.220 19.710 2049.280 ;
        RECT 259.510 2049.220 259.830 2049.280 ;
      LAYER via ;
        RECT 19.420 2049.220 19.680 2049.480 ;
        RECT 259.540 2049.220 259.800 2049.480 ;
      LAYER met2 ;
        RECT 19.410 2052.395 19.690 2052.765 ;
        RECT 19.480 2049.510 19.620 2052.395 ;
        RECT 19.420 2049.190 19.680 2049.510 ;
        RECT 259.540 2049.190 259.800 2049.510 ;
        RECT 259.600 1014.405 259.740 2049.190 ;
        RECT 259.530 1014.035 259.810 1014.405 ;
        RECT 259.530 1011.315 259.810 1011.685 ;
        RECT 259.600 262.325 259.740 1011.315 ;
        RECT 2607.830 272.155 2608.110 272.525 ;
        RECT 2607.900 262.325 2608.040 272.155 ;
        RECT 259.530 261.955 259.810 262.325 ;
        RECT 2607.830 261.955 2608.110 262.325 ;
      LAYER via2 ;
        RECT 19.410 2052.440 19.690 2052.720 ;
        RECT 259.530 1014.080 259.810 1014.360 ;
        RECT 259.530 1011.360 259.810 1011.640 ;
        RECT 2607.830 272.200 2608.110 272.480 ;
        RECT 259.530 262.000 259.810 262.280 ;
        RECT 2607.830 262.000 2608.110 262.280 ;
      LAYER met3 ;
        RECT -4.800 2052.730 2.400 2053.180 ;
        RECT 19.385 2052.730 19.715 2052.745 ;
        RECT -4.800 2052.430 19.715 2052.730 ;
        RECT -4.800 2051.980 2.400 2052.430 ;
        RECT 19.385 2052.415 19.715 2052.430 ;
        RECT 259.505 1014.370 259.835 1014.385 ;
        RECT 259.505 1014.055 260.050 1014.370 ;
        RECT 259.750 1011.665 260.050 1014.055 ;
        RECT 259.505 1011.350 260.050 1011.665 ;
        RECT 259.505 1011.335 259.835 1011.350 ;
        RECT 2606.000 275.000 2610.000 275.600 ;
        RECT 2607.590 272.505 2607.890 275.000 ;
        RECT 2607.590 272.190 2608.135 272.505 ;
        RECT 2607.805 272.175 2608.135 272.190 ;
        RECT 259.505 262.290 259.835 262.305 ;
        RECT 2607.805 262.290 2608.135 262.305 ;
        RECT 259.505 261.990 2608.135 262.290 ;
        RECT 259.505 261.975 259.835 261.990 ;
        RECT 2607.805 261.975 2608.135 261.990 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2728.790 669.360 2729.110 669.420 ;
        RECT 2900.830 669.360 2901.150 669.420 ;
        RECT 2728.790 669.220 2901.150 669.360 ;
        RECT 2728.790 669.160 2729.110 669.220 ;
        RECT 2900.830 669.160 2901.150 669.220 ;
      LAYER via ;
        RECT 2728.820 669.160 2729.080 669.420 ;
        RECT 2900.860 669.160 2901.120 669.420 ;
      LAYER met2 ;
        RECT 1449.090 3265.515 1449.370 3265.885 ;
        RECT 2728.810 3265.515 2729.090 3265.885 ;
        RECT 1449.160 3260.000 1449.300 3265.515 ;
        RECT 1449.050 3256.000 1449.330 3260.000 ;
        RECT 2728.880 669.450 2729.020 3265.515 ;
        RECT 2728.820 669.130 2729.080 669.450 ;
        RECT 2900.860 669.130 2901.120 669.450 ;
        RECT 2900.920 664.885 2901.060 669.130 ;
        RECT 2900.850 664.515 2901.130 664.885 ;
      LAYER via2 ;
        RECT 1449.090 3265.560 1449.370 3265.840 ;
        RECT 2728.810 3265.560 2729.090 3265.840 ;
        RECT 2900.850 664.560 2901.130 664.840 ;
      LAYER met3 ;
        RECT 1449.065 3265.850 1449.395 3265.865 ;
        RECT 2728.785 3265.850 2729.115 3265.865 ;
        RECT 1449.065 3265.550 2729.115 3265.850 ;
        RECT 1449.065 3265.535 1449.395 3265.550 ;
        RECT 2728.785 3265.535 2729.115 3265.550 ;
        RECT 2900.825 664.850 2901.155 664.865 ;
        RECT 2917.600 664.850 2924.800 665.300 ;
        RECT 2900.825 664.550 2924.800 664.850 ;
        RECT 2900.825 664.535 2901.155 664.550 ;
        RECT 2917.600 664.100 2924.800 664.550 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 1801.220 20.630 1801.280 ;
        RECT 65.850 1801.220 66.170 1801.280 ;
        RECT 20.310 1801.080 66.170 1801.220 ;
        RECT 20.310 1801.020 20.630 1801.080 ;
        RECT 65.850 1801.020 66.170 1801.080 ;
        RECT 65.850 1345.280 66.170 1345.340 ;
        RECT 296.770 1345.280 297.090 1345.340 ;
        RECT 65.850 1345.140 297.090 1345.280 ;
        RECT 65.850 1345.080 66.170 1345.140 ;
        RECT 296.770 1345.080 297.090 1345.140 ;
      LAYER via ;
        RECT 20.340 1801.020 20.600 1801.280 ;
        RECT 65.880 1801.020 66.140 1801.280 ;
        RECT 65.880 1345.080 66.140 1345.340 ;
        RECT 296.800 1345.080 297.060 1345.340 ;
      LAYER met2 ;
        RECT 20.330 1801.475 20.610 1801.845 ;
        RECT 20.400 1801.310 20.540 1801.475 ;
        RECT 20.340 1800.990 20.600 1801.310 ;
        RECT 65.880 1800.990 66.140 1801.310 ;
        RECT 65.940 1345.370 66.080 1800.990 ;
        RECT 65.880 1345.050 66.140 1345.370 ;
        RECT 296.800 1345.050 297.060 1345.370 ;
        RECT 296.860 1341.485 297.000 1345.050 ;
        RECT 296.790 1341.115 297.070 1341.485 ;
      LAYER via2 ;
        RECT 20.330 1801.520 20.610 1801.800 ;
        RECT 296.790 1341.160 297.070 1341.440 ;
      LAYER met3 ;
        RECT -4.800 1801.810 2.400 1802.260 ;
        RECT 20.305 1801.810 20.635 1801.825 ;
        RECT -4.800 1801.510 20.635 1801.810 ;
        RECT -4.800 1801.060 2.400 1801.510 ;
        RECT 20.305 1801.495 20.635 1801.510 ;
        RECT 296.765 1341.450 297.095 1341.465 ;
        RECT 310.000 1341.450 314.000 1341.840 ;
        RECT 296.765 1341.240 314.000 1341.450 ;
        RECT 296.765 1341.150 310.500 1341.240 ;
        RECT 296.765 1341.135 297.095 1341.150 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1548.260 16.030 1548.320 ;
        RECT 44.690 1548.260 45.010 1548.320 ;
        RECT 15.710 1548.120 45.010 1548.260 ;
        RECT 15.710 1548.060 16.030 1548.120 ;
        RECT 44.690 1548.060 45.010 1548.120 ;
        RECT 44.690 254.220 45.010 254.280 ;
        RECT 1699.310 254.220 1699.630 254.280 ;
        RECT 44.690 254.080 1699.630 254.220 ;
        RECT 44.690 254.020 45.010 254.080 ;
        RECT 1699.310 254.020 1699.630 254.080 ;
      LAYER via ;
        RECT 15.740 1548.060 16.000 1548.320 ;
        RECT 44.720 1548.060 44.980 1548.320 ;
        RECT 44.720 254.020 44.980 254.280 ;
        RECT 1699.340 254.020 1699.600 254.280 ;
      LAYER met2 ;
        RECT 15.730 1549.875 16.010 1550.245 ;
        RECT 15.800 1548.350 15.940 1549.875 ;
        RECT 15.740 1548.030 16.000 1548.350 ;
        RECT 44.720 1548.030 44.980 1548.350 ;
        RECT 44.780 254.310 44.920 1548.030 ;
        RECT 1699.290 260.000 1699.570 264.000 ;
        RECT 1699.400 254.310 1699.540 260.000 ;
        RECT 44.720 253.990 44.980 254.310 ;
        RECT 1699.340 253.990 1699.600 254.310 ;
      LAYER via2 ;
        RECT 15.730 1549.920 16.010 1550.200 ;
      LAYER met3 ;
        RECT -4.800 1550.210 2.400 1550.660 ;
        RECT 15.705 1550.210 16.035 1550.225 ;
        RECT -4.800 1549.910 16.035 1550.210 ;
        RECT -4.800 1549.460 2.400 1549.910 ;
        RECT 15.705 1549.895 16.035 1549.910 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 53.045 1303.985 54.135 1304.155 ;
      LAYER mcon ;
        RECT 53.965 1303.985 54.135 1304.155 ;
      LAYER met1 ;
        RECT 230.530 3261.520 230.850 3261.580 ;
        RECT 319.310 3261.520 319.630 3261.580 ;
        RECT 230.530 3261.380 319.630 3261.520 ;
        RECT 230.530 3261.320 230.850 3261.380 ;
        RECT 319.310 3261.320 319.630 3261.380 ;
        RECT 16.630 1304.140 16.950 1304.200 ;
        RECT 52.985 1304.140 53.275 1304.185 ;
        RECT 16.630 1304.000 53.275 1304.140 ;
        RECT 16.630 1303.940 16.950 1304.000 ;
        RECT 52.985 1303.955 53.275 1304.000 ;
        RECT 53.905 1304.140 54.195 1304.185 ;
        RECT 230.530 1304.140 230.850 1304.200 ;
        RECT 53.905 1304.000 230.850 1304.140 ;
        RECT 53.905 1303.955 54.195 1304.000 ;
        RECT 230.530 1303.940 230.850 1304.000 ;
      LAYER via ;
        RECT 230.560 3261.320 230.820 3261.580 ;
        RECT 319.340 3261.320 319.600 3261.580 ;
        RECT 16.660 1303.940 16.920 1304.200 ;
        RECT 230.560 1303.940 230.820 1304.200 ;
      LAYER met2 ;
        RECT 230.560 3261.290 230.820 3261.610 ;
        RECT 319.340 3261.290 319.600 3261.610 ;
        RECT 230.620 1304.230 230.760 3261.290 ;
        RECT 319.400 3260.000 319.540 3261.290 ;
        RECT 319.290 3256.000 319.570 3260.000 ;
        RECT 16.660 1303.910 16.920 1304.230 ;
        RECT 230.560 1303.910 230.820 1304.230 ;
        RECT 16.720 1298.645 16.860 1303.910 ;
        RECT 230.620 1303.615 230.760 1303.910 ;
        RECT 16.650 1298.275 16.930 1298.645 ;
      LAYER via2 ;
        RECT 16.650 1298.320 16.930 1298.600 ;
      LAYER met3 ;
        RECT -4.800 1298.610 2.400 1299.060 ;
        RECT 16.625 1298.610 16.955 1298.625 ;
        RECT -4.800 1298.310 16.955 1298.610 ;
        RECT -4.800 1297.860 2.400 1298.310 ;
        RECT 16.625 1298.295 16.955 1298.310 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 265.490 2946.680 265.810 2946.740 ;
        RECT 296.770 2946.680 297.090 2946.740 ;
        RECT 265.490 2946.540 297.090 2946.680 ;
        RECT 265.490 2946.480 265.810 2946.540 ;
        RECT 296.770 2946.480 297.090 2946.540 ;
        RECT 19.850 1052.200 20.170 1052.260 ;
        RECT 265.490 1052.200 265.810 1052.260 ;
        RECT 19.850 1052.060 265.810 1052.200 ;
        RECT 19.850 1052.000 20.170 1052.060 ;
        RECT 265.490 1052.000 265.810 1052.060 ;
      LAYER via ;
        RECT 265.520 2946.480 265.780 2946.740 ;
        RECT 296.800 2946.480 297.060 2946.740 ;
        RECT 19.880 1052.000 20.140 1052.260 ;
        RECT 265.520 1052.000 265.780 1052.260 ;
      LAYER met2 ;
        RECT 296.790 2947.275 297.070 2947.645 ;
        RECT 296.860 2946.770 297.000 2947.275 ;
        RECT 265.520 2946.450 265.780 2946.770 ;
        RECT 296.800 2946.450 297.060 2946.770 ;
        RECT 265.580 1052.290 265.720 2946.450 ;
        RECT 19.880 1051.970 20.140 1052.290 ;
        RECT 265.520 1051.970 265.780 1052.290 ;
        RECT 19.940 1047.045 20.080 1051.970 ;
        RECT 19.870 1046.675 20.150 1047.045 ;
      LAYER via2 ;
        RECT 296.790 2947.320 297.070 2947.600 ;
        RECT 19.870 1046.720 20.150 1047.000 ;
      LAYER met3 ;
        RECT 296.765 2947.610 297.095 2947.625 ;
        RECT 310.000 2947.610 314.000 2948.000 ;
        RECT 296.765 2947.400 314.000 2947.610 ;
        RECT 296.765 2947.310 310.500 2947.400 ;
        RECT 296.765 2947.295 297.095 2947.310 ;
        RECT -4.800 1047.010 2.400 1047.460 ;
        RECT 19.845 1047.010 20.175 1047.025 ;
        RECT -4.800 1046.710 20.175 1047.010 ;
        RECT -4.800 1046.260 2.400 1046.710 ;
        RECT 19.845 1046.695 20.175 1046.710 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 793.800 20.630 793.860 ;
        RECT 265.490 793.800 265.810 793.860 ;
        RECT 20.310 793.660 265.810 793.800 ;
        RECT 20.310 793.600 20.630 793.660 ;
        RECT 265.490 793.600 265.810 793.660 ;
        RECT 265.490 255.240 265.810 255.300 ;
        RECT 698.350 255.240 698.670 255.300 ;
        RECT 265.490 255.100 698.670 255.240 ;
        RECT 265.490 255.040 265.810 255.100 ;
        RECT 698.350 255.040 698.670 255.100 ;
      LAYER via ;
        RECT 20.340 793.600 20.600 793.860 ;
        RECT 265.520 793.600 265.780 793.860 ;
        RECT 265.520 255.040 265.780 255.300 ;
        RECT 698.380 255.040 698.640 255.300 ;
      LAYER met2 ;
        RECT 20.330 795.755 20.610 796.125 ;
        RECT 20.400 793.890 20.540 795.755 ;
        RECT 20.340 793.570 20.600 793.890 ;
        RECT 265.520 793.570 265.780 793.890 ;
        RECT 265.580 255.330 265.720 793.570 ;
        RECT 698.330 260.000 698.610 264.000 ;
        RECT 698.440 255.330 698.580 260.000 ;
        RECT 265.520 255.010 265.780 255.330 ;
        RECT 698.380 255.010 698.640 255.330 ;
      LAYER via2 ;
        RECT 20.330 795.800 20.610 796.080 ;
      LAYER met3 ;
        RECT -4.800 796.090 2.400 796.540 ;
        RECT 20.305 796.090 20.635 796.105 ;
        RECT -4.800 795.790 20.635 796.090 ;
        RECT -4.800 795.340 2.400 795.790 ;
        RECT 20.305 795.775 20.635 795.790 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 86.090 1511.200 86.410 1511.260 ;
        RECT 296.770 1511.200 297.090 1511.260 ;
        RECT 86.090 1511.060 297.090 1511.200 ;
        RECT 86.090 1511.000 86.410 1511.060 ;
        RECT 296.770 1511.000 297.090 1511.060 ;
        RECT 20.310 544.920 20.630 544.980 ;
        RECT 86.090 544.920 86.410 544.980 ;
        RECT 20.310 544.780 86.410 544.920 ;
        RECT 20.310 544.720 20.630 544.780 ;
        RECT 86.090 544.720 86.410 544.780 ;
      LAYER via ;
        RECT 86.120 1511.000 86.380 1511.260 ;
        RECT 296.800 1511.000 297.060 1511.260 ;
        RECT 20.340 544.720 20.600 544.980 ;
        RECT 86.120 544.720 86.380 544.980 ;
      LAYER met2 ;
        RECT 86.120 1510.970 86.380 1511.290 ;
        RECT 296.790 1511.115 297.070 1511.485 ;
        RECT 296.800 1510.970 297.060 1511.115 ;
        RECT 86.180 545.010 86.320 1510.970 ;
        RECT 20.340 544.690 20.600 545.010 ;
        RECT 86.120 544.690 86.380 545.010 ;
        RECT 20.400 544.525 20.540 544.690 ;
        RECT 20.330 544.155 20.610 544.525 ;
      LAYER via2 ;
        RECT 296.790 1511.160 297.070 1511.440 ;
        RECT 20.330 544.200 20.610 544.480 ;
      LAYER met3 ;
        RECT 296.765 1511.450 297.095 1511.465 ;
        RECT 310.000 1511.450 314.000 1511.840 ;
        RECT 296.765 1511.240 314.000 1511.450 ;
        RECT 296.765 1511.150 310.500 1511.240 ;
        RECT 296.765 1511.135 297.095 1511.150 ;
        RECT -4.800 544.490 2.400 544.940 ;
        RECT 20.305 544.490 20.635 544.505 ;
        RECT -4.800 544.190 20.635 544.490 ;
        RECT -4.800 543.740 2.400 544.190 ;
        RECT 20.305 544.175 20.635 544.190 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 120.590 3091.520 120.910 3091.580 ;
        RECT 296.770 3091.520 297.090 3091.580 ;
        RECT 120.590 3091.380 297.090 3091.520 ;
        RECT 120.590 3091.320 120.910 3091.380 ;
        RECT 296.770 3091.320 297.090 3091.380 ;
        RECT 15.250 296.720 15.570 296.780 ;
        RECT 120.590 296.720 120.910 296.780 ;
        RECT 15.250 296.580 120.910 296.720 ;
        RECT 15.250 296.520 15.570 296.580 ;
        RECT 120.590 296.520 120.910 296.580 ;
      LAYER via ;
        RECT 120.620 3091.320 120.880 3091.580 ;
        RECT 296.800 3091.320 297.060 3091.580 ;
        RECT 15.280 296.520 15.540 296.780 ;
        RECT 120.620 296.520 120.880 296.780 ;
      LAYER met2 ;
        RECT 296.790 3095.515 297.070 3095.885 ;
        RECT 296.860 3091.610 297.000 3095.515 ;
        RECT 120.620 3091.290 120.880 3091.610 ;
        RECT 296.800 3091.290 297.060 3091.610 ;
        RECT 120.680 296.810 120.820 3091.290 ;
        RECT 15.280 296.490 15.540 296.810 ;
        RECT 120.620 296.490 120.880 296.810 ;
        RECT 15.340 292.925 15.480 296.490 ;
        RECT 15.270 292.555 15.550 292.925 ;
      LAYER via2 ;
        RECT 296.790 3095.560 297.070 3095.840 ;
        RECT 15.270 292.600 15.550 292.880 ;
      LAYER met3 ;
        RECT 296.765 3095.850 297.095 3095.865 ;
        RECT 310.000 3095.850 314.000 3096.240 ;
        RECT 296.765 3095.640 314.000 3095.850 ;
        RECT 296.765 3095.550 310.500 3095.640 ;
        RECT 296.765 3095.535 297.095 3095.550 ;
        RECT -4.800 292.890 2.400 293.340 ;
        RECT 15.245 292.890 15.575 292.905 ;
        RECT -4.800 292.590 15.575 292.890 ;
        RECT -4.800 292.140 2.400 292.590 ;
        RECT 15.245 292.575 15.575 292.590 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2657.510 2124.475 2657.790 2124.845 ;
        RECT 2657.580 2101.045 2657.720 2124.475 ;
        RECT 2657.510 2100.675 2657.790 2101.045 ;
        RECT 2657.510 1641.675 2657.790 1642.045 ;
        RECT 2657.580 1640.005 2657.720 1641.675 ;
        RECT 2657.510 1639.635 2657.790 1640.005 ;
        RECT 17.110 47.755 17.390 48.125 ;
        RECT 17.180 42.005 17.320 47.755 ;
        RECT 17.110 41.635 17.390 42.005 ;
      LAYER via2 ;
        RECT 2657.510 2124.520 2657.790 2124.800 ;
        RECT 2657.510 2100.720 2657.790 2101.000 ;
        RECT 2657.510 1641.720 2657.790 1642.000 ;
        RECT 2657.510 1639.680 2657.790 1639.960 ;
        RECT 17.110 47.800 17.390 48.080 ;
        RECT 17.110 41.680 17.390 41.960 ;
      LAYER met3 ;
        RECT 2606.000 2198.040 2610.000 2198.640 ;
        RECT 2609.430 2194.850 2609.730 2198.040 ;
        RECT 2657.230 2194.850 2657.610 2194.860 ;
        RECT 2609.430 2194.550 2657.610 2194.850 ;
        RECT 2657.230 2194.540 2657.610 2194.550 ;
        RECT 2657.485 2124.820 2657.815 2124.825 ;
        RECT 2657.230 2124.810 2657.815 2124.820 ;
        RECT 2657.230 2124.510 2658.040 2124.810 ;
        RECT 2657.230 2124.500 2657.815 2124.510 ;
        RECT 2657.485 2124.495 2657.815 2124.500 ;
        RECT 2657.485 2101.020 2657.815 2101.025 ;
        RECT 2657.230 2101.010 2657.815 2101.020 ;
        RECT 2657.030 2100.710 2657.815 2101.010 ;
        RECT 2657.230 2100.700 2657.815 2100.710 ;
        RECT 2657.485 2100.695 2657.815 2100.700 ;
        RECT 2657.485 1642.020 2657.815 1642.025 ;
        RECT 2657.230 1642.010 2657.815 1642.020 ;
        RECT 2657.230 1641.710 2658.040 1642.010 ;
        RECT 2657.230 1641.700 2657.815 1641.710 ;
        RECT 2657.485 1641.695 2657.815 1641.700 ;
        RECT 2657.485 1639.970 2657.815 1639.985 ;
        RECT 2658.150 1639.970 2658.530 1639.980 ;
        RECT 2657.485 1639.670 2658.530 1639.970 ;
        RECT 2657.485 1639.655 2657.815 1639.670 ;
        RECT 2658.150 1639.660 2658.530 1639.670 ;
        RECT 17.085 48.090 17.415 48.105 ;
        RECT 2657.230 48.090 2657.610 48.100 ;
        RECT 17.085 47.790 2657.610 48.090 ;
        RECT 17.085 47.775 17.415 47.790 ;
        RECT 2657.230 47.780 2657.610 47.790 ;
        RECT -4.800 41.970 2.400 42.420 ;
        RECT 17.085 41.970 17.415 41.985 ;
        RECT -4.800 41.670 17.415 41.970 ;
        RECT -4.800 41.220 2.400 41.670 ;
        RECT 17.085 41.655 17.415 41.670 ;
      LAYER via3 ;
        RECT 2657.260 2194.540 2657.580 2194.860 ;
        RECT 2657.260 2124.500 2657.580 2124.820 ;
        RECT 2657.260 2100.700 2657.580 2101.020 ;
        RECT 2657.260 1641.700 2657.580 1642.020 ;
        RECT 2658.180 1639.660 2658.500 1639.980 ;
        RECT 2657.260 47.780 2657.580 48.100 ;
      LAYER met4 ;
        RECT 2657.255 2194.535 2657.585 2194.865 ;
        RECT 2657.270 2124.825 2657.570 2194.535 ;
        RECT 2657.255 2124.495 2657.585 2124.825 ;
        RECT 2657.255 2100.695 2657.585 2101.025 ;
        RECT 2657.270 1642.025 2657.570 2100.695 ;
        RECT 2657.255 1641.695 2657.585 1642.025 ;
        RECT 2658.175 1639.655 2658.505 1639.985 ;
        RECT 2658.190 1616.850 2658.490 1639.655 ;
        RECT 2657.270 1616.550 2658.490 1616.850 ;
        RECT 2657.270 48.105 2657.570 1616.550 ;
        RECT 2657.255 47.775 2657.585 48.105 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2901.770 899.115 2902.050 899.485 ;
        RECT 2901.840 813.805 2901.980 899.115 ;
        RECT 2901.770 813.435 2902.050 813.805 ;
      LAYER via2 ;
        RECT 2901.770 899.160 2902.050 899.440 ;
        RECT 2901.770 813.480 2902.050 813.760 ;
      LAYER met3 ;
        RECT 2901.745 899.450 2902.075 899.465 ;
        RECT 2917.600 899.450 2924.800 899.900 ;
        RECT 2901.745 899.150 2924.800 899.450 ;
        RECT 2901.745 899.135 2902.075 899.150 ;
        RECT 2917.600 898.700 2924.800 899.150 ;
        RECT 310.000 813.560 314.000 814.160 ;
        RECT 2626.870 813.770 2627.250 813.780 ;
        RECT 2901.745 813.770 2902.075 813.785 ;
        RECT 309.390 811.050 309.770 811.060 ;
        RECT 310.350 811.050 310.650 813.560 ;
        RECT 2626.870 813.470 2902.075 813.770 ;
        RECT 2626.870 813.460 2627.250 813.470 ;
        RECT 2901.745 813.455 2902.075 813.470 ;
        RECT 309.390 810.750 310.650 811.050 ;
        RECT 309.390 810.740 309.770 810.750 ;
      LAYER via3 ;
        RECT 309.420 810.740 309.740 811.060 ;
        RECT 2626.900 813.460 2627.220 813.780 ;
      LAYER met4 ;
        RECT 2626.895 813.455 2627.225 813.785 ;
        RECT 2626.910 811.490 2627.210 813.455 ;
        RECT 308.990 810.310 310.170 811.490 ;
        RECT 2626.470 810.310 2627.650 811.490 ;
      LAYER met5 ;
        RECT 348.340 813.500 404.220 815.100 ;
        RECT 348.340 811.700 349.940 813.500 ;
        RECT 308.780 810.100 349.940 811.700 ;
        RECT 402.620 798.100 404.220 813.500 ;
        RECT 414.580 813.500 485.180 815.100 ;
        RECT 414.580 798.100 416.180 813.500 ;
        RECT 483.580 811.700 485.180 813.500 ;
        RECT 482.660 810.100 485.180 811.700 ;
        RECT 543.380 813.500 581.780 815.100 ;
        RECT 482.660 801.500 484.260 810.100 ;
        RECT 543.380 808.300 544.980 813.500 ;
        RECT 580.180 811.700 581.780 813.500 ;
        RECT 529.580 806.700 544.980 808.300 ;
        RECT 579.260 810.100 581.780 811.700 ;
        RECT 639.980 813.500 678.380 815.100 ;
        RECT 529.580 801.500 531.180 806.700 ;
        RECT 482.660 799.900 531.180 801.500 ;
        RECT 579.260 801.500 580.860 810.100 ;
        RECT 639.980 808.300 641.580 813.500 ;
        RECT 676.780 811.700 678.380 813.500 ;
        RECT 626.180 806.700 641.580 808.300 ;
        RECT 675.860 810.100 678.380 811.700 ;
        RECT 736.580 813.500 786.940 815.100 ;
        RECT 626.180 801.500 627.780 806.700 ;
        RECT 579.260 799.900 627.780 801.500 ;
        RECT 675.860 801.500 677.460 810.100 ;
        RECT 736.580 808.300 738.180 813.500 ;
        RECT 722.780 806.700 738.180 808.300 ;
        RECT 785.340 808.300 786.940 813.500 ;
        RECT 806.500 813.500 855.940 815.100 ;
        RECT 806.500 808.300 808.100 813.500 ;
        RECT 785.340 806.700 808.100 808.300 ;
        RECT 854.340 808.300 855.940 813.500 ;
        RECT 903.100 813.500 952.540 815.100 ;
        RECT 903.100 808.300 904.700 813.500 ;
        RECT 854.340 806.700 904.700 808.300 ;
        RECT 950.940 808.300 952.540 813.500 ;
        RECT 999.700 813.500 1049.140 815.100 ;
        RECT 999.700 808.300 1001.300 813.500 ;
        RECT 950.940 806.700 1001.300 808.300 ;
        RECT 1047.540 808.300 1049.140 813.500 ;
        RECT 1096.300 813.500 1145.740 815.100 ;
        RECT 1096.300 808.300 1097.900 813.500 ;
        RECT 1047.540 806.700 1097.900 808.300 ;
        RECT 1144.140 808.300 1145.740 813.500 ;
        RECT 1192.900 813.500 1242.340 815.100 ;
        RECT 1192.900 808.300 1194.500 813.500 ;
        RECT 1144.140 806.700 1194.500 808.300 ;
        RECT 1240.740 808.300 1242.340 813.500 ;
        RECT 1289.500 813.500 1338.940 815.100 ;
        RECT 1289.500 808.300 1291.100 813.500 ;
        RECT 1240.740 806.700 1291.100 808.300 ;
        RECT 1337.340 808.300 1338.940 813.500 ;
        RECT 1386.100 813.500 1435.540 815.100 ;
        RECT 1386.100 808.300 1387.700 813.500 ;
        RECT 1337.340 806.700 1387.700 808.300 ;
        RECT 1433.940 808.300 1435.540 813.500 ;
        RECT 1482.700 813.500 1532.140 815.100 ;
        RECT 1482.700 808.300 1484.300 813.500 ;
        RECT 1433.940 806.700 1484.300 808.300 ;
        RECT 1530.540 808.300 1532.140 813.500 ;
        RECT 1579.300 813.500 1628.740 815.100 ;
        RECT 1579.300 808.300 1580.900 813.500 ;
        RECT 1530.540 806.700 1580.900 808.300 ;
        RECT 1627.140 808.300 1628.740 813.500 ;
        RECT 1675.900 813.500 1725.340 815.100 ;
        RECT 1675.900 808.300 1677.500 813.500 ;
        RECT 1627.140 806.700 1677.500 808.300 ;
        RECT 1723.740 808.300 1725.340 813.500 ;
        RECT 1772.500 813.500 1821.940 815.100 ;
        RECT 1772.500 808.300 1774.100 813.500 ;
        RECT 1723.740 806.700 1774.100 808.300 ;
        RECT 1820.340 808.300 1821.940 813.500 ;
        RECT 1869.100 813.500 1918.540 815.100 ;
        RECT 1869.100 808.300 1870.700 813.500 ;
        RECT 1820.340 806.700 1870.700 808.300 ;
        RECT 1916.940 808.300 1918.540 813.500 ;
        RECT 1965.700 813.500 2015.140 815.100 ;
        RECT 1965.700 808.300 1967.300 813.500 ;
        RECT 1916.940 806.700 1967.300 808.300 ;
        RECT 2013.540 808.300 2015.140 813.500 ;
        RECT 2062.300 813.500 2111.740 815.100 ;
        RECT 2062.300 808.300 2063.900 813.500 ;
        RECT 2013.540 806.700 2063.900 808.300 ;
        RECT 2110.140 808.300 2111.740 813.500 ;
        RECT 2158.900 813.500 2208.340 815.100 ;
        RECT 2158.900 808.300 2160.500 813.500 ;
        RECT 2110.140 806.700 2160.500 808.300 ;
        RECT 2206.740 808.300 2208.340 813.500 ;
        RECT 2255.500 813.500 2304.940 815.100 ;
        RECT 2255.500 808.300 2257.100 813.500 ;
        RECT 2206.740 806.700 2257.100 808.300 ;
        RECT 2303.340 808.300 2304.940 813.500 ;
        RECT 2352.100 813.500 2401.540 815.100 ;
        RECT 2352.100 808.300 2353.700 813.500 ;
        RECT 2303.340 806.700 2353.700 808.300 ;
        RECT 2399.940 808.300 2401.540 813.500 ;
        RECT 2448.700 813.500 2525.740 815.100 ;
        RECT 2448.700 808.300 2450.300 813.500 ;
        RECT 2399.940 806.700 2450.300 808.300 ;
        RECT 2524.140 808.300 2525.740 813.500 ;
        RECT 2545.300 813.500 2574.500 815.100 ;
        RECT 2545.300 808.300 2546.900 813.500 ;
        RECT 2572.900 811.700 2574.500 813.500 ;
        RECT 2572.900 810.100 2627.860 811.700 ;
        RECT 2524.140 806.700 2546.900 808.300 ;
        RECT 722.780 801.500 724.380 806.700 ;
        RECT 675.860 799.900 724.380 801.500 ;
        RECT 402.620 796.500 416.180 798.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2435.310 3267.980 2435.630 3268.040 ;
        RECT 2694.290 3267.980 2694.610 3268.040 ;
        RECT 2435.310 3267.840 2694.610 3267.980 ;
        RECT 2435.310 3267.780 2435.630 3267.840 ;
        RECT 2694.290 3267.780 2694.610 3267.840 ;
        RECT 2694.290 1138.560 2694.610 1138.620 ;
        RECT 2900.830 1138.560 2901.150 1138.620 ;
        RECT 2694.290 1138.420 2901.150 1138.560 ;
        RECT 2694.290 1138.360 2694.610 1138.420 ;
        RECT 2900.830 1138.360 2901.150 1138.420 ;
      LAYER via ;
        RECT 2435.340 3267.780 2435.600 3268.040 ;
        RECT 2694.320 3267.780 2694.580 3268.040 ;
        RECT 2694.320 1138.360 2694.580 1138.620 ;
        RECT 2900.860 1138.360 2901.120 1138.620 ;
      LAYER met2 ;
        RECT 2435.340 3267.750 2435.600 3268.070 ;
        RECT 2694.320 3267.750 2694.580 3268.070 ;
        RECT 2435.400 3260.000 2435.540 3267.750 ;
        RECT 2435.290 3256.000 2435.570 3260.000 ;
        RECT 2694.380 1138.650 2694.520 3267.750 ;
        RECT 2694.320 1138.330 2694.580 1138.650 ;
        RECT 2900.860 1138.330 2901.120 1138.650 ;
        RECT 2900.920 1134.085 2901.060 1138.330 ;
        RECT 2900.850 1133.715 2901.130 1134.085 ;
      LAYER via2 ;
        RECT 2900.850 1133.760 2901.130 1134.040 ;
      LAYER met3 ;
        RECT 2900.825 1134.050 2901.155 1134.065 ;
        RECT 2917.600 1134.050 2924.800 1134.500 ;
        RECT 2900.825 1133.750 2924.800 1134.050 ;
        RECT 2900.825 1133.735 2901.155 1133.750 ;
        RECT 2917.600 1133.300 2924.800 1133.750 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 861.725 3253.205 861.895 3256.435 ;
      LAYER mcon ;
        RECT 861.725 3256.265 861.895 3256.435 ;
      LAYER met1 ;
        RECT 861.650 3256.420 861.970 3256.480 ;
        RECT 861.455 3256.280 861.970 3256.420 ;
        RECT 861.650 3256.220 861.970 3256.280 ;
        RECT 861.665 3253.360 861.955 3253.405 ;
        RECT 2763.290 3253.360 2763.610 3253.420 ;
        RECT 861.665 3253.220 2763.610 3253.360 ;
        RECT 861.665 3253.175 861.955 3253.220 ;
        RECT 2763.290 3253.160 2763.610 3253.220 ;
        RECT 2763.290 1373.160 2763.610 1373.220 ;
        RECT 2900.830 1373.160 2901.150 1373.220 ;
        RECT 2763.290 1373.020 2901.150 1373.160 ;
        RECT 2763.290 1372.960 2763.610 1373.020 ;
        RECT 2900.830 1372.960 2901.150 1373.020 ;
      LAYER via ;
        RECT 861.680 3256.220 861.940 3256.480 ;
        RECT 2763.320 3253.160 2763.580 3253.420 ;
        RECT 2763.320 1372.960 2763.580 1373.220 ;
        RECT 2900.860 1372.960 2901.120 1373.220 ;
      LAYER met2 ;
        RECT 862.090 3256.930 862.370 3260.000 ;
        RECT 861.740 3256.790 862.370 3256.930 ;
        RECT 861.740 3256.510 861.880 3256.790 ;
        RECT 861.680 3256.190 861.940 3256.510 ;
        RECT 862.090 3256.000 862.370 3256.790 ;
        RECT 2763.320 3253.130 2763.580 3253.450 ;
        RECT 2763.380 1373.250 2763.520 3253.130 ;
        RECT 2763.320 1372.930 2763.580 1373.250 ;
        RECT 2900.860 1372.930 2901.120 1373.250 ;
        RECT 2900.920 1368.685 2901.060 1372.930 ;
        RECT 2900.850 1368.315 2901.130 1368.685 ;
      LAYER via2 ;
        RECT 2900.850 1368.360 2901.130 1368.640 ;
      LAYER met3 ;
        RECT 2900.825 1368.650 2901.155 1368.665 ;
        RECT 2917.600 1368.650 2924.800 1369.100 ;
        RECT 2900.825 1368.350 2924.800 1368.650 ;
        RECT 2900.825 1368.335 2901.155 1368.350 ;
        RECT 2917.600 1367.900 2924.800 1368.350 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2549.390 3271.040 2549.710 3271.100 ;
        RECT 2660.250 3271.040 2660.570 3271.100 ;
        RECT 2549.390 3270.900 2660.570 3271.040 ;
        RECT 2549.390 3270.840 2549.710 3270.900 ;
        RECT 2660.250 3270.840 2660.570 3270.900 ;
        RECT 2660.250 1607.760 2660.570 1607.820 ;
        RECT 2900.830 1607.760 2901.150 1607.820 ;
        RECT 2660.250 1607.620 2901.150 1607.760 ;
        RECT 2660.250 1607.560 2660.570 1607.620 ;
        RECT 2900.830 1607.560 2901.150 1607.620 ;
      LAYER via ;
        RECT 2549.420 3270.840 2549.680 3271.100 ;
        RECT 2660.280 3270.840 2660.540 3271.100 ;
        RECT 2660.280 1607.560 2660.540 1607.820 ;
        RECT 2900.860 1607.560 2901.120 1607.820 ;
      LAYER met2 ;
        RECT 2549.420 3270.810 2549.680 3271.130 ;
        RECT 2660.280 3270.810 2660.540 3271.130 ;
        RECT 2549.480 3260.000 2549.620 3270.810 ;
        RECT 2549.370 3256.000 2549.650 3260.000 ;
        RECT 2660.340 1607.850 2660.480 3270.810 ;
        RECT 2660.280 1607.530 2660.540 1607.850 ;
        RECT 2900.860 1607.530 2901.120 1607.850 ;
        RECT 2900.920 1603.285 2901.060 1607.530 ;
        RECT 2900.850 1602.915 2901.130 1603.285 ;
      LAYER via2 ;
        RECT 2900.850 1602.960 2901.130 1603.240 ;
      LAYER met3 ;
        RECT 2900.825 1603.250 2901.155 1603.265 ;
        RECT 2917.600 1603.250 2924.800 1603.700 ;
        RECT 2900.825 1602.950 2924.800 1603.250 ;
        RECT 2900.825 1602.935 2901.155 1602.950 ;
        RECT 2917.600 1602.500 2924.800 1602.950 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2849.845 1836.765 2850.935 1836.935 ;
        RECT 2849.845 1835.405 2850.015 1836.765 ;
        RECT 2850.765 1835.405 2850.935 1836.765 ;
      LAYER met1 ;
        RECT 2749.490 1835.560 2749.810 1835.620 ;
        RECT 2849.785 1835.560 2850.075 1835.605 ;
        RECT 2749.490 1835.420 2850.075 1835.560 ;
        RECT 2749.490 1835.360 2749.810 1835.420 ;
        RECT 2849.785 1835.375 2850.075 1835.420 ;
        RECT 2850.705 1835.560 2850.995 1835.605 ;
        RECT 2900.830 1835.560 2901.150 1835.620 ;
        RECT 2850.705 1835.420 2901.150 1835.560 ;
        RECT 2850.705 1835.375 2850.995 1835.420 ;
        RECT 2900.830 1835.360 2901.150 1835.420 ;
        RECT 1528.190 251.500 1528.510 251.560 ;
        RECT 2749.490 251.500 2749.810 251.560 ;
        RECT 1528.190 251.360 2749.810 251.500 ;
        RECT 1528.190 251.300 1528.510 251.360 ;
        RECT 2749.490 251.300 2749.810 251.360 ;
      LAYER via ;
        RECT 2749.520 1835.360 2749.780 1835.620 ;
        RECT 2900.860 1835.360 2901.120 1835.620 ;
        RECT 1528.220 251.300 1528.480 251.560 ;
        RECT 2749.520 251.300 2749.780 251.560 ;
      LAYER met2 ;
        RECT 2900.850 1837.515 2901.130 1837.885 ;
        RECT 2900.920 1835.650 2901.060 1837.515 ;
        RECT 2749.520 1835.330 2749.780 1835.650 ;
        RECT 2900.860 1835.330 2901.120 1835.650 ;
        RECT 1528.170 260.000 1528.450 264.000 ;
        RECT 1528.280 251.590 1528.420 260.000 ;
        RECT 2749.580 251.590 2749.720 1835.330 ;
        RECT 1528.220 251.270 1528.480 251.590 ;
        RECT 2749.520 251.270 2749.780 251.590 ;
      LAYER via2 ;
        RECT 2900.850 1837.560 2901.130 1837.840 ;
      LAYER met3 ;
        RECT 2900.825 1837.850 2901.155 1837.865 ;
        RECT 2917.600 1837.850 2924.800 1838.300 ;
        RECT 2900.825 1837.550 2924.800 1837.850 ;
        RECT 2900.825 1837.535 2901.155 1837.550 ;
        RECT 2917.600 1837.100 2924.800 1837.550 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2092.150 3273.420 2092.470 3273.480 ;
        RECT 2701.190 3273.420 2701.510 3273.480 ;
        RECT 2092.150 3273.280 2701.510 3273.420 ;
        RECT 2092.150 3273.220 2092.470 3273.280 ;
        RECT 2701.190 3273.220 2701.510 3273.280 ;
        RECT 2701.190 2076.960 2701.510 2077.020 ;
        RECT 2900.830 2076.960 2901.150 2077.020 ;
        RECT 2701.190 2076.820 2901.150 2076.960 ;
        RECT 2701.190 2076.760 2701.510 2076.820 ;
        RECT 2900.830 2076.760 2901.150 2076.820 ;
      LAYER via ;
        RECT 2092.180 3273.220 2092.440 3273.480 ;
        RECT 2701.220 3273.220 2701.480 3273.480 ;
        RECT 2701.220 2076.760 2701.480 2077.020 ;
        RECT 2900.860 2076.760 2901.120 2077.020 ;
      LAYER met2 ;
        RECT 2092.180 3273.190 2092.440 3273.510 ;
        RECT 2701.220 3273.190 2701.480 3273.510 ;
        RECT 2092.240 3260.000 2092.380 3273.190 ;
        RECT 2092.130 3256.000 2092.410 3260.000 ;
        RECT 2701.280 2077.050 2701.420 3273.190 ;
        RECT 2701.220 2076.730 2701.480 2077.050 ;
        RECT 2900.860 2076.730 2901.120 2077.050 ;
        RECT 2900.920 2072.485 2901.060 2076.730 ;
        RECT 2900.850 2072.115 2901.130 2072.485 ;
      LAYER via2 ;
        RECT 2900.850 2072.160 2901.130 2072.440 ;
      LAYER met3 ;
        RECT 2900.825 2072.450 2901.155 2072.465 ;
        RECT 2917.600 2072.450 2924.800 2072.900 ;
        RECT 2900.825 2072.150 2924.800 2072.450 ;
        RECT 2900.825 2072.135 2901.155 2072.150 ;
        RECT 2917.600 2071.700 2924.800 2072.150 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2687.390 2304.760 2687.710 2304.820 ;
        RECT 2900.830 2304.760 2901.150 2304.820 ;
        RECT 2687.390 2304.620 2901.150 2304.760 ;
        RECT 2687.390 2304.560 2687.710 2304.620 ;
        RECT 2900.830 2304.560 2901.150 2304.620 ;
        RECT 813.350 240.280 813.670 240.340 ;
        RECT 2687.390 240.280 2687.710 240.340 ;
        RECT 813.350 240.140 2687.710 240.280 ;
        RECT 813.350 240.080 813.670 240.140 ;
        RECT 2687.390 240.080 2687.710 240.140 ;
      LAYER via ;
        RECT 2687.420 2304.560 2687.680 2304.820 ;
        RECT 2900.860 2304.560 2901.120 2304.820 ;
        RECT 813.380 240.080 813.640 240.340 ;
        RECT 2687.420 240.080 2687.680 240.340 ;
      LAYER met2 ;
        RECT 2900.850 2306.715 2901.130 2307.085 ;
        RECT 2900.920 2304.850 2901.060 2306.715 ;
        RECT 2687.420 2304.530 2687.680 2304.850 ;
        RECT 2900.860 2304.530 2901.120 2304.850 ;
        RECT 813.330 260.000 813.610 264.000 ;
        RECT 813.440 240.370 813.580 260.000 ;
        RECT 2687.480 240.370 2687.620 2304.530 ;
        RECT 813.380 240.050 813.640 240.370 ;
        RECT 2687.420 240.050 2687.680 240.370 ;
      LAYER via2 ;
        RECT 2900.850 2306.760 2901.130 2307.040 ;
      LAYER met3 ;
        RECT 2900.825 2307.050 2901.155 2307.065 ;
        RECT 2917.600 2307.050 2924.800 2307.500 ;
        RECT 2900.825 2306.750 2924.800 2307.050 ;
        RECT 2900.825 2306.735 2901.155 2306.750 ;
        RECT 2917.600 2306.300 2924.800 2306.750 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2708.090 124.000 2708.410 124.060 ;
        RECT 2900.830 124.000 2901.150 124.060 ;
        RECT 2708.090 123.860 2901.150 124.000 ;
        RECT 2708.090 123.800 2708.410 123.860 ;
        RECT 2900.830 123.800 2901.150 123.860 ;
      LAYER via ;
        RECT 2708.120 123.800 2708.380 124.060 ;
        RECT 2900.860 123.800 2901.120 124.060 ;
      LAYER met2 ;
        RECT 719.490 3258.290 719.770 3260.000 ;
        RECT 720.450 3258.290 720.730 3258.405 ;
        RECT 719.490 3258.150 720.730 3258.290 ;
        RECT 719.490 3256.000 719.770 3258.150 ;
        RECT 720.450 3258.035 720.730 3258.150 ;
        RECT 2708.110 3249.875 2708.390 3250.245 ;
        RECT 2708.180 124.090 2708.320 3249.875 ;
        RECT 2708.120 123.770 2708.380 124.090 ;
        RECT 2900.860 123.770 2901.120 124.090 ;
        RECT 2900.920 117.485 2901.060 123.770 ;
        RECT 2900.850 117.115 2901.130 117.485 ;
      LAYER via2 ;
        RECT 720.450 3258.080 720.730 3258.360 ;
        RECT 2708.110 3249.920 2708.390 3250.200 ;
        RECT 2900.850 117.160 2901.130 117.440 ;
      LAYER met3 ;
        RECT 720.425 3258.380 720.755 3258.385 ;
        RECT 720.425 3258.370 721.010 3258.380 ;
        RECT 720.425 3258.070 721.210 3258.370 ;
        RECT 720.425 3258.060 721.010 3258.070 ;
        RECT 720.425 3258.055 720.755 3258.060 ;
        RECT 720.630 3250.210 721.010 3250.220 ;
        RECT 2708.085 3250.210 2708.415 3250.225 ;
        RECT 720.630 3249.910 2708.415 3250.210 ;
        RECT 720.630 3249.900 721.010 3249.910 ;
        RECT 2708.085 3249.895 2708.415 3249.910 ;
        RECT 2900.825 117.450 2901.155 117.465 ;
        RECT 2917.600 117.450 2924.800 117.900 ;
        RECT 2900.825 117.150 2924.800 117.450 ;
        RECT 2900.825 117.135 2901.155 117.150 ;
        RECT 2917.600 116.700 2924.800 117.150 ;
      LAYER via3 ;
        RECT 720.660 3258.060 720.980 3258.380 ;
        RECT 720.660 3249.900 720.980 3250.220 ;
      LAYER met4 ;
        RECT 720.655 3258.055 720.985 3258.385 ;
        RECT 720.670 3250.225 720.970 3258.055 ;
        RECT 720.655 3249.895 720.985 3250.225 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 605.965 3252.525 606.135 3256.435 ;
      LAYER mcon ;
        RECT 605.965 3256.265 606.135 3256.435 ;
      LAYER met1 ;
        RECT 605.890 3256.420 606.210 3256.480 ;
        RECT 605.695 3256.280 606.210 3256.420 ;
        RECT 605.890 3256.220 606.210 3256.280 ;
        RECT 605.905 3252.680 606.195 3252.725 ;
        RECT 2680.490 3252.680 2680.810 3252.740 ;
        RECT 605.905 3252.540 2680.810 3252.680 ;
        RECT 605.905 3252.495 606.195 3252.540 ;
        RECT 2680.490 3252.480 2680.810 3252.540 ;
        RECT 2680.490 2470.000 2680.810 2470.060 ;
        RECT 2900.830 2470.000 2901.150 2470.060 ;
        RECT 2680.490 2469.860 2901.150 2470.000 ;
        RECT 2680.490 2469.800 2680.810 2469.860 ;
        RECT 2900.830 2469.800 2901.150 2469.860 ;
      LAYER via ;
        RECT 605.920 3256.220 606.180 3256.480 ;
        RECT 2680.520 3252.480 2680.780 3252.740 ;
        RECT 2680.520 2469.800 2680.780 2470.060 ;
        RECT 2900.860 2469.800 2901.120 2470.060 ;
      LAYER met2 ;
        RECT 604.490 3256.930 604.770 3260.000 ;
        RECT 604.490 3256.790 606.120 3256.930 ;
        RECT 604.490 3256.000 604.770 3256.790 ;
        RECT 605.980 3256.510 606.120 3256.790 ;
        RECT 605.920 3256.190 606.180 3256.510 ;
        RECT 2680.520 3252.450 2680.780 3252.770 ;
        RECT 2680.580 2470.090 2680.720 3252.450 ;
        RECT 2680.520 2469.770 2680.780 2470.090 ;
        RECT 2900.860 2469.770 2901.120 2470.090 ;
        RECT 2900.920 2463.485 2901.060 2469.770 ;
        RECT 2900.850 2463.115 2901.130 2463.485 ;
      LAYER via2 ;
        RECT 2900.850 2463.160 2901.130 2463.440 ;
      LAYER met3 ;
        RECT 2900.825 2463.450 2901.155 2463.465 ;
        RECT 2917.600 2463.450 2924.800 2463.900 ;
        RECT 2900.825 2463.150 2924.800 2463.450 ;
        RECT 2900.825 2463.135 2901.155 2463.150 ;
        RECT 2917.600 2462.700 2924.800 2463.150 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2859.890 2698.140 2860.210 2698.200 ;
        RECT 2900.830 2698.140 2901.150 2698.200 ;
        RECT 2859.890 2698.000 2901.150 2698.140 ;
        RECT 2859.890 2697.940 2860.210 2698.000 ;
        RECT 2900.830 2697.940 2901.150 2698.000 ;
        RECT 941.230 240.620 941.550 240.680 ;
        RECT 2859.890 240.620 2860.210 240.680 ;
        RECT 941.230 240.480 2860.210 240.620 ;
        RECT 941.230 240.420 941.550 240.480 ;
        RECT 2859.890 240.420 2860.210 240.480 ;
      LAYER via ;
        RECT 2859.920 2697.940 2860.180 2698.200 ;
        RECT 2900.860 2697.940 2901.120 2698.200 ;
        RECT 941.260 240.420 941.520 240.680 ;
        RECT 2859.920 240.420 2860.180 240.680 ;
      LAYER met2 ;
        RECT 2859.920 2697.910 2860.180 2698.230 ;
        RECT 2900.860 2698.085 2901.120 2698.230 ;
        RECT 941.210 260.000 941.490 264.000 ;
        RECT 941.320 240.710 941.460 260.000 ;
        RECT 2859.980 240.710 2860.120 2697.910 ;
        RECT 2900.850 2697.715 2901.130 2698.085 ;
        RECT 941.260 240.390 941.520 240.710 ;
        RECT 2859.920 240.390 2860.180 240.710 ;
      LAYER via2 ;
        RECT 2900.850 2697.760 2901.130 2698.040 ;
      LAYER met3 ;
        RECT 2900.825 2698.050 2901.155 2698.065 ;
        RECT 2917.600 2698.050 2924.800 2698.500 ;
        RECT 2900.825 2697.750 2924.800 2698.050 ;
        RECT 2900.825 2697.735 2901.155 2697.750 ;
        RECT 2917.600 2697.300 2924.800 2697.750 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2735.690 2932.740 2736.010 2932.800 ;
        RECT 2900.830 2932.740 2901.150 2932.800 ;
        RECT 2735.690 2932.600 2901.150 2932.740 ;
        RECT 2735.690 2932.540 2736.010 2932.600 ;
        RECT 2900.830 2932.540 2901.150 2932.600 ;
        RECT 2085.710 254.220 2086.030 254.280 ;
        RECT 2735.690 254.220 2736.010 254.280 ;
        RECT 2085.710 254.080 2736.010 254.220 ;
        RECT 2085.710 254.020 2086.030 254.080 ;
        RECT 2735.690 254.020 2736.010 254.080 ;
      LAYER via ;
        RECT 2735.720 2932.540 2735.980 2932.800 ;
        RECT 2900.860 2932.540 2901.120 2932.800 ;
        RECT 2085.740 254.020 2086.000 254.280 ;
        RECT 2735.720 254.020 2735.980 254.280 ;
      LAYER met2 ;
        RECT 2735.720 2932.510 2735.980 2932.830 ;
        RECT 2900.860 2932.685 2901.120 2932.830 ;
        RECT 2085.690 260.000 2085.970 264.000 ;
        RECT 2085.800 254.310 2085.940 260.000 ;
        RECT 2735.780 254.310 2735.920 2932.510 ;
        RECT 2900.850 2932.315 2901.130 2932.685 ;
        RECT 2085.740 253.990 2086.000 254.310 ;
        RECT 2735.720 253.990 2735.980 254.310 ;
      LAYER via2 ;
        RECT 2900.850 2932.360 2901.130 2932.640 ;
      LAYER met3 ;
        RECT 2900.825 2932.650 2901.155 2932.665 ;
        RECT 2917.600 2932.650 2924.800 2933.100 ;
        RECT 2900.825 2932.350 2924.800 2932.650 ;
        RECT 2900.825 2932.335 2901.155 2932.350 ;
        RECT 2917.600 2931.900 2924.800 2932.350 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2673.590 3167.340 2673.910 3167.400 ;
        RECT 2900.830 3167.340 2901.150 3167.400 ;
        RECT 2673.590 3167.200 2901.150 3167.340 ;
        RECT 2673.590 3167.140 2673.910 3167.200 ;
        RECT 2900.830 3167.140 2901.150 3167.200 ;
        RECT 2171.270 254.900 2171.590 254.960 ;
        RECT 2673.590 254.900 2673.910 254.960 ;
        RECT 2171.270 254.760 2673.910 254.900 ;
        RECT 2171.270 254.700 2171.590 254.760 ;
        RECT 2673.590 254.700 2673.910 254.760 ;
      LAYER via ;
        RECT 2673.620 3167.140 2673.880 3167.400 ;
        RECT 2900.860 3167.140 2901.120 3167.400 ;
        RECT 2171.300 254.700 2171.560 254.960 ;
        RECT 2673.620 254.700 2673.880 254.960 ;
      LAYER met2 ;
        RECT 2673.620 3167.110 2673.880 3167.430 ;
        RECT 2900.860 3167.285 2901.120 3167.430 ;
        RECT 2171.250 260.000 2171.530 264.000 ;
        RECT 2171.360 254.990 2171.500 260.000 ;
        RECT 2673.680 254.990 2673.820 3167.110 ;
        RECT 2900.850 3166.915 2901.130 3167.285 ;
        RECT 2171.300 254.670 2171.560 254.990 ;
        RECT 2673.620 254.670 2673.880 254.990 ;
      LAYER via2 ;
        RECT 2900.850 3166.960 2901.130 3167.240 ;
      LAYER met3 ;
        RECT 2900.825 3167.250 2901.155 3167.265 ;
        RECT 2917.600 3167.250 2924.800 3167.700 ;
        RECT 2900.825 3166.950 2924.800 3167.250 ;
        RECT 2900.825 3166.935 2901.155 3166.950 ;
        RECT 2917.600 3166.500 2924.800 3166.950 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2729.250 3401.940 2729.570 3402.000 ;
        RECT 2900.830 3401.940 2901.150 3402.000 ;
        RECT 2729.250 3401.800 2901.150 3401.940 ;
        RECT 2729.250 3401.740 2729.570 3401.800 ;
        RECT 2900.830 3401.740 2901.150 3401.800 ;
        RECT 2615.170 2035.480 2615.490 2035.540 ;
        RECT 2729.250 2035.480 2729.570 2035.540 ;
        RECT 2615.170 2035.340 2729.570 2035.480 ;
        RECT 2615.170 2035.280 2615.490 2035.340 ;
        RECT 2729.250 2035.280 2729.570 2035.340 ;
      LAYER via ;
        RECT 2729.280 3401.740 2729.540 3402.000 ;
        RECT 2900.860 3401.740 2901.120 3402.000 ;
        RECT 2615.200 2035.280 2615.460 2035.540 ;
        RECT 2729.280 2035.280 2729.540 2035.540 ;
      LAYER met2 ;
        RECT 2729.280 3401.710 2729.540 3402.030 ;
        RECT 2900.860 3401.885 2901.120 3402.030 ;
        RECT 2729.340 2035.570 2729.480 3401.710 ;
        RECT 2900.850 3401.515 2901.130 3401.885 ;
        RECT 2615.200 2035.250 2615.460 2035.570 ;
        RECT 2729.280 2035.250 2729.540 2035.570 ;
        RECT 2615.260 2029.645 2615.400 2035.250 ;
        RECT 2615.190 2029.275 2615.470 2029.645 ;
      LAYER via2 ;
        RECT 2900.850 3401.560 2901.130 3401.840 ;
        RECT 2615.190 2029.320 2615.470 2029.600 ;
      LAYER met3 ;
        RECT 2900.825 3401.850 2901.155 3401.865 ;
        RECT 2917.600 3401.850 2924.800 3402.300 ;
        RECT 2900.825 3401.550 2924.800 3401.850 ;
        RECT 2900.825 3401.535 2901.155 3401.550 ;
        RECT 2917.600 3401.100 2924.800 3401.550 ;
        RECT 2606.000 2029.610 2610.000 2030.000 ;
        RECT 2615.165 2029.610 2615.495 2029.625 ;
        RECT 2606.000 2029.400 2615.495 2029.610 ;
        RECT 2609.580 2029.310 2615.495 2029.400 ;
        RECT 2615.165 2029.295 2615.495 2029.310 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2753.170 3464.160 2753.490 3464.220 ;
        RECT 2757.770 3464.160 2758.090 3464.220 ;
        RECT 2753.170 3464.020 2758.090 3464.160 ;
        RECT 2753.170 3463.960 2753.490 3464.020 ;
        RECT 2757.770 3463.960 2758.090 3464.020 ;
        RECT 2701.650 3432.540 2701.970 3432.600 ;
        RECT 2753.170 3432.540 2753.490 3432.600 ;
        RECT 2701.650 3432.400 2753.490 3432.540 ;
        RECT 2701.650 3432.340 2701.970 3432.400 ;
        RECT 2753.170 3432.340 2753.490 3432.400 ;
        RECT 2615.170 3070.440 2615.490 3070.500 ;
        RECT 2701.650 3070.440 2701.970 3070.500 ;
        RECT 2615.170 3070.300 2701.970 3070.440 ;
        RECT 2615.170 3070.240 2615.490 3070.300 ;
        RECT 2701.650 3070.240 2701.970 3070.300 ;
      LAYER via ;
        RECT 2753.200 3463.960 2753.460 3464.220 ;
        RECT 2757.800 3463.960 2758.060 3464.220 ;
        RECT 2701.680 3432.340 2701.940 3432.600 ;
        RECT 2753.200 3432.340 2753.460 3432.600 ;
        RECT 2615.200 3070.240 2615.460 3070.500 ;
        RECT 2701.680 3070.240 2701.940 3070.500 ;
      LAYER met2 ;
        RECT 2757.190 3517.600 2757.750 3524.800 ;
        RECT 2757.400 3517.370 2757.540 3517.600 ;
        RECT 2757.400 3517.230 2758.000 3517.370 ;
        RECT 2757.860 3464.250 2758.000 3517.230 ;
        RECT 2753.200 3463.930 2753.460 3464.250 ;
        RECT 2757.800 3463.930 2758.060 3464.250 ;
        RECT 2753.260 3432.630 2753.400 3463.930 ;
        RECT 2701.680 3432.310 2701.940 3432.630 ;
        RECT 2753.200 3432.310 2753.460 3432.630 ;
        RECT 2701.740 3070.530 2701.880 3432.310 ;
        RECT 2615.200 3070.210 2615.460 3070.530 ;
        RECT 2701.680 3070.210 2701.940 3070.530 ;
        RECT 2615.260 3065.965 2615.400 3070.210 ;
        RECT 2615.190 3065.595 2615.470 3065.965 ;
      LAYER via2 ;
        RECT 2615.190 3065.640 2615.470 3065.920 ;
      LAYER met3 ;
        RECT 2606.000 3065.930 2610.000 3066.320 ;
        RECT 2615.165 3065.930 2615.495 3065.945 ;
        RECT 2606.000 3065.720 2615.495 3065.930 ;
        RECT 2609.580 3065.630 2615.495 3065.720 ;
        RECT 2615.165 3065.615 2615.495 3065.630 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2428.870 3464.160 2429.190 3464.220 ;
        RECT 2433.470 3464.160 2433.790 3464.220 ;
        RECT 2428.870 3464.020 2433.790 3464.160 ;
        RECT 2428.870 3463.960 2429.190 3464.020 ;
        RECT 2433.470 3463.960 2433.790 3464.020 ;
        RECT 2428.870 3367.600 2429.190 3367.660 ;
        RECT 2429.790 3367.600 2430.110 3367.660 ;
        RECT 2428.870 3367.460 2430.110 3367.600 ;
        RECT 2428.870 3367.400 2429.190 3367.460 ;
        RECT 2429.790 3367.400 2430.110 3367.460 ;
        RECT 304.130 3308.440 304.450 3308.500 ;
        RECT 2429.790 3308.440 2430.110 3308.500 ;
        RECT 304.130 3308.300 2430.110 3308.440 ;
        RECT 304.130 3308.240 304.450 3308.300 ;
        RECT 2429.790 3308.240 2430.110 3308.300 ;
      LAYER via ;
        RECT 2428.900 3463.960 2429.160 3464.220 ;
        RECT 2433.500 3463.960 2433.760 3464.220 ;
        RECT 2428.900 3367.400 2429.160 3367.660 ;
        RECT 2429.820 3367.400 2430.080 3367.660 ;
        RECT 304.160 3308.240 304.420 3308.500 ;
        RECT 2429.820 3308.240 2430.080 3308.500 ;
      LAYER met2 ;
        RECT 2432.890 3517.600 2433.450 3524.800 ;
        RECT 2433.100 3517.370 2433.240 3517.600 ;
        RECT 2433.100 3517.230 2433.700 3517.370 ;
        RECT 2433.560 3464.250 2433.700 3517.230 ;
        RECT 2428.900 3463.930 2429.160 3464.250 ;
        RECT 2433.500 3463.930 2433.760 3464.250 ;
        RECT 2428.960 3415.370 2429.100 3463.930 ;
        RECT 2428.960 3415.230 2430.020 3415.370 ;
        RECT 2429.880 3367.690 2430.020 3415.230 ;
        RECT 2428.900 3367.370 2429.160 3367.690 ;
        RECT 2429.820 3367.370 2430.080 3367.690 ;
        RECT 2428.960 3318.810 2429.100 3367.370 ;
        RECT 2428.960 3318.670 2430.020 3318.810 ;
        RECT 2429.880 3308.530 2430.020 3318.670 ;
        RECT 304.160 3308.210 304.420 3308.530 ;
        RECT 2429.820 3308.210 2430.080 3308.530 ;
        RECT 304.220 2568.205 304.360 3308.210 ;
        RECT 304.150 2567.835 304.430 2568.205 ;
      LAYER via2 ;
        RECT 304.150 2567.880 304.430 2568.160 ;
      LAYER met3 ;
        RECT 304.125 2568.170 304.455 2568.185 ;
        RECT 310.000 2568.170 314.000 2568.560 ;
        RECT 304.125 2567.960 314.000 2568.170 ;
        RECT 304.125 2567.870 310.500 2567.960 ;
        RECT 304.125 2567.855 304.455 2567.870 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2108.590 3517.600 2109.150 3524.800 ;
        RECT 2108.800 3501.845 2108.940 3517.600 ;
        RECT 2108.730 3501.475 2109.010 3501.845 ;
        RECT 341.370 260.000 341.650 264.000 ;
        RECT 341.480 255.525 341.620 260.000 ;
        RECT 341.410 255.155 341.690 255.525 ;
      LAYER via2 ;
        RECT 2108.730 3501.520 2109.010 3501.800 ;
        RECT 341.410 255.200 341.690 255.480 ;
      LAYER met3 ;
        RECT 267.990 3501.810 268.370 3501.820 ;
        RECT 2108.705 3501.810 2109.035 3501.825 ;
        RECT 267.990 3501.510 2109.035 3501.810 ;
        RECT 267.990 3501.500 268.370 3501.510 ;
        RECT 2108.705 3501.495 2109.035 3501.510 ;
        RECT 267.990 255.490 268.370 255.500 ;
        RECT 341.385 255.490 341.715 255.505 ;
        RECT 267.990 255.190 341.715 255.490 ;
        RECT 267.990 255.180 268.370 255.190 ;
        RECT 341.385 255.175 341.715 255.190 ;
      LAYER via3 ;
        RECT 268.020 3501.500 268.340 3501.820 ;
        RECT 268.020 255.180 268.340 255.500 ;
      LAYER met4 ;
        RECT 268.015 3501.495 268.345 3501.825 ;
        RECT 268.030 255.505 268.330 3501.495 ;
        RECT 268.015 255.175 268.345 255.505 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1783.830 3517.600 1784.390 3524.800 ;
        RECT 1784.040 3502.525 1784.180 3517.600 ;
        RECT 1783.970 3502.155 1784.250 3502.525 ;
        RECT 555.730 260.000 556.010 264.000 ;
        RECT 555.840 247.365 555.980 260.000 ;
        RECT 555.770 246.995 556.050 247.365 ;
      LAYER via2 ;
        RECT 1783.970 3502.200 1784.250 3502.480 ;
        RECT 555.770 247.040 556.050 247.320 ;
      LAYER met3 ;
        RECT 253.270 3502.490 253.650 3502.500 ;
        RECT 1783.945 3502.490 1784.275 3502.505 ;
        RECT 253.270 3502.190 1784.275 3502.490 ;
        RECT 253.270 3502.180 253.650 3502.190 ;
        RECT 1783.945 3502.175 1784.275 3502.190 ;
        RECT 253.270 247.330 253.650 247.340 ;
        RECT 555.745 247.330 556.075 247.345 ;
        RECT 253.270 247.030 556.075 247.330 ;
        RECT 253.270 247.020 253.650 247.030 ;
        RECT 555.745 247.015 556.075 247.030 ;
      LAYER via3 ;
        RECT 253.300 3502.180 253.620 3502.500 ;
        RECT 253.300 247.020 253.620 247.340 ;
      LAYER met4 ;
        RECT 253.295 3502.175 253.625 3502.505 ;
        RECT 253.310 247.345 253.610 3502.175 ;
        RECT 253.295 247.015 253.625 247.345 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1459.650 3502.920 1459.970 3502.980 ;
        RECT 1600.870 3502.920 1601.190 3502.980 ;
        RECT 1459.650 3502.780 1601.190 3502.920 ;
        RECT 1459.650 3502.720 1459.970 3502.780 ;
        RECT 1600.870 3502.720 1601.190 3502.780 ;
      LAYER via ;
        RECT 1459.680 3502.720 1459.940 3502.980 ;
        RECT 1600.900 3502.720 1601.160 3502.980 ;
      LAYER met2 ;
        RECT 1459.530 3517.600 1460.090 3524.800 ;
        RECT 1459.740 3503.010 1459.880 3517.600 ;
        RECT 1459.680 3502.690 1459.940 3503.010 ;
        RECT 1600.900 3502.690 1601.160 3503.010 ;
        RECT 1600.960 3258.970 1601.100 3502.690 ;
        RECT 1605.450 3258.970 1605.730 3260.000 ;
        RECT 1600.960 3258.830 1605.730 3258.970 ;
        RECT 1605.450 3256.000 1605.730 3258.830 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 271.470 724.780 271.790 724.840 ;
        RECT 296.770 724.780 297.090 724.840 ;
        RECT 271.470 724.640 297.090 724.780 ;
        RECT 271.470 724.580 271.790 724.640 ;
        RECT 296.770 724.580 297.090 724.640 ;
        RECT 271.470 262.040 271.790 262.100 ;
        RECT 2901.750 262.040 2902.070 262.100 ;
        RECT 271.470 261.900 2902.070 262.040 ;
        RECT 271.470 261.840 271.790 261.900 ;
        RECT 2901.750 261.840 2902.070 261.900 ;
      LAYER via ;
        RECT 271.500 724.580 271.760 724.840 ;
        RECT 296.800 724.580 297.060 724.840 ;
        RECT 271.500 261.840 271.760 262.100 ;
        RECT 2901.780 261.840 2902.040 262.100 ;
      LAYER met2 ;
        RECT 296.790 727.755 297.070 728.125 ;
        RECT 296.860 724.870 297.000 727.755 ;
        RECT 271.500 724.550 271.760 724.870 ;
        RECT 296.800 724.550 297.060 724.870 ;
        RECT 271.560 262.130 271.700 724.550 ;
        RECT 2901.770 351.715 2902.050 352.085 ;
        RECT 2901.840 262.130 2901.980 351.715 ;
        RECT 271.500 261.810 271.760 262.130 ;
        RECT 2901.780 261.810 2902.040 262.130 ;
      LAYER via2 ;
        RECT 296.790 727.800 297.070 728.080 ;
        RECT 2901.770 351.760 2902.050 352.040 ;
      LAYER met3 ;
        RECT 296.765 728.090 297.095 728.105 ;
        RECT 310.000 728.090 314.000 728.480 ;
        RECT 296.765 727.880 314.000 728.090 ;
        RECT 296.765 727.790 310.500 727.880 ;
        RECT 296.765 727.775 297.095 727.790 ;
        RECT 2901.745 352.050 2902.075 352.065 ;
        RECT 2917.600 352.050 2924.800 352.500 ;
        RECT 2901.745 351.750 2924.800 352.050 ;
        RECT 2901.745 351.735 2902.075 351.750 ;
        RECT 2917.600 351.300 2924.800 351.750 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 314.325 313.225 314.495 337.875 ;
      LAYER mcon ;
        RECT 314.325 337.705 314.495 337.875 ;
      LAYER met1 ;
        RECT 286.190 3503.600 286.510 3503.660 ;
        RECT 1135.350 3503.600 1135.670 3503.660 ;
        RECT 286.190 3503.460 1135.670 3503.600 ;
        RECT 286.190 3503.400 286.510 3503.460 ;
        RECT 1135.350 3503.400 1135.670 3503.460 ;
        RECT 278.830 761.160 279.150 761.220 ;
        RECT 286.190 761.160 286.510 761.220 ;
        RECT 278.830 761.020 286.510 761.160 ;
        RECT 278.830 760.960 279.150 761.020 ;
        RECT 286.190 760.960 286.510 761.020 ;
        RECT 278.830 483.040 279.150 483.100 ;
        RECT 311.030 483.040 311.350 483.100 ;
        RECT 278.830 482.900 311.350 483.040 ;
        RECT 278.830 482.840 279.150 482.900 ;
        RECT 311.030 482.840 311.350 482.900 ;
        RECT 303.210 386.140 303.530 386.200 ;
        RECT 311.030 386.140 311.350 386.200 ;
        RECT 303.210 386.000 311.350 386.140 ;
        RECT 303.210 385.940 303.530 386.000 ;
        RECT 311.030 385.940 311.350 386.000 ;
        RECT 303.210 358.260 303.530 358.320 ;
        RECT 314.250 358.260 314.570 358.320 ;
        RECT 303.210 358.120 314.570 358.260 ;
        RECT 303.210 358.060 303.530 358.120 ;
        RECT 314.250 358.060 314.570 358.120 ;
        RECT 314.250 337.860 314.570 337.920 ;
        RECT 314.250 337.720 314.765 337.860 ;
        RECT 314.250 337.660 314.570 337.720 ;
        RECT 314.250 313.380 314.570 313.440 ;
        RECT 314.055 313.240 314.570 313.380 ;
        RECT 314.250 313.180 314.570 313.240 ;
        RECT 314.250 253.880 314.570 253.940 ;
        RECT 1742.550 253.880 1742.870 253.940 ;
        RECT 314.250 253.740 1742.870 253.880 ;
        RECT 314.250 253.680 314.570 253.740 ;
        RECT 1742.550 253.680 1742.870 253.740 ;
      LAYER via ;
        RECT 286.220 3503.400 286.480 3503.660 ;
        RECT 1135.380 3503.400 1135.640 3503.660 ;
        RECT 278.860 760.960 279.120 761.220 ;
        RECT 286.220 760.960 286.480 761.220 ;
        RECT 278.860 482.840 279.120 483.100 ;
        RECT 311.060 482.840 311.320 483.100 ;
        RECT 303.240 385.940 303.500 386.200 ;
        RECT 311.060 385.940 311.320 386.200 ;
        RECT 303.240 358.060 303.500 358.320 ;
        RECT 314.280 358.060 314.540 358.320 ;
        RECT 314.280 337.660 314.540 337.920 ;
        RECT 314.280 313.180 314.540 313.440 ;
        RECT 314.280 253.680 314.540 253.940 ;
        RECT 1742.580 253.680 1742.840 253.940 ;
      LAYER met2 ;
        RECT 1135.230 3517.600 1135.790 3524.800 ;
        RECT 1135.440 3503.690 1135.580 3517.600 ;
        RECT 286.220 3503.370 286.480 3503.690 ;
        RECT 1135.380 3503.370 1135.640 3503.690 ;
        RECT 286.280 761.250 286.420 3503.370 ;
        RECT 278.860 760.930 279.120 761.250 ;
        RECT 286.220 760.930 286.480 761.250 ;
        RECT 278.920 483.130 279.060 760.930 ;
        RECT 278.860 482.810 279.120 483.130 ;
        RECT 311.060 482.810 311.320 483.130 ;
        RECT 311.120 386.230 311.260 482.810 ;
        RECT 303.240 385.910 303.500 386.230 ;
        RECT 311.060 385.910 311.320 386.230 ;
        RECT 303.300 358.350 303.440 385.910 ;
        RECT 303.240 358.030 303.500 358.350 ;
        RECT 314.280 358.030 314.540 358.350 ;
        RECT 314.340 337.950 314.480 358.030 ;
        RECT 314.280 337.630 314.540 337.950 ;
        RECT 314.280 313.150 314.540 313.470 ;
        RECT 314.340 253.970 314.480 313.150 ;
        RECT 1742.530 260.000 1742.810 264.000 ;
        RECT 1742.640 253.970 1742.780 260.000 ;
        RECT 314.280 253.650 314.540 253.970 ;
        RECT 1742.580 253.650 1742.840 253.970 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 313.790 3503.940 314.110 3504.000 ;
        RECT 810.590 3503.940 810.910 3504.000 ;
        RECT 313.790 3503.800 810.910 3503.940 ;
        RECT 313.790 3503.740 314.110 3503.800 ;
        RECT 810.590 3503.740 810.910 3503.800 ;
      LAYER via ;
        RECT 313.820 3503.740 314.080 3504.000 ;
        RECT 810.620 3503.740 810.880 3504.000 ;
      LAYER met2 ;
        RECT 810.470 3517.600 811.030 3524.800 ;
        RECT 810.680 3504.030 810.820 3517.600 ;
        RECT 313.820 3503.710 314.080 3504.030 ;
        RECT 810.620 3503.710 810.880 3504.030 ;
        RECT 313.350 485.930 313.630 486.045 ;
        RECT 313.880 485.930 314.020 3503.710 ;
        RECT 313.350 485.790 314.020 485.930 ;
        RECT 313.350 485.675 313.630 485.790 ;
        RECT 598.050 260.000 598.330 264.000 ;
        RECT 598.160 246.685 598.300 260.000 ;
        RECT 598.090 246.315 598.370 246.685 ;
      LAYER via2 ;
        RECT 313.350 485.720 313.630 486.000 ;
        RECT 598.090 246.360 598.370 246.640 ;
      LAYER met3 ;
        RECT 285.470 486.010 285.850 486.020 ;
        RECT 313.325 486.010 313.655 486.025 ;
        RECT 285.470 485.710 313.655 486.010 ;
        RECT 285.470 485.700 285.850 485.710 ;
        RECT 313.325 485.695 313.655 485.710 ;
        RECT 326.870 246.650 327.250 246.660 ;
        RECT 598.065 246.650 598.395 246.665 ;
        RECT 326.870 246.350 598.395 246.650 ;
        RECT 326.870 246.340 327.250 246.350 ;
        RECT 598.065 246.335 598.395 246.350 ;
      LAYER via3 ;
        RECT 285.500 485.700 285.820 486.020 ;
        RECT 326.900 246.340 327.220 246.660 ;
      LAYER met4 ;
        RECT 285.495 485.695 285.825 486.025 ;
        RECT 285.510 270.890 285.810 485.695 ;
        RECT 285.070 269.710 286.250 270.890 ;
        RECT 326.470 266.310 327.650 267.490 ;
        RECT 326.910 246.665 327.210 266.310 ;
        RECT 326.895 246.335 327.225 246.665 ;
      LAYER met5 ;
        RECT 284.860 269.500 327.860 271.100 ;
        RECT 326.260 266.100 327.860 269.500 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 3504.280 255.230 3504.340 ;
        RECT 486.290 3504.280 486.610 3504.340 ;
        RECT 254.910 3504.140 486.610 3504.280 ;
        RECT 254.910 3504.080 255.230 3504.140 ;
        RECT 486.290 3504.080 486.610 3504.140 ;
        RECT 254.910 247.760 255.230 247.820 ;
        RECT 912.710 247.760 913.030 247.820 ;
        RECT 254.910 247.620 913.030 247.760 ;
        RECT 254.910 247.560 255.230 247.620 ;
        RECT 912.710 247.560 913.030 247.620 ;
      LAYER via ;
        RECT 254.940 3504.080 255.200 3504.340 ;
        RECT 486.320 3504.080 486.580 3504.340 ;
        RECT 254.940 247.560 255.200 247.820 ;
        RECT 912.740 247.560 913.000 247.820 ;
      LAYER met2 ;
        RECT 486.170 3517.600 486.730 3524.800 ;
        RECT 486.380 3504.370 486.520 3517.600 ;
        RECT 254.940 3504.050 255.200 3504.370 ;
        RECT 486.320 3504.050 486.580 3504.370 ;
        RECT 255.000 247.850 255.140 3504.050 ;
        RECT 912.690 260.000 912.970 264.000 ;
        RECT 912.800 247.850 912.940 260.000 ;
        RECT 254.940 247.530 255.200 247.850 ;
        RECT 912.740 247.530 913.000 247.850 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.870 3517.600 162.430 3524.800 ;
        RECT 162.080 3501.845 162.220 3517.600 ;
        RECT 162.010 3501.475 162.290 3501.845 ;
        RECT 2385.610 260.000 2385.890 264.000 ;
        RECT 2385.720 241.245 2385.860 260.000 ;
        RECT 2385.650 240.875 2385.930 241.245 ;
      LAYER via2 ;
        RECT 162.010 3501.520 162.290 3501.800 ;
        RECT 2385.650 240.920 2385.930 241.200 ;
      LAYER met3 ;
        RECT 161.985 3501.810 162.315 3501.825 ;
        RECT 244.070 3501.810 244.450 3501.820 ;
        RECT 161.985 3501.510 244.450 3501.810 ;
        RECT 161.985 3501.495 162.315 3501.510 ;
        RECT 244.070 3501.500 244.450 3501.510 ;
        RECT 244.070 241.210 244.450 241.220 ;
        RECT 2385.625 241.210 2385.955 241.225 ;
        RECT 244.070 240.910 2385.955 241.210 ;
        RECT 244.070 240.900 244.450 240.910 ;
        RECT 2385.625 240.895 2385.955 240.910 ;
      LAYER via3 ;
        RECT 244.100 3501.500 244.420 3501.820 ;
        RECT 244.100 240.900 244.420 241.220 ;
      LAYER met4 ;
        RECT 244.095 3501.495 244.425 3501.825 ;
        RECT 244.110 241.225 244.410 3501.495 ;
        RECT 244.095 240.895 244.425 241.225 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3388.000 17.410 3388.060 ;
        RECT 2616.550 3388.000 2616.870 3388.060 ;
        RECT 17.090 3387.860 2616.870 3388.000 ;
        RECT 17.090 3387.800 17.410 3387.860 ;
        RECT 2616.550 3387.800 2616.870 3387.860 ;
      LAYER via ;
        RECT 17.120 3387.800 17.380 3388.060 ;
        RECT 2616.580 3387.800 2616.840 3388.060 ;
      LAYER met2 ;
        RECT 17.110 3393.355 17.390 3393.725 ;
        RECT 17.180 3388.090 17.320 3393.355 ;
        RECT 17.120 3387.770 17.380 3388.090 ;
        RECT 2616.580 3387.770 2616.840 3388.090 ;
        RECT 2616.640 2262.205 2616.780 3387.770 ;
        RECT 2616.570 2261.835 2616.850 2262.205 ;
      LAYER via2 ;
        RECT 17.110 3393.400 17.390 3393.680 ;
        RECT 2616.570 2261.880 2616.850 2262.160 ;
      LAYER met3 ;
        RECT -4.800 3393.690 2.400 3394.140 ;
        RECT 17.085 3393.690 17.415 3393.705 ;
        RECT -4.800 3393.390 17.415 3393.690 ;
        RECT -4.800 3392.940 2.400 3393.390 ;
        RECT 17.085 3393.375 17.415 3393.390 ;
        RECT 2606.000 2262.170 2610.000 2262.560 ;
        RECT 2616.545 2262.170 2616.875 2262.185 ;
        RECT 2606.000 2261.960 2616.875 2262.170 ;
        RECT 2609.580 2261.870 2616.875 2261.960 ;
        RECT 2616.545 2261.855 2616.875 2261.870 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 3139.800 16.950 3139.860 ;
        RECT 65.850 3139.800 66.170 3139.860 ;
        RECT 16.630 3139.660 66.170 3139.800 ;
        RECT 16.630 3139.600 16.950 3139.660 ;
        RECT 65.850 3139.600 66.170 3139.660 ;
        RECT 65.850 2235.400 66.170 2235.460 ;
        RECT 296.770 2235.400 297.090 2235.460 ;
        RECT 65.850 2235.260 297.090 2235.400 ;
        RECT 65.850 2235.200 66.170 2235.260 ;
        RECT 296.770 2235.200 297.090 2235.260 ;
      LAYER via ;
        RECT 16.660 3139.600 16.920 3139.860 ;
        RECT 65.880 3139.600 66.140 3139.860 ;
        RECT 65.880 2235.200 66.140 2235.460 ;
        RECT 296.800 2235.200 297.060 2235.460 ;
      LAYER met2 ;
        RECT 16.650 3141.755 16.930 3142.125 ;
        RECT 16.720 3139.890 16.860 3141.755 ;
        RECT 16.660 3139.570 16.920 3139.890 ;
        RECT 65.880 3139.570 66.140 3139.890 ;
        RECT 65.940 2235.490 66.080 3139.570 ;
        RECT 65.880 2235.170 66.140 2235.490 ;
        RECT 296.800 2235.170 297.060 2235.490 ;
        RECT 296.860 2229.565 297.000 2235.170 ;
        RECT 296.790 2229.195 297.070 2229.565 ;
      LAYER via2 ;
        RECT 16.650 3141.800 16.930 3142.080 ;
        RECT 296.790 2229.240 297.070 2229.520 ;
      LAYER met3 ;
        RECT -4.800 3142.090 2.400 3142.540 ;
        RECT 16.625 3142.090 16.955 3142.105 ;
        RECT -4.800 3141.790 16.955 3142.090 ;
        RECT -4.800 3141.340 2.400 3141.790 ;
        RECT 16.625 3141.775 16.955 3141.790 ;
        RECT 296.765 2229.530 297.095 2229.545 ;
        RECT 310.000 2229.530 314.000 2229.920 ;
        RECT 296.765 2229.320 314.000 2229.530 ;
        RECT 296.765 2229.230 310.500 2229.320 ;
        RECT 296.765 2229.215 297.095 2229.230 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2884.460 15.110 2884.520 ;
        RECT 92.990 2884.460 93.310 2884.520 ;
        RECT 14.790 2884.320 93.310 2884.460 ;
        RECT 14.790 2884.260 15.110 2884.320 ;
        RECT 92.990 2884.260 93.310 2884.320 ;
        RECT 92.990 254.560 93.310 254.620 ;
        RECT 798.630 254.560 798.950 254.620 ;
        RECT 92.990 254.420 798.950 254.560 ;
        RECT 92.990 254.360 93.310 254.420 ;
        RECT 798.630 254.360 798.950 254.420 ;
      LAYER via ;
        RECT 14.820 2884.260 15.080 2884.520 ;
        RECT 93.020 2884.260 93.280 2884.520 ;
        RECT 93.020 254.360 93.280 254.620 ;
        RECT 798.660 254.360 798.920 254.620 ;
      LAYER met2 ;
        RECT 14.810 2890.835 15.090 2891.205 ;
        RECT 14.880 2884.550 15.020 2890.835 ;
        RECT 14.820 2884.230 15.080 2884.550 ;
        RECT 93.020 2884.230 93.280 2884.550 ;
        RECT 93.080 254.650 93.220 2884.230 ;
        RECT 798.610 260.000 798.890 264.000 ;
        RECT 798.720 254.650 798.860 260.000 ;
        RECT 93.020 254.330 93.280 254.650 ;
        RECT 798.660 254.330 798.920 254.650 ;
      LAYER via2 ;
        RECT 14.810 2890.880 15.090 2891.160 ;
      LAYER met3 ;
        RECT -4.800 2891.170 2.400 2891.620 ;
        RECT 14.785 2891.170 15.115 2891.185 ;
        RECT -4.800 2890.870 15.115 2891.170 ;
        RECT -4.800 2890.420 2.400 2890.870 ;
        RECT 14.785 2890.855 15.115 2890.870 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 731.545 3253.205 731.715 3256.435 ;
      LAYER mcon ;
        RECT 731.545 3256.265 731.715 3256.435 ;
      LAYER met1 ;
        RECT 731.470 3256.420 731.790 3256.480 ;
        RECT 731.275 3256.280 731.790 3256.420 ;
        RECT 731.470 3256.220 731.790 3256.280 ;
        RECT 162.450 3253.360 162.770 3253.420 ;
        RECT 731.485 3253.360 731.775 3253.405 ;
        RECT 162.450 3253.220 731.775 3253.360 ;
        RECT 162.450 3253.160 162.770 3253.220 ;
        RECT 731.485 3253.175 731.775 3253.220 ;
        RECT 19.390 2642.720 19.710 2642.780 ;
        RECT 162.450 2642.720 162.770 2642.780 ;
        RECT 19.390 2642.580 162.770 2642.720 ;
        RECT 19.390 2642.520 19.710 2642.580 ;
        RECT 162.450 2642.520 162.770 2642.580 ;
      LAYER via ;
        RECT 731.500 3256.220 731.760 3256.480 ;
        RECT 162.480 3253.160 162.740 3253.420 ;
        RECT 19.420 2642.520 19.680 2642.780 ;
        RECT 162.480 2642.520 162.740 2642.780 ;
      LAYER met2 ;
        RECT 733.290 3256.930 733.570 3260.000 ;
        RECT 731.560 3256.790 733.570 3256.930 ;
        RECT 731.560 3256.510 731.700 3256.790 ;
        RECT 731.500 3256.190 731.760 3256.510 ;
        RECT 733.290 3256.000 733.570 3256.790 ;
        RECT 162.480 3253.130 162.740 3253.450 ;
        RECT 162.540 2642.810 162.680 3253.130 ;
        RECT 19.420 2642.490 19.680 2642.810 ;
        RECT 162.480 2642.490 162.740 2642.810 ;
        RECT 19.480 2639.605 19.620 2642.490 ;
        RECT 19.410 2639.235 19.690 2639.605 ;
      LAYER via2 ;
        RECT 19.410 2639.280 19.690 2639.560 ;
      LAYER met3 ;
        RECT -4.800 2639.570 2.400 2640.020 ;
        RECT 19.385 2639.570 19.715 2639.585 ;
        RECT -4.800 2639.270 19.715 2639.570 ;
        RECT -4.800 2638.820 2.400 2639.270 ;
        RECT 19.385 2639.255 19.715 2639.270 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2387.720 20.630 2387.780 ;
        RECT 251.690 2387.720 252.010 2387.780 ;
        RECT 20.310 2387.580 252.010 2387.720 ;
        RECT 20.310 2387.520 20.630 2387.580 ;
        RECT 251.690 2387.520 252.010 2387.580 ;
        RECT 251.690 253.540 252.010 253.600 ;
        RECT 855.670 253.540 855.990 253.600 ;
        RECT 251.690 253.400 855.990 253.540 ;
        RECT 251.690 253.340 252.010 253.400 ;
        RECT 855.670 253.340 855.990 253.400 ;
      LAYER via ;
        RECT 20.340 2387.520 20.600 2387.780 ;
        RECT 251.720 2387.520 251.980 2387.780 ;
        RECT 251.720 253.340 251.980 253.600 ;
        RECT 855.700 253.340 855.960 253.600 ;
      LAYER met2 ;
        RECT 20.330 2387.635 20.610 2388.005 ;
        RECT 20.340 2387.490 20.600 2387.635 ;
        RECT 251.720 2387.490 251.980 2387.810 ;
        RECT 251.780 253.630 251.920 2387.490 ;
        RECT 855.650 260.000 855.930 264.000 ;
        RECT 855.760 253.630 855.900 260.000 ;
        RECT 251.720 253.310 251.980 253.630 ;
        RECT 855.700 253.310 855.960 253.630 ;
      LAYER via2 ;
        RECT 20.330 2387.680 20.610 2387.960 ;
      LAYER met3 ;
        RECT -4.800 2387.970 2.400 2388.420 ;
        RECT 20.305 2387.970 20.635 2387.985 ;
        RECT -4.800 2387.670 20.635 2387.970 ;
        RECT -4.800 2387.220 2.400 2387.670 ;
        RECT 20.305 2387.655 20.635 2387.670 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 2132.380 20.170 2132.440 ;
        RECT 73.210 2132.380 73.530 2132.440 ;
        RECT 19.850 2132.240 73.530 2132.380 ;
        RECT 19.850 2132.180 20.170 2132.240 ;
        RECT 73.210 2132.180 73.530 2132.240 ;
        RECT 73.210 1531.600 73.530 1531.660 ;
        RECT 296.770 1531.600 297.090 1531.660 ;
        RECT 73.210 1531.460 297.090 1531.600 ;
        RECT 73.210 1531.400 73.530 1531.460 ;
        RECT 296.770 1531.400 297.090 1531.460 ;
      LAYER via ;
        RECT 19.880 2132.180 20.140 2132.440 ;
        RECT 73.240 2132.180 73.500 2132.440 ;
        RECT 73.240 1531.400 73.500 1531.660 ;
        RECT 296.800 1531.400 297.060 1531.660 ;
      LAYER met2 ;
        RECT 19.870 2136.035 20.150 2136.405 ;
        RECT 19.940 2132.470 20.080 2136.035 ;
        RECT 19.880 2132.150 20.140 2132.470 ;
        RECT 73.240 2132.150 73.500 2132.470 ;
        RECT 73.300 1531.690 73.440 2132.150 ;
        RECT 73.240 1531.370 73.500 1531.690 ;
        RECT 296.790 1531.515 297.070 1531.885 ;
        RECT 296.800 1531.370 297.060 1531.515 ;
      LAYER via2 ;
        RECT 19.870 2136.080 20.150 2136.360 ;
        RECT 296.790 1531.560 297.070 1531.840 ;
      LAYER met3 ;
        RECT -4.800 2136.370 2.400 2136.820 ;
        RECT 19.845 2136.370 20.175 2136.385 ;
        RECT -4.800 2136.070 20.175 2136.370 ;
        RECT -4.800 2135.620 2.400 2136.070 ;
        RECT 19.845 2136.055 20.175 2136.070 ;
        RECT 296.765 1531.850 297.095 1531.865 ;
        RECT 310.000 1531.850 314.000 1532.240 ;
        RECT 296.765 1531.640 314.000 1531.850 ;
        RECT 296.765 1531.550 310.500 1531.640 ;
        RECT 296.765 1531.535 297.095 1531.550 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 3163.600 2615.490 3163.660 ;
        RECT 2818.490 3163.600 2818.810 3163.660 ;
        RECT 2615.170 3163.460 2818.810 3163.600 ;
        RECT 2615.170 3163.400 2615.490 3163.460 ;
        RECT 2818.490 3163.400 2818.810 3163.460 ;
        RECT 2818.490 593.200 2818.810 593.260 ;
        RECT 2900.830 593.200 2901.150 593.260 ;
        RECT 2818.490 593.060 2901.150 593.200 ;
        RECT 2818.490 593.000 2818.810 593.060 ;
        RECT 2900.830 593.000 2901.150 593.060 ;
      LAYER via ;
        RECT 2615.200 3163.400 2615.460 3163.660 ;
        RECT 2818.520 3163.400 2818.780 3163.660 ;
        RECT 2818.520 593.000 2818.780 593.260 ;
        RECT 2900.860 593.000 2901.120 593.260 ;
      LAYER met2 ;
        RECT 2615.190 3170.315 2615.470 3170.685 ;
        RECT 2615.260 3163.690 2615.400 3170.315 ;
        RECT 2615.200 3163.370 2615.460 3163.690 ;
        RECT 2818.520 3163.370 2818.780 3163.690 ;
        RECT 2818.580 593.290 2818.720 3163.370 ;
        RECT 2818.520 592.970 2818.780 593.290 ;
        RECT 2900.860 592.970 2901.120 593.290 ;
        RECT 2900.920 586.685 2901.060 592.970 ;
        RECT 2900.850 586.315 2901.130 586.685 ;
      LAYER via2 ;
        RECT 2615.190 3170.360 2615.470 3170.640 ;
        RECT 2900.850 586.360 2901.130 586.640 ;
      LAYER met3 ;
        RECT 2606.000 3170.650 2610.000 3171.040 ;
        RECT 2615.165 3170.650 2615.495 3170.665 ;
        RECT 2606.000 3170.440 2615.495 3170.650 ;
        RECT 2609.580 3170.350 2615.495 3170.440 ;
        RECT 2615.165 3170.335 2615.495 3170.350 ;
        RECT 2900.825 586.650 2901.155 586.665 ;
        RECT 2917.600 586.650 2924.800 587.100 ;
        RECT 2900.825 586.350 2924.800 586.650 ;
        RECT 2900.825 586.335 2901.155 586.350 ;
        RECT 2917.600 585.900 2924.800 586.350 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1124.385 3254.225 1124.555 3255.075 ;
        RECT 1159.345 3254.225 1159.515 3255.755 ;
        RECT 1207.185 3253.885 1207.355 3255.755 ;
        RECT 1218.225 3253.885 1218.395 3256.435 ;
      LAYER mcon ;
        RECT 1218.225 3256.265 1218.395 3256.435 ;
        RECT 1159.345 3255.585 1159.515 3255.755 ;
        RECT 1124.385 3254.905 1124.555 3255.075 ;
        RECT 1207.185 3255.585 1207.355 3255.755 ;
      LAYER met1 ;
        RECT 1218.150 3256.420 1218.470 3256.480 ;
        RECT 1217.955 3256.280 1218.470 3256.420 ;
        RECT 1218.150 3256.220 1218.470 3256.280 ;
        RECT 1159.285 3255.740 1159.575 3255.785 ;
        RECT 1207.125 3255.740 1207.415 3255.785 ;
        RECT 1159.285 3255.600 1207.415 3255.740 ;
        RECT 1159.285 3255.555 1159.575 3255.600 ;
        RECT 1207.125 3255.555 1207.415 3255.600 ;
        RECT 1124.325 3255.060 1124.615 3255.105 ;
        RECT 1028.720 3254.920 1124.615 3255.060 ;
        RECT 169.350 3254.380 169.670 3254.440 ;
        RECT 1028.720 3254.380 1028.860 3254.920 ;
        RECT 1124.325 3254.875 1124.615 3254.920 ;
        RECT 169.350 3254.240 1028.860 3254.380 ;
        RECT 1124.325 3254.380 1124.615 3254.425 ;
        RECT 1159.285 3254.380 1159.575 3254.425 ;
        RECT 1124.325 3254.240 1159.575 3254.380 ;
        RECT 169.350 3254.180 169.670 3254.240 ;
        RECT 1124.325 3254.195 1124.615 3254.240 ;
        RECT 1159.285 3254.195 1159.575 3254.240 ;
        RECT 1207.125 3254.040 1207.415 3254.085 ;
        RECT 1218.165 3254.040 1218.455 3254.085 ;
        RECT 1207.125 3253.900 1218.455 3254.040 ;
        RECT 1207.125 3253.855 1207.415 3253.900 ;
        RECT 1218.165 3253.855 1218.455 3253.900 ;
        RECT 19.850 1890.640 20.170 1890.700 ;
        RECT 169.350 1890.640 169.670 1890.700 ;
        RECT 19.850 1890.500 169.670 1890.640 ;
        RECT 19.850 1890.440 20.170 1890.500 ;
        RECT 169.350 1890.440 169.670 1890.500 ;
      LAYER via ;
        RECT 1218.180 3256.220 1218.440 3256.480 ;
        RECT 169.380 3254.180 169.640 3254.440 ;
        RECT 19.880 1890.440 20.140 1890.700 ;
        RECT 169.380 1890.440 169.640 1890.700 ;
      LAYER met2 ;
        RECT 1219.970 3256.930 1220.250 3260.000 ;
        RECT 1218.240 3256.790 1220.250 3256.930 ;
        RECT 1218.240 3256.510 1218.380 3256.790 ;
        RECT 1218.180 3256.190 1218.440 3256.510 ;
        RECT 1219.970 3256.000 1220.250 3256.790 ;
        RECT 169.380 3254.150 169.640 3254.470 ;
        RECT 169.440 1890.730 169.580 3254.150 ;
        RECT 19.880 1890.410 20.140 1890.730 ;
        RECT 169.380 1890.410 169.640 1890.730 ;
        RECT 19.940 1885.485 20.080 1890.410 ;
        RECT 19.870 1885.115 20.150 1885.485 ;
      LAYER via2 ;
        RECT 19.870 1885.160 20.150 1885.440 ;
      LAYER met3 ;
        RECT -4.800 1885.450 2.400 1885.900 ;
        RECT 19.845 1885.450 20.175 1885.465 ;
        RECT -4.800 1885.150 20.175 1885.450 ;
        RECT -4.800 1884.700 2.400 1885.150 ;
        RECT 19.845 1885.135 20.175 1885.150 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.330 1633.515 20.610 1633.885 ;
        RECT 20.400 1629.125 20.540 1633.515 ;
        RECT 20.330 1628.755 20.610 1629.125 ;
        RECT 159.710 1628.755 159.990 1629.125 ;
        RECT 159.780 1594.445 159.920 1628.755 ;
        RECT 159.710 1594.075 159.990 1594.445 ;
        RECT 174.430 1545.115 174.710 1545.485 ;
        RECT 174.500 1498.565 174.640 1545.115 ;
        RECT 174.430 1498.195 174.710 1498.565 ;
        RECT 176.270 1448.555 176.550 1448.925 ;
        RECT 176.340 1402.005 176.480 1448.555 ;
        RECT 176.270 1401.635 176.550 1402.005 ;
        RECT 174.430 1351.995 174.710 1352.365 ;
        RECT 174.500 1305.445 174.640 1351.995 ;
        RECT 174.430 1305.075 174.710 1305.445 ;
        RECT 176.270 1296.915 176.550 1297.285 ;
        RECT 176.340 1250.365 176.480 1296.915 ;
        RECT 176.270 1249.995 176.550 1250.365 ;
        RECT 176.270 1200.355 176.550 1200.725 ;
        RECT 176.340 1153.805 176.480 1200.355 ;
        RECT 176.270 1153.435 176.550 1153.805 ;
        RECT 177.190 1141.875 177.470 1142.245 ;
        RECT 177.260 1112.325 177.400 1141.875 ;
        RECT 177.190 1111.955 177.470 1112.325 ;
      LAYER via2 ;
        RECT 20.330 1633.560 20.610 1633.840 ;
        RECT 20.330 1628.800 20.610 1629.080 ;
        RECT 159.710 1628.800 159.990 1629.080 ;
        RECT 159.710 1594.120 159.990 1594.400 ;
        RECT 174.430 1545.160 174.710 1545.440 ;
        RECT 174.430 1498.240 174.710 1498.520 ;
        RECT 176.270 1448.600 176.550 1448.880 ;
        RECT 176.270 1401.680 176.550 1401.960 ;
        RECT 174.430 1352.040 174.710 1352.320 ;
        RECT 174.430 1305.120 174.710 1305.400 ;
        RECT 176.270 1296.960 176.550 1297.240 ;
        RECT 176.270 1250.040 176.550 1250.320 ;
        RECT 176.270 1200.400 176.550 1200.680 ;
        RECT 176.270 1153.480 176.550 1153.760 ;
        RECT 177.190 1141.920 177.470 1142.200 ;
        RECT 177.190 1112.000 177.470 1112.280 ;
      LAYER met3 ;
        RECT -4.800 1633.850 2.400 1634.300 ;
        RECT 20.305 1633.850 20.635 1633.865 ;
        RECT -4.800 1633.550 20.635 1633.850 ;
        RECT -4.800 1633.100 2.400 1633.550 ;
        RECT 20.305 1633.535 20.635 1633.550 ;
        RECT 20.305 1629.090 20.635 1629.105 ;
        RECT 159.685 1629.090 160.015 1629.105 ;
        RECT 20.305 1628.790 160.015 1629.090 ;
        RECT 20.305 1628.775 20.635 1628.790 ;
        RECT 159.685 1628.775 160.015 1628.790 ;
        RECT 159.685 1594.410 160.015 1594.425 ;
        RECT 175.070 1594.410 175.450 1594.420 ;
        RECT 159.685 1594.110 175.450 1594.410 ;
        RECT 159.685 1594.095 160.015 1594.110 ;
        RECT 175.070 1594.100 175.450 1594.110 ;
        RECT 175.070 1560.410 175.450 1560.420 ;
        RECT 174.190 1560.110 175.450 1560.410 ;
        RECT 174.190 1559.060 174.490 1560.110 ;
        RECT 175.070 1560.100 175.450 1560.110 ;
        RECT 174.150 1558.740 174.530 1559.060 ;
        RECT 174.405 1545.460 174.735 1545.465 ;
        RECT 174.150 1545.450 174.735 1545.460 ;
        RECT 174.150 1545.150 174.960 1545.450 ;
        RECT 174.150 1545.140 174.735 1545.150 ;
        RECT 174.405 1545.135 174.735 1545.140 ;
        RECT 174.405 1498.530 174.735 1498.545 ;
        RECT 173.270 1498.230 174.735 1498.530 ;
        RECT 173.270 1497.860 173.570 1498.230 ;
        RECT 174.405 1498.215 174.735 1498.230 ;
        RECT 173.230 1497.540 173.610 1497.860 ;
        RECT 173.230 1463.540 173.610 1463.860 ;
        RECT 173.270 1463.170 173.570 1463.540 ;
        RECT 175.990 1463.170 176.370 1463.180 ;
        RECT 173.270 1462.870 176.370 1463.170 ;
        RECT 175.990 1462.860 176.370 1462.870 ;
        RECT 176.245 1448.900 176.575 1448.905 ;
        RECT 175.990 1448.890 176.575 1448.900 ;
        RECT 175.990 1448.590 176.800 1448.890 ;
        RECT 175.990 1448.580 176.575 1448.590 ;
        RECT 176.245 1448.575 176.575 1448.580 ;
        RECT 176.245 1401.970 176.575 1401.985 ;
        RECT 175.110 1401.670 176.575 1401.970 ;
        RECT 175.110 1401.300 175.410 1401.670 ;
        RECT 176.245 1401.655 176.575 1401.670 ;
        RECT 175.070 1400.980 175.450 1401.300 ;
        RECT 175.070 1367.290 175.450 1367.300 ;
        RECT 174.190 1366.990 175.450 1367.290 ;
        RECT 174.190 1365.940 174.490 1366.990 ;
        RECT 175.070 1366.980 175.450 1366.990 ;
        RECT 174.150 1365.620 174.530 1365.940 ;
        RECT 174.405 1352.340 174.735 1352.345 ;
        RECT 174.150 1352.330 174.735 1352.340 ;
        RECT 173.950 1352.030 174.735 1352.330 ;
        RECT 174.150 1352.020 174.735 1352.030 ;
        RECT 174.405 1352.015 174.735 1352.020 ;
        RECT 174.405 1305.410 174.735 1305.425 ;
        RECT 175.070 1305.410 175.450 1305.420 ;
        RECT 174.405 1305.110 175.450 1305.410 ;
        RECT 174.405 1305.095 174.735 1305.110 ;
        RECT 175.070 1305.100 175.450 1305.110 ;
        RECT 175.070 1304.050 175.450 1304.060 ;
        RECT 175.990 1304.050 176.370 1304.060 ;
        RECT 175.070 1303.750 176.370 1304.050 ;
        RECT 175.070 1303.740 175.450 1303.750 ;
        RECT 175.990 1303.740 176.370 1303.750 ;
        RECT 176.245 1297.260 176.575 1297.265 ;
        RECT 175.990 1297.250 176.575 1297.260 ;
        RECT 175.990 1296.950 176.800 1297.250 ;
        RECT 175.990 1296.940 176.575 1296.950 ;
        RECT 176.245 1296.935 176.575 1296.940 ;
        RECT 176.245 1250.330 176.575 1250.345 ;
        RECT 176.030 1250.015 176.575 1250.330 ;
        RECT 176.030 1249.660 176.330 1250.015 ;
        RECT 175.990 1249.340 176.370 1249.660 ;
        RECT 175.990 1221.460 176.370 1221.780 ;
        RECT 176.030 1220.410 176.330 1221.460 ;
        RECT 176.910 1220.410 177.290 1220.420 ;
        RECT 176.030 1220.110 177.290 1220.410 ;
        RECT 176.910 1220.100 177.290 1220.110 ;
        RECT 176.245 1200.690 176.575 1200.705 ;
        RECT 176.910 1200.690 177.290 1200.700 ;
        RECT 176.245 1200.390 177.290 1200.690 ;
        RECT 176.245 1200.375 176.575 1200.390 ;
        RECT 176.910 1200.380 177.290 1200.390 ;
        RECT 176.245 1153.770 176.575 1153.785 ;
        RECT 176.030 1153.455 176.575 1153.770 ;
        RECT 176.030 1153.100 176.330 1153.455 ;
        RECT 175.990 1152.780 176.370 1153.100 ;
        RECT 175.990 1142.210 176.370 1142.220 ;
        RECT 177.165 1142.210 177.495 1142.225 ;
        RECT 175.990 1141.910 177.495 1142.210 ;
        RECT 175.990 1141.900 176.370 1141.910 ;
        RECT 177.165 1141.895 177.495 1141.910 ;
        RECT 177.165 1112.290 177.495 1112.305 ;
        RECT 177.830 1112.290 178.210 1112.300 ;
        RECT 177.165 1111.990 178.210 1112.290 ;
        RECT 177.165 1111.975 177.495 1111.990 ;
        RECT 177.830 1111.980 178.210 1111.990 ;
        RECT 177.830 1110.930 178.210 1110.940 ;
        RECT 192.550 1110.930 192.930 1110.940 ;
        RECT 177.830 1110.630 192.930 1110.930 ;
        RECT 177.830 1110.620 178.210 1110.630 ;
        RECT 192.550 1110.620 192.930 1110.630 ;
        RECT 285.470 1062.650 285.850 1062.660 ;
        RECT 308.470 1062.650 308.850 1062.660 ;
        RECT 285.470 1062.350 308.850 1062.650 ;
        RECT 285.470 1062.340 285.850 1062.350 ;
        RECT 308.470 1062.340 308.850 1062.350 ;
        RECT 2612.150 1059.930 2612.530 1059.940 ;
        RECT 2609.430 1059.630 2612.530 1059.930 ;
        RECT 2609.430 1057.600 2609.730 1059.630 ;
        RECT 2612.150 1059.620 2612.530 1059.630 ;
        RECT 2606.000 1057.000 2610.000 1057.600 ;
      LAYER via3 ;
        RECT 175.100 1594.100 175.420 1594.420 ;
        RECT 175.100 1560.100 175.420 1560.420 ;
        RECT 174.180 1558.740 174.500 1559.060 ;
        RECT 174.180 1545.140 174.500 1545.460 ;
        RECT 173.260 1497.540 173.580 1497.860 ;
        RECT 173.260 1463.540 173.580 1463.860 ;
        RECT 176.020 1462.860 176.340 1463.180 ;
        RECT 176.020 1448.580 176.340 1448.900 ;
        RECT 175.100 1400.980 175.420 1401.300 ;
        RECT 175.100 1366.980 175.420 1367.300 ;
        RECT 174.180 1365.620 174.500 1365.940 ;
        RECT 174.180 1352.020 174.500 1352.340 ;
        RECT 175.100 1305.100 175.420 1305.420 ;
        RECT 175.100 1303.740 175.420 1304.060 ;
        RECT 176.020 1303.740 176.340 1304.060 ;
        RECT 176.020 1296.940 176.340 1297.260 ;
        RECT 176.020 1249.340 176.340 1249.660 ;
        RECT 176.020 1221.460 176.340 1221.780 ;
        RECT 176.940 1220.100 177.260 1220.420 ;
        RECT 176.940 1200.380 177.260 1200.700 ;
        RECT 176.020 1152.780 176.340 1153.100 ;
        RECT 176.020 1141.900 176.340 1142.220 ;
        RECT 177.860 1111.980 178.180 1112.300 ;
        RECT 177.860 1110.620 178.180 1110.940 ;
        RECT 192.580 1110.620 192.900 1110.940 ;
        RECT 285.500 1062.340 285.820 1062.660 ;
        RECT 308.500 1062.340 308.820 1062.660 ;
        RECT 2612.180 1059.620 2612.500 1059.940 ;
      LAYER met4 ;
        RECT 175.095 1594.095 175.425 1594.425 ;
        RECT 175.110 1560.425 175.410 1594.095 ;
        RECT 175.095 1560.095 175.425 1560.425 ;
        RECT 174.175 1558.735 174.505 1559.065 ;
        RECT 174.190 1545.465 174.490 1558.735 ;
        RECT 174.175 1545.135 174.505 1545.465 ;
        RECT 173.255 1497.535 173.585 1497.865 ;
        RECT 173.270 1463.865 173.570 1497.535 ;
        RECT 173.255 1463.535 173.585 1463.865 ;
        RECT 176.015 1462.855 176.345 1463.185 ;
        RECT 176.030 1448.905 176.330 1462.855 ;
        RECT 176.015 1448.575 176.345 1448.905 ;
        RECT 175.095 1400.975 175.425 1401.305 ;
        RECT 175.110 1367.305 175.410 1400.975 ;
        RECT 175.095 1366.975 175.425 1367.305 ;
        RECT 174.175 1365.615 174.505 1365.945 ;
        RECT 174.190 1352.345 174.490 1365.615 ;
        RECT 174.175 1352.015 174.505 1352.345 ;
        RECT 175.095 1305.095 175.425 1305.425 ;
        RECT 175.110 1304.065 175.410 1305.095 ;
        RECT 175.095 1303.735 175.425 1304.065 ;
        RECT 176.015 1303.735 176.345 1304.065 ;
        RECT 176.030 1297.265 176.330 1303.735 ;
        RECT 176.015 1296.935 176.345 1297.265 ;
        RECT 176.015 1249.335 176.345 1249.665 ;
        RECT 176.030 1221.785 176.330 1249.335 ;
        RECT 176.015 1221.455 176.345 1221.785 ;
        RECT 176.935 1220.095 177.265 1220.425 ;
        RECT 176.950 1200.705 177.250 1220.095 ;
        RECT 176.935 1200.375 177.265 1200.705 ;
        RECT 176.015 1152.775 176.345 1153.105 ;
        RECT 176.030 1142.225 176.330 1152.775 ;
        RECT 176.015 1141.895 176.345 1142.225 ;
        RECT 177.855 1111.975 178.185 1112.305 ;
        RECT 177.870 1110.945 178.170 1111.975 ;
        RECT 177.855 1110.615 178.185 1110.945 ;
        RECT 192.575 1110.615 192.905 1110.945 ;
        RECT 192.590 1066.490 192.890 1110.615 ;
        RECT 192.150 1065.310 193.330 1066.490 ;
        RECT 285.070 1061.910 286.250 1063.090 ;
        RECT 308.495 1062.335 308.825 1062.665 ;
        RECT 308.510 1059.690 308.810 1062.335 ;
        RECT 2611.750 1061.910 2612.930 1063.090 ;
        RECT 2612.190 1059.945 2612.490 1061.910 ;
        RECT 308.070 1058.510 309.250 1059.690 ;
        RECT 2612.175 1059.615 2612.505 1059.945 ;
      LAYER met5 ;
        RECT 367.660 1085.500 408.820 1087.100 ;
        RECT 191.940 1065.100 228.500 1066.700 ;
        RECT 226.900 1063.300 228.500 1065.100 ;
        RECT 254.500 1065.100 276.340 1066.700 ;
        RECT 254.500 1063.300 256.100 1065.100 ;
        RECT 226.900 1061.700 256.100 1063.300 ;
        RECT 274.740 1063.300 276.340 1065.100 ;
        RECT 323.500 1065.100 355.460 1066.700 ;
        RECT 274.740 1061.700 286.460 1063.300 ;
        RECT 323.500 1059.900 325.100 1065.100 ;
        RECT 307.860 1058.300 325.100 1059.900 ;
        RECT 353.860 1059.900 355.460 1065.100 ;
        RECT 367.660 1063.300 369.260 1085.500 ;
        RECT 407.220 1083.700 408.820 1085.500 ;
        RECT 407.220 1082.100 414.340 1083.700 ;
        RECT 412.740 1073.500 414.340 1082.100 ;
        RECT 364.900 1061.700 369.260 1063.300 ;
        RECT 411.820 1071.900 414.340 1073.500 ;
        RECT 411.820 1063.300 413.420 1071.900 ;
        RECT 444.020 1065.100 449.300 1066.700 ;
        RECT 444.020 1063.300 445.620 1065.100 ;
        RECT 411.820 1061.700 445.620 1063.300 ;
        RECT 364.900 1059.900 366.500 1061.700 ;
        RECT 353.860 1058.300 366.500 1059.900 ;
        RECT 447.700 1059.900 449.300 1065.100 ;
        RECT 495.540 1065.100 545.900 1066.700 ;
        RECT 495.540 1059.900 497.140 1065.100 ;
        RECT 447.700 1058.300 497.140 1059.900 ;
        RECT 544.300 1059.900 545.900 1065.100 ;
        RECT 592.140 1065.100 642.500 1066.700 ;
        RECT 592.140 1059.900 593.740 1065.100 ;
        RECT 544.300 1058.300 593.740 1059.900 ;
        RECT 640.900 1059.900 642.500 1065.100 ;
        RECT 688.740 1065.100 739.100 1066.700 ;
        RECT 688.740 1059.900 690.340 1065.100 ;
        RECT 640.900 1058.300 690.340 1059.900 ;
        RECT 737.500 1059.900 739.100 1065.100 ;
        RECT 785.340 1065.100 835.700 1066.700 ;
        RECT 785.340 1059.900 786.940 1065.100 ;
        RECT 737.500 1058.300 786.940 1059.900 ;
        RECT 834.100 1059.900 835.700 1065.100 ;
        RECT 881.940 1065.100 932.300 1066.700 ;
        RECT 881.940 1059.900 883.540 1065.100 ;
        RECT 834.100 1058.300 883.540 1059.900 ;
        RECT 930.700 1059.900 932.300 1065.100 ;
        RECT 978.540 1059.900 981.060 1066.700 ;
        RECT 1026.380 1065.100 1077.660 1066.700 ;
        RECT 1026.380 1059.900 1027.980 1065.100 ;
        RECT 930.700 1058.300 1027.980 1059.900 ;
        RECT 1076.060 1059.900 1077.660 1065.100 ;
        RECT 1122.980 1065.100 1174.260 1066.700 ;
        RECT 1122.980 1059.900 1124.580 1065.100 ;
        RECT 1076.060 1058.300 1124.580 1059.900 ;
        RECT 1172.660 1059.900 1174.260 1065.100 ;
        RECT 1219.580 1065.100 1270.860 1066.700 ;
        RECT 1219.580 1059.900 1221.180 1065.100 ;
        RECT 1172.660 1058.300 1221.180 1059.900 ;
        RECT 1269.260 1059.900 1270.860 1065.100 ;
        RECT 1316.180 1065.100 1367.460 1066.700 ;
        RECT 1316.180 1059.900 1317.780 1065.100 ;
        RECT 1269.260 1058.300 1317.780 1059.900 ;
        RECT 1365.860 1059.900 1367.460 1065.100 ;
        RECT 1412.780 1065.100 1464.060 1066.700 ;
        RECT 1412.780 1059.900 1414.380 1065.100 ;
        RECT 1365.860 1058.300 1414.380 1059.900 ;
        RECT 1462.460 1059.900 1464.060 1065.100 ;
        RECT 1509.380 1065.100 1560.660 1066.700 ;
        RECT 1509.380 1059.900 1510.980 1065.100 ;
        RECT 1462.460 1058.300 1510.980 1059.900 ;
        RECT 1559.060 1059.900 1560.660 1065.100 ;
        RECT 1605.980 1065.100 1657.260 1066.700 ;
        RECT 1605.980 1059.900 1607.580 1065.100 ;
        RECT 1559.060 1058.300 1607.580 1059.900 ;
        RECT 1655.660 1059.900 1657.260 1065.100 ;
        RECT 1702.580 1065.100 1753.860 1066.700 ;
        RECT 1702.580 1059.900 1704.180 1065.100 ;
        RECT 1655.660 1058.300 1704.180 1059.900 ;
        RECT 1752.260 1059.900 1753.860 1065.100 ;
        RECT 1799.180 1065.100 1850.460 1066.700 ;
        RECT 1799.180 1059.900 1800.780 1065.100 ;
        RECT 1752.260 1058.300 1800.780 1059.900 ;
        RECT 1848.860 1059.900 1850.460 1065.100 ;
        RECT 1895.780 1065.100 1947.060 1066.700 ;
        RECT 1895.780 1059.900 1897.380 1065.100 ;
        RECT 1848.860 1058.300 1897.380 1059.900 ;
        RECT 1945.460 1059.900 1947.060 1065.100 ;
        RECT 1992.380 1065.100 2043.660 1066.700 ;
        RECT 1992.380 1059.900 1993.980 1065.100 ;
        RECT 1945.460 1058.300 1993.980 1059.900 ;
        RECT 2042.060 1059.900 2043.660 1065.100 ;
        RECT 2088.980 1065.100 2140.260 1066.700 ;
        RECT 2088.980 1059.900 2090.580 1065.100 ;
        RECT 2042.060 1058.300 2090.580 1059.900 ;
        RECT 2138.660 1059.900 2140.260 1065.100 ;
        RECT 2185.580 1065.100 2236.860 1066.700 ;
        RECT 2185.580 1059.900 2187.180 1065.100 ;
        RECT 2138.660 1058.300 2187.180 1059.900 ;
        RECT 2235.260 1059.900 2236.860 1065.100 ;
        RECT 2282.180 1065.100 2333.460 1066.700 ;
        RECT 2282.180 1059.900 2283.780 1065.100 ;
        RECT 2235.260 1058.300 2283.780 1059.900 ;
        RECT 2331.860 1059.900 2333.460 1065.100 ;
        RECT 2378.780 1065.100 2430.060 1066.700 ;
        RECT 2378.780 1059.900 2380.380 1065.100 ;
        RECT 2331.860 1058.300 2380.380 1059.900 ;
        RECT 2428.460 1059.900 2430.060 1065.100 ;
        RECT 2449.620 1065.100 2546.900 1066.700 ;
        RECT 2449.620 1059.900 2451.220 1065.100 ;
        RECT 2545.300 1063.300 2546.900 1065.100 ;
        RECT 2545.300 1061.700 2613.140 1063.300 ;
        RECT 2428.460 1058.300 2451.220 1059.900 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1052.165 3253.545 1052.335 3255.415 ;
        RECT 1100.465 3253.545 1100.635 3255.415 ;
        RECT 1125.305 3253.715 1125.475 3255.075 ;
        RECT 1124.845 3253.545 1125.475 3253.715 ;
        RECT 1242.145 3253.545 1242.315 3254.395 ;
        RECT 1269.285 3254.225 1269.915 3254.395 ;
        RECT 1304.245 3253.885 1304.415 3255.075 ;
        RECT 1352.085 3254.225 1352.255 3255.075 ;
        RECT 1365.885 3254.225 1366.515 3254.395 ;
        RECT 1400.845 3253.885 1401.015 3255.075 ;
        RECT 1424.765 3253.885 1424.935 3255.075 ;
        RECT 1560.005 3254.055 1560.175 3254.395 ;
        RECT 1594.045 3254.225 1594.215 3255.075 ;
        RECT 1559.085 3253.885 1560.175 3254.055 ;
        RECT 1641.885 3253.885 1642.055 3255.075 ;
        RECT 1661.665 3253.885 1661.835 3256.435 ;
      LAYER mcon ;
        RECT 1661.665 3256.265 1661.835 3256.435 ;
        RECT 1052.165 3255.245 1052.335 3255.415 ;
        RECT 1100.465 3255.245 1100.635 3255.415 ;
        RECT 1125.305 3254.905 1125.475 3255.075 ;
        RECT 1304.245 3254.905 1304.415 3255.075 ;
        RECT 1242.145 3254.225 1242.315 3254.395 ;
        RECT 1269.745 3254.225 1269.915 3254.395 ;
        RECT 1352.085 3254.905 1352.255 3255.075 ;
        RECT 1400.845 3254.905 1401.015 3255.075 ;
        RECT 1366.345 3254.225 1366.515 3254.395 ;
        RECT 1424.765 3254.905 1424.935 3255.075 ;
        RECT 1594.045 3254.905 1594.215 3255.075 ;
        RECT 1560.005 3254.225 1560.175 3254.395 ;
        RECT 1641.885 3254.905 1642.055 3255.075 ;
      LAYER met1 ;
        RECT 1661.590 3256.420 1661.910 3256.480 ;
        RECT 1661.395 3256.280 1661.910 3256.420 ;
        RECT 1661.590 3256.220 1661.910 3256.280 ;
        RECT 1052.105 3255.400 1052.395 3255.445 ;
        RECT 1100.405 3255.400 1100.695 3255.445 ;
        RECT 1052.105 3255.260 1100.695 3255.400 ;
        RECT 1052.105 3255.215 1052.395 3255.260 ;
        RECT 1100.405 3255.215 1100.695 3255.260 ;
        RECT 1125.245 3255.060 1125.535 3255.105 ;
        RECT 1304.185 3255.060 1304.475 3255.105 ;
        RECT 1352.025 3255.060 1352.315 3255.105 ;
        RECT 1125.245 3254.920 1219.300 3255.060 ;
        RECT 1125.245 3254.875 1125.535 3254.920 ;
        RECT 161.990 3253.700 162.310 3253.760 ;
        RECT 1052.105 3253.700 1052.395 3253.745 ;
        RECT 161.990 3253.560 1052.395 3253.700 ;
        RECT 161.990 3253.500 162.310 3253.560 ;
        RECT 1052.105 3253.515 1052.395 3253.560 ;
        RECT 1100.405 3253.700 1100.695 3253.745 ;
        RECT 1124.785 3253.700 1125.075 3253.745 ;
        RECT 1100.405 3253.560 1125.075 3253.700 ;
        RECT 1219.160 3253.700 1219.300 3254.920 ;
        RECT 1304.185 3254.920 1352.315 3255.060 ;
        RECT 1304.185 3254.875 1304.475 3254.920 ;
        RECT 1352.025 3254.875 1352.315 3254.920 ;
        RECT 1400.785 3255.060 1401.075 3255.105 ;
        RECT 1424.705 3255.060 1424.995 3255.105 ;
        RECT 1400.785 3254.920 1424.995 3255.060 ;
        RECT 1400.785 3254.875 1401.075 3254.920 ;
        RECT 1424.705 3254.875 1424.995 3254.920 ;
        RECT 1593.985 3255.060 1594.275 3255.105 ;
        RECT 1641.825 3255.060 1642.115 3255.105 ;
        RECT 1593.985 3254.920 1642.115 3255.060 ;
        RECT 1593.985 3254.875 1594.275 3254.920 ;
        RECT 1641.825 3254.875 1642.115 3254.920 ;
        RECT 1242.085 3254.380 1242.375 3254.425 ;
        RECT 1269.225 3254.380 1269.515 3254.425 ;
        RECT 1242.085 3254.240 1269.515 3254.380 ;
        RECT 1242.085 3254.195 1242.375 3254.240 ;
        RECT 1269.225 3254.195 1269.515 3254.240 ;
        RECT 1269.685 3254.380 1269.975 3254.425 ;
        RECT 1352.025 3254.380 1352.315 3254.425 ;
        RECT 1365.825 3254.380 1366.115 3254.425 ;
        RECT 1269.685 3254.240 1273.580 3254.380 ;
        RECT 1269.685 3254.195 1269.975 3254.240 ;
        RECT 1273.440 3254.040 1273.580 3254.240 ;
        RECT 1352.025 3254.240 1366.115 3254.380 ;
        RECT 1352.025 3254.195 1352.315 3254.240 ;
        RECT 1365.825 3254.195 1366.115 3254.240 ;
        RECT 1366.285 3254.380 1366.575 3254.425 ;
        RECT 1559.945 3254.380 1560.235 3254.425 ;
        RECT 1593.985 3254.380 1594.275 3254.425 ;
        RECT 1366.285 3254.240 1370.180 3254.380 ;
        RECT 1366.285 3254.195 1366.575 3254.240 ;
        RECT 1304.185 3254.040 1304.475 3254.085 ;
        RECT 1273.440 3253.900 1304.475 3254.040 ;
        RECT 1370.040 3254.040 1370.180 3254.240 ;
        RECT 1462.960 3254.240 1511.400 3254.380 ;
        RECT 1400.785 3254.040 1401.075 3254.085 ;
        RECT 1370.040 3253.900 1401.075 3254.040 ;
        RECT 1304.185 3253.855 1304.475 3253.900 ;
        RECT 1400.785 3253.855 1401.075 3253.900 ;
        RECT 1424.705 3254.040 1424.995 3254.085 ;
        RECT 1462.960 3254.040 1463.100 3254.240 ;
        RECT 1424.705 3253.900 1463.100 3254.040 ;
        RECT 1511.260 3254.040 1511.400 3254.240 ;
        RECT 1559.945 3254.240 1594.275 3254.380 ;
        RECT 1559.945 3254.195 1560.235 3254.240 ;
        RECT 1593.985 3254.195 1594.275 3254.240 ;
        RECT 1559.025 3254.040 1559.315 3254.085 ;
        RECT 1511.260 3253.900 1559.315 3254.040 ;
        RECT 1424.705 3253.855 1424.995 3253.900 ;
        RECT 1559.025 3253.855 1559.315 3253.900 ;
        RECT 1641.825 3254.040 1642.115 3254.085 ;
        RECT 1661.605 3254.040 1661.895 3254.085 ;
        RECT 1641.825 3253.900 1661.895 3254.040 ;
        RECT 1641.825 3253.855 1642.115 3253.900 ;
        RECT 1661.605 3253.855 1661.895 3253.900 ;
        RECT 1242.085 3253.700 1242.375 3253.745 ;
        RECT 1219.160 3253.560 1242.375 3253.700 ;
        RECT 1100.405 3253.515 1100.695 3253.560 ;
        RECT 1124.785 3253.515 1125.075 3253.560 ;
        RECT 1242.085 3253.515 1242.375 3253.560 ;
        RECT 19.850 1386.760 20.170 1386.820 ;
        RECT 161.990 1386.760 162.310 1386.820 ;
        RECT 19.850 1386.620 162.310 1386.760 ;
        RECT 19.850 1386.560 20.170 1386.620 ;
        RECT 161.990 1386.560 162.310 1386.620 ;
      LAYER via ;
        RECT 1661.620 3256.220 1661.880 3256.480 ;
        RECT 162.020 3253.500 162.280 3253.760 ;
        RECT 19.880 1386.560 20.140 1386.820 ;
        RECT 162.020 1386.560 162.280 1386.820 ;
      LAYER met2 ;
        RECT 1663.410 3256.930 1663.690 3260.000 ;
        RECT 1661.680 3256.790 1663.690 3256.930 ;
        RECT 1661.680 3256.510 1661.820 3256.790 ;
        RECT 1661.620 3256.190 1661.880 3256.510 ;
        RECT 1663.410 3256.000 1663.690 3256.790 ;
        RECT 162.020 3253.470 162.280 3253.790 ;
        RECT 162.080 1386.850 162.220 3253.470 ;
        RECT 19.880 1386.530 20.140 1386.850 ;
        RECT 162.020 1386.530 162.280 1386.850 ;
        RECT 19.940 1382.285 20.080 1386.530 ;
        RECT 19.870 1381.915 20.150 1382.285 ;
      LAYER via2 ;
        RECT 19.870 1381.960 20.150 1382.240 ;
      LAYER met3 ;
        RECT -4.800 1382.250 2.400 1382.700 ;
        RECT 19.845 1382.250 20.175 1382.265 ;
        RECT -4.800 1381.950 20.175 1382.250 ;
        RECT -4.800 1381.500 2.400 1381.950 ;
        RECT 19.845 1381.935 20.175 1381.950 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1028.705 3254.735 1028.875 3255.755 ;
        RECT 1028.245 3254.565 1028.875 3254.735 ;
      LAYER mcon ;
        RECT 1028.705 3255.585 1028.875 3255.755 ;
      LAYER met1 ;
        RECT 1118.330 3256.220 1118.650 3256.480 ;
        RECT 1028.645 3255.740 1028.935 3255.785 ;
        RECT 1118.420 3255.740 1118.560 3256.220 ;
        RECT 1028.645 3255.600 1118.560 3255.740 ;
        RECT 1028.645 3255.555 1028.935 3255.600 ;
        RECT 272.390 3254.720 272.710 3254.780 ;
        RECT 1028.185 3254.720 1028.475 3254.765 ;
        RECT 272.390 3254.580 1028.475 3254.720 ;
        RECT 272.390 3254.520 272.710 3254.580 ;
        RECT 1028.185 3254.535 1028.475 3254.580 ;
        RECT 20.310 1131.420 20.630 1131.480 ;
        RECT 272.390 1131.420 272.710 1131.480 ;
        RECT 20.310 1131.280 272.710 1131.420 ;
        RECT 20.310 1131.220 20.630 1131.280 ;
        RECT 272.390 1131.220 272.710 1131.280 ;
      LAYER via ;
        RECT 1118.360 3256.220 1118.620 3256.480 ;
        RECT 272.420 3254.520 272.680 3254.780 ;
        RECT 20.340 1131.220 20.600 1131.480 ;
        RECT 272.420 1131.220 272.680 1131.480 ;
      LAYER met2 ;
        RECT 1119.690 3256.930 1119.970 3260.000 ;
        RECT 1118.420 3256.790 1119.970 3256.930 ;
        RECT 1118.420 3256.510 1118.560 3256.790 ;
        RECT 1118.360 3256.190 1118.620 3256.510 ;
        RECT 1119.690 3256.000 1119.970 3256.790 ;
        RECT 272.420 3254.490 272.680 3254.810 ;
        RECT 272.480 1131.510 272.620 3254.490 ;
        RECT 20.340 1131.365 20.600 1131.510 ;
        RECT 20.330 1130.995 20.610 1131.365 ;
        RECT 272.420 1131.190 272.680 1131.510 ;
      LAYER via2 ;
        RECT 20.330 1131.040 20.610 1131.320 ;
      LAYER met3 ;
        RECT -4.800 1131.330 2.400 1131.780 ;
        RECT 20.305 1131.330 20.635 1131.345 ;
        RECT -4.800 1131.030 20.635 1131.330 ;
        RECT -4.800 1130.580 2.400 1131.030 ;
        RECT 20.305 1131.015 20.635 1131.030 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 79.190 3257.780 79.510 3257.840 ;
        RECT 531.830 3257.780 532.150 3257.840 ;
        RECT 79.190 3257.640 532.150 3257.780 ;
        RECT 79.190 3257.580 79.510 3257.640 ;
        RECT 531.830 3257.580 532.150 3257.640 ;
        RECT 20.310 883.220 20.630 883.280 ;
        RECT 79.190 883.220 79.510 883.280 ;
        RECT 20.310 883.080 79.510 883.220 ;
        RECT 20.310 883.020 20.630 883.080 ;
        RECT 79.190 883.020 79.510 883.080 ;
      LAYER via ;
        RECT 79.220 3257.580 79.480 3257.840 ;
        RECT 531.860 3257.580 532.120 3257.840 ;
        RECT 20.340 883.020 20.600 883.280 ;
        RECT 79.220 883.020 79.480 883.280 ;
      LAYER met2 ;
        RECT 79.220 3257.550 79.480 3257.870 ;
        RECT 531.860 3257.610 532.120 3257.870 ;
        RECT 533.650 3257.610 533.930 3260.000 ;
        RECT 531.860 3257.550 533.930 3257.610 ;
        RECT 79.280 883.310 79.420 3257.550 ;
        RECT 531.920 3257.470 533.930 3257.550 ;
        RECT 533.650 3256.000 533.930 3257.470 ;
        RECT 20.340 882.990 20.600 883.310 ;
        RECT 79.220 882.990 79.480 883.310 ;
        RECT 20.400 879.765 20.540 882.990 ;
        RECT 20.330 879.395 20.610 879.765 ;
      LAYER via2 ;
        RECT 20.330 879.440 20.610 879.720 ;
      LAYER met3 ;
        RECT -4.800 879.730 2.400 880.180 ;
        RECT 20.305 879.730 20.635 879.745 ;
        RECT -4.800 879.430 20.635 879.730 ;
        RECT -4.800 878.980 2.400 879.430 ;
        RECT 20.305 879.415 20.635 879.430 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.330 634.595 20.610 634.965 ;
        RECT 20.400 628.165 20.540 634.595 ;
        RECT 20.330 627.795 20.610 628.165 ;
      LAYER via2 ;
        RECT 20.330 634.640 20.610 634.920 ;
        RECT 20.330 627.840 20.610 628.120 ;
      LAYER met3 ;
        RECT 301.110 1188.450 301.490 1188.460 ;
        RECT 308.470 1188.450 308.850 1188.460 ;
        RECT 301.110 1188.150 308.850 1188.450 ;
        RECT 301.110 1188.140 301.490 1188.150 ;
        RECT 308.470 1188.140 308.850 1188.150 ;
        RECT 156.670 1185.050 157.050 1185.060 ;
        RECT 159.430 1185.050 159.810 1185.060 ;
        RECT 156.670 1184.750 159.810 1185.050 ;
        RECT 156.670 1184.740 157.050 1184.750 ;
        RECT 159.430 1184.740 159.810 1184.750 ;
        RECT 2606.630 1184.740 2607.010 1185.060 ;
        RECT 2606.670 1184.080 2606.970 1184.740 ;
        RECT 2606.000 1183.480 2610.000 1184.080 ;
        RECT 20.305 634.930 20.635 634.945 ;
        RECT 156.670 634.930 157.050 634.940 ;
        RECT 20.305 634.630 157.050 634.930 ;
        RECT 20.305 634.615 20.635 634.630 ;
        RECT 156.670 634.620 157.050 634.630 ;
        RECT -4.800 628.130 2.400 628.580 ;
        RECT 20.305 628.130 20.635 628.145 ;
        RECT -4.800 627.830 20.635 628.130 ;
        RECT -4.800 627.380 2.400 627.830 ;
        RECT 20.305 627.815 20.635 627.830 ;
      LAYER via3 ;
        RECT 301.140 1188.140 301.460 1188.460 ;
        RECT 308.500 1188.140 308.820 1188.460 ;
        RECT 156.700 1184.740 157.020 1185.060 ;
        RECT 159.460 1184.740 159.780 1185.060 ;
        RECT 2606.660 1184.740 2606.980 1185.060 ;
        RECT 156.700 634.620 157.020 634.940 ;
      LAYER met4 ;
        RECT 159.030 1187.710 160.210 1188.890 ;
        RECT 300.710 1187.710 301.890 1188.890 ;
        RECT 308.495 1188.135 308.825 1188.465 ;
        RECT 159.470 1185.065 159.770 1187.710 ;
        RECT 308.510 1185.490 308.810 1188.135 ;
        RECT 156.695 1184.735 157.025 1185.065 ;
        RECT 159.455 1184.735 159.785 1185.065 ;
        RECT 156.710 634.945 157.010 1184.735 ;
        RECT 308.070 1184.310 309.250 1185.490 ;
        RECT 2606.230 1184.310 2607.410 1185.490 ;
        RECT 156.695 634.615 157.025 634.945 ;
      LAYER met5 ;
        RECT 348.340 1190.900 408.820 1192.500 ;
        RECT 158.820 1187.500 302.100 1189.100 ;
        RECT 348.340 1185.700 349.940 1190.900 ;
        RECT 407.220 1189.100 408.820 1190.900 ;
        RECT 516.700 1190.900 566.140 1192.500 ;
        RECT 407.220 1187.500 497.140 1189.100 ;
        RECT 307.860 1184.100 349.940 1185.700 ;
        RECT 495.540 1185.700 497.140 1187.500 ;
        RECT 516.700 1185.700 518.300 1190.900 ;
        RECT 495.540 1184.100 518.300 1185.700 ;
        RECT 564.540 1185.700 566.140 1190.900 ;
        RECT 613.300 1190.900 662.740 1192.500 ;
        RECT 613.300 1185.700 614.900 1190.900 ;
        RECT 564.540 1184.100 614.900 1185.700 ;
        RECT 661.140 1185.700 662.740 1190.900 ;
        RECT 709.900 1190.900 759.340 1192.500 ;
        RECT 709.900 1185.700 711.500 1190.900 ;
        RECT 661.140 1184.100 711.500 1185.700 ;
        RECT 757.740 1185.700 759.340 1190.900 ;
        RECT 806.500 1190.900 855.940 1192.500 ;
        RECT 806.500 1185.700 808.100 1190.900 ;
        RECT 757.740 1184.100 808.100 1185.700 ;
        RECT 854.340 1185.700 855.940 1190.900 ;
        RECT 903.100 1190.900 952.540 1192.500 ;
        RECT 903.100 1185.700 904.700 1190.900 ;
        RECT 854.340 1184.100 904.700 1185.700 ;
        RECT 950.940 1185.700 952.540 1190.900 ;
        RECT 999.700 1190.900 1049.140 1192.500 ;
        RECT 999.700 1185.700 1001.300 1190.900 ;
        RECT 950.940 1184.100 1001.300 1185.700 ;
        RECT 1047.540 1185.700 1049.140 1190.900 ;
        RECT 1096.300 1190.900 1145.740 1192.500 ;
        RECT 1096.300 1185.700 1097.900 1190.900 ;
        RECT 1047.540 1184.100 1097.900 1185.700 ;
        RECT 1144.140 1185.700 1145.740 1190.900 ;
        RECT 1192.900 1190.900 1242.340 1192.500 ;
        RECT 1192.900 1185.700 1194.500 1190.900 ;
        RECT 1144.140 1184.100 1194.500 1185.700 ;
        RECT 1240.740 1185.700 1242.340 1190.900 ;
        RECT 1289.500 1190.900 1338.940 1192.500 ;
        RECT 1289.500 1185.700 1291.100 1190.900 ;
        RECT 1240.740 1184.100 1291.100 1185.700 ;
        RECT 1337.340 1185.700 1338.940 1190.900 ;
        RECT 1386.100 1190.900 1435.540 1192.500 ;
        RECT 1386.100 1185.700 1387.700 1190.900 ;
        RECT 1337.340 1184.100 1387.700 1185.700 ;
        RECT 1433.940 1185.700 1435.540 1190.900 ;
        RECT 1482.700 1190.900 1532.140 1192.500 ;
        RECT 1482.700 1185.700 1484.300 1190.900 ;
        RECT 1433.940 1184.100 1484.300 1185.700 ;
        RECT 1530.540 1185.700 1532.140 1190.900 ;
        RECT 1579.300 1190.900 1628.740 1192.500 ;
        RECT 1579.300 1185.700 1580.900 1190.900 ;
        RECT 1530.540 1184.100 1580.900 1185.700 ;
        RECT 1627.140 1185.700 1628.740 1190.900 ;
        RECT 1675.900 1190.900 1725.340 1192.500 ;
        RECT 1675.900 1185.700 1677.500 1190.900 ;
        RECT 1627.140 1184.100 1677.500 1185.700 ;
        RECT 1723.740 1185.700 1725.340 1190.900 ;
        RECT 1772.500 1190.900 1821.940 1192.500 ;
        RECT 1772.500 1185.700 1774.100 1190.900 ;
        RECT 1723.740 1184.100 1774.100 1185.700 ;
        RECT 1820.340 1185.700 1821.940 1190.900 ;
        RECT 1869.100 1190.900 1918.540 1192.500 ;
        RECT 1869.100 1185.700 1870.700 1190.900 ;
        RECT 1820.340 1184.100 1870.700 1185.700 ;
        RECT 1916.940 1185.700 1918.540 1190.900 ;
        RECT 1965.700 1190.900 2015.140 1192.500 ;
        RECT 1965.700 1185.700 1967.300 1190.900 ;
        RECT 1916.940 1184.100 1967.300 1185.700 ;
        RECT 2013.540 1185.700 2015.140 1190.900 ;
        RECT 2062.300 1190.900 2111.740 1192.500 ;
        RECT 2062.300 1185.700 2063.900 1190.900 ;
        RECT 2013.540 1184.100 2063.900 1185.700 ;
        RECT 2110.140 1185.700 2111.740 1190.900 ;
        RECT 2158.900 1190.900 2208.340 1192.500 ;
        RECT 2158.900 1185.700 2160.500 1190.900 ;
        RECT 2110.140 1184.100 2160.500 1185.700 ;
        RECT 2206.740 1185.700 2208.340 1190.900 ;
        RECT 2255.500 1190.900 2304.940 1192.500 ;
        RECT 2255.500 1185.700 2257.100 1190.900 ;
        RECT 2206.740 1184.100 2257.100 1185.700 ;
        RECT 2303.340 1185.700 2304.940 1190.900 ;
        RECT 2352.100 1190.900 2381.300 1192.500 ;
        RECT 2352.100 1185.700 2353.700 1190.900 ;
        RECT 2379.700 1189.100 2381.300 1190.900 ;
        RECT 2448.700 1190.900 2477.900 1192.500 ;
        RECT 2379.700 1187.500 2429.140 1189.100 ;
        RECT 2303.340 1184.100 2353.700 1185.700 ;
        RECT 2427.540 1185.700 2429.140 1187.500 ;
        RECT 2448.700 1185.700 2450.300 1190.900 ;
        RECT 2476.300 1189.100 2477.900 1190.900 ;
        RECT 2545.300 1190.900 2574.500 1192.500 ;
        RECT 2476.300 1187.500 2525.740 1189.100 ;
        RECT 2427.540 1184.100 2450.300 1185.700 ;
        RECT 2524.140 1185.700 2525.740 1187.500 ;
        RECT 2545.300 1185.700 2546.900 1190.900 ;
        RECT 2524.140 1184.100 2546.900 1185.700 ;
        RECT 2572.900 1185.700 2574.500 1190.900 ;
        RECT 2572.900 1184.100 2607.620 1185.700 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 134.390 1801.220 134.710 1801.280 ;
        RECT 296.770 1801.220 297.090 1801.280 ;
        RECT 134.390 1801.080 297.090 1801.220 ;
        RECT 134.390 1801.020 134.710 1801.080 ;
        RECT 296.770 1801.020 297.090 1801.080 ;
        RECT 17.550 379.340 17.870 379.400 ;
        RECT 134.390 379.340 134.710 379.400 ;
        RECT 17.550 379.200 134.710 379.340 ;
        RECT 17.550 379.140 17.870 379.200 ;
        RECT 134.390 379.140 134.710 379.200 ;
      LAYER via ;
        RECT 134.420 1801.020 134.680 1801.280 ;
        RECT 296.800 1801.020 297.060 1801.280 ;
        RECT 17.580 379.140 17.840 379.400 ;
        RECT 134.420 379.140 134.680 379.400 ;
      LAYER met2 ;
        RECT 296.790 1806.235 297.070 1806.605 ;
        RECT 296.860 1801.310 297.000 1806.235 ;
        RECT 134.420 1800.990 134.680 1801.310 ;
        RECT 296.800 1800.990 297.060 1801.310 ;
        RECT 134.480 379.430 134.620 1800.990 ;
        RECT 17.580 379.110 17.840 379.430 ;
        RECT 134.420 379.110 134.680 379.430 ;
        RECT 17.640 376.565 17.780 379.110 ;
        RECT 17.570 376.195 17.850 376.565 ;
      LAYER via2 ;
        RECT 296.790 1806.280 297.070 1806.560 ;
        RECT 17.570 376.240 17.850 376.520 ;
      LAYER met3 ;
        RECT 296.765 1806.570 297.095 1806.585 ;
        RECT 310.000 1806.570 314.000 1806.960 ;
        RECT 296.765 1806.360 314.000 1806.570 ;
        RECT 296.765 1806.270 310.500 1806.360 ;
        RECT 296.765 1806.255 297.095 1806.270 ;
        RECT -4.800 376.530 2.400 376.980 ;
        RECT 17.545 376.530 17.875 376.545 ;
        RECT -4.800 376.230 17.875 376.530 ;
        RECT -4.800 375.780 2.400 376.230 ;
        RECT 17.545 376.215 17.875 376.230 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 3125.860 2615.490 3125.920 ;
        RECT 2657.950 3125.860 2658.270 3125.920 ;
        RECT 2615.170 3125.720 2658.270 3125.860 ;
        RECT 2615.170 3125.660 2615.490 3125.720 ;
        RECT 2657.950 3125.660 2658.270 3125.720 ;
      LAYER via ;
        RECT 2615.200 3125.660 2615.460 3125.920 ;
        RECT 2657.980 3125.660 2658.240 3125.920 ;
      LAYER met2 ;
        RECT 2615.190 3128.155 2615.470 3128.525 ;
        RECT 2615.260 3125.950 2615.400 3128.155 ;
        RECT 2615.200 3125.630 2615.460 3125.950 ;
        RECT 2657.980 3125.630 2658.240 3125.950 ;
        RECT 2658.040 517.325 2658.180 3125.630 ;
        RECT 2657.970 516.955 2658.250 517.325 ;
        RECT 15.730 130.715 16.010 131.085 ;
        RECT 15.800 125.645 15.940 130.715 ;
        RECT 15.730 125.275 16.010 125.645 ;
      LAYER via2 ;
        RECT 2615.190 3128.200 2615.470 3128.480 ;
        RECT 2657.970 517.000 2658.250 517.280 ;
        RECT 15.730 130.760 16.010 131.040 ;
        RECT 15.730 125.320 16.010 125.600 ;
      LAYER met3 ;
        RECT 2606.000 3128.490 2610.000 3128.880 ;
        RECT 2615.165 3128.490 2615.495 3128.505 ;
        RECT 2606.000 3128.280 2615.495 3128.490 ;
        RECT 2609.580 3128.190 2615.495 3128.280 ;
        RECT 2615.165 3128.175 2615.495 3128.190 ;
        RECT 2657.945 517.300 2658.275 517.305 ;
        RECT 2657.945 517.290 2658.530 517.300 ;
        RECT 2657.720 516.990 2658.530 517.290 ;
        RECT 2657.945 516.980 2658.530 516.990 ;
        RECT 2657.945 516.975 2658.275 516.980 ;
        RECT 15.705 131.050 16.035 131.065 ;
        RECT 2658.150 131.050 2658.530 131.060 ;
        RECT 15.705 130.750 2658.530 131.050 ;
        RECT 15.705 130.735 16.035 130.750 ;
        RECT 2658.150 130.740 2658.530 130.750 ;
        RECT -4.800 125.610 2.400 126.060 ;
        RECT 15.705 125.610 16.035 125.625 ;
        RECT -4.800 125.310 16.035 125.610 ;
        RECT -4.800 124.860 2.400 125.310 ;
        RECT 15.705 125.295 16.035 125.310 ;
      LAYER via3 ;
        RECT 2658.180 516.980 2658.500 517.300 ;
        RECT 2658.180 130.740 2658.500 131.060 ;
      LAYER met4 ;
        RECT 2658.175 516.975 2658.505 517.305 ;
        RECT 2658.190 131.065 2658.490 516.975 ;
        RECT 2658.175 130.735 2658.505 131.065 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1707.130 3256.220 1707.450 3256.480 ;
        RECT 1707.220 3253.700 1707.360 3256.220 ;
        RECT 2790.890 3253.700 2791.210 3253.760 ;
        RECT 1707.220 3253.560 2791.210 3253.700 ;
        RECT 2790.890 3253.500 2791.210 3253.560 ;
        RECT 2790.890 827.800 2791.210 827.860 ;
        RECT 2900.830 827.800 2901.150 827.860 ;
        RECT 2790.890 827.660 2901.150 827.800 ;
        RECT 2790.890 827.600 2791.210 827.660 ;
        RECT 2900.830 827.600 2901.150 827.660 ;
      LAYER via ;
        RECT 1707.160 3256.220 1707.420 3256.480 ;
        RECT 2790.920 3253.500 2791.180 3253.760 ;
        RECT 2790.920 827.600 2791.180 827.860 ;
        RECT 2900.860 827.600 2901.120 827.860 ;
      LAYER met2 ;
        RECT 1705.730 3256.930 1706.010 3260.000 ;
        RECT 1705.730 3256.790 1707.360 3256.930 ;
        RECT 1705.730 3256.000 1706.010 3256.790 ;
        RECT 1707.220 3256.510 1707.360 3256.790 ;
        RECT 1707.160 3256.190 1707.420 3256.510 ;
        RECT 2790.920 3253.470 2791.180 3253.790 ;
        RECT 2790.980 827.890 2791.120 3253.470 ;
        RECT 2790.920 827.570 2791.180 827.890 ;
        RECT 2900.860 827.570 2901.120 827.890 ;
        RECT 2900.920 821.285 2901.060 827.570 ;
        RECT 2900.850 820.915 2901.130 821.285 ;
      LAYER via2 ;
        RECT 2900.850 820.960 2901.130 821.240 ;
      LAYER met3 ;
        RECT 2900.825 821.250 2901.155 821.265 ;
        RECT 2917.600 821.250 2924.800 821.700 ;
        RECT 2900.825 820.950 2924.800 821.250 ;
        RECT 2900.825 820.935 2901.155 820.950 ;
        RECT 2917.600 820.500 2924.800 820.950 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1518.340 2615.490 1518.400 ;
        RECT 2715.450 1518.340 2715.770 1518.400 ;
        RECT 2615.170 1518.200 2715.770 1518.340 ;
        RECT 2615.170 1518.140 2615.490 1518.200 ;
        RECT 2715.450 1518.140 2715.770 1518.200 ;
        RECT 2715.450 1062.400 2715.770 1062.460 ;
        RECT 2900.830 1062.400 2901.150 1062.460 ;
        RECT 2715.450 1062.260 2901.150 1062.400 ;
        RECT 2715.450 1062.200 2715.770 1062.260 ;
        RECT 2900.830 1062.200 2901.150 1062.260 ;
      LAYER via ;
        RECT 2615.200 1518.140 2615.460 1518.400 ;
        RECT 2715.480 1518.140 2715.740 1518.400 ;
        RECT 2715.480 1062.200 2715.740 1062.460 ;
        RECT 2900.860 1062.200 2901.120 1062.460 ;
      LAYER met2 ;
        RECT 2615.190 1521.995 2615.470 1522.365 ;
        RECT 2615.260 1518.430 2615.400 1521.995 ;
        RECT 2615.200 1518.110 2615.460 1518.430 ;
        RECT 2715.480 1518.110 2715.740 1518.430 ;
        RECT 2715.540 1062.490 2715.680 1518.110 ;
        RECT 2715.480 1062.170 2715.740 1062.490 ;
        RECT 2900.860 1062.170 2901.120 1062.490 ;
        RECT 2900.920 1055.885 2901.060 1062.170 ;
        RECT 2900.850 1055.515 2901.130 1055.885 ;
      LAYER via2 ;
        RECT 2615.190 1522.040 2615.470 1522.320 ;
        RECT 2900.850 1055.560 2901.130 1055.840 ;
      LAYER met3 ;
        RECT 2606.000 1522.330 2610.000 1522.720 ;
        RECT 2615.165 1522.330 2615.495 1522.345 ;
        RECT 2606.000 1522.120 2615.495 1522.330 ;
        RECT 2609.580 1522.030 2615.495 1522.120 ;
        RECT 2615.165 1522.015 2615.495 1522.030 ;
        RECT 2900.825 1055.850 2901.155 1055.865 ;
        RECT 2917.600 1055.850 2924.800 1056.300 ;
        RECT 2900.825 1055.550 2924.800 1055.850 ;
        RECT 2900.825 1055.535 2901.155 1055.550 ;
        RECT 2917.600 1055.100 2924.800 1055.550 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 310.000 1679.880 314.000 1680.480 ;
        RECT 309.390 1677.370 309.770 1677.380 ;
        RECT 310.350 1677.370 310.650 1679.880 ;
        RECT 309.390 1677.070 310.650 1677.370 ;
        RECT 309.390 1677.060 309.770 1677.070 ;
        RECT 2620.430 1671.250 2620.810 1671.260 ;
        RECT 2654.470 1671.250 2654.850 1671.260 ;
        RECT 2620.430 1670.950 2654.850 1671.250 ;
        RECT 2620.430 1670.940 2620.810 1670.950 ;
        RECT 2654.470 1670.940 2654.850 1670.950 ;
        RECT 2660.910 1290.450 2661.290 1290.460 ;
        RECT 2917.600 1290.450 2924.800 1290.900 ;
        RECT 2660.910 1290.150 2924.800 1290.450 ;
        RECT 2660.910 1290.140 2661.290 1290.150 ;
        RECT 2917.600 1289.700 2924.800 1290.150 ;
      LAYER via3 ;
        RECT 309.420 1677.060 309.740 1677.380 ;
        RECT 2620.460 1670.940 2620.780 1671.260 ;
        RECT 2654.500 1670.940 2654.820 1671.260 ;
        RECT 2660.940 1290.140 2661.260 1290.460 ;
      LAYER met4 ;
        RECT 309.415 1677.055 309.745 1677.385 ;
        RECT 309.430 1675.090 309.730 1677.055 ;
        RECT 308.990 1673.910 310.170 1675.090 ;
        RECT 2620.030 1673.910 2621.210 1675.090 ;
        RECT 2660.510 1673.910 2661.690 1675.090 ;
        RECT 2620.470 1671.265 2620.770 1673.910 ;
        RECT 2620.455 1670.935 2620.785 1671.265 ;
        RECT 2654.070 1670.510 2655.250 1671.690 ;
        RECT 2660.950 1290.465 2661.250 1673.910 ;
        RECT 2660.935 1290.135 2661.265 1290.465 ;
      LAYER met5 ;
        RECT 361.220 1677.100 366.500 1678.700 ;
        RECT 361.220 1675.300 362.820 1677.100 ;
        RECT 308.780 1673.700 362.820 1675.300 ;
        RECT 364.900 1675.300 366.500 1677.100 ;
        RECT 446.780 1677.100 498.060 1678.700 ;
        RECT 364.900 1673.700 369.260 1675.300 ;
        RECT 367.660 1671.900 369.260 1673.700 ;
        RECT 446.780 1671.900 448.380 1677.100 ;
        RECT 367.660 1670.300 448.380 1671.900 ;
        RECT 496.460 1671.900 498.060 1677.100 ;
        RECT 543.380 1677.100 594.660 1678.700 ;
        RECT 543.380 1671.900 544.980 1677.100 ;
        RECT 593.060 1675.300 594.660 1677.100 ;
        RECT 2558.180 1677.100 2609.460 1678.700 ;
        RECT 593.060 1673.700 641.580 1675.300 ;
        RECT 496.460 1670.300 544.980 1671.900 ;
        RECT 639.980 1671.900 641.580 1673.700 ;
        RECT 690.580 1673.700 738.180 1675.300 ;
        RECT 690.580 1671.900 692.180 1673.700 ;
        RECT 639.980 1670.300 692.180 1671.900 ;
        RECT 736.580 1671.900 738.180 1673.700 ;
        RECT 787.180 1673.700 834.780 1675.300 ;
        RECT 787.180 1671.900 788.780 1673.700 ;
        RECT 736.580 1670.300 788.780 1671.900 ;
        RECT 833.180 1671.900 834.780 1673.700 ;
        RECT 883.780 1673.700 931.380 1675.300 ;
        RECT 883.780 1671.900 885.380 1673.700 ;
        RECT 833.180 1670.300 885.380 1671.900 ;
        RECT 929.780 1671.900 931.380 1673.700 ;
        RECT 980.380 1673.700 1027.980 1675.300 ;
        RECT 980.380 1671.900 981.980 1673.700 ;
        RECT 929.780 1670.300 981.980 1671.900 ;
        RECT 1026.380 1671.900 1027.980 1673.700 ;
        RECT 1076.980 1673.700 1124.580 1675.300 ;
        RECT 1076.980 1671.900 1078.580 1673.700 ;
        RECT 1026.380 1670.300 1078.580 1671.900 ;
        RECT 1122.980 1671.900 1124.580 1673.700 ;
        RECT 1173.580 1673.700 1221.180 1675.300 ;
        RECT 1173.580 1671.900 1175.180 1673.700 ;
        RECT 1122.980 1670.300 1175.180 1671.900 ;
        RECT 1219.580 1671.900 1221.180 1673.700 ;
        RECT 1270.180 1673.700 1317.780 1675.300 ;
        RECT 1270.180 1671.900 1271.780 1673.700 ;
        RECT 1219.580 1670.300 1271.780 1671.900 ;
        RECT 1316.180 1671.900 1317.780 1673.700 ;
        RECT 1366.780 1673.700 1414.380 1675.300 ;
        RECT 1366.780 1671.900 1368.380 1673.700 ;
        RECT 1316.180 1670.300 1368.380 1671.900 ;
        RECT 1412.780 1671.900 1414.380 1673.700 ;
        RECT 1463.380 1673.700 1510.980 1675.300 ;
        RECT 1463.380 1671.900 1464.980 1673.700 ;
        RECT 1412.780 1670.300 1464.980 1671.900 ;
        RECT 1509.380 1671.900 1510.980 1673.700 ;
        RECT 1559.980 1673.700 1607.580 1675.300 ;
        RECT 1559.980 1671.900 1561.580 1673.700 ;
        RECT 1509.380 1670.300 1561.580 1671.900 ;
        RECT 1605.980 1671.900 1607.580 1673.700 ;
        RECT 1656.580 1673.700 1704.180 1675.300 ;
        RECT 1656.580 1671.900 1658.180 1673.700 ;
        RECT 1605.980 1670.300 1658.180 1671.900 ;
        RECT 1702.580 1671.900 1704.180 1673.700 ;
        RECT 1753.180 1673.700 1800.780 1675.300 ;
        RECT 1753.180 1671.900 1754.780 1673.700 ;
        RECT 1702.580 1670.300 1754.780 1671.900 ;
        RECT 1799.180 1671.900 1800.780 1673.700 ;
        RECT 1849.780 1673.700 1897.380 1675.300 ;
        RECT 1849.780 1671.900 1851.380 1673.700 ;
        RECT 1799.180 1670.300 1851.380 1671.900 ;
        RECT 1895.780 1671.900 1897.380 1673.700 ;
        RECT 1946.380 1673.700 1993.980 1675.300 ;
        RECT 1946.380 1671.900 1947.980 1673.700 ;
        RECT 1895.780 1670.300 1947.980 1671.900 ;
        RECT 1992.380 1671.900 1993.980 1673.700 ;
        RECT 2042.980 1673.700 2090.580 1675.300 ;
        RECT 2042.980 1671.900 2044.580 1673.700 ;
        RECT 1992.380 1670.300 2044.580 1671.900 ;
        RECT 2088.980 1671.900 2090.580 1673.700 ;
        RECT 2139.580 1673.700 2187.180 1675.300 ;
        RECT 2139.580 1671.900 2141.180 1673.700 ;
        RECT 2088.980 1670.300 2141.180 1671.900 ;
        RECT 2185.580 1671.900 2187.180 1673.700 ;
        RECT 2236.180 1673.700 2283.780 1675.300 ;
        RECT 2236.180 1671.900 2237.780 1673.700 ;
        RECT 2185.580 1670.300 2237.780 1671.900 ;
        RECT 2282.180 1671.900 2283.780 1673.700 ;
        RECT 2332.780 1673.700 2380.380 1675.300 ;
        RECT 2332.780 1671.900 2334.380 1673.700 ;
        RECT 2282.180 1670.300 2334.380 1671.900 ;
        RECT 2378.780 1671.900 2380.380 1673.700 ;
        RECT 2429.380 1673.700 2476.980 1675.300 ;
        RECT 2429.380 1671.900 2430.980 1673.700 ;
        RECT 2378.780 1670.300 2430.980 1671.900 ;
        RECT 2475.380 1671.900 2476.980 1673.700 ;
        RECT 2558.180 1671.900 2559.780 1677.100 ;
        RECT 2607.860 1675.300 2609.460 1677.100 ;
        RECT 2607.860 1673.700 2621.420 1675.300 ;
        RECT 2654.780 1673.700 2661.900 1675.300 ;
        RECT 2654.780 1672.580 2656.380 1673.700 ;
        RECT 2475.380 1670.300 2559.780 1671.900 ;
        RECT 2653.860 1670.980 2656.380 1672.580 ;
        RECT 2653.860 1670.300 2655.460 1670.980 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2149.190 3264.240 2149.510 3264.300 ;
        RECT 2652.890 3264.240 2653.210 3264.300 ;
        RECT 2149.190 3264.100 2653.210 3264.240 ;
        RECT 2149.190 3264.040 2149.510 3264.100 ;
        RECT 2652.890 3264.040 2653.210 3264.100 ;
        RECT 2652.890 1531.600 2653.210 1531.660 ;
        RECT 2900.830 1531.600 2901.150 1531.660 ;
        RECT 2652.890 1531.460 2901.150 1531.600 ;
        RECT 2652.890 1531.400 2653.210 1531.460 ;
        RECT 2900.830 1531.400 2901.150 1531.460 ;
      LAYER via ;
        RECT 2149.220 3264.040 2149.480 3264.300 ;
        RECT 2652.920 3264.040 2653.180 3264.300 ;
        RECT 2652.920 1531.400 2653.180 1531.660 ;
        RECT 2900.860 1531.400 2901.120 1531.660 ;
      LAYER met2 ;
        RECT 2149.220 3264.010 2149.480 3264.330 ;
        RECT 2652.920 3264.010 2653.180 3264.330 ;
        RECT 2149.280 3260.000 2149.420 3264.010 ;
        RECT 2149.170 3256.000 2149.450 3260.000 ;
        RECT 2652.980 1531.690 2653.120 3264.010 ;
        RECT 2652.920 1531.370 2653.180 1531.690 ;
        RECT 2900.860 1531.370 2901.120 1531.690 ;
        RECT 2900.920 1525.085 2901.060 1531.370 ;
        RECT 2900.850 1524.715 2901.130 1525.085 ;
      LAYER via2 ;
        RECT 2900.850 1524.760 2901.130 1525.040 ;
      LAYER met3 ;
        RECT 2900.825 1525.050 2901.155 1525.065 ;
        RECT 2917.600 1525.050 2924.800 1525.500 ;
        RECT 2900.825 1524.750 2924.800 1525.050 ;
        RECT 2900.825 1524.735 2901.155 1524.750 ;
        RECT 2917.600 1524.300 2924.800 1524.750 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2653.350 1759.740 2653.670 1759.800 ;
        RECT 2900.830 1759.740 2901.150 1759.800 ;
        RECT 2653.350 1759.600 2901.150 1759.740 ;
        RECT 2653.350 1759.540 2653.670 1759.600 ;
        RECT 2900.830 1759.540 2901.150 1759.600 ;
        RECT 955.950 254.560 956.270 254.620 ;
        RECT 2653.350 254.560 2653.670 254.620 ;
        RECT 955.950 254.420 2653.670 254.560 ;
        RECT 955.950 254.360 956.270 254.420 ;
        RECT 2653.350 254.360 2653.670 254.420 ;
      LAYER via ;
        RECT 2653.380 1759.540 2653.640 1759.800 ;
        RECT 2900.860 1759.540 2901.120 1759.800 ;
        RECT 955.980 254.360 956.240 254.620 ;
        RECT 2653.380 254.360 2653.640 254.620 ;
      LAYER met2 ;
        RECT 2653.380 1759.510 2653.640 1759.830 ;
        RECT 2900.860 1759.685 2901.120 1759.830 ;
        RECT 955.930 260.000 956.210 264.000 ;
        RECT 956.040 254.650 956.180 260.000 ;
        RECT 2653.440 254.650 2653.580 1759.510 ;
        RECT 2900.850 1759.315 2901.130 1759.685 ;
        RECT 955.980 254.330 956.240 254.650 ;
        RECT 2653.380 254.330 2653.640 254.650 ;
      LAYER via2 ;
        RECT 2900.850 1759.360 2901.130 1759.640 ;
      LAYER met3 ;
        RECT 2900.825 1759.650 2901.155 1759.665 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2900.825 1759.350 2924.800 1759.650 ;
        RECT 2900.825 1759.335 2901.155 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2729.250 1994.340 2729.570 1994.400 ;
        RECT 2900.830 1994.340 2901.150 1994.400 ;
        RECT 2729.250 1994.200 2901.150 1994.340 ;
        RECT 2729.250 1994.140 2729.570 1994.200 ;
        RECT 2900.830 1994.140 2901.150 1994.200 ;
        RECT 1727.830 248.440 1728.150 248.500 ;
        RECT 2729.250 248.440 2729.570 248.500 ;
        RECT 1727.830 248.300 2729.570 248.440 ;
        RECT 1727.830 248.240 1728.150 248.300 ;
        RECT 2729.250 248.240 2729.570 248.300 ;
      LAYER via ;
        RECT 2729.280 1994.140 2729.540 1994.400 ;
        RECT 2900.860 1994.140 2901.120 1994.400 ;
        RECT 1727.860 248.240 1728.120 248.500 ;
        RECT 2729.280 248.240 2729.540 248.500 ;
      LAYER met2 ;
        RECT 2729.280 1994.110 2729.540 1994.430 ;
        RECT 2900.860 1994.285 2901.120 1994.430 ;
        RECT 1727.810 260.000 1728.090 264.000 ;
        RECT 1727.920 248.530 1728.060 260.000 ;
        RECT 2729.340 248.530 2729.480 1994.110 ;
        RECT 2900.850 1993.915 2901.130 1994.285 ;
        RECT 1727.860 248.210 1728.120 248.530 ;
        RECT 2729.280 248.210 2729.540 248.530 ;
      LAYER via2 ;
        RECT 2900.850 1993.960 2901.130 1994.240 ;
      LAYER met3 ;
        RECT 2900.825 1994.250 2901.155 1994.265 ;
        RECT 2917.600 1994.250 2924.800 1994.700 ;
        RECT 2900.825 1993.950 2924.800 1994.250 ;
        RECT 2900.825 1993.935 2901.155 1993.950 ;
        RECT 2917.600 1993.500 2924.800 1993.950 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 404.870 3278.180 405.190 3278.240 ;
        RECT 2687.850 3278.180 2688.170 3278.240 ;
        RECT 404.870 3278.040 2688.170 3278.180 ;
        RECT 404.870 3277.980 405.190 3278.040 ;
        RECT 2687.850 3277.980 2688.170 3278.040 ;
        RECT 2687.850 2235.400 2688.170 2235.460 ;
        RECT 2900.830 2235.400 2901.150 2235.460 ;
        RECT 2687.850 2235.260 2901.150 2235.400 ;
        RECT 2687.850 2235.200 2688.170 2235.260 ;
        RECT 2900.830 2235.200 2901.150 2235.260 ;
      LAYER via ;
        RECT 404.900 3277.980 405.160 3278.240 ;
        RECT 2687.880 3277.980 2688.140 3278.240 ;
        RECT 2687.880 2235.200 2688.140 2235.460 ;
        RECT 2900.860 2235.200 2901.120 2235.460 ;
      LAYER met2 ;
        RECT 404.900 3277.950 405.160 3278.270 ;
        RECT 2687.880 3277.950 2688.140 3278.270 ;
        RECT 404.960 3260.000 405.100 3277.950 ;
        RECT 404.850 3256.000 405.130 3260.000 ;
        RECT 2687.940 2235.490 2688.080 3277.950 ;
        RECT 2687.880 2235.170 2688.140 2235.490 ;
        RECT 2900.860 2235.170 2901.120 2235.490 ;
        RECT 2900.920 2228.885 2901.060 2235.170 ;
        RECT 2900.850 2228.515 2901.130 2228.885 ;
      LAYER via2 ;
        RECT 2900.850 2228.560 2901.130 2228.840 ;
      LAYER met3 ;
        RECT 2900.825 2228.850 2901.155 2228.865 ;
        RECT 2917.600 2228.850 2924.800 2229.300 ;
        RECT 2900.825 2228.550 2924.800 2228.850 ;
        RECT 2900.825 2228.535 2901.155 2228.550 ;
        RECT 2917.600 2228.100 2924.800 2228.550 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 633.105 48.365 633.275 66.555 ;
      LAYER mcon ;
        RECT 633.105 66.385 633.275 66.555 ;
      LAYER met1 ;
        RECT 633.045 66.540 633.335 66.585 ;
        RECT 1538.770 66.540 1539.090 66.600 ;
        RECT 633.045 66.400 1539.090 66.540 ;
        RECT 633.045 66.355 633.335 66.400 ;
        RECT 1538.770 66.340 1539.090 66.400 ;
        RECT 633.030 48.520 633.350 48.580 ;
        RECT 632.835 48.380 633.350 48.520 ;
        RECT 633.030 48.320 633.350 48.380 ;
      LAYER via ;
        RECT 1538.800 66.340 1539.060 66.600 ;
        RECT 633.060 48.320 633.320 48.580 ;
      LAYER met2 ;
        RECT 1541.970 260.170 1542.250 264.000 ;
        RECT 1538.860 260.030 1542.250 260.170 ;
        RECT 1538.860 66.630 1539.000 260.030 ;
        RECT 1541.970 260.000 1542.250 260.030 ;
        RECT 1538.800 66.310 1539.060 66.630 ;
        RECT 633.060 48.290 633.320 48.610 ;
        RECT 633.120 2.400 633.260 48.290 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2448.725 257.465 2448.895 261.375 ;
        RECT 2497.945 257.805 2498.115 261.375 ;
        RECT 2545.785 257.975 2545.955 261.375 ;
        RECT 2545.325 257.805 2545.955 257.975 ;
      LAYER mcon ;
        RECT 2448.725 261.205 2448.895 261.375 ;
        RECT 2497.945 261.205 2498.115 261.375 ;
        RECT 2545.785 261.205 2545.955 261.375 ;
      LAYER met1 ;
        RECT 2615.170 986.920 2615.490 986.980 ;
        RECT 2652.890 986.920 2653.210 986.980 ;
        RECT 2615.170 986.780 2653.210 986.920 ;
        RECT 2615.170 986.720 2615.490 986.780 ;
        RECT 2652.890 986.720 2653.210 986.780 ;
        RECT 2652.890 261.700 2653.210 261.760 ;
        RECT 2597.780 261.560 2653.210 261.700 ;
        RECT 2448.665 261.360 2448.955 261.405 ;
        RECT 2497.885 261.360 2498.175 261.405 ;
        RECT 2448.665 261.220 2498.175 261.360 ;
        RECT 2448.665 261.175 2448.955 261.220 ;
        RECT 2497.885 261.175 2498.175 261.220 ;
        RECT 2545.725 261.360 2546.015 261.405 ;
        RECT 2597.780 261.360 2597.920 261.560 ;
        RECT 2652.890 261.500 2653.210 261.560 ;
        RECT 2545.725 261.220 2597.920 261.360 ;
        RECT 2545.725 261.175 2546.015 261.220 ;
        RECT 2497.885 257.960 2498.175 258.005 ;
        RECT 2545.265 257.960 2545.555 258.005 ;
        RECT 2497.885 257.820 2545.555 257.960 ;
        RECT 2497.885 257.775 2498.175 257.820 ;
        RECT 2545.265 257.775 2545.555 257.820 ;
        RECT 2421.510 257.620 2421.830 257.680 ;
        RECT 2448.665 257.620 2448.955 257.665 ;
        RECT 2421.510 257.480 2448.955 257.620 ;
        RECT 2421.510 257.420 2421.830 257.480 ;
        RECT 2448.665 257.435 2448.955 257.480 ;
        RECT 2417.370 17.920 2417.690 17.980 ;
        RECT 2421.510 17.920 2421.830 17.980 ;
        RECT 2417.370 17.780 2421.830 17.920 ;
        RECT 2417.370 17.720 2417.690 17.780 ;
        RECT 2421.510 17.720 2421.830 17.780 ;
      LAYER via ;
        RECT 2615.200 986.720 2615.460 986.980 ;
        RECT 2652.920 986.720 2653.180 986.980 ;
        RECT 2652.920 261.500 2653.180 261.760 ;
        RECT 2421.540 257.420 2421.800 257.680 ;
        RECT 2417.400 17.720 2417.660 17.980 ;
        RECT 2421.540 17.720 2421.800 17.980 ;
      LAYER met2 ;
        RECT 2615.190 992.955 2615.470 993.325 ;
        RECT 2615.260 987.010 2615.400 992.955 ;
        RECT 2615.200 986.690 2615.460 987.010 ;
        RECT 2652.920 986.690 2653.180 987.010 ;
        RECT 2652.980 261.790 2653.120 986.690 ;
        RECT 2652.920 261.470 2653.180 261.790 ;
        RECT 2421.540 257.390 2421.800 257.710 ;
        RECT 2421.600 18.010 2421.740 257.390 ;
        RECT 2417.400 17.690 2417.660 18.010 ;
        RECT 2421.540 17.690 2421.800 18.010 ;
        RECT 2417.460 2.400 2417.600 17.690 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
      LAYER via2 ;
        RECT 2615.190 993.000 2615.470 993.280 ;
      LAYER met3 ;
        RECT 2606.000 993.290 2610.000 993.680 ;
        RECT 2615.165 993.290 2615.495 993.305 ;
        RECT 2606.000 993.080 2615.495 993.290 ;
        RECT 2609.580 992.990 2615.495 993.080 ;
        RECT 2615.165 992.975 2615.495 992.990 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2449.185 257.805 2449.355 261.715 ;
        RECT 2498.405 257.125 2498.575 261.715 ;
        RECT 2545.325 258.315 2545.495 261.715 ;
        RECT 2597.305 261.545 2598.395 261.715 ;
        RECT 2598.225 261.205 2598.395 261.545 ;
        RECT 2544.865 258.145 2545.495 258.315 ;
        RECT 2544.865 257.125 2545.035 258.145 ;
      LAYER mcon ;
        RECT 2449.185 261.545 2449.355 261.715 ;
        RECT 2498.405 261.545 2498.575 261.715 ;
        RECT 2545.325 261.545 2545.495 261.715 ;
      LAYER met1 ;
        RECT 2615.170 586.740 2615.490 586.800 ;
        RECT 2645.530 586.740 2645.850 586.800 ;
        RECT 2615.170 586.600 2645.850 586.740 ;
        RECT 2615.170 586.540 2615.490 586.600 ;
        RECT 2645.530 586.540 2645.850 586.600 ;
        RECT 2449.125 261.700 2449.415 261.745 ;
        RECT 2498.345 261.700 2498.635 261.745 ;
        RECT 2449.125 261.560 2498.635 261.700 ;
        RECT 2449.125 261.515 2449.415 261.560 ;
        RECT 2498.345 261.515 2498.635 261.560 ;
        RECT 2545.265 261.700 2545.555 261.745 ;
        RECT 2597.245 261.700 2597.535 261.745 ;
        RECT 2545.265 261.560 2597.535 261.700 ;
        RECT 2545.265 261.515 2545.555 261.560 ;
        RECT 2597.245 261.515 2597.535 261.560 ;
        RECT 2598.165 261.360 2598.455 261.405 ;
        RECT 2645.530 261.360 2645.850 261.420 ;
        RECT 2598.165 261.220 2645.850 261.360 ;
        RECT 2598.165 261.175 2598.455 261.220 ;
        RECT 2645.530 261.160 2645.850 261.220 ;
        RECT 2435.310 257.960 2435.630 258.020 ;
        RECT 2449.125 257.960 2449.415 258.005 ;
        RECT 2435.310 257.820 2449.415 257.960 ;
        RECT 2435.310 257.760 2435.630 257.820 ;
        RECT 2449.125 257.775 2449.415 257.820 ;
        RECT 2498.345 257.280 2498.635 257.325 ;
        RECT 2544.805 257.280 2545.095 257.325 ;
        RECT 2498.345 257.140 2545.095 257.280 ;
        RECT 2498.345 257.095 2498.635 257.140 ;
        RECT 2544.805 257.095 2545.095 257.140 ;
      LAYER via ;
        RECT 2615.200 586.540 2615.460 586.800 ;
        RECT 2645.560 586.540 2645.820 586.800 ;
        RECT 2645.560 261.160 2645.820 261.420 ;
        RECT 2435.340 257.760 2435.600 258.020 ;
      LAYER met2 ;
        RECT 2615.190 591.755 2615.470 592.125 ;
        RECT 2615.260 586.830 2615.400 591.755 ;
        RECT 2615.200 586.510 2615.460 586.830 ;
        RECT 2645.560 586.510 2645.820 586.830 ;
        RECT 2645.620 261.450 2645.760 586.510 ;
        RECT 2645.560 261.130 2645.820 261.450 ;
        RECT 2435.340 257.730 2435.600 258.050 ;
        RECT 2435.400 19.450 2435.540 257.730 ;
        RECT 2434.940 19.310 2435.540 19.450 ;
        RECT 2434.940 2.400 2435.080 19.310 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
      LAYER via2 ;
        RECT 2615.190 591.800 2615.470 592.080 ;
      LAYER met3 ;
        RECT 2606.000 592.090 2610.000 592.480 ;
        RECT 2615.165 592.090 2615.495 592.105 ;
        RECT 2606.000 591.880 2615.495 592.090 ;
        RECT 2609.580 591.790 2615.495 591.880 ;
        RECT 2615.165 591.775 2615.495 591.790 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.810 3258.970 877.090 3260.000 ;
        RECT 878.230 3258.970 878.510 3259.085 ;
        RECT 876.810 3258.830 878.510 3258.970 ;
        RECT 876.810 3256.000 877.090 3258.830 ;
        RECT 878.230 3258.715 878.510 3258.830 ;
        RECT 2452.810 15.115 2453.090 15.485 ;
        RECT 2452.880 2.400 2453.020 15.115 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
      LAYER via2 ;
        RECT 878.230 3258.760 878.510 3259.040 ;
        RECT 2452.810 15.160 2453.090 15.440 ;
      LAYER met3 ;
        RECT 878.205 3259.050 878.535 3259.065 ;
        RECT 2636.070 3259.050 2636.450 3259.060 ;
        RECT 878.205 3258.750 2636.450 3259.050 ;
        RECT 878.205 3258.735 878.535 3258.750 ;
        RECT 2636.070 3258.740 2636.450 3258.750 ;
        RECT 2452.785 15.450 2453.115 15.465 ;
        RECT 2455.750 15.450 2456.130 15.460 ;
        RECT 2452.785 15.150 2456.130 15.450 ;
        RECT 2452.785 15.135 2453.115 15.150 ;
        RECT 2455.750 15.140 2456.130 15.150 ;
      LAYER via3 ;
        RECT 2636.100 3258.740 2636.420 3259.060 ;
        RECT 2455.780 15.140 2456.100 15.460 ;
      LAYER met4 ;
        RECT 2636.095 3258.735 2636.425 3259.065 ;
        RECT 2636.110 19.290 2636.410 3258.735 ;
        RECT 2455.350 18.110 2456.530 19.290 ;
        RECT 2635.670 18.110 2636.850 19.290 ;
        RECT 2455.790 15.465 2456.090 18.110 ;
        RECT 2455.775 15.135 2456.105 15.465 ;
      LAYER met5 ;
        RECT 2455.140 17.900 2637.060 19.500 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2511.745 20.145 2511.915 21.335 ;
        RECT 2546.245 20.485 2546.415 21.335 ;
        RECT 2589.025 17.765 2589.195 19.975 ;
        RECT 2597.305 19.805 2598.395 19.975 ;
        RECT 2597.305 17.765 2597.475 19.805 ;
        RECT 2598.225 19.465 2598.395 19.805 ;
        RECT 2607.885 19.465 2608.055 20.655 ;
        RECT 2624.905 18.445 2625.075 20.655 ;
      LAYER mcon ;
        RECT 2511.745 21.165 2511.915 21.335 ;
        RECT 2546.245 21.165 2546.415 21.335 ;
        RECT 2607.885 20.485 2608.055 20.655 ;
        RECT 2589.025 19.805 2589.195 19.975 ;
        RECT 2624.905 20.485 2625.075 20.655 ;
      LAYER met1 ;
        RECT 2277.990 3274.100 2278.310 3274.160 ;
        RECT 2636.330 3274.100 2636.650 3274.160 ;
        RECT 2277.990 3273.960 2636.650 3274.100 ;
        RECT 2277.990 3273.900 2278.310 3273.960 ;
        RECT 2636.330 3273.900 2636.650 3273.960 ;
        RECT 2511.685 21.320 2511.975 21.365 ;
        RECT 2546.185 21.320 2546.475 21.365 ;
        RECT 2511.685 21.180 2546.475 21.320 ;
        RECT 2511.685 21.135 2511.975 21.180 ;
        RECT 2546.185 21.135 2546.475 21.180 ;
        RECT 2546.185 20.640 2546.475 20.685 ;
        RECT 2607.825 20.640 2608.115 20.685 ;
        RECT 2624.845 20.640 2625.135 20.685 ;
        RECT 2546.185 20.500 2563.880 20.640 ;
        RECT 2546.185 20.455 2546.475 20.500 ;
        RECT 2470.730 20.300 2471.050 20.360 ;
        RECT 2511.685 20.300 2511.975 20.345 ;
        RECT 2470.730 20.160 2511.975 20.300 ;
        RECT 2470.730 20.100 2471.050 20.160 ;
        RECT 2511.685 20.115 2511.975 20.160 ;
        RECT 2563.740 19.960 2563.880 20.500 ;
        RECT 2607.825 20.500 2625.135 20.640 ;
        RECT 2607.825 20.455 2608.115 20.500 ;
        RECT 2624.845 20.455 2625.135 20.500 ;
        RECT 2588.965 19.960 2589.255 20.005 ;
        RECT 2563.740 19.820 2589.255 19.960 ;
        RECT 2588.965 19.775 2589.255 19.820 ;
        RECT 2598.165 19.620 2598.455 19.665 ;
        RECT 2607.825 19.620 2608.115 19.665 ;
        RECT 2598.165 19.480 2608.115 19.620 ;
        RECT 2598.165 19.435 2598.455 19.480 ;
        RECT 2607.825 19.435 2608.115 19.480 ;
        RECT 2624.845 18.600 2625.135 18.645 ;
        RECT 2636.330 18.600 2636.650 18.660 ;
        RECT 2624.845 18.460 2636.650 18.600 ;
        RECT 2624.845 18.415 2625.135 18.460 ;
        RECT 2636.330 18.400 2636.650 18.460 ;
        RECT 2588.965 17.920 2589.255 17.965 ;
        RECT 2597.245 17.920 2597.535 17.965 ;
        RECT 2588.965 17.780 2597.535 17.920 ;
        RECT 2588.965 17.735 2589.255 17.780 ;
        RECT 2597.245 17.735 2597.535 17.780 ;
      LAYER via ;
        RECT 2278.020 3273.900 2278.280 3274.160 ;
        RECT 2636.360 3273.900 2636.620 3274.160 ;
        RECT 2470.760 20.100 2471.020 20.360 ;
        RECT 2636.360 18.400 2636.620 18.660 ;
      LAYER met2 ;
        RECT 2278.020 3273.870 2278.280 3274.190 ;
        RECT 2636.360 3273.870 2636.620 3274.190 ;
        RECT 2278.080 3260.000 2278.220 3273.870 ;
        RECT 2277.970 3256.000 2278.250 3260.000 ;
        RECT 2470.760 20.070 2471.020 20.390 ;
        RECT 2470.820 2.400 2470.960 20.070 ;
        RECT 2636.420 18.690 2636.560 3273.870 ;
        RECT 2636.360 18.370 2636.620 18.690 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2597.765 17.765 2597.935 19.635 ;
      LAYER mcon ;
        RECT 2597.765 19.465 2597.935 19.635 ;
      LAYER met1 ;
        RECT 1748.990 3273.080 1749.310 3273.140 ;
        RECT 2649.670 3273.080 2649.990 3273.140 ;
        RECT 1748.990 3272.940 2649.990 3273.080 ;
        RECT 1748.990 3272.880 1749.310 3272.940 ;
        RECT 2649.670 3272.880 2649.990 3272.940 ;
        RECT 2488.670 19.620 2488.990 19.680 ;
        RECT 2597.705 19.620 2597.995 19.665 ;
        RECT 2488.670 19.480 2597.995 19.620 ;
        RECT 2488.670 19.420 2488.990 19.480 ;
        RECT 2597.705 19.435 2597.995 19.480 ;
        RECT 2597.705 17.920 2597.995 17.965 ;
        RECT 2649.670 17.920 2649.990 17.980 ;
        RECT 2597.705 17.780 2649.990 17.920 ;
        RECT 2597.705 17.735 2597.995 17.780 ;
        RECT 2649.670 17.720 2649.990 17.780 ;
      LAYER via ;
        RECT 1749.020 3272.880 1749.280 3273.140 ;
        RECT 2649.700 3272.880 2649.960 3273.140 ;
        RECT 2488.700 19.420 2488.960 19.680 ;
        RECT 2649.700 17.720 2649.960 17.980 ;
      LAYER met2 ;
        RECT 1749.020 3272.850 1749.280 3273.170 ;
        RECT 2649.700 3272.850 2649.960 3273.170 ;
        RECT 1749.080 3260.000 1749.220 3272.850 ;
        RECT 1748.970 3256.000 1749.250 3260.000 ;
        RECT 2488.700 19.390 2488.960 19.710 ;
        RECT 2488.760 2.400 2488.900 19.390 ;
        RECT 2649.760 18.010 2649.900 3272.850 ;
        RECT 2649.700 17.690 2649.960 18.010 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2504.845 144.925 2505.015 193.035 ;
        RECT 2504.845 48.365 2505.015 96.475 ;
      LAYER mcon ;
        RECT 2504.845 192.865 2505.015 193.035 ;
        RECT 2504.845 96.305 2505.015 96.475 ;
      LAYER met1 ;
        RECT 2300.070 244.020 2300.390 244.080 ;
        RECT 2304.210 244.020 2304.530 244.080 ;
        RECT 2300.070 243.880 2304.530 244.020 ;
        RECT 2300.070 243.820 2300.390 243.880 ;
        RECT 2304.210 243.820 2304.530 243.880 ;
        RECT 2304.210 217.160 2304.530 217.220 ;
        RECT 2505.230 217.160 2505.550 217.220 ;
        RECT 2304.210 217.020 2505.550 217.160 ;
        RECT 2304.210 216.960 2304.530 217.020 ;
        RECT 2505.230 216.960 2505.550 217.020 ;
        RECT 2504.770 193.020 2505.090 193.080 ;
        RECT 2504.575 192.880 2505.090 193.020 ;
        RECT 2504.770 192.820 2505.090 192.880 ;
        RECT 2504.770 145.080 2505.090 145.140 ;
        RECT 2504.575 144.940 2505.090 145.080 ;
        RECT 2504.770 144.880 2505.090 144.940 ;
        RECT 2504.770 96.460 2505.090 96.520 ;
        RECT 2504.575 96.320 2505.090 96.460 ;
        RECT 2504.770 96.260 2505.090 96.320 ;
        RECT 2504.770 48.520 2505.090 48.580 ;
        RECT 2504.575 48.380 2505.090 48.520 ;
        RECT 2504.770 48.320 2505.090 48.380 ;
      LAYER via ;
        RECT 2300.100 243.820 2300.360 244.080 ;
        RECT 2304.240 243.820 2304.500 244.080 ;
        RECT 2304.240 216.960 2304.500 217.220 ;
        RECT 2505.260 216.960 2505.520 217.220 ;
        RECT 2504.800 192.820 2505.060 193.080 ;
        RECT 2504.800 144.880 2505.060 145.140 ;
        RECT 2504.800 96.260 2505.060 96.520 ;
        RECT 2504.800 48.320 2505.060 48.580 ;
      LAYER met2 ;
        RECT 2300.050 260.000 2300.330 264.000 ;
        RECT 2300.160 244.110 2300.300 260.000 ;
        RECT 2300.100 243.790 2300.360 244.110 ;
        RECT 2304.240 243.790 2304.500 244.110 ;
        RECT 2304.300 217.250 2304.440 243.790 ;
        RECT 2304.240 216.930 2304.500 217.250 ;
        RECT 2505.260 216.930 2505.520 217.250 ;
        RECT 2505.320 193.530 2505.460 216.930 ;
        RECT 2504.860 193.390 2505.460 193.530 ;
        RECT 2504.860 193.110 2505.000 193.390 ;
        RECT 2504.800 192.790 2505.060 193.110 ;
        RECT 2504.800 144.850 2505.060 145.170 ;
        RECT 2504.860 96.550 2505.000 144.850 ;
        RECT 2504.800 96.230 2505.060 96.550 ;
        RECT 2504.800 48.290 2505.060 48.610 ;
        RECT 2504.860 14.180 2505.000 48.290 ;
        RECT 2504.860 14.040 2505.920 14.180 ;
        RECT 2505.780 13.840 2505.920 14.040 ;
        RECT 2505.780 13.700 2506.380 13.840 ;
        RECT 2506.240 2.400 2506.380 13.700 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 267.330 1297.340 267.650 1297.400 ;
        RECT 296.770 1297.340 297.090 1297.400 ;
        RECT 267.330 1297.200 297.090 1297.340 ;
        RECT 267.330 1297.140 267.650 1297.200 ;
        RECT 296.770 1297.140 297.090 1297.200 ;
      LAYER via ;
        RECT 267.360 1297.140 267.620 1297.400 ;
        RECT 296.800 1297.140 297.060 1297.400 ;
      LAYER met2 ;
        RECT 296.790 1298.955 297.070 1299.325 ;
        RECT 296.860 1297.430 297.000 1298.955 ;
        RECT 267.360 1297.110 267.620 1297.430 ;
        RECT 296.800 1297.110 297.060 1297.430 ;
        RECT 267.420 16.845 267.560 1297.110 ;
        RECT 267.350 16.475 267.630 16.845 ;
        RECT 2524.110 16.475 2524.390 16.845 ;
        RECT 2524.180 2.400 2524.320 16.475 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
      LAYER via2 ;
        RECT 296.790 1299.000 297.070 1299.280 ;
        RECT 267.350 16.520 267.630 16.800 ;
        RECT 2524.110 16.520 2524.390 16.800 ;
      LAYER met3 ;
        RECT 296.765 1299.290 297.095 1299.305 ;
        RECT 310.000 1299.290 314.000 1299.680 ;
        RECT 296.765 1299.080 314.000 1299.290 ;
        RECT 296.765 1298.990 310.500 1299.080 ;
        RECT 296.765 1298.975 297.095 1298.990 ;
        RECT 267.325 16.810 267.655 16.825 ;
        RECT 2524.085 16.810 2524.415 16.825 ;
        RECT 267.325 16.510 2524.415 16.810 ;
        RECT 267.325 16.495 267.655 16.510 ;
        RECT 2524.085 16.495 2524.415 16.510 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1352.760 2615.490 1352.820 ;
        RECT 2666.690 1352.760 2667.010 1352.820 ;
        RECT 2615.170 1352.620 2667.010 1352.760 ;
        RECT 2615.170 1352.560 2615.490 1352.620 ;
        RECT 2666.690 1352.560 2667.010 1352.620 ;
        RECT 2545.710 257.960 2546.030 258.020 ;
        RECT 2666.690 257.960 2667.010 258.020 ;
        RECT 2545.710 257.820 2667.010 257.960 ;
        RECT 2545.710 257.760 2546.030 257.820 ;
        RECT 2666.690 257.760 2667.010 257.820 ;
        RECT 2542.030 20.640 2542.350 20.700 ;
        RECT 2545.710 20.640 2546.030 20.700 ;
        RECT 2542.030 20.500 2546.030 20.640 ;
        RECT 2542.030 20.440 2542.350 20.500 ;
        RECT 2545.710 20.440 2546.030 20.500 ;
      LAYER via ;
        RECT 2615.200 1352.560 2615.460 1352.820 ;
        RECT 2666.720 1352.560 2666.980 1352.820 ;
        RECT 2545.740 257.760 2546.000 258.020 ;
        RECT 2666.720 257.760 2666.980 258.020 ;
        RECT 2542.060 20.440 2542.320 20.700 ;
        RECT 2545.740 20.440 2546.000 20.700 ;
      LAYER met2 ;
        RECT 2615.190 1353.355 2615.470 1353.725 ;
        RECT 2615.260 1352.850 2615.400 1353.355 ;
        RECT 2615.200 1352.530 2615.460 1352.850 ;
        RECT 2666.720 1352.530 2666.980 1352.850 ;
        RECT 2666.780 258.050 2666.920 1352.530 ;
        RECT 2545.740 257.730 2546.000 258.050 ;
        RECT 2666.720 257.730 2666.980 258.050 ;
        RECT 2545.800 20.730 2545.940 257.730 ;
        RECT 2542.060 20.410 2542.320 20.730 ;
        RECT 2545.740 20.410 2546.000 20.730 ;
        RECT 2542.120 2.400 2542.260 20.410 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1353.400 2615.470 1353.680 ;
      LAYER met3 ;
        RECT 2606.000 1353.690 2610.000 1354.080 ;
        RECT 2615.165 1353.690 2615.495 1353.705 ;
        RECT 2606.000 1353.480 2615.495 1353.690 ;
        RECT 2609.580 1353.390 2615.495 1353.480 ;
        RECT 2615.165 1353.375 2615.495 1353.390 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2646.065 15.725 2646.235 20.655 ;
      LAYER mcon ;
        RECT 2646.065 20.485 2646.235 20.655 ;
      LAYER met1 ;
        RECT 2420.590 3274.780 2420.910 3274.840 ;
        RECT 2670.830 3274.780 2671.150 3274.840 ;
        RECT 2420.590 3274.640 2671.150 3274.780 ;
        RECT 2420.590 3274.580 2420.910 3274.640 ;
        RECT 2670.830 3274.580 2671.150 3274.640 ;
        RECT 2646.005 20.640 2646.295 20.685 ;
        RECT 2670.830 20.640 2671.150 20.700 ;
        RECT 2646.005 20.500 2671.150 20.640 ;
        RECT 2646.005 20.455 2646.295 20.500 ;
        RECT 2670.830 20.440 2671.150 20.500 ;
        RECT 2646.005 15.880 2646.295 15.925 ;
        RECT 2560.060 15.740 2646.295 15.880 ;
        RECT 2560.060 15.600 2560.200 15.740 ;
        RECT 2646.005 15.695 2646.295 15.740 ;
        RECT 2559.970 15.340 2560.290 15.600 ;
      LAYER via ;
        RECT 2420.620 3274.580 2420.880 3274.840 ;
        RECT 2670.860 3274.580 2671.120 3274.840 ;
        RECT 2670.860 20.440 2671.120 20.700 ;
        RECT 2560.000 15.340 2560.260 15.600 ;
      LAYER met2 ;
        RECT 2420.620 3274.550 2420.880 3274.870 ;
        RECT 2670.860 3274.550 2671.120 3274.870 ;
        RECT 2420.680 3260.000 2420.820 3274.550 ;
        RECT 2420.570 3256.000 2420.850 3260.000 ;
        RECT 2670.920 20.730 2671.060 3274.550 ;
        RECT 2670.860 20.410 2671.120 20.730 ;
        RECT 2560.000 15.310 2560.260 15.630 ;
        RECT 2560.060 2.400 2560.200 15.310 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 303.745 15.385 303.915 17.255 ;
        RECT 351.585 15.385 351.755 17.595 ;
        RECT 2560.045 14.025 2560.215 17.595 ;
      LAYER mcon ;
        RECT 351.585 17.425 351.755 17.595 ;
        RECT 303.745 17.085 303.915 17.255 ;
        RECT 2560.045 17.425 2560.215 17.595 ;
      LAYER met1 ;
        RECT 259.970 1127.680 260.290 1127.740 ;
        RECT 296.770 1127.680 297.090 1127.740 ;
        RECT 259.970 1127.540 297.090 1127.680 ;
        RECT 259.970 1127.480 260.290 1127.540 ;
        RECT 296.770 1127.480 297.090 1127.540 ;
        RECT 351.525 17.580 351.815 17.625 ;
        RECT 2559.985 17.580 2560.275 17.625 ;
        RECT 351.525 17.440 2560.275 17.580 ;
        RECT 351.525 17.395 351.815 17.440 ;
        RECT 2559.985 17.395 2560.275 17.440 ;
        RECT 259.970 17.240 260.290 17.300 ;
        RECT 303.685 17.240 303.975 17.285 ;
        RECT 259.970 17.100 303.975 17.240 ;
        RECT 259.970 17.040 260.290 17.100 ;
        RECT 303.685 17.055 303.975 17.100 ;
        RECT 303.685 15.540 303.975 15.585 ;
        RECT 351.525 15.540 351.815 15.585 ;
        RECT 303.685 15.400 351.815 15.540 ;
        RECT 303.685 15.355 303.975 15.400 ;
        RECT 351.525 15.355 351.815 15.400 ;
        RECT 2559.985 14.180 2560.275 14.225 ;
        RECT 2577.910 14.180 2578.230 14.240 ;
        RECT 2559.985 14.040 2578.230 14.180 ;
        RECT 2559.985 13.995 2560.275 14.040 ;
        RECT 2577.910 13.980 2578.230 14.040 ;
      LAYER via ;
        RECT 260.000 1127.480 260.260 1127.740 ;
        RECT 296.800 1127.480 297.060 1127.740 ;
        RECT 260.000 17.040 260.260 17.300 ;
        RECT 2577.940 13.980 2578.200 14.240 ;
      LAYER met2 ;
        RECT 296.790 1130.315 297.070 1130.685 ;
        RECT 296.860 1127.770 297.000 1130.315 ;
        RECT 260.000 1127.450 260.260 1127.770 ;
        RECT 296.800 1127.450 297.060 1127.770 ;
        RECT 260.060 17.330 260.200 1127.450 ;
        RECT 260.000 17.010 260.260 17.330 ;
        RECT 2577.940 13.950 2578.200 14.270 ;
        RECT 2578.000 2.400 2578.140 13.950 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
      LAYER via2 ;
        RECT 296.790 1130.360 297.070 1130.640 ;
      LAYER met3 ;
        RECT 296.765 1130.650 297.095 1130.665 ;
        RECT 310.000 1130.650 314.000 1131.040 ;
        RECT 296.765 1130.440 314.000 1130.650 ;
        RECT 296.765 1130.350 310.500 1130.440 ;
        RECT 296.765 1130.335 297.095 1130.350 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 297.305 17.425 297.475 19.975 ;
      LAYER mcon ;
        RECT 297.305 19.805 297.475 19.975 ;
      LAYER met1 ;
        RECT 267.790 2159.920 268.110 2159.980 ;
        RECT 296.770 2159.920 297.090 2159.980 ;
        RECT 267.790 2159.780 297.090 2159.920 ;
        RECT 267.790 2159.720 268.110 2159.780 ;
        RECT 296.770 2159.720 297.090 2159.780 ;
        RECT 297.245 19.960 297.535 20.005 ;
        RECT 811.510 19.960 811.830 20.020 ;
        RECT 297.245 19.820 811.830 19.960 ;
        RECT 297.245 19.775 297.535 19.820 ;
        RECT 811.510 19.760 811.830 19.820 ;
        RECT 267.790 17.580 268.110 17.640 ;
        RECT 297.245 17.580 297.535 17.625 ;
        RECT 267.790 17.440 297.535 17.580 ;
        RECT 267.790 17.380 268.110 17.440 ;
        RECT 297.245 17.395 297.535 17.440 ;
      LAYER via ;
        RECT 267.820 2159.720 268.080 2159.980 ;
        RECT 296.800 2159.720 297.060 2159.980 ;
        RECT 811.540 19.760 811.800 20.020 ;
        RECT 267.820 17.380 268.080 17.640 ;
      LAYER met2 ;
        RECT 296.790 2165.275 297.070 2165.645 ;
        RECT 296.860 2160.010 297.000 2165.275 ;
        RECT 267.820 2159.690 268.080 2160.010 ;
        RECT 296.800 2159.690 297.060 2160.010 ;
        RECT 267.880 17.670 268.020 2159.690 ;
        RECT 811.540 19.730 811.800 20.050 ;
        RECT 267.820 17.350 268.080 17.670 ;
        RECT 811.600 2.400 811.740 19.730 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 296.790 2165.320 297.070 2165.600 ;
      LAYER met3 ;
        RECT 296.765 2165.610 297.095 2165.625 ;
        RECT 310.000 2165.610 314.000 2166.000 ;
        RECT 296.765 2165.400 314.000 2165.610 ;
        RECT 296.765 2165.310 310.500 2165.400 ;
        RECT 296.765 2165.295 297.095 2165.310 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 86.260 358.730 86.320 ;
        RECT 2594.470 86.260 2594.790 86.320 ;
        RECT 358.410 86.120 2594.790 86.260 ;
        RECT 358.410 86.060 358.730 86.120 ;
        RECT 2594.470 86.060 2594.790 86.120 ;
        RECT 2594.470 2.960 2594.790 3.020 ;
        RECT 2595.390 2.960 2595.710 3.020 ;
        RECT 2594.470 2.820 2595.710 2.960 ;
        RECT 2594.470 2.760 2594.790 2.820 ;
        RECT 2595.390 2.760 2595.710 2.820 ;
      LAYER via ;
        RECT 358.440 86.060 358.700 86.320 ;
        RECT 2594.500 86.060 2594.760 86.320 ;
        RECT 2594.500 2.760 2594.760 3.020 ;
        RECT 2595.420 2.760 2595.680 3.020 ;
      LAYER met2 ;
        RECT 355.170 260.170 355.450 264.000 ;
        RECT 355.170 260.030 358.640 260.170 ;
        RECT 355.170 260.000 355.450 260.030 ;
        RECT 358.500 86.350 358.640 260.030 ;
        RECT 358.440 86.030 358.700 86.350 ;
        RECT 2594.500 86.030 2594.760 86.350 ;
        RECT 2594.560 3.050 2594.700 86.030 ;
        RECT 2594.500 2.730 2594.760 3.050 ;
        RECT 2595.420 2.730 2595.680 3.050 ;
        RECT 2595.480 2.400 2595.620 2.730 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 257.745 1015.325 257.915 1097.095 ;
        RECT 257.745 966.025 257.915 980.135 ;
        RECT 256.825 193.205 256.995 241.315 ;
        RECT 258.205 144.925 258.375 192.695 ;
        RECT 258.205 96.645 258.375 111.095 ;
      LAYER mcon ;
        RECT 257.745 1096.925 257.915 1097.095 ;
        RECT 257.745 979.965 257.915 980.135 ;
        RECT 256.825 241.145 256.995 241.315 ;
        RECT 258.205 192.525 258.375 192.695 ;
        RECT 258.205 110.925 258.375 111.095 ;
      LAYER met1 ;
        RECT 258.130 1104.220 258.450 1104.280 ;
        RECT 296.770 1104.220 297.090 1104.280 ;
        RECT 258.130 1104.080 297.090 1104.220 ;
        RECT 258.130 1104.020 258.450 1104.080 ;
        RECT 296.770 1104.020 297.090 1104.080 ;
        RECT 257.670 1097.080 257.990 1097.140 ;
        RECT 257.475 1096.940 257.990 1097.080 ;
        RECT 257.670 1096.880 257.990 1096.940 ;
        RECT 257.670 1015.480 257.990 1015.540 ;
        RECT 257.475 1015.340 257.990 1015.480 ;
        RECT 257.670 1015.280 257.990 1015.340 ;
        RECT 257.670 980.120 257.990 980.180 ;
        RECT 257.475 979.980 257.990 980.120 ;
        RECT 257.670 979.920 257.990 979.980 ;
        RECT 257.670 966.180 257.990 966.240 ;
        RECT 257.475 966.040 257.990 966.180 ;
        RECT 257.670 965.980 257.990 966.040 ;
        RECT 256.750 931.500 257.070 931.560 ;
        RECT 257.670 931.500 257.990 931.560 ;
        RECT 256.750 931.360 257.990 931.500 ;
        RECT 256.750 931.300 257.070 931.360 ;
        RECT 257.670 931.300 257.990 931.360 ;
        RECT 256.750 903.960 257.070 904.020 ;
        RECT 257.670 903.960 257.990 904.020 ;
        RECT 256.750 903.820 257.990 903.960 ;
        RECT 256.750 903.760 257.070 903.820 ;
        RECT 257.670 903.760 257.990 903.820 ;
        RECT 256.750 845.480 257.070 845.540 ;
        RECT 258.130 845.480 258.450 845.540 ;
        RECT 256.750 845.340 258.450 845.480 ;
        RECT 256.750 845.280 257.070 845.340 ;
        RECT 258.130 845.280 258.450 845.340 ;
        RECT 256.750 738.380 257.070 738.440 ;
        RECT 258.130 738.380 258.450 738.440 ;
        RECT 256.750 738.240 258.450 738.380 ;
        RECT 256.750 738.180 257.070 738.240 ;
        RECT 258.130 738.180 258.450 738.240 ;
        RECT 256.750 689.760 257.070 689.820 ;
        RECT 258.130 689.760 258.450 689.820 ;
        RECT 256.750 689.620 258.450 689.760 ;
        RECT 256.750 689.560 257.070 689.620 ;
        RECT 258.130 689.560 258.450 689.620 ;
        RECT 256.750 642.160 257.070 642.220 ;
        RECT 258.130 642.160 258.450 642.220 ;
        RECT 256.750 642.020 258.450 642.160 ;
        RECT 256.750 641.960 257.070 642.020 ;
        RECT 258.130 641.960 258.450 642.020 ;
        RECT 256.750 593.200 257.070 593.260 ;
        RECT 258.130 593.200 258.450 593.260 ;
        RECT 256.750 593.060 258.450 593.200 ;
        RECT 256.750 593.000 257.070 593.060 ;
        RECT 258.130 593.000 258.450 593.060 ;
        RECT 256.750 545.260 257.070 545.320 ;
        RECT 258.130 545.260 258.450 545.320 ;
        RECT 256.750 545.120 258.450 545.260 ;
        RECT 256.750 545.060 257.070 545.120 ;
        RECT 258.130 545.060 258.450 545.120 ;
        RECT 256.750 496.640 257.070 496.700 ;
        RECT 258.130 496.640 258.450 496.700 ;
        RECT 256.750 496.500 258.450 496.640 ;
        RECT 256.750 496.440 257.070 496.500 ;
        RECT 258.130 496.440 258.450 496.500 ;
        RECT 256.750 448.700 257.070 448.760 ;
        RECT 258.130 448.700 258.450 448.760 ;
        RECT 256.750 448.560 258.450 448.700 ;
        RECT 256.750 448.500 257.070 448.560 ;
        RECT 258.130 448.500 258.450 448.560 ;
        RECT 256.750 400.080 257.070 400.140 ;
        RECT 258.130 400.080 258.450 400.140 ;
        RECT 256.750 399.940 258.450 400.080 ;
        RECT 256.750 399.880 257.070 399.940 ;
        RECT 258.130 399.880 258.450 399.940 ;
        RECT 256.750 352.140 257.070 352.200 ;
        RECT 258.130 352.140 258.450 352.200 ;
        RECT 256.750 352.000 258.450 352.140 ;
        RECT 256.750 351.940 257.070 352.000 ;
        RECT 258.130 351.940 258.450 352.000 ;
        RECT 256.750 303.520 257.070 303.580 ;
        RECT 258.130 303.520 258.450 303.580 ;
        RECT 256.750 303.380 258.450 303.520 ;
        RECT 256.750 303.320 257.070 303.380 ;
        RECT 258.130 303.320 258.450 303.380 ;
        RECT 256.750 255.240 257.070 255.300 ;
        RECT 258.130 255.240 258.450 255.300 ;
        RECT 256.750 255.100 258.450 255.240 ;
        RECT 256.750 255.040 257.070 255.100 ;
        RECT 258.130 255.040 258.450 255.100 ;
        RECT 256.750 241.300 257.070 241.360 ;
        RECT 256.555 241.160 257.070 241.300 ;
        RECT 256.750 241.100 257.070 241.160 ;
        RECT 256.765 193.360 257.055 193.405 ;
        RECT 258.130 193.360 258.450 193.420 ;
        RECT 256.765 193.220 258.450 193.360 ;
        RECT 256.765 193.175 257.055 193.220 ;
        RECT 258.130 193.160 258.450 193.220 ;
        RECT 258.130 192.680 258.450 192.740 ;
        RECT 257.935 192.540 258.450 192.680 ;
        RECT 258.130 192.480 258.450 192.540 ;
        RECT 258.145 145.080 258.435 145.125 ;
        RECT 258.590 145.080 258.910 145.140 ;
        RECT 258.145 144.940 258.910 145.080 ;
        RECT 258.145 144.895 258.435 144.940 ;
        RECT 258.590 144.880 258.910 144.940 ;
        RECT 258.130 111.080 258.450 111.140 ;
        RECT 257.935 110.940 258.450 111.080 ;
        RECT 258.130 110.880 258.450 110.940 ;
        RECT 258.130 96.800 258.450 96.860 ;
        RECT 257.935 96.660 258.450 96.800 ;
        RECT 258.130 96.600 258.450 96.660 ;
        RECT 258.590 32.200 258.910 32.260 ;
        RECT 2613.330 32.200 2613.650 32.260 ;
        RECT 258.590 32.060 2613.650 32.200 ;
        RECT 258.590 32.000 258.910 32.060 ;
        RECT 2613.330 32.000 2613.650 32.060 ;
      LAYER via ;
        RECT 258.160 1104.020 258.420 1104.280 ;
        RECT 296.800 1104.020 297.060 1104.280 ;
        RECT 257.700 1096.880 257.960 1097.140 ;
        RECT 257.700 1015.280 257.960 1015.540 ;
        RECT 257.700 979.920 257.960 980.180 ;
        RECT 257.700 965.980 257.960 966.240 ;
        RECT 256.780 931.300 257.040 931.560 ;
        RECT 257.700 931.300 257.960 931.560 ;
        RECT 256.780 903.760 257.040 904.020 ;
        RECT 257.700 903.760 257.960 904.020 ;
        RECT 256.780 845.280 257.040 845.540 ;
        RECT 258.160 845.280 258.420 845.540 ;
        RECT 256.780 738.180 257.040 738.440 ;
        RECT 258.160 738.180 258.420 738.440 ;
        RECT 256.780 689.560 257.040 689.820 ;
        RECT 258.160 689.560 258.420 689.820 ;
        RECT 256.780 641.960 257.040 642.220 ;
        RECT 258.160 641.960 258.420 642.220 ;
        RECT 256.780 593.000 257.040 593.260 ;
        RECT 258.160 593.000 258.420 593.260 ;
        RECT 256.780 545.060 257.040 545.320 ;
        RECT 258.160 545.060 258.420 545.320 ;
        RECT 256.780 496.440 257.040 496.700 ;
        RECT 258.160 496.440 258.420 496.700 ;
        RECT 256.780 448.500 257.040 448.760 ;
        RECT 258.160 448.500 258.420 448.760 ;
        RECT 256.780 399.880 257.040 400.140 ;
        RECT 258.160 399.880 258.420 400.140 ;
        RECT 256.780 351.940 257.040 352.200 ;
        RECT 258.160 351.940 258.420 352.200 ;
        RECT 256.780 303.320 257.040 303.580 ;
        RECT 258.160 303.320 258.420 303.580 ;
        RECT 256.780 255.040 257.040 255.300 ;
        RECT 258.160 255.040 258.420 255.300 ;
        RECT 256.780 241.100 257.040 241.360 ;
        RECT 258.160 193.160 258.420 193.420 ;
        RECT 258.160 192.480 258.420 192.740 ;
        RECT 258.620 144.880 258.880 145.140 ;
        RECT 258.160 110.880 258.420 111.140 ;
        RECT 258.160 96.600 258.420 96.860 ;
        RECT 258.620 32.000 258.880 32.260 ;
        RECT 2613.360 32.000 2613.620 32.260 ;
      LAYER met2 ;
        RECT 296.790 1108.555 297.070 1108.925 ;
        RECT 296.860 1104.310 297.000 1108.555 ;
        RECT 258.160 1104.220 258.420 1104.310 ;
        RECT 257.760 1104.080 258.420 1104.220 ;
        RECT 257.760 1097.170 257.900 1104.080 ;
        RECT 258.160 1103.990 258.420 1104.080 ;
        RECT 296.800 1103.990 297.060 1104.310 ;
        RECT 257.700 1096.850 257.960 1097.170 ;
        RECT 257.700 1015.250 257.960 1015.570 ;
        RECT 257.760 980.210 257.900 1015.250 ;
        RECT 257.700 979.890 257.960 980.210 ;
        RECT 257.700 966.125 257.960 966.270 ;
        RECT 256.770 965.755 257.050 966.125 ;
        RECT 257.690 965.755 257.970 966.125 ;
        RECT 256.840 931.590 256.980 965.755 ;
        RECT 256.780 931.270 257.040 931.590 ;
        RECT 257.700 931.270 257.960 931.590 ;
        RECT 257.760 904.050 257.900 931.270 ;
        RECT 256.780 903.730 257.040 904.050 ;
        RECT 257.700 903.730 257.960 904.050 ;
        RECT 256.840 855.965 256.980 903.730 ;
        RECT 256.770 855.595 257.050 855.965 ;
        RECT 258.150 855.595 258.430 855.965 ;
        RECT 258.220 845.570 258.360 855.595 ;
        RECT 256.780 845.250 257.040 845.570 ;
        RECT 258.160 845.250 258.420 845.570 ;
        RECT 256.840 738.470 256.980 845.250 ;
        RECT 256.780 738.150 257.040 738.470 ;
        RECT 258.160 738.150 258.420 738.470 ;
        RECT 258.220 689.850 258.360 738.150 ;
        RECT 256.780 689.530 257.040 689.850 ;
        RECT 258.160 689.530 258.420 689.850 ;
        RECT 256.840 642.250 256.980 689.530 ;
        RECT 256.780 641.930 257.040 642.250 ;
        RECT 258.160 641.930 258.420 642.250 ;
        RECT 258.220 593.290 258.360 641.930 ;
        RECT 256.780 592.970 257.040 593.290 ;
        RECT 258.160 592.970 258.420 593.290 ;
        RECT 256.840 545.350 256.980 592.970 ;
        RECT 256.780 545.030 257.040 545.350 ;
        RECT 258.160 545.030 258.420 545.350 ;
        RECT 258.220 496.730 258.360 545.030 ;
        RECT 256.780 496.410 257.040 496.730 ;
        RECT 258.160 496.410 258.420 496.730 ;
        RECT 256.840 448.790 256.980 496.410 ;
        RECT 256.780 448.470 257.040 448.790 ;
        RECT 258.160 448.470 258.420 448.790 ;
        RECT 258.220 400.170 258.360 448.470 ;
        RECT 256.780 399.850 257.040 400.170 ;
        RECT 258.160 399.850 258.420 400.170 ;
        RECT 256.840 352.230 256.980 399.850 ;
        RECT 256.780 351.910 257.040 352.230 ;
        RECT 258.160 351.910 258.420 352.230 ;
        RECT 258.220 303.610 258.360 351.910 ;
        RECT 256.780 303.290 257.040 303.610 ;
        RECT 258.160 303.290 258.420 303.610 ;
        RECT 256.840 255.525 256.980 303.290 ;
        RECT 256.770 255.155 257.050 255.525 ;
        RECT 258.150 255.155 258.430 255.525 ;
        RECT 256.780 255.010 257.040 255.155 ;
        RECT 258.160 255.010 258.420 255.155 ;
        RECT 256.840 241.390 256.980 255.010 ;
        RECT 256.780 241.070 257.040 241.390 ;
        RECT 258.160 193.130 258.420 193.450 ;
        RECT 258.220 192.770 258.360 193.130 ;
        RECT 258.160 192.450 258.420 192.770 ;
        RECT 258.620 144.850 258.880 145.170 ;
        RECT 258.680 144.570 258.820 144.850 ;
        RECT 258.220 144.430 258.820 144.570 ;
        RECT 258.220 111.170 258.360 144.430 ;
        RECT 258.160 110.850 258.420 111.170 ;
        RECT 258.160 96.570 258.420 96.890 ;
        RECT 258.220 47.330 258.360 96.570 ;
        RECT 258.220 47.190 258.820 47.330 ;
        RECT 258.680 32.290 258.820 47.190 ;
        RECT 258.620 31.970 258.880 32.290 ;
        RECT 2613.360 31.970 2613.620 32.290 ;
        RECT 2613.420 2.400 2613.560 31.970 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
      LAYER via2 ;
        RECT 296.790 1108.600 297.070 1108.880 ;
        RECT 256.770 965.800 257.050 966.080 ;
        RECT 257.690 965.800 257.970 966.080 ;
        RECT 256.770 855.640 257.050 855.920 ;
        RECT 258.150 855.640 258.430 855.920 ;
        RECT 256.770 255.200 257.050 255.480 ;
        RECT 258.150 255.200 258.430 255.480 ;
      LAYER met3 ;
        RECT 296.765 1108.890 297.095 1108.905 ;
        RECT 310.000 1108.890 314.000 1109.280 ;
        RECT 296.765 1108.680 314.000 1108.890 ;
        RECT 296.765 1108.590 310.500 1108.680 ;
        RECT 296.765 1108.575 297.095 1108.590 ;
        RECT 256.745 966.090 257.075 966.105 ;
        RECT 257.665 966.090 257.995 966.105 ;
        RECT 256.745 965.790 257.995 966.090 ;
        RECT 256.745 965.775 257.075 965.790 ;
        RECT 257.665 965.775 257.995 965.790 ;
        RECT 256.745 855.930 257.075 855.945 ;
        RECT 258.125 855.930 258.455 855.945 ;
        RECT 256.745 855.630 258.455 855.930 ;
        RECT 256.745 855.615 257.075 855.630 ;
        RECT 258.125 855.615 258.455 855.630 ;
        RECT 256.745 255.490 257.075 255.505 ;
        RECT 258.125 255.490 258.455 255.505 ;
        RECT 256.745 255.190 258.455 255.490 ;
        RECT 256.745 255.175 257.075 255.190 ;
        RECT 258.125 255.175 258.455 255.190 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2428.870 244.020 2429.190 244.080 ;
        RECT 2434.390 244.020 2434.710 244.080 ;
        RECT 2428.870 243.880 2434.710 244.020 ;
        RECT 2428.870 243.820 2429.190 243.880 ;
        RECT 2434.390 243.820 2434.710 243.880 ;
        RECT 2434.390 45.120 2434.710 45.180 ;
        RECT 2631.270 45.120 2631.590 45.180 ;
        RECT 2434.390 44.980 2631.590 45.120 ;
        RECT 2434.390 44.920 2434.710 44.980 ;
        RECT 2631.270 44.920 2631.590 44.980 ;
      LAYER via ;
        RECT 2428.900 243.820 2429.160 244.080 ;
        RECT 2434.420 243.820 2434.680 244.080 ;
        RECT 2434.420 44.920 2434.680 45.180 ;
        RECT 2631.300 44.920 2631.560 45.180 ;
      LAYER met2 ;
        RECT 2428.850 260.000 2429.130 264.000 ;
        RECT 2428.960 244.110 2429.100 260.000 ;
        RECT 2428.900 243.790 2429.160 244.110 ;
        RECT 2434.420 243.790 2434.680 244.110 ;
        RECT 2434.480 45.210 2434.620 243.790 ;
        RECT 2434.420 44.890 2434.680 45.210 ;
        RECT 2631.300 44.890 2631.560 45.210 ;
        RECT 2631.360 2.400 2631.500 44.890 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 65.520 2573.630 65.580 ;
        RECT 2643.230 65.520 2643.550 65.580 ;
        RECT 2573.310 65.380 2643.550 65.520 ;
        RECT 2573.310 65.320 2573.630 65.380 ;
        RECT 2643.230 65.320 2643.550 65.380 ;
        RECT 2643.230 37.980 2643.550 38.040 ;
        RECT 2649.210 37.980 2649.530 38.040 ;
        RECT 2643.230 37.840 2649.530 37.980 ;
        RECT 2643.230 37.780 2643.550 37.840 ;
        RECT 2649.210 37.780 2649.530 37.840 ;
      LAYER via ;
        RECT 2573.340 65.320 2573.600 65.580 ;
        RECT 2643.260 65.320 2643.520 65.580 ;
        RECT 2643.260 37.780 2643.520 38.040 ;
        RECT 2649.240 37.780 2649.500 38.040 ;
      LAYER met2 ;
        RECT 2571.450 260.170 2571.730 264.000 ;
        RECT 2571.450 260.030 2573.540 260.170 ;
        RECT 2571.450 260.000 2571.730 260.030 ;
        RECT 2573.400 65.610 2573.540 260.030 ;
        RECT 2573.340 65.290 2573.600 65.610 ;
        RECT 2643.260 65.290 2643.520 65.610 ;
        RECT 2643.320 38.070 2643.460 65.290 ;
        RECT 2643.260 37.750 2643.520 38.070 ;
        RECT 2649.240 37.750 2649.500 38.070 ;
        RECT 2649.300 2.400 2649.440 37.750 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 906.750 3260.075 907.030 3260.445 ;
        RECT 905.330 3259.650 905.610 3260.000 ;
        RECT 906.820 3259.650 906.960 3260.075 ;
        RECT 905.330 3259.510 906.960 3259.650 ;
        RECT 905.330 3256.000 905.610 3259.510 ;
        RECT 2667.170 19.875 2667.450 20.245 ;
        RECT 2667.240 2.400 2667.380 19.875 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
      LAYER via2 ;
        RECT 906.750 3260.120 907.030 3260.400 ;
        RECT 2667.170 19.920 2667.450 20.200 ;
      LAYER met3 ;
        RECT 906.725 3260.410 907.055 3260.425 ;
        RECT 907.390 3260.410 907.770 3260.420 ;
        RECT 906.725 3260.110 907.770 3260.410 ;
        RECT 906.725 3260.095 907.055 3260.110 ;
        RECT 907.390 3260.100 907.770 3260.110 ;
        RECT 907.390 3250.890 907.770 3250.900 ;
        RECT 2663.670 3250.890 2664.050 3250.900 ;
        RECT 907.390 3250.590 2664.050 3250.890 ;
        RECT 907.390 3250.580 907.770 3250.590 ;
        RECT 2663.670 3250.580 2664.050 3250.590 ;
        RECT 2663.670 20.210 2664.050 20.220 ;
        RECT 2667.145 20.210 2667.475 20.225 ;
        RECT 2663.670 19.910 2667.475 20.210 ;
        RECT 2663.670 19.900 2664.050 19.910 ;
        RECT 2667.145 19.895 2667.475 19.910 ;
      LAYER via3 ;
        RECT 907.420 3260.100 907.740 3260.420 ;
        RECT 907.420 3250.580 907.740 3250.900 ;
        RECT 2663.700 3250.580 2664.020 3250.900 ;
        RECT 2663.700 19.900 2664.020 20.220 ;
      LAYER met4 ;
        RECT 907.415 3260.095 907.745 3260.425 ;
        RECT 907.430 3250.905 907.730 3260.095 ;
        RECT 907.415 3250.575 907.745 3250.905 ;
        RECT 2663.695 3250.575 2664.025 3250.905 ;
        RECT 2663.710 20.225 2664.010 3250.575 ;
        RECT 2663.695 19.895 2664.025 20.225 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 266.870 1166.440 267.190 1166.500 ;
        RECT 296.770 1166.440 297.090 1166.500 ;
        RECT 266.870 1166.300 297.090 1166.440 ;
        RECT 266.870 1166.240 267.190 1166.300 ;
        RECT 296.770 1166.240 297.090 1166.300 ;
        RECT 266.870 31.860 267.190 31.920 ;
        RECT 2684.630 31.860 2684.950 31.920 ;
        RECT 266.870 31.720 2684.950 31.860 ;
        RECT 266.870 31.660 267.190 31.720 ;
        RECT 2684.630 31.660 2684.950 31.720 ;
      LAYER via ;
        RECT 266.900 1166.240 267.160 1166.500 ;
        RECT 296.800 1166.240 297.060 1166.500 ;
        RECT 266.900 31.660 267.160 31.920 ;
        RECT 2684.660 31.660 2684.920 31.920 ;
      LAYER met2 ;
        RECT 296.790 1172.475 297.070 1172.845 ;
        RECT 296.860 1166.530 297.000 1172.475 ;
        RECT 266.900 1166.210 267.160 1166.530 ;
        RECT 296.800 1166.210 297.060 1166.530 ;
        RECT 266.960 31.950 267.100 1166.210 ;
        RECT 266.900 31.630 267.160 31.950 ;
        RECT 2684.660 31.630 2684.920 31.950 ;
        RECT 2684.720 2.400 2684.860 31.630 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
      LAYER via2 ;
        RECT 296.790 1172.520 297.070 1172.800 ;
      LAYER met3 ;
        RECT 296.765 1172.810 297.095 1172.825 ;
        RECT 310.000 1172.810 314.000 1173.200 ;
        RECT 296.765 1172.600 314.000 1172.810 ;
        RECT 296.765 1172.510 310.500 1172.600 ;
        RECT 296.765 1172.495 297.095 1172.510 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 713.070 244.020 713.390 244.080 ;
        RECT 717.210 244.020 717.530 244.080 ;
        RECT 713.070 243.880 717.530 244.020 ;
        RECT 713.070 243.820 713.390 243.880 ;
        RECT 717.210 243.820 717.530 243.880 ;
        RECT 717.210 93.400 717.530 93.460 ;
        RECT 2698.430 93.400 2698.750 93.460 ;
        RECT 717.210 93.260 2698.750 93.400 ;
        RECT 717.210 93.200 717.530 93.260 ;
        RECT 2698.430 93.200 2698.750 93.260 ;
      LAYER via ;
        RECT 713.100 243.820 713.360 244.080 ;
        RECT 717.240 243.820 717.500 244.080 ;
        RECT 717.240 93.200 717.500 93.460 ;
        RECT 2698.460 93.200 2698.720 93.460 ;
      LAYER met2 ;
        RECT 713.050 260.000 713.330 264.000 ;
        RECT 713.160 244.110 713.300 260.000 ;
        RECT 713.100 243.790 713.360 244.110 ;
        RECT 717.240 243.790 717.500 244.110 ;
        RECT 717.300 93.490 717.440 243.790 ;
        RECT 717.240 93.170 717.500 93.490 ;
        RECT 2698.460 93.170 2698.720 93.490 ;
        RECT 2698.520 17.410 2698.660 93.170 ;
        RECT 2698.520 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2714.990 17.920 2715.310 17.980 ;
        RECT 2720.510 17.920 2720.830 17.980 ;
        RECT 2714.990 17.780 2720.830 17.920 ;
        RECT 2714.990 17.720 2715.310 17.780 ;
        RECT 2720.510 17.720 2720.830 17.780 ;
      LAYER via ;
        RECT 2715.020 17.720 2715.280 17.980 ;
        RECT 2720.540 17.720 2720.800 17.980 ;
      LAYER met2 ;
        RECT 1934.850 3267.555 1935.130 3267.925 ;
        RECT 2715.010 3267.555 2715.290 3267.925 ;
        RECT 1934.920 3260.000 1935.060 3267.555 ;
        RECT 1934.810 3256.000 1935.090 3260.000 ;
        RECT 2715.080 18.010 2715.220 3267.555 ;
        RECT 2715.020 17.690 2715.280 18.010 ;
        RECT 2720.540 17.690 2720.800 18.010 ;
        RECT 2720.600 2.400 2720.740 17.690 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
      LAYER via2 ;
        RECT 1934.850 3267.600 1935.130 3267.880 ;
        RECT 2715.010 3267.600 2715.290 3267.880 ;
      LAYER met3 ;
        RECT 1934.825 3267.890 1935.155 3267.905 ;
        RECT 2714.985 3267.890 2715.315 3267.905 ;
        RECT 1934.825 3267.590 2715.315 3267.890 ;
        RECT 1934.825 3267.575 1935.155 3267.590 ;
        RECT 2714.985 3267.575 2715.315 3267.590 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1944.950 100.880 1945.270 100.940 ;
        RECT 2732.470 100.880 2732.790 100.940 ;
        RECT 1944.950 100.740 2732.790 100.880 ;
        RECT 1944.950 100.680 1945.270 100.740 ;
        RECT 2732.470 100.680 2732.790 100.740 ;
        RECT 2732.470 37.980 2732.790 38.040 ;
        RECT 2738.450 37.980 2738.770 38.040 ;
        RECT 2732.470 37.840 2738.770 37.980 ;
        RECT 2732.470 37.780 2732.790 37.840 ;
        RECT 2738.450 37.780 2738.770 37.840 ;
      LAYER via ;
        RECT 1944.980 100.680 1945.240 100.940 ;
        RECT 2732.500 100.680 2732.760 100.940 ;
        RECT 2732.500 37.780 2732.760 38.040 ;
        RECT 2738.480 37.780 2738.740 38.040 ;
      LAYER met2 ;
        RECT 1942.170 260.170 1942.450 264.000 ;
        RECT 1942.170 260.030 1945.180 260.170 ;
        RECT 1942.170 260.000 1942.450 260.030 ;
        RECT 1945.040 100.970 1945.180 260.030 ;
        RECT 1944.980 100.650 1945.240 100.970 ;
        RECT 2732.500 100.650 2732.760 100.970 ;
        RECT 2732.560 38.070 2732.700 100.650 ;
        RECT 2732.500 37.750 2732.760 38.070 ;
        RECT 2738.480 37.750 2738.740 38.070 ;
        RECT 2738.540 2.400 2738.680 37.750 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 469.270 241.640 469.590 241.700 ;
        RECT 475.710 241.640 476.030 241.700 ;
        RECT 469.270 241.500 476.030 241.640 ;
        RECT 469.270 241.440 469.590 241.500 ;
        RECT 475.710 241.440 476.030 241.500 ;
        RECT 475.710 203.560 476.030 203.620 ;
        RECT 2753.170 203.560 2753.490 203.620 ;
        RECT 475.710 203.420 2753.490 203.560 ;
        RECT 475.710 203.360 476.030 203.420 ;
        RECT 2753.170 203.360 2753.490 203.420 ;
        RECT 2753.170 62.120 2753.490 62.180 ;
        RECT 2755.930 62.120 2756.250 62.180 ;
        RECT 2753.170 61.980 2756.250 62.120 ;
        RECT 2753.170 61.920 2753.490 61.980 ;
        RECT 2755.930 61.920 2756.250 61.980 ;
      LAYER via ;
        RECT 469.300 241.440 469.560 241.700 ;
        RECT 475.740 241.440 476.000 241.700 ;
        RECT 475.740 203.360 476.000 203.620 ;
        RECT 2753.200 203.360 2753.460 203.620 ;
        RECT 2753.200 61.920 2753.460 62.180 ;
        RECT 2755.960 61.920 2756.220 62.180 ;
      LAYER met2 ;
        RECT 469.250 260.000 469.530 264.000 ;
        RECT 469.360 241.730 469.500 260.000 ;
        RECT 469.300 241.410 469.560 241.730 ;
        RECT 475.740 241.410 476.000 241.730 ;
        RECT 475.800 203.650 475.940 241.410 ;
        RECT 475.740 203.330 476.000 203.650 ;
        RECT 2753.200 203.330 2753.460 203.650 ;
        RECT 2753.260 62.210 2753.400 203.330 ;
        RECT 2753.200 61.890 2753.460 62.210 ;
        RECT 2755.960 61.890 2756.220 62.210 ;
        RECT 2756.020 2.400 2756.160 61.890 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 253.070 2967.080 253.390 2967.140 ;
        RECT 296.770 2967.080 297.090 2967.140 ;
        RECT 253.070 2966.940 297.090 2967.080 ;
        RECT 253.070 2966.880 253.390 2966.940 ;
        RECT 296.770 2966.880 297.090 2966.940 ;
      LAYER via ;
        RECT 253.100 2966.880 253.360 2967.140 ;
        RECT 296.800 2966.880 297.060 2967.140 ;
      LAYER met2 ;
        RECT 296.790 2969.035 297.070 2969.405 ;
        RECT 296.860 2967.170 297.000 2969.035 ;
        RECT 253.100 2966.850 253.360 2967.170 ;
        RECT 296.800 2966.850 297.060 2967.170 ;
        RECT 253.160 19.565 253.300 2966.850 ;
        RECT 253.090 19.195 253.370 19.565 ;
        RECT 829.470 19.195 829.750 19.565 ;
        RECT 829.540 2.400 829.680 19.195 ;
        RECT 829.330 -4.800 829.890 2.400 ;
      LAYER via2 ;
        RECT 296.790 2969.080 297.070 2969.360 ;
        RECT 253.090 19.240 253.370 19.520 ;
        RECT 829.470 19.240 829.750 19.520 ;
      LAYER met3 ;
        RECT 296.765 2969.370 297.095 2969.385 ;
        RECT 310.000 2969.370 314.000 2969.760 ;
        RECT 296.765 2969.160 314.000 2969.370 ;
        RECT 296.765 2969.070 310.500 2969.160 ;
        RECT 296.765 2969.055 297.095 2969.070 ;
        RECT 253.065 19.530 253.395 19.545 ;
        RECT 829.445 19.530 829.775 19.545 ;
        RECT 253.065 19.230 829.775 19.530 ;
        RECT 253.065 19.215 253.395 19.230 ;
        RECT 829.445 19.215 829.775 19.230 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 272.390 897.160 272.710 897.220 ;
        RECT 296.770 897.160 297.090 897.220 ;
        RECT 272.390 897.020 297.090 897.160 ;
        RECT 272.390 896.960 272.710 897.020 ;
        RECT 296.770 896.960 297.090 897.020 ;
        RECT 272.390 31.520 272.710 31.580 ;
        RECT 2773.870 31.520 2774.190 31.580 ;
        RECT 272.390 31.380 2774.190 31.520 ;
        RECT 272.390 31.320 272.710 31.380 ;
        RECT 2773.870 31.320 2774.190 31.380 ;
      LAYER via ;
        RECT 272.420 896.960 272.680 897.220 ;
        RECT 296.800 896.960 297.060 897.220 ;
        RECT 272.420 31.320 272.680 31.580 ;
        RECT 2773.900 31.320 2774.160 31.580 ;
      LAYER met2 ;
        RECT 296.790 897.755 297.070 898.125 ;
        RECT 296.860 897.250 297.000 897.755 ;
        RECT 272.420 896.930 272.680 897.250 ;
        RECT 296.800 896.930 297.060 897.250 ;
        RECT 272.480 31.610 272.620 896.930 ;
        RECT 272.420 31.290 272.680 31.610 ;
        RECT 2773.900 31.290 2774.160 31.610 ;
        RECT 2773.960 2.400 2774.100 31.290 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
      LAYER via2 ;
        RECT 296.790 897.800 297.070 898.080 ;
      LAYER met3 ;
        RECT 296.765 898.090 297.095 898.105 ;
        RECT 310.000 898.090 314.000 898.480 ;
        RECT 296.765 897.880 314.000 898.090 ;
        RECT 296.765 897.790 310.500 897.880 ;
        RECT 296.765 897.775 297.095 897.790 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 260.430 2415.260 260.750 2415.320 ;
        RECT 296.770 2415.260 297.090 2415.320 ;
        RECT 260.430 2415.120 297.090 2415.260 ;
        RECT 260.430 2415.060 260.750 2415.120 ;
        RECT 296.770 2415.060 297.090 2415.120 ;
        RECT 260.430 31.180 260.750 31.240 ;
        RECT 2791.810 31.180 2792.130 31.240 ;
        RECT 260.430 31.040 2792.130 31.180 ;
        RECT 260.430 30.980 260.750 31.040 ;
        RECT 2791.810 30.980 2792.130 31.040 ;
      LAYER via ;
        RECT 260.460 2415.060 260.720 2415.320 ;
        RECT 296.800 2415.060 297.060 2415.320 ;
        RECT 260.460 30.980 260.720 31.240 ;
        RECT 2791.840 30.980 2792.100 31.240 ;
      LAYER met2 ;
        RECT 296.790 2419.595 297.070 2419.965 ;
        RECT 296.860 2415.350 297.000 2419.595 ;
        RECT 260.460 2415.030 260.720 2415.350 ;
        RECT 296.800 2415.030 297.060 2415.350 ;
        RECT 260.520 31.270 260.660 2415.030 ;
        RECT 260.460 30.950 260.720 31.270 ;
        RECT 2791.840 30.950 2792.100 31.270 ;
        RECT 2791.900 2.400 2792.040 30.950 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
      LAYER via2 ;
        RECT 296.790 2419.640 297.070 2419.920 ;
      LAYER met3 ;
        RECT 296.765 2419.930 297.095 2419.945 ;
        RECT 310.000 2419.930 314.000 2420.320 ;
        RECT 296.765 2419.720 314.000 2419.930 ;
        RECT 296.765 2419.630 310.500 2419.720 ;
        RECT 296.765 2419.615 297.095 2419.630 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.770 30.755 2810.050 31.125 ;
        RECT 2809.840 2.400 2809.980 30.755 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
      LAYER via2 ;
        RECT 2809.770 30.800 2810.050 31.080 ;
      LAYER met3 ;
        RECT 310.000 2313.640 314.000 2314.240 ;
        RECT 246.830 2311.810 247.210 2311.820 ;
        RECT 310.350 2311.810 310.650 2313.640 ;
        RECT 246.830 2311.510 310.650 2311.810 ;
        RECT 246.830 2311.500 247.210 2311.510 ;
        RECT 246.830 31.090 247.210 31.100 ;
        RECT 2809.745 31.090 2810.075 31.105 ;
        RECT 246.830 30.790 2810.075 31.090 ;
        RECT 246.830 30.780 247.210 30.790 ;
        RECT 2809.745 30.775 2810.075 30.790 ;
      LAYER via3 ;
        RECT 246.860 2311.500 247.180 2311.820 ;
        RECT 246.860 30.780 247.180 31.100 ;
      LAYER met4 ;
        RECT 246.855 2311.495 247.185 2311.825 ;
        RECT 246.870 31.105 247.170 2311.495 ;
        RECT 246.855 30.775 247.185 31.105 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2711.385 1690.565 2712.475 1690.735 ;
      LAYER mcon ;
        RECT 2712.305 1690.565 2712.475 1690.735 ;
      LAYER met1 ;
        RECT 2615.170 1690.720 2615.490 1690.780 ;
        RECT 2711.325 1690.720 2711.615 1690.765 ;
        RECT 2615.170 1690.580 2711.615 1690.720 ;
        RECT 2615.170 1690.520 2615.490 1690.580 ;
        RECT 2711.325 1690.535 2711.615 1690.580 ;
        RECT 2712.245 1690.720 2712.535 1690.765 ;
        RECT 2822.170 1690.720 2822.490 1690.780 ;
        RECT 2712.245 1690.580 2822.490 1690.720 ;
        RECT 2712.245 1690.535 2712.535 1690.580 ;
        RECT 2822.170 1690.520 2822.490 1690.580 ;
        RECT 2822.170 62.120 2822.490 62.180 ;
        RECT 2827.690 62.120 2828.010 62.180 ;
        RECT 2822.170 61.980 2828.010 62.120 ;
        RECT 2822.170 61.920 2822.490 61.980 ;
        RECT 2827.690 61.920 2828.010 61.980 ;
      LAYER via ;
        RECT 2615.200 1690.520 2615.460 1690.780 ;
        RECT 2822.200 1690.520 2822.460 1690.780 ;
        RECT 2822.200 61.920 2822.460 62.180 ;
        RECT 2827.720 61.920 2827.980 62.180 ;
      LAYER met2 ;
        RECT 2615.190 1690.635 2615.470 1691.005 ;
        RECT 2615.200 1690.490 2615.460 1690.635 ;
        RECT 2822.200 1690.490 2822.460 1690.810 ;
        RECT 2822.260 62.210 2822.400 1690.490 ;
        RECT 2822.200 61.890 2822.460 62.210 ;
        RECT 2827.720 61.890 2827.980 62.210 ;
        RECT 2827.780 2.400 2827.920 61.890 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1690.680 2615.470 1690.960 ;
      LAYER met3 ;
        RECT 2606.000 1690.970 2610.000 1691.360 ;
        RECT 2615.165 1690.970 2615.495 1690.985 ;
        RECT 2606.000 1690.760 2615.495 1690.970 ;
        RECT 2609.580 1690.670 2615.495 1690.760 ;
        RECT 2615.165 1690.655 2615.495 1690.670 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 251.230 959.380 251.550 959.440 ;
        RECT 296.770 959.380 297.090 959.440 ;
        RECT 251.230 959.240 297.090 959.380 ;
        RECT 251.230 959.180 251.550 959.240 ;
        RECT 296.770 959.180 297.090 959.240 ;
        RECT 251.230 30.840 251.550 30.900 ;
        RECT 2845.170 30.840 2845.490 30.900 ;
        RECT 251.230 30.700 2845.490 30.840 ;
        RECT 251.230 30.640 251.550 30.700 ;
        RECT 2845.170 30.640 2845.490 30.700 ;
      LAYER via ;
        RECT 251.260 959.180 251.520 959.440 ;
        RECT 296.800 959.180 297.060 959.440 ;
        RECT 251.260 30.640 251.520 30.900 ;
        RECT 2845.200 30.640 2845.460 30.900 ;
      LAYER met2 ;
        RECT 296.790 960.315 297.070 960.685 ;
        RECT 296.860 959.470 297.000 960.315 ;
        RECT 251.260 959.150 251.520 959.470 ;
        RECT 296.800 959.150 297.060 959.470 ;
        RECT 251.320 30.930 251.460 959.150 ;
        RECT 251.260 30.610 251.520 30.930 ;
        RECT 2845.200 30.610 2845.460 30.930 ;
        RECT 2845.260 2.400 2845.400 30.610 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
      LAYER via2 ;
        RECT 296.790 960.360 297.070 960.640 ;
      LAYER met3 ;
        RECT 296.765 960.650 297.095 960.665 ;
        RECT 310.000 960.650 314.000 961.040 ;
        RECT 296.765 960.440 314.000 960.650 ;
        RECT 296.765 960.350 310.500 960.440 ;
        RECT 296.765 960.335 297.095 960.350 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 484.400 2615.490 484.460 ;
        RECT 2646.450 484.400 2646.770 484.460 ;
        RECT 2615.170 484.260 2646.770 484.400 ;
        RECT 2615.170 484.200 2615.490 484.260 ;
        RECT 2646.450 484.200 2646.770 484.260 ;
        RECT 2646.450 17.580 2646.770 17.640 ;
        RECT 2863.110 17.580 2863.430 17.640 ;
        RECT 2646.450 17.440 2863.430 17.580 ;
        RECT 2646.450 17.380 2646.770 17.440 ;
        RECT 2863.110 17.380 2863.430 17.440 ;
      LAYER via ;
        RECT 2615.200 484.200 2615.460 484.460 ;
        RECT 2646.480 484.200 2646.740 484.460 ;
        RECT 2646.480 17.380 2646.740 17.640 ;
        RECT 2863.140 17.380 2863.400 17.640 ;
      LAYER met2 ;
        RECT 2615.190 485.675 2615.470 486.045 ;
        RECT 2615.260 484.490 2615.400 485.675 ;
        RECT 2615.200 484.170 2615.460 484.490 ;
        RECT 2646.480 484.170 2646.740 484.490 ;
        RECT 2646.540 17.670 2646.680 484.170 ;
        RECT 2646.480 17.350 2646.740 17.670 ;
        RECT 2863.140 17.350 2863.400 17.670 ;
        RECT 2863.200 2.400 2863.340 17.350 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
      LAYER via2 ;
        RECT 2615.190 485.720 2615.470 486.000 ;
      LAYER met3 ;
        RECT 2606.000 486.010 2610.000 486.400 ;
        RECT 2615.165 486.010 2615.495 486.025 ;
        RECT 2606.000 485.800 2615.495 486.010 ;
        RECT 2609.580 485.710 2615.495 485.800 ;
        RECT 2615.165 485.695 2615.495 485.710 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2684.200 2615.490 2684.260 ;
        RECT 2804.690 2684.200 2805.010 2684.260 ;
        RECT 2615.170 2684.060 2805.010 2684.200 ;
        RECT 2615.170 2684.000 2615.490 2684.060 ;
        RECT 2804.690 2684.000 2805.010 2684.060 ;
        RECT 2881.050 17.240 2881.370 17.300 ;
        RECT 2820.420 17.100 2881.370 17.240 ;
        RECT 2804.690 16.560 2805.010 16.620 ;
        RECT 2820.420 16.560 2820.560 17.100 ;
        RECT 2881.050 17.040 2881.370 17.100 ;
        RECT 2804.690 16.420 2820.560 16.560 ;
        RECT 2804.690 16.360 2805.010 16.420 ;
      LAYER via ;
        RECT 2615.200 2684.000 2615.460 2684.260 ;
        RECT 2804.720 2684.000 2804.980 2684.260 ;
        RECT 2804.720 16.360 2804.980 16.620 ;
        RECT 2881.080 17.040 2881.340 17.300 ;
      LAYER met2 ;
        RECT 2615.190 2684.795 2615.470 2685.165 ;
        RECT 2615.260 2684.290 2615.400 2684.795 ;
        RECT 2615.200 2683.970 2615.460 2684.290 ;
        RECT 2804.720 2683.970 2804.980 2684.290 ;
        RECT 2804.780 16.650 2804.920 2683.970 ;
        RECT 2881.080 17.010 2881.340 17.330 ;
        RECT 2804.720 16.330 2804.980 16.650 ;
        RECT 2881.140 2.400 2881.280 17.010 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2684.840 2615.470 2685.120 ;
      LAYER met3 ;
        RECT 2606.000 2685.130 2610.000 2685.520 ;
        RECT 2615.165 2685.130 2615.495 2685.145 ;
        RECT 2606.000 2684.920 2615.495 2685.130 ;
        RECT 2609.580 2684.830 2615.495 2684.920 ;
        RECT 2615.165 2684.815 2615.495 2684.830 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2898.070 2.960 2898.390 3.020 ;
        RECT 2898.990 2.960 2899.310 3.020 ;
        RECT 2898.070 2.820 2899.310 2.960 ;
        RECT 2898.070 2.760 2898.390 2.820 ;
        RECT 2898.990 2.760 2899.310 2.820 ;
      LAYER via ;
        RECT 2898.100 2.760 2898.360 3.020 ;
        RECT 2899.020 2.760 2899.280 3.020 ;
      LAYER met2 ;
        RECT 2898.090 57.955 2898.370 58.325 ;
        RECT 2898.160 3.050 2898.300 57.955 ;
        RECT 2898.100 2.730 2898.360 3.050 ;
        RECT 2899.020 2.730 2899.280 3.050 ;
        RECT 2899.080 2.400 2899.220 2.730 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 2898.090 58.000 2898.370 58.280 ;
      LAYER met3 ;
        RECT 303.870 3075.450 304.250 3075.460 ;
        RECT 310.000 3075.450 314.000 3075.840 ;
        RECT 303.870 3075.240 314.000 3075.450 ;
        RECT 303.870 3075.150 310.500 3075.240 ;
        RECT 303.870 3075.140 304.250 3075.150 ;
        RECT 303.870 58.290 304.250 58.300 ;
        RECT 2898.065 58.290 2898.395 58.305 ;
        RECT 303.870 57.990 2898.395 58.290 ;
        RECT 303.870 57.980 304.250 57.990 ;
        RECT 2898.065 57.975 2898.395 57.990 ;
      LAYER via3 ;
        RECT 303.900 3075.140 304.220 3075.460 ;
        RECT 303.900 57.980 304.220 58.300 ;
      LAYER met4 ;
        RECT 303.895 3075.135 304.225 3075.465 ;
        RECT 303.910 58.305 304.210 3075.135 ;
        RECT 303.895 57.975 304.225 58.305 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 846.930 2.960 847.250 3.020 ;
        RECT 848.310 2.960 848.630 3.020 ;
        RECT 846.930 2.820 848.630 2.960 ;
        RECT 846.930 2.760 847.250 2.820 ;
        RECT 848.310 2.760 848.630 2.820 ;
      LAYER via ;
        RECT 846.960 2.760 847.220 3.020 ;
        RECT 848.340 2.760 848.600 3.020 ;
      LAYER met2 ;
        RECT 2564.130 3275.035 2564.410 3275.405 ;
        RECT 2564.200 3260.000 2564.340 3275.035 ;
        RECT 2564.090 3256.000 2564.370 3260.000 ;
        RECT 848.330 251.075 848.610 251.445 ;
        RECT 848.400 3.050 848.540 251.075 ;
        RECT 846.960 2.730 847.220 3.050 ;
        RECT 848.340 2.730 848.600 3.050 ;
        RECT 847.020 2.400 847.160 2.730 ;
        RECT 846.810 -4.800 847.370 2.400 ;
      LAYER via2 ;
        RECT 2564.130 3275.080 2564.410 3275.360 ;
        RECT 848.330 251.120 848.610 251.400 ;
      LAYER met3 ;
        RECT 2564.105 3275.370 2564.435 3275.385 ;
        RECT 2664.590 3275.370 2664.970 3275.380 ;
        RECT 2564.105 3275.070 2664.970 3275.370 ;
        RECT 2564.105 3275.055 2564.435 3275.070 ;
        RECT 2664.590 3275.060 2664.970 3275.070 ;
        RECT 848.305 251.410 848.635 251.425 ;
        RECT 2664.590 251.410 2664.970 251.420 ;
        RECT 848.305 251.110 2664.970 251.410 ;
        RECT 848.305 251.095 848.635 251.110 ;
        RECT 2664.590 251.100 2664.970 251.110 ;
      LAYER via3 ;
        RECT 2664.620 3275.060 2664.940 3275.380 ;
        RECT 2664.620 251.100 2664.940 251.420 ;
      LAYER met4 ;
        RECT 2664.615 3275.055 2664.945 3275.385 ;
        RECT 2664.630 251.425 2664.930 3275.055 ;
        RECT 2664.615 251.095 2664.945 251.425 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.010 190.300 869.330 190.360 ;
        RECT 966.070 190.300 966.390 190.360 ;
        RECT 869.010 190.160 966.390 190.300 ;
        RECT 869.010 190.100 869.330 190.160 ;
        RECT 966.070 190.100 966.390 190.160 ;
        RECT 864.870 20.640 865.190 20.700 ;
        RECT 869.010 20.640 869.330 20.700 ;
        RECT 864.870 20.500 869.330 20.640 ;
        RECT 864.870 20.440 865.190 20.500 ;
        RECT 869.010 20.440 869.330 20.500 ;
      LAYER via ;
        RECT 869.040 190.100 869.300 190.360 ;
        RECT 966.100 190.100 966.360 190.360 ;
        RECT 864.900 20.440 865.160 20.700 ;
        RECT 869.040 20.440 869.300 20.700 ;
      LAYER met2 ;
        RECT 969.730 260.170 970.010 264.000 ;
        RECT 966.160 260.030 970.010 260.170 ;
        RECT 966.160 190.390 966.300 260.030 ;
        RECT 969.730 260.000 970.010 260.030 ;
        RECT 869.040 190.070 869.300 190.390 ;
        RECT 966.100 190.070 966.360 190.390 ;
        RECT 869.100 20.730 869.240 190.070 ;
        RECT 864.900 20.410 865.160 20.730 ;
        RECT 869.040 20.410 869.300 20.730 ;
        RECT 864.960 2.400 865.100 20.410 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.350 79.460 882.670 79.520 ;
        RECT 924.670 79.460 924.990 79.520 ;
        RECT 882.350 79.320 924.990 79.460 ;
        RECT 882.350 79.260 882.670 79.320 ;
        RECT 924.670 79.260 924.990 79.320 ;
      LAYER via ;
        RECT 882.380 79.260 882.640 79.520 ;
        RECT 924.700 79.260 924.960 79.520 ;
      LAYER met2 ;
        RECT 927.410 260.170 927.690 264.000 ;
        RECT 924.760 260.030 927.690 260.170 ;
        RECT 924.760 79.550 924.900 260.030 ;
        RECT 927.410 260.000 927.690 260.030 ;
        RECT 882.380 79.230 882.640 79.550 ;
        RECT 924.700 79.230 924.960 79.550 ;
        RECT 882.440 15.370 882.580 79.230 ;
        RECT 882.440 15.230 883.040 15.370 ;
        RECT 882.900 2.400 883.040 15.230 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 378.265 3254.905 378.435 3255.755 ;
        RECT 393.445 3254.905 393.615 3255.755 ;
        RECT 603.665 3254.905 603.835 3256.775 ;
        RECT 627.585 3255.585 627.755 3256.775 ;
        RECT 628.045 3255.245 628.215 3256.435 ;
        RECT 675.885 3254.905 676.055 3256.435 ;
        RECT 966.145 3254.905 966.315 3255.755 ;
      LAYER mcon ;
        RECT 603.665 3256.605 603.835 3256.775 ;
        RECT 378.265 3255.585 378.435 3255.755 ;
        RECT 393.445 3255.585 393.615 3255.755 ;
        RECT 627.585 3256.605 627.755 3256.775 ;
        RECT 628.045 3256.265 628.215 3256.435 ;
        RECT 675.885 3256.265 676.055 3256.435 ;
        RECT 966.145 3255.585 966.315 3255.755 ;
      LAYER met1 ;
        RECT 603.605 3256.760 603.895 3256.805 ;
        RECT 627.525 3256.760 627.815 3256.805 ;
        RECT 603.605 3256.620 627.815 3256.760 ;
        RECT 603.605 3256.575 603.895 3256.620 ;
        RECT 627.525 3256.575 627.815 3256.620 ;
        RECT 627.985 3256.420 628.275 3256.465 ;
        RECT 675.825 3256.420 676.115 3256.465 ;
        RECT 627.985 3256.280 676.115 3256.420 ;
        RECT 627.985 3256.235 628.275 3256.280 ;
        RECT 675.825 3256.235 676.115 3256.280 ;
        RECT 1063.130 3256.220 1063.450 3256.480 ;
        RECT 1063.220 3256.080 1063.360 3256.220 ;
        RECT 1028.260 3255.940 1063.360 3256.080 ;
        RECT 378.205 3255.740 378.495 3255.785 ;
        RECT 278.920 3255.600 378.495 3255.740 ;
        RECT 253.530 3255.400 253.850 3255.460 ;
        RECT 278.920 3255.400 279.060 3255.600 ;
        RECT 378.205 3255.555 378.495 3255.600 ;
        RECT 393.385 3255.740 393.675 3255.785 ;
        RECT 393.385 3255.600 472.720 3255.740 ;
        RECT 393.385 3255.555 393.675 3255.600 ;
        RECT 253.530 3255.260 279.060 3255.400 ;
        RECT 253.530 3255.200 253.850 3255.260 ;
        RECT 378.205 3255.060 378.495 3255.105 ;
        RECT 393.385 3255.060 393.675 3255.105 ;
        RECT 378.205 3254.920 393.675 3255.060 ;
        RECT 472.580 3255.060 472.720 3255.600 ;
        RECT 520.880 3255.600 569.320 3255.740 ;
        RECT 520.880 3255.060 521.020 3255.600 ;
        RECT 472.580 3254.920 521.020 3255.060 ;
        RECT 569.180 3255.060 569.320 3255.600 ;
        RECT 627.525 3255.555 627.815 3255.785 ;
        RECT 966.085 3255.740 966.375 3255.785 ;
        RECT 1028.260 3255.740 1028.400 3255.940 ;
        RECT 714.080 3255.600 762.520 3255.740 ;
        RECT 627.600 3255.400 627.740 3255.555 ;
        RECT 627.985 3255.400 628.275 3255.445 ;
        RECT 627.600 3255.260 628.275 3255.400 ;
        RECT 627.985 3255.215 628.275 3255.260 ;
        RECT 603.605 3255.060 603.895 3255.105 ;
        RECT 569.180 3254.920 603.895 3255.060 ;
        RECT 378.205 3254.875 378.495 3254.920 ;
        RECT 393.385 3254.875 393.675 3254.920 ;
        RECT 603.605 3254.875 603.895 3254.920 ;
        RECT 675.825 3255.060 676.115 3255.105 ;
        RECT 714.080 3255.060 714.220 3255.600 ;
        RECT 675.825 3254.920 714.220 3255.060 ;
        RECT 762.380 3255.060 762.520 3255.600 ;
        RECT 810.680 3255.600 859.120 3255.740 ;
        RECT 810.680 3255.060 810.820 3255.600 ;
        RECT 762.380 3254.920 810.820 3255.060 ;
        RECT 858.980 3255.060 859.120 3255.600 ;
        RECT 966.085 3255.600 1028.400 3255.740 ;
        RECT 966.085 3255.555 966.375 3255.600 ;
        RECT 907.280 3255.260 931.800 3255.400 ;
        RECT 907.280 3255.060 907.420 3255.260 ;
        RECT 858.980 3254.920 907.420 3255.060 ;
        RECT 931.660 3255.060 931.800 3255.260 ;
        RECT 966.085 3255.060 966.375 3255.105 ;
        RECT 931.660 3254.920 966.375 3255.060 ;
        RECT 675.825 3254.875 676.115 3254.920 ;
        RECT 966.085 3254.875 966.375 3254.920 ;
        RECT 253.530 251.840 253.850 251.900 ;
        RECT 897.530 251.840 897.850 251.900 ;
        RECT 253.530 251.700 897.850 251.840 ;
        RECT 253.530 251.640 253.850 251.700 ;
        RECT 897.530 251.640 897.850 251.700 ;
        RECT 897.530 20.640 897.850 20.700 ;
        RECT 900.750 20.640 901.070 20.700 ;
        RECT 897.530 20.500 901.070 20.640 ;
        RECT 897.530 20.440 897.850 20.500 ;
        RECT 900.750 20.440 901.070 20.500 ;
      LAYER via ;
        RECT 1063.160 3256.220 1063.420 3256.480 ;
        RECT 253.560 3255.200 253.820 3255.460 ;
        RECT 253.560 251.640 253.820 251.900 ;
        RECT 897.560 251.640 897.820 251.900 ;
        RECT 897.560 20.440 897.820 20.700 ;
        RECT 900.780 20.440 901.040 20.700 ;
      LAYER met2 ;
        RECT 1062.650 3256.930 1062.930 3260.000 ;
        RECT 1062.650 3256.790 1063.360 3256.930 ;
        RECT 1062.650 3256.000 1062.930 3256.790 ;
        RECT 1063.220 3256.510 1063.360 3256.790 ;
        RECT 1063.160 3256.190 1063.420 3256.510 ;
        RECT 253.560 3255.170 253.820 3255.490 ;
        RECT 253.620 251.930 253.760 3255.170 ;
        RECT 253.560 251.610 253.820 251.930 ;
        RECT 897.560 251.610 897.820 251.930 ;
        RECT 897.620 20.730 897.760 251.610 ;
        RECT 897.560 20.410 897.820 20.730 ;
        RECT 900.780 20.410 901.040 20.730 ;
        RECT 900.840 2.400 900.980 20.410 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 225.930 2794.700 226.250 2794.760 ;
        RECT 296.770 2794.700 297.090 2794.760 ;
        RECT 225.930 2794.560 297.090 2794.700 ;
        RECT 225.930 2794.500 226.250 2794.560 ;
        RECT 296.770 2794.500 297.090 2794.560 ;
        RECT 225.930 24.720 226.250 24.780 ;
        RECT 918.690 24.720 919.010 24.780 ;
        RECT 225.930 24.580 919.010 24.720 ;
        RECT 225.930 24.520 226.250 24.580 ;
        RECT 918.690 24.520 919.010 24.580 ;
      LAYER via ;
        RECT 225.960 2794.500 226.220 2794.760 ;
        RECT 296.800 2794.500 297.060 2794.760 ;
        RECT 225.960 24.520 226.220 24.780 ;
        RECT 918.720 24.520 918.980 24.780 ;
      LAYER met2 ;
        RECT 296.790 2800.395 297.070 2800.765 ;
        RECT 296.860 2794.790 297.000 2800.395 ;
        RECT 225.960 2794.470 226.220 2794.790 ;
        RECT 296.800 2794.470 297.060 2794.790 ;
        RECT 226.020 24.810 226.160 2794.470 ;
        RECT 225.960 24.490 226.220 24.810 ;
        RECT 918.720 24.490 918.980 24.810 ;
        RECT 918.780 2.400 918.920 24.490 ;
        RECT 918.570 -4.800 919.130 2.400 ;
      LAYER via2 ;
        RECT 296.790 2800.440 297.070 2800.720 ;
      LAYER met3 ;
        RECT 296.765 2800.730 297.095 2800.745 ;
        RECT 310.000 2800.730 314.000 2801.120 ;
        RECT 296.765 2800.520 314.000 2800.730 ;
        RECT 296.765 2800.430 310.500 2800.520 ;
        RECT 296.765 2800.415 297.095 2800.430 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 931.645 48.365 931.815 96.475 ;
      LAYER mcon ;
        RECT 931.645 96.305 931.815 96.475 ;
      LAYER met1 ;
        RECT 498.710 244.020 499.030 244.080 ;
        RECT 503.310 244.020 503.630 244.080 ;
        RECT 498.710 243.880 503.630 244.020 ;
        RECT 498.710 243.820 499.030 243.880 ;
        RECT 503.310 243.820 503.630 243.880 ;
        RECT 503.310 121.960 503.630 122.020 ;
        RECT 931.570 121.960 931.890 122.020 ;
        RECT 503.310 121.820 931.890 121.960 ;
        RECT 503.310 121.760 503.630 121.820 ;
        RECT 931.570 121.760 931.890 121.820 ;
        RECT 931.570 96.460 931.890 96.520 ;
        RECT 931.375 96.320 931.890 96.460 ;
        RECT 931.570 96.260 931.890 96.320 ;
        RECT 931.585 48.520 931.875 48.565 ;
        RECT 936.170 48.520 936.490 48.580 ;
        RECT 931.585 48.380 936.490 48.520 ;
        RECT 931.585 48.335 931.875 48.380 ;
        RECT 936.170 48.320 936.490 48.380 ;
      LAYER via ;
        RECT 498.740 243.820 499.000 244.080 ;
        RECT 503.340 243.820 503.600 244.080 ;
        RECT 503.340 121.760 503.600 122.020 ;
        RECT 931.600 121.760 931.860 122.020 ;
        RECT 931.600 96.260 931.860 96.520 ;
        RECT 936.200 48.320 936.460 48.580 ;
      LAYER met2 ;
        RECT 498.690 260.000 498.970 264.000 ;
        RECT 498.800 244.110 498.940 260.000 ;
        RECT 498.740 243.790 499.000 244.110 ;
        RECT 503.340 243.790 503.600 244.110 ;
        RECT 503.400 122.050 503.540 243.790 ;
        RECT 503.340 121.730 503.600 122.050 ;
        RECT 931.600 121.730 931.860 122.050 ;
        RECT 931.660 96.550 931.800 121.730 ;
        RECT 931.600 96.230 931.860 96.550 ;
        RECT 936.200 48.290 936.460 48.610 ;
        RECT 936.260 2.400 936.400 48.290 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 353.350 3274.100 353.670 3274.160 ;
        RECT 690.990 3274.100 691.310 3274.160 ;
        RECT 353.350 3273.960 691.310 3274.100 ;
        RECT 353.350 3273.900 353.670 3273.960 ;
        RECT 690.990 3273.900 691.310 3273.960 ;
        RECT 306.890 3260.840 307.210 3260.900 ;
        RECT 353.350 3260.840 353.670 3260.900 ;
        RECT 306.890 3260.700 353.670 3260.840 ;
        RECT 306.890 3260.640 307.210 3260.700 ;
        RECT 353.350 3260.640 353.670 3260.700 ;
        RECT 268.250 382.740 268.570 382.800 ;
        RECT 306.890 382.740 307.210 382.800 ;
        RECT 268.250 382.600 307.210 382.740 ;
        RECT 268.250 382.540 268.570 382.600 ;
        RECT 306.890 382.540 307.210 382.600 ;
        RECT 268.250 43.760 268.570 43.820 ;
        RECT 954.110 43.760 954.430 43.820 ;
        RECT 268.250 43.620 954.430 43.760 ;
        RECT 268.250 43.560 268.570 43.620 ;
        RECT 954.110 43.560 954.430 43.620 ;
      LAYER via ;
        RECT 353.380 3273.900 353.640 3274.160 ;
        RECT 691.020 3273.900 691.280 3274.160 ;
        RECT 306.920 3260.640 307.180 3260.900 ;
        RECT 353.380 3260.640 353.640 3260.900 ;
        RECT 268.280 382.540 268.540 382.800 ;
        RECT 306.920 382.540 307.180 382.800 ;
        RECT 268.280 43.560 268.540 43.820 ;
        RECT 954.140 43.560 954.400 43.820 ;
      LAYER met2 ;
        RECT 353.380 3273.870 353.640 3274.190 ;
        RECT 691.020 3273.870 691.280 3274.190 ;
        RECT 353.440 3260.930 353.580 3273.870 ;
        RECT 306.920 3260.610 307.180 3260.930 ;
        RECT 353.380 3260.610 353.640 3260.930 ;
        RECT 306.980 382.830 307.120 3260.610 ;
        RECT 691.080 3260.000 691.220 3273.870 ;
        RECT 690.970 3256.000 691.250 3260.000 ;
        RECT 268.280 382.510 268.540 382.830 ;
        RECT 306.920 382.510 307.180 382.830 ;
        RECT 268.340 43.850 268.480 382.510 ;
        RECT 268.280 43.530 268.540 43.850 ;
        RECT 954.140 43.530 954.400 43.850 ;
        RECT 954.200 2.400 954.340 43.530 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 972.585 145.265 972.755 193.035 ;
        RECT 972.585 48.365 972.755 96.475 ;
      LAYER mcon ;
        RECT 972.585 192.865 972.755 193.035 ;
        RECT 972.585 96.305 972.755 96.475 ;
      LAYER met1 ;
        RECT 2615.170 291.960 2615.490 292.020 ;
        RECT 2645.990 291.960 2646.310 292.020 ;
        RECT 2615.170 291.820 2646.310 291.960 ;
        RECT 2615.170 291.760 2615.490 291.820 ;
        RECT 2645.990 291.760 2646.310 291.820 ;
        RECT 972.510 251.840 972.830 251.900 ;
        RECT 2645.990 251.840 2646.310 251.900 ;
        RECT 972.510 251.700 2646.310 251.840 ;
        RECT 972.510 251.640 972.830 251.700 ;
        RECT 2645.990 251.640 2646.310 251.700 ;
        RECT 972.510 193.020 972.830 193.080 ;
        RECT 972.315 192.880 972.830 193.020 ;
        RECT 972.510 192.820 972.830 192.880 ;
        RECT 972.510 145.420 972.830 145.480 ;
        RECT 972.315 145.280 972.830 145.420 ;
        RECT 972.510 145.220 972.830 145.280 ;
        RECT 971.590 144.740 971.910 144.800 ;
        RECT 972.510 144.740 972.830 144.800 ;
        RECT 971.590 144.600 972.830 144.740 ;
        RECT 971.590 144.540 971.910 144.600 ;
        RECT 972.510 144.540 972.830 144.600 ;
        RECT 972.510 96.460 972.830 96.520 ;
        RECT 972.315 96.320 972.830 96.460 ;
        RECT 972.510 96.260 972.830 96.320 ;
        RECT 972.510 48.520 972.830 48.580 ;
        RECT 972.315 48.380 972.830 48.520 ;
        RECT 972.510 48.320 972.830 48.380 ;
      LAYER via ;
        RECT 2615.200 291.760 2615.460 292.020 ;
        RECT 2646.020 291.760 2646.280 292.020 ;
        RECT 972.540 251.640 972.800 251.900 ;
        RECT 2646.020 251.640 2646.280 251.900 ;
        RECT 972.540 192.820 972.800 193.080 ;
        RECT 972.540 145.220 972.800 145.480 ;
        RECT 971.620 144.540 971.880 144.800 ;
        RECT 972.540 144.540 972.800 144.800 ;
        RECT 972.540 96.260 972.800 96.520 ;
        RECT 972.540 48.320 972.800 48.580 ;
      LAYER met2 ;
        RECT 2615.190 295.275 2615.470 295.645 ;
        RECT 2615.260 292.050 2615.400 295.275 ;
        RECT 2615.200 291.730 2615.460 292.050 ;
        RECT 2646.020 291.730 2646.280 292.050 ;
        RECT 2646.080 251.930 2646.220 291.730 ;
        RECT 972.540 251.610 972.800 251.930 ;
        RECT 2646.020 251.610 2646.280 251.930 ;
        RECT 972.600 241.130 972.740 251.610 ;
        RECT 972.600 240.990 973.200 241.130 ;
        RECT 973.060 194.325 973.200 240.990 ;
        RECT 972.990 193.955 973.270 194.325 ;
        RECT 972.530 193.275 972.810 193.645 ;
        RECT 972.600 193.110 972.740 193.275 ;
        RECT 972.540 192.790 972.800 193.110 ;
        RECT 972.540 145.190 972.800 145.510 ;
        RECT 972.600 144.830 972.740 145.190 ;
        RECT 971.620 144.510 971.880 144.830 ;
        RECT 972.540 144.510 972.800 144.830 ;
        RECT 971.680 97.085 971.820 144.510 ;
        RECT 971.610 96.715 971.890 97.085 ;
        RECT 972.530 96.715 972.810 97.085 ;
        RECT 972.600 96.550 972.740 96.715 ;
        RECT 972.540 96.230 972.800 96.550 ;
        RECT 972.540 48.290 972.800 48.610 ;
        RECT 972.600 14.010 972.740 48.290 ;
        RECT 972.600 13.870 973.200 14.010 ;
        RECT 973.060 13.330 973.200 13.870 ;
        RECT 972.140 13.190 973.200 13.330 ;
        RECT 972.140 2.400 972.280 13.190 ;
        RECT 971.930 -4.800 972.490 2.400 ;
      LAYER via2 ;
        RECT 2615.190 295.320 2615.470 295.600 ;
        RECT 972.990 194.000 973.270 194.280 ;
        RECT 972.530 193.320 972.810 193.600 ;
        RECT 971.610 96.760 971.890 97.040 ;
        RECT 972.530 96.760 972.810 97.040 ;
      LAYER met3 ;
        RECT 2606.000 295.610 2610.000 296.000 ;
        RECT 2615.165 295.610 2615.495 295.625 ;
        RECT 2606.000 295.400 2615.495 295.610 ;
        RECT 2609.580 295.310 2615.495 295.400 ;
        RECT 2615.165 295.295 2615.495 295.310 ;
        RECT 972.965 194.290 973.295 194.305 ;
        RECT 971.830 193.990 973.295 194.290 ;
        RECT 971.830 193.610 972.130 193.990 ;
        RECT 972.965 193.975 973.295 193.990 ;
        RECT 972.505 193.610 972.835 193.625 ;
        RECT 971.830 193.310 972.835 193.610 ;
        RECT 972.505 193.295 972.835 193.310 ;
        RECT 971.585 97.050 971.915 97.065 ;
        RECT 972.505 97.050 972.835 97.065 ;
        RECT 971.585 96.750 972.835 97.050 ;
        RECT 971.585 96.735 971.915 96.750 ;
        RECT 972.505 96.735 972.835 96.750 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.670 20.640 648.990 20.700 ;
        RECT 650.970 20.640 651.290 20.700 ;
        RECT 648.670 20.500 651.290 20.640 ;
        RECT 648.670 20.440 648.990 20.500 ;
        RECT 650.970 20.440 651.290 20.500 ;
      LAYER via ;
        RECT 648.700 20.440 648.960 20.700 ;
        RECT 651.000 20.440 651.260 20.700 ;
      LAYER met2 ;
        RECT 2133.570 3257.610 2133.850 3257.725 ;
        RECT 2135.370 3257.610 2135.650 3260.000 ;
        RECT 2133.570 3257.470 2135.650 3257.610 ;
        RECT 2133.570 3257.355 2133.850 3257.470 ;
        RECT 2135.370 3256.000 2135.650 3257.470 ;
        RECT 648.690 245.635 648.970 246.005 ;
        RECT 648.760 20.730 648.900 245.635 ;
        RECT 648.700 20.410 648.960 20.730 ;
        RECT 651.000 20.410 651.260 20.730 ;
        RECT 651.060 2.400 651.200 20.410 ;
        RECT 650.850 -4.800 651.410 2.400 ;
      LAYER via2 ;
        RECT 2133.570 3257.400 2133.850 3257.680 ;
        RECT 648.690 245.680 648.970 245.960 ;
      LAYER met3 ;
        RECT 271.670 3257.690 272.050 3257.700 ;
        RECT 2133.545 3257.690 2133.875 3257.705 ;
        RECT 271.670 3257.390 2133.875 3257.690 ;
        RECT 271.670 3257.380 272.050 3257.390 ;
        RECT 2133.545 3257.375 2133.875 3257.390 ;
        RECT 271.670 245.970 272.050 245.980 ;
        RECT 648.665 245.970 648.995 245.985 ;
        RECT 271.670 245.670 648.995 245.970 ;
        RECT 271.670 245.660 272.050 245.670 ;
        RECT 648.665 245.655 648.995 245.670 ;
      LAYER via3 ;
        RECT 271.700 3257.380 272.020 3257.700 ;
        RECT 271.700 245.660 272.020 245.980 ;
      LAYER met4 ;
        RECT 271.695 3257.375 272.025 3257.705 ;
        RECT 271.710 245.985 272.010 3257.375 ;
        RECT 271.695 245.655 272.025 245.985 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2617.930 1159.300 2618.250 1159.360 ;
        RECT 2660.250 1159.300 2660.570 1159.360 ;
        RECT 2617.930 1159.160 2660.570 1159.300 ;
        RECT 2617.930 1159.100 2618.250 1159.160 ;
        RECT 2660.250 1159.100 2660.570 1159.160 ;
        RECT 993.210 252.180 993.530 252.240 ;
        RECT 2660.250 252.180 2660.570 252.240 ;
        RECT 993.210 252.040 2660.570 252.180 ;
        RECT 993.210 251.980 993.530 252.040 ;
        RECT 2660.250 251.980 2660.570 252.040 ;
        RECT 989.990 20.640 990.310 20.700 ;
        RECT 993.210 20.640 993.530 20.700 ;
        RECT 989.990 20.500 993.530 20.640 ;
        RECT 989.990 20.440 990.310 20.500 ;
        RECT 993.210 20.440 993.530 20.500 ;
      LAYER via ;
        RECT 2617.960 1159.100 2618.220 1159.360 ;
        RECT 2660.280 1159.100 2660.540 1159.360 ;
        RECT 993.240 251.980 993.500 252.240 ;
        RECT 2660.280 251.980 2660.540 252.240 ;
        RECT 990.020 20.440 990.280 20.700 ;
        RECT 993.240 20.440 993.500 20.700 ;
      LAYER met2 ;
        RECT 2617.950 1162.955 2618.230 1163.325 ;
        RECT 2618.020 1159.390 2618.160 1162.955 ;
        RECT 2617.960 1159.070 2618.220 1159.390 ;
        RECT 2660.280 1159.070 2660.540 1159.390 ;
        RECT 2660.340 252.270 2660.480 1159.070 ;
        RECT 993.240 251.950 993.500 252.270 ;
        RECT 2660.280 251.950 2660.540 252.270 ;
        RECT 993.300 20.730 993.440 251.950 ;
        RECT 990.020 20.410 990.280 20.730 ;
        RECT 993.240 20.410 993.500 20.730 ;
        RECT 990.080 2.400 990.220 20.410 ;
        RECT 989.870 -4.800 990.430 2.400 ;
      LAYER via2 ;
        RECT 2617.950 1163.000 2618.230 1163.280 ;
      LAYER met3 ;
        RECT 2606.000 1163.290 2610.000 1163.680 ;
        RECT 2617.925 1163.290 2618.255 1163.305 ;
        RECT 2606.000 1163.080 2618.255 1163.290 ;
        RECT 2609.580 1162.990 2618.255 1163.080 ;
        RECT 2617.925 1162.975 2618.255 1162.990 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.930 24.720 1008.250 24.780 ;
        RECT 1966.570 24.720 1966.890 24.780 ;
        RECT 1007.930 24.580 1966.890 24.720 ;
        RECT 1007.930 24.520 1008.250 24.580 ;
        RECT 1966.570 24.520 1966.890 24.580 ;
      LAYER via ;
        RECT 1007.960 24.520 1008.220 24.780 ;
        RECT 1966.600 24.520 1966.860 24.780 ;
      LAYER met2 ;
        RECT 1970.690 260.170 1970.970 264.000 ;
        RECT 1966.660 260.030 1970.970 260.170 ;
        RECT 1966.660 24.810 1966.800 260.030 ;
        RECT 1970.690 260.000 1970.970 260.030 ;
        RECT 1007.960 24.490 1008.220 24.810 ;
        RECT 1966.600 24.490 1966.860 24.810 ;
        RECT 1008.020 2.960 1008.160 24.490 ;
        RECT 1007.560 2.820 1008.160 2.960 ;
        RECT 1007.560 2.400 1007.700 2.820 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 244.020 527.550 244.080 ;
        RECT 530.910 244.020 531.230 244.080 ;
        RECT 527.230 243.880 531.230 244.020 ;
        RECT 527.230 243.820 527.550 243.880 ;
        RECT 530.910 243.820 531.230 243.880 ;
        RECT 530.910 25.740 531.230 25.800 ;
        RECT 1025.410 25.740 1025.730 25.800 ;
        RECT 530.910 25.600 1025.730 25.740 ;
        RECT 530.910 25.540 531.230 25.600 ;
        RECT 1025.410 25.540 1025.730 25.600 ;
      LAYER via ;
        RECT 527.260 243.820 527.520 244.080 ;
        RECT 530.940 243.820 531.200 244.080 ;
        RECT 530.940 25.540 531.200 25.800 ;
        RECT 1025.440 25.540 1025.700 25.800 ;
      LAYER met2 ;
        RECT 527.210 260.000 527.490 264.000 ;
        RECT 527.320 244.110 527.460 260.000 ;
        RECT 527.260 243.790 527.520 244.110 ;
        RECT 530.940 243.790 531.200 244.110 ;
        RECT 531.000 25.830 531.140 243.790 ;
        RECT 530.940 25.510 531.200 25.830 ;
        RECT 1025.440 25.510 1025.700 25.830 ;
        RECT 1025.500 2.400 1025.640 25.510 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.350 15.540 1043.670 15.600 ;
        RECT 1048.410 15.540 1048.730 15.600 ;
        RECT 1043.350 15.400 1048.730 15.540 ;
        RECT 1043.350 15.340 1043.670 15.400 ;
        RECT 1048.410 15.340 1048.730 15.400 ;
      LAYER via ;
        RECT 1043.380 15.340 1043.640 15.600 ;
        RECT 1048.440 15.340 1048.700 15.600 ;
      LAYER met2 ;
        RECT 1048.430 251.755 1048.710 252.125 ;
        RECT 1048.500 15.630 1048.640 251.755 ;
        RECT 1043.380 15.310 1043.640 15.630 ;
        RECT 1048.440 15.310 1048.700 15.630 ;
        RECT 1043.440 2.400 1043.580 15.310 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
      LAYER via2 ;
        RECT 1048.430 251.800 1048.710 252.080 ;
      LAYER met3 ;
        RECT 2672.870 3087.010 2673.250 3087.020 ;
        RECT 2606.000 3086.120 2610.000 3086.720 ;
        RECT 2646.230 3086.710 2673.250 3087.010 ;
        RECT 2609.430 3085.650 2609.730 3086.120 ;
        RECT 2646.230 3085.650 2646.530 3086.710 ;
        RECT 2672.870 3086.700 2673.250 3086.710 ;
        RECT 2609.430 3085.350 2646.530 3085.650 ;
        RECT 1048.405 252.090 1048.735 252.105 ;
        RECT 2672.870 252.090 2673.250 252.100 ;
        RECT 1048.405 251.790 2673.250 252.090 ;
        RECT 1048.405 251.775 1048.735 251.790 ;
        RECT 2672.870 251.780 2673.250 251.790 ;
      LAYER via3 ;
        RECT 2672.900 3086.700 2673.220 3087.020 ;
        RECT 2672.900 251.780 2673.220 252.100 ;
      LAYER met4 ;
        RECT 2672.895 3086.695 2673.225 3087.025 ;
        RECT 2672.910 252.105 2673.210 3086.695 ;
        RECT 2672.895 251.775 2673.225 252.105 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1960.000 2615.490 1960.060 ;
        RECT 2665.770 1960.000 2666.090 1960.060 ;
        RECT 2615.170 1959.860 2666.090 1960.000 ;
        RECT 2615.170 1959.800 2615.490 1959.860 ;
        RECT 2665.770 1959.800 2666.090 1959.860 ;
        RECT 1062.210 252.520 1062.530 252.580 ;
        RECT 2665.770 252.520 2666.090 252.580 ;
        RECT 1062.210 252.380 2666.090 252.520 ;
        RECT 1062.210 252.320 1062.530 252.380 ;
        RECT 2665.770 252.320 2666.090 252.380 ;
      LAYER via ;
        RECT 2615.200 1959.800 2615.460 1960.060 ;
        RECT 2665.800 1959.800 2666.060 1960.060 ;
        RECT 1062.240 252.320 1062.500 252.580 ;
        RECT 2665.800 252.320 2666.060 252.580 ;
      LAYER met2 ;
        RECT 2615.190 1965.355 2615.470 1965.725 ;
        RECT 2615.260 1960.090 2615.400 1965.355 ;
        RECT 2615.200 1959.770 2615.460 1960.090 ;
        RECT 2665.800 1959.770 2666.060 1960.090 ;
        RECT 2665.860 252.610 2666.000 1959.770 ;
        RECT 1062.240 252.290 1062.500 252.610 ;
        RECT 2665.800 252.290 2666.060 252.610 ;
        RECT 1062.300 14.010 1062.440 252.290 ;
        RECT 1061.840 13.870 1062.440 14.010 ;
        RECT 1061.840 13.330 1061.980 13.870 ;
        RECT 1061.380 13.190 1061.980 13.330 ;
        RECT 1061.380 2.400 1061.520 13.190 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1965.400 2615.470 1965.680 ;
      LAYER met3 ;
        RECT 2606.000 1965.690 2610.000 1966.080 ;
        RECT 2615.165 1965.690 2615.495 1965.705 ;
        RECT 2606.000 1965.480 2615.495 1965.690 ;
        RECT 2609.580 1965.390 2615.495 1965.480 ;
        RECT 2615.165 1965.375 2615.495 1965.390 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2611.030 2387.720 2611.350 2387.780 ;
        RECT 2665.310 2387.720 2665.630 2387.780 ;
        RECT 2611.030 2387.580 2665.630 2387.720 ;
        RECT 2611.030 2387.520 2611.350 2387.580 ;
        RECT 2665.310 2387.520 2665.630 2387.580 ;
        RECT 1082.910 252.860 1083.230 252.920 ;
        RECT 2665.310 252.860 2665.630 252.920 ;
        RECT 1082.910 252.720 2665.630 252.860 ;
        RECT 1082.910 252.660 1083.230 252.720 ;
        RECT 2665.310 252.660 2665.630 252.720 ;
        RECT 1079.230 20.640 1079.550 20.700 ;
        RECT 1082.910 20.640 1083.230 20.700 ;
        RECT 1079.230 20.500 1083.230 20.640 ;
        RECT 1079.230 20.440 1079.550 20.500 ;
        RECT 1082.910 20.440 1083.230 20.500 ;
      LAYER via ;
        RECT 2611.060 2387.520 2611.320 2387.780 ;
        RECT 2665.340 2387.520 2665.600 2387.780 ;
        RECT 1082.940 252.660 1083.200 252.920 ;
        RECT 2665.340 252.660 2665.600 252.920 ;
        RECT 1079.260 20.440 1079.520 20.700 ;
        RECT 1082.940 20.440 1083.200 20.700 ;
      LAYER met2 ;
        RECT 2611.050 2388.315 2611.330 2388.685 ;
        RECT 2611.120 2387.810 2611.260 2388.315 ;
        RECT 2611.060 2387.490 2611.320 2387.810 ;
        RECT 2665.340 2387.490 2665.600 2387.810 ;
        RECT 2665.400 252.950 2665.540 2387.490 ;
        RECT 1082.940 252.630 1083.200 252.950 ;
        RECT 2665.340 252.630 2665.600 252.950 ;
        RECT 1083.000 20.730 1083.140 252.630 ;
        RECT 1079.260 20.410 1079.520 20.730 ;
        RECT 1082.940 20.410 1083.200 20.730 ;
        RECT 1079.320 2.400 1079.460 20.410 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
      LAYER via2 ;
        RECT 2611.050 2388.360 2611.330 2388.640 ;
      LAYER met3 ;
        RECT 2606.000 2388.650 2610.000 2389.040 ;
        RECT 2611.025 2388.650 2611.355 2388.665 ;
        RECT 2606.000 2388.440 2611.355 2388.650 ;
        RECT 2609.580 2388.350 2611.355 2388.440 ;
        RECT 2611.025 2388.335 2611.355 2388.350 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 3273.760 372.530 3273.820 ;
        RECT 933.870 3273.760 934.190 3273.820 ;
        RECT 372.210 3273.620 934.190 3273.760 ;
        RECT 372.210 3273.560 372.530 3273.620 ;
        RECT 933.870 3273.560 934.190 3273.620 ;
        RECT 226.850 3267.980 227.170 3268.040 ;
        RECT 372.210 3267.980 372.530 3268.040 ;
        RECT 226.850 3267.840 372.530 3267.980 ;
        RECT 226.850 3267.780 227.170 3267.840 ;
        RECT 372.210 3267.780 372.530 3267.840 ;
        RECT 226.850 61.780 227.170 61.840 ;
        RECT 1096.250 61.780 1096.570 61.840 ;
        RECT 226.850 61.640 1096.570 61.780 ;
        RECT 226.850 61.580 227.170 61.640 ;
        RECT 1096.250 61.580 1096.570 61.640 ;
      LAYER via ;
        RECT 372.240 3273.560 372.500 3273.820 ;
        RECT 933.900 3273.560 934.160 3273.820 ;
        RECT 226.880 3267.780 227.140 3268.040 ;
        RECT 372.240 3267.780 372.500 3268.040 ;
        RECT 226.880 61.580 227.140 61.840 ;
        RECT 1096.280 61.580 1096.540 61.840 ;
      LAYER met2 ;
        RECT 372.240 3273.530 372.500 3273.850 ;
        RECT 933.900 3273.530 934.160 3273.850 ;
        RECT 372.300 3268.070 372.440 3273.530 ;
        RECT 226.880 3267.750 227.140 3268.070 ;
        RECT 372.240 3267.750 372.500 3268.070 ;
        RECT 226.940 61.870 227.080 3267.750 ;
        RECT 933.960 3260.000 934.100 3273.530 ;
        RECT 933.850 3256.000 934.130 3260.000 ;
        RECT 226.880 61.550 227.140 61.870 ;
        RECT 1096.280 61.550 1096.540 61.870 ;
        RECT 1096.340 16.050 1096.480 61.550 ;
        RECT 1096.340 15.910 1096.940 16.050 ;
        RECT 1096.800 2.400 1096.940 15.910 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 305.050 142.020 305.370 142.080 ;
        RECT 1110.970 142.020 1111.290 142.080 ;
        RECT 305.050 141.880 1111.290 142.020 ;
        RECT 305.050 141.820 305.370 141.880 ;
        RECT 1110.970 141.820 1111.290 141.880 ;
        RECT 1110.970 2.960 1111.290 3.020 ;
        RECT 1114.650 2.960 1114.970 3.020 ;
        RECT 1110.970 2.820 1114.970 2.960 ;
        RECT 1110.970 2.760 1111.290 2.820 ;
        RECT 1114.650 2.760 1114.970 2.820 ;
      LAYER via ;
        RECT 305.080 141.820 305.340 142.080 ;
        RECT 1111.000 141.820 1111.260 142.080 ;
        RECT 1111.000 2.760 1111.260 3.020 ;
        RECT 1114.680 2.760 1114.940 3.020 ;
      LAYER met2 ;
        RECT 305.070 1848.395 305.350 1848.765 ;
        RECT 305.140 142.110 305.280 1848.395 ;
        RECT 305.080 141.790 305.340 142.110 ;
        RECT 1111.000 141.790 1111.260 142.110 ;
        RECT 1111.060 3.050 1111.200 141.790 ;
        RECT 1111.000 2.730 1111.260 3.050 ;
        RECT 1114.680 2.730 1114.940 3.050 ;
        RECT 1114.740 2.400 1114.880 2.730 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
      LAYER via2 ;
        RECT 305.070 1848.440 305.350 1848.720 ;
      LAYER met3 ;
        RECT 305.045 1848.730 305.375 1848.745 ;
        RECT 310.000 1848.730 314.000 1849.120 ;
        RECT 305.045 1848.520 314.000 1848.730 ;
        RECT 305.045 1848.430 310.500 1848.520 ;
        RECT 305.045 1848.415 305.375 1848.430 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 148.140 1138.430 148.200 ;
        RECT 2624.370 148.140 2624.690 148.200 ;
        RECT 1138.110 148.000 2624.690 148.140 ;
        RECT 1138.110 147.940 1138.430 148.000 ;
        RECT 2624.370 147.940 2624.690 148.000 ;
        RECT 1132.590 20.640 1132.910 20.700 ;
        RECT 1138.110 20.640 1138.430 20.700 ;
        RECT 1132.590 20.500 1138.430 20.640 ;
        RECT 1132.590 20.440 1132.910 20.500 ;
        RECT 1138.110 20.440 1138.430 20.500 ;
      LAYER via ;
        RECT 1138.140 147.940 1138.400 148.200 ;
        RECT 2624.400 147.940 2624.660 148.200 ;
        RECT 1132.620 20.440 1132.880 20.700 ;
        RECT 1138.140 20.440 1138.400 20.700 ;
      LAYER met2 ;
        RECT 2624.390 1141.195 2624.670 1141.565 ;
        RECT 2624.460 148.230 2624.600 1141.195 ;
        RECT 1138.140 147.910 1138.400 148.230 ;
        RECT 2624.400 147.910 2624.660 148.230 ;
        RECT 1138.200 20.730 1138.340 147.910 ;
        RECT 1132.620 20.410 1132.880 20.730 ;
        RECT 1138.140 20.410 1138.400 20.730 ;
        RECT 1132.680 2.400 1132.820 20.410 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
      LAYER via2 ;
        RECT 2624.390 1141.240 2624.670 1141.520 ;
      LAYER met3 ;
        RECT 2606.000 1141.530 2610.000 1141.920 ;
        RECT 2624.365 1141.530 2624.695 1141.545 ;
        RECT 2606.000 1141.320 2624.695 1141.530 ;
        RECT 2609.580 1141.230 2624.695 1141.320 ;
        RECT 2624.365 1141.215 2624.695 1141.230 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 314.250 3291.440 314.570 3291.500 ;
        RECT 833.590 3291.440 833.910 3291.500 ;
        RECT 314.250 3291.300 833.910 3291.440 ;
        RECT 314.250 3291.240 314.570 3291.300 ;
        RECT 833.590 3291.240 833.910 3291.300 ;
        RECT 259.050 500.040 259.370 500.100 ;
        RECT 314.250 500.040 314.570 500.100 ;
        RECT 259.050 499.900 314.570 500.040 ;
        RECT 259.050 499.840 259.370 499.900 ;
        RECT 314.250 499.840 314.570 499.900 ;
        RECT 259.050 61.440 259.370 61.500 ;
        RECT 1150.530 61.440 1150.850 61.500 ;
        RECT 259.050 61.300 1150.850 61.440 ;
        RECT 259.050 61.240 259.370 61.300 ;
        RECT 1150.530 61.240 1150.850 61.300 ;
      LAYER via ;
        RECT 314.280 3291.240 314.540 3291.500 ;
        RECT 833.620 3291.240 833.880 3291.500 ;
        RECT 259.080 499.840 259.340 500.100 ;
        RECT 314.280 499.840 314.540 500.100 ;
        RECT 259.080 61.240 259.340 61.500 ;
        RECT 1150.560 61.240 1150.820 61.500 ;
      LAYER met2 ;
        RECT 314.280 3291.210 314.540 3291.530 ;
        RECT 833.620 3291.210 833.880 3291.530 ;
        RECT 314.340 500.130 314.480 3291.210 ;
        RECT 833.680 3260.000 833.820 3291.210 ;
        RECT 833.570 3256.000 833.850 3260.000 ;
        RECT 259.080 499.810 259.340 500.130 ;
        RECT 314.280 499.810 314.540 500.130 ;
        RECT 259.140 61.530 259.280 499.810 ;
        RECT 259.080 61.210 259.340 61.530 ;
        RECT 1150.560 61.210 1150.820 61.530 ;
        RECT 1150.620 2.400 1150.760 61.210 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 245.250 2056.560 245.570 2056.620 ;
        RECT 296.770 2056.560 297.090 2056.620 ;
        RECT 245.250 2056.420 297.090 2056.560 ;
        RECT 245.250 2056.360 245.570 2056.420 ;
        RECT 296.770 2056.360 297.090 2056.420 ;
        RECT 245.250 30.160 245.570 30.220 ;
        RECT 668.910 30.160 669.230 30.220 ;
        RECT 245.250 30.020 669.230 30.160 ;
        RECT 245.250 29.960 245.570 30.020 ;
        RECT 668.910 29.960 669.230 30.020 ;
      LAYER via ;
        RECT 245.280 2056.360 245.540 2056.620 ;
        RECT 296.800 2056.360 297.060 2056.620 ;
        RECT 245.280 29.960 245.540 30.220 ;
        RECT 668.940 29.960 669.200 30.220 ;
      LAYER met2 ;
        RECT 296.790 2060.555 297.070 2060.925 ;
        RECT 296.860 2056.650 297.000 2060.555 ;
        RECT 245.280 2056.330 245.540 2056.650 ;
        RECT 296.800 2056.330 297.060 2056.650 ;
        RECT 245.340 30.250 245.480 2056.330 ;
        RECT 245.280 29.930 245.540 30.250 ;
        RECT 668.940 29.930 669.200 30.250 ;
        RECT 669.000 2.400 669.140 29.930 ;
        RECT 668.790 -4.800 669.350 2.400 ;
      LAYER via2 ;
        RECT 296.790 2060.600 297.070 2060.880 ;
      LAYER met3 ;
        RECT 296.765 2060.890 297.095 2060.905 ;
        RECT 310.000 2060.890 314.000 2061.280 ;
        RECT 296.765 2060.680 314.000 2060.890 ;
        RECT 296.765 2060.590 310.500 2060.680 ;
        RECT 296.765 2060.575 297.095 2060.590 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1084.750 244.020 1085.070 244.080 ;
        RECT 1089.810 244.020 1090.130 244.080 ;
        RECT 1084.750 243.880 1090.130 244.020 ;
        RECT 1084.750 243.820 1085.070 243.880 ;
        RECT 1089.810 243.820 1090.130 243.880 ;
        RECT 1089.810 226.340 1090.130 226.400 ;
        RECT 1166.170 226.340 1166.490 226.400 ;
        RECT 1089.810 226.200 1166.490 226.340 ;
        RECT 1089.810 226.140 1090.130 226.200 ;
        RECT 1166.170 226.140 1166.490 226.200 ;
        RECT 1166.170 62.120 1166.490 62.180 ;
        RECT 1168.470 62.120 1168.790 62.180 ;
        RECT 1166.170 61.980 1168.790 62.120 ;
        RECT 1166.170 61.920 1166.490 61.980 ;
        RECT 1168.470 61.920 1168.790 61.980 ;
      LAYER via ;
        RECT 1084.780 243.820 1085.040 244.080 ;
        RECT 1089.840 243.820 1090.100 244.080 ;
        RECT 1089.840 226.140 1090.100 226.400 ;
        RECT 1166.200 226.140 1166.460 226.400 ;
        RECT 1166.200 61.920 1166.460 62.180 ;
        RECT 1168.500 61.920 1168.760 62.180 ;
      LAYER met2 ;
        RECT 1084.730 260.000 1085.010 264.000 ;
        RECT 1084.840 244.110 1084.980 260.000 ;
        RECT 1084.780 243.790 1085.040 244.110 ;
        RECT 1089.840 243.790 1090.100 244.110 ;
        RECT 1089.900 226.430 1090.040 243.790 ;
        RECT 1089.840 226.110 1090.100 226.430 ;
        RECT 1166.200 226.110 1166.460 226.430 ;
        RECT 1166.260 62.210 1166.400 226.110 ;
        RECT 1166.200 61.890 1166.460 62.210 ;
        RECT 1168.500 61.890 1168.760 62.210 ;
        RECT 1168.560 2.400 1168.700 61.890 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.970 141.595 1186.250 141.965 ;
        RECT 1186.040 2.400 1186.180 141.595 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 1185.970 141.640 1186.250 141.920 ;
      LAYER met3 ;
        RECT 2606.000 3150.250 2610.000 3150.640 ;
        RECT 2622.270 3150.250 2622.650 3150.260 ;
        RECT 2606.000 3150.040 2622.650 3150.250 ;
        RECT 2609.580 3149.950 2622.650 3150.040 ;
        RECT 2622.270 3149.940 2622.650 3149.950 ;
        RECT 1185.945 141.930 1186.275 141.945 ;
        RECT 2622.270 141.930 2622.650 141.940 ;
        RECT 1185.945 141.630 2622.650 141.930 ;
        RECT 1185.945 141.615 1186.275 141.630 ;
        RECT 2622.270 141.620 2622.650 141.630 ;
      LAYER via3 ;
        RECT 2622.300 3149.940 2622.620 3150.260 ;
        RECT 2622.300 141.620 2622.620 141.940 ;
      LAYER met4 ;
        RECT 2622.295 3149.935 2622.625 3150.265 ;
        RECT 2622.310 141.945 2622.610 3149.935 ;
        RECT 2622.295 141.615 2622.625 141.945 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1711.460 2615.490 1711.520 ;
        RECT 2658.870 1711.460 2659.190 1711.520 ;
        RECT 2615.170 1711.320 2659.190 1711.460 ;
        RECT 2615.170 1711.260 2615.490 1711.320 ;
        RECT 2658.870 1711.260 2659.190 1711.320 ;
        RECT 1207.110 253.200 1207.430 253.260 ;
        RECT 2658.870 253.200 2659.190 253.260 ;
        RECT 1207.110 253.060 2659.190 253.200 ;
        RECT 1207.110 253.000 1207.430 253.060 ;
        RECT 2658.870 253.000 2659.190 253.060 ;
        RECT 1203.890 20.640 1204.210 20.700 ;
        RECT 1207.110 20.640 1207.430 20.700 ;
        RECT 1203.890 20.500 1207.430 20.640 ;
        RECT 1203.890 20.440 1204.210 20.500 ;
        RECT 1207.110 20.440 1207.430 20.500 ;
      LAYER via ;
        RECT 2615.200 1711.260 2615.460 1711.520 ;
        RECT 2658.900 1711.260 2659.160 1711.520 ;
        RECT 1207.140 253.000 1207.400 253.260 ;
        RECT 2658.900 253.000 2659.160 253.260 ;
        RECT 1203.920 20.440 1204.180 20.700 ;
        RECT 1207.140 20.440 1207.400 20.700 ;
      LAYER met2 ;
        RECT 2615.190 1712.395 2615.470 1712.765 ;
        RECT 2615.260 1711.550 2615.400 1712.395 ;
        RECT 2615.200 1711.230 2615.460 1711.550 ;
        RECT 2658.900 1711.230 2659.160 1711.550 ;
        RECT 2658.960 253.290 2659.100 1711.230 ;
        RECT 1207.140 252.970 1207.400 253.290 ;
        RECT 2658.900 252.970 2659.160 253.290 ;
        RECT 1207.200 20.730 1207.340 252.970 ;
        RECT 1203.920 20.410 1204.180 20.730 ;
        RECT 1207.140 20.410 1207.400 20.730 ;
        RECT 1203.980 2.400 1204.120 20.410 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1712.440 2615.470 1712.720 ;
      LAYER met3 ;
        RECT 2606.000 1712.730 2610.000 1713.120 ;
        RECT 2615.165 1712.730 2615.495 1712.745 ;
        RECT 2606.000 1712.520 2615.495 1712.730 ;
        RECT 2609.580 1712.430 2615.495 1712.520 ;
        RECT 2615.165 1712.415 2615.495 1712.430 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 223.630 490.180 223.950 490.240 ;
        RECT 296.770 490.180 297.090 490.240 ;
        RECT 223.630 490.040 297.090 490.180 ;
        RECT 223.630 489.980 223.950 490.040 ;
        RECT 296.770 489.980 297.090 490.040 ;
        RECT 223.630 61.100 223.950 61.160 ;
        RECT 1221.830 61.100 1222.150 61.160 ;
        RECT 223.630 60.960 1222.150 61.100 ;
        RECT 223.630 60.900 223.950 60.960 ;
        RECT 1221.830 60.900 1222.150 60.960 ;
      LAYER via ;
        RECT 223.660 489.980 223.920 490.240 ;
        RECT 296.800 489.980 297.060 490.240 ;
        RECT 223.660 60.900 223.920 61.160 ;
        RECT 1221.860 60.900 1222.120 61.160 ;
      LAYER met2 ;
        RECT 296.790 495.195 297.070 495.565 ;
        RECT 296.860 490.270 297.000 495.195 ;
        RECT 223.660 489.950 223.920 490.270 ;
        RECT 296.800 489.950 297.060 490.270 ;
        RECT 223.720 61.190 223.860 489.950 ;
        RECT 223.660 60.870 223.920 61.190 ;
        RECT 1221.860 60.870 1222.120 61.190 ;
        RECT 1221.920 2.400 1222.060 60.870 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
      LAYER via2 ;
        RECT 296.790 495.240 297.070 495.520 ;
      LAYER met3 ;
        RECT 296.765 495.530 297.095 495.545 ;
        RECT 310.000 495.530 314.000 495.920 ;
        RECT 296.765 495.320 314.000 495.530 ;
        RECT 296.765 495.230 310.500 495.320 ;
        RECT 296.765 495.215 297.095 495.230 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2643.060 2615.490 2643.120 ;
        RECT 2664.850 2643.060 2665.170 2643.120 ;
        RECT 2615.170 2642.920 2665.170 2643.060 ;
        RECT 2615.170 2642.860 2615.490 2642.920 ;
        RECT 2664.850 2642.860 2665.170 2642.920 ;
        RECT 1241.610 237.900 1241.930 237.960 ;
        RECT 2664.850 237.900 2665.170 237.960 ;
        RECT 1241.610 237.760 2665.170 237.900 ;
        RECT 1241.610 237.700 1241.930 237.760 ;
        RECT 2664.850 237.700 2665.170 237.760 ;
        RECT 1239.770 14.180 1240.090 14.240 ;
        RECT 1241.610 14.180 1241.930 14.240 ;
        RECT 1239.770 14.040 1241.930 14.180 ;
        RECT 1239.770 13.980 1240.090 14.040 ;
        RECT 1241.610 13.980 1241.930 14.040 ;
      LAYER via ;
        RECT 2615.200 2642.860 2615.460 2643.120 ;
        RECT 2664.880 2642.860 2665.140 2643.120 ;
        RECT 1241.640 237.700 1241.900 237.960 ;
        RECT 2664.880 237.700 2665.140 237.960 ;
        RECT 1239.800 13.980 1240.060 14.240 ;
        RECT 1241.640 13.980 1241.900 14.240 ;
      LAYER met2 ;
        RECT 2615.200 2643.005 2615.460 2643.150 ;
        RECT 2615.190 2642.635 2615.470 2643.005 ;
        RECT 2664.880 2642.830 2665.140 2643.150 ;
        RECT 2664.940 237.990 2665.080 2642.830 ;
        RECT 1241.640 237.670 1241.900 237.990 ;
        RECT 2664.880 237.670 2665.140 237.990 ;
        RECT 1241.700 14.270 1241.840 237.670 ;
        RECT 1239.800 13.950 1240.060 14.270 ;
        RECT 1241.640 13.950 1241.900 14.270 ;
        RECT 1239.860 2.400 1240.000 13.950 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2642.680 2615.470 2642.960 ;
      LAYER met3 ;
        RECT 2606.000 2642.970 2610.000 2643.360 ;
        RECT 2615.165 2642.970 2615.495 2642.985 ;
        RECT 2606.000 2642.760 2615.495 2642.970 ;
        RECT 2609.580 2642.670 2615.495 2642.760 ;
        RECT 2615.165 2642.655 2615.495 2642.670 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1257.250 20.640 1257.570 20.700 ;
        RECT 1262.310 20.640 1262.630 20.700 ;
        RECT 1257.250 20.500 1262.630 20.640 ;
        RECT 1257.250 20.440 1257.570 20.500 ;
        RECT 1262.310 20.440 1262.630 20.500 ;
      LAYER via ;
        RECT 1257.280 20.440 1257.540 20.700 ;
        RECT 1262.340 20.440 1262.600 20.700 ;
      LAYER met2 ;
        RECT 1820.770 3266.195 1821.050 3266.565 ;
        RECT 1820.840 3260.000 1820.980 3266.195 ;
        RECT 1820.730 3256.000 1821.010 3260.000 ;
        RECT 1262.330 230.675 1262.610 231.045 ;
        RECT 1262.400 20.730 1262.540 230.675 ;
        RECT 1257.280 20.410 1257.540 20.730 ;
        RECT 1262.340 20.410 1262.600 20.730 ;
        RECT 1257.340 2.400 1257.480 20.410 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
      LAYER via2 ;
        RECT 1820.770 3266.240 1821.050 3266.520 ;
        RECT 1262.330 230.720 1262.610 231.000 ;
      LAYER met3 ;
        RECT 1820.745 3266.530 1821.075 3266.545 ;
        RECT 2608.470 3266.530 2608.850 3266.540 ;
        RECT 1820.745 3266.230 2608.850 3266.530 ;
        RECT 1820.745 3266.215 1821.075 3266.230 ;
        RECT 2608.470 3266.220 2608.850 3266.230 ;
        RECT 1262.305 231.010 1262.635 231.025 ;
        RECT 2608.470 231.010 2608.850 231.020 ;
        RECT 1262.305 230.710 2608.850 231.010 ;
        RECT 1262.305 230.695 1262.635 230.710 ;
        RECT 2608.470 230.700 2608.850 230.710 ;
      LAYER via3 ;
        RECT 2608.500 3266.220 2608.820 3266.540 ;
        RECT 2608.500 230.700 2608.820 231.020 ;
      LAYER met4 ;
        RECT 2608.495 3266.215 2608.825 3266.545 ;
        RECT 2608.510 231.025 2608.810 3266.215 ;
        RECT 2608.495 230.695 2608.825 231.025 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 252.610 2394.520 252.930 2394.580 ;
        RECT 296.770 2394.520 297.090 2394.580 ;
        RECT 252.610 2394.380 297.090 2394.520 ;
        RECT 252.610 2394.320 252.930 2394.380 ;
        RECT 296.770 2394.320 297.090 2394.380 ;
        RECT 252.610 33.900 252.930 33.960 ;
        RECT 1275.190 33.900 1275.510 33.960 ;
        RECT 252.610 33.760 1275.510 33.900 ;
        RECT 252.610 33.700 252.930 33.760 ;
        RECT 1275.190 33.700 1275.510 33.760 ;
      LAYER via ;
        RECT 252.640 2394.320 252.900 2394.580 ;
        RECT 296.800 2394.320 297.060 2394.580 ;
        RECT 252.640 33.700 252.900 33.960 ;
        RECT 1275.220 33.700 1275.480 33.960 ;
      LAYER met2 ;
        RECT 296.790 2397.835 297.070 2398.205 ;
        RECT 296.860 2394.610 297.000 2397.835 ;
        RECT 252.640 2394.290 252.900 2394.610 ;
        RECT 296.800 2394.290 297.060 2394.610 ;
        RECT 252.700 33.990 252.840 2394.290 ;
        RECT 252.640 33.670 252.900 33.990 ;
        RECT 1275.220 33.670 1275.480 33.990 ;
        RECT 1275.280 2.400 1275.420 33.670 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
      LAYER via2 ;
        RECT 296.790 2397.880 297.070 2398.160 ;
      LAYER met3 ;
        RECT 296.765 2398.170 297.095 2398.185 ;
        RECT 310.000 2398.170 314.000 2398.560 ;
        RECT 296.765 2397.960 314.000 2398.170 ;
        RECT 296.765 2397.870 310.500 2397.960 ;
        RECT 296.765 2397.855 297.095 2397.870 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1290.445 48.365 1290.615 96.475 ;
      LAYER mcon ;
        RECT 1290.445 96.305 1290.615 96.475 ;
      LAYER met1 ;
        RECT 1261.850 145.080 1262.170 145.140 ;
        RECT 1290.370 145.080 1290.690 145.140 ;
        RECT 1261.850 144.940 1290.690 145.080 ;
        RECT 1261.850 144.880 1262.170 144.940 ;
        RECT 1290.370 144.880 1290.690 144.940 ;
        RECT 1290.370 96.460 1290.690 96.520 ;
        RECT 1290.175 96.320 1290.690 96.460 ;
        RECT 1290.370 96.260 1290.690 96.320 ;
        RECT 1290.370 48.520 1290.690 48.580 ;
        RECT 1290.175 48.380 1290.690 48.520 ;
        RECT 1290.370 48.320 1290.690 48.380 ;
        RECT 1290.370 14.180 1290.690 14.240 ;
        RECT 1290.370 14.040 1293.360 14.180 ;
        RECT 1290.370 13.980 1290.690 14.040 ;
        RECT 1293.220 13.900 1293.360 14.040 ;
        RECT 1293.130 13.640 1293.450 13.900 ;
      LAYER via ;
        RECT 1261.880 144.880 1262.140 145.140 ;
        RECT 1290.400 144.880 1290.660 145.140 ;
        RECT 1290.400 96.260 1290.660 96.520 ;
        RECT 1290.400 48.320 1290.660 48.580 ;
        RECT 1290.400 13.980 1290.660 14.240 ;
        RECT 1293.160 13.640 1293.420 13.900 ;
      LAYER met2 ;
        RECT 312.890 2752.115 313.170 2752.485 ;
        RECT 312.960 2728.685 313.100 2752.115 ;
        RECT 312.890 2728.315 313.170 2728.685 ;
        RECT 312.890 2558.315 313.170 2558.685 ;
        RECT 312.960 2517.885 313.100 2558.315 ;
        RECT 312.890 2517.515 313.170 2517.885 ;
        RECT 312.890 2480.795 313.170 2481.165 ;
        RECT 312.960 2456.685 313.100 2480.795 ;
        RECT 312.890 2456.315 313.170 2456.685 ;
        RECT 312.430 2225.115 312.710 2225.485 ;
        RECT 312.500 2201.685 312.640 2225.115 ;
        RECT 312.430 2201.315 312.710 2201.685 ;
        RECT 312.890 2150.315 313.170 2150.685 ;
        RECT 312.960 2113.285 313.100 2150.315 ;
        RECT 312.890 2112.915 313.170 2113.285 ;
        RECT 312.890 1038.515 313.170 1038.885 ;
        RECT 312.960 1000.805 313.100 1038.515 ;
        RECT 312.890 1000.435 313.170 1000.805 ;
        RECT 315.190 191.915 315.470 192.285 ;
        RECT 315.260 155.565 315.400 191.915 ;
        RECT 315.190 155.195 315.470 155.565 ;
        RECT 1261.870 155.195 1262.150 155.565 ;
        RECT 1261.940 145.170 1262.080 155.195 ;
        RECT 1261.880 144.850 1262.140 145.170 ;
        RECT 1290.400 144.850 1290.660 145.170 ;
        RECT 1290.460 96.550 1290.600 144.850 ;
        RECT 1290.400 96.230 1290.660 96.550 ;
        RECT 1290.400 48.290 1290.660 48.610 ;
        RECT 1290.460 14.270 1290.600 48.290 ;
        RECT 1290.400 13.950 1290.660 14.270 ;
        RECT 1293.160 13.610 1293.420 13.930 ;
        RECT 1293.220 2.400 1293.360 13.610 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
      LAYER via2 ;
        RECT 312.890 2752.160 313.170 2752.440 ;
        RECT 312.890 2728.360 313.170 2728.640 ;
        RECT 312.890 2558.360 313.170 2558.640 ;
        RECT 312.890 2517.560 313.170 2517.840 ;
        RECT 312.890 2480.840 313.170 2481.120 ;
        RECT 312.890 2456.360 313.170 2456.640 ;
        RECT 312.430 2225.160 312.710 2225.440 ;
        RECT 312.430 2201.360 312.710 2201.640 ;
        RECT 312.890 2150.360 313.170 2150.640 ;
        RECT 312.890 2112.960 313.170 2113.240 ;
        RECT 312.890 1038.560 313.170 1038.840 ;
        RECT 312.890 1000.480 313.170 1000.760 ;
        RECT 315.190 191.960 315.470 192.240 ;
        RECT 315.190 155.240 315.470 155.520 ;
        RECT 1261.870 155.240 1262.150 155.520 ;
      LAYER met3 ;
        RECT 313.070 2759.620 313.450 2759.940 ;
        RECT 313.110 2758.960 313.410 2759.620 ;
        RECT 310.000 2758.360 314.000 2758.960 ;
        RECT 312.865 2752.460 313.195 2752.465 ;
        RECT 312.865 2752.450 313.450 2752.460 ;
        RECT 312.865 2752.150 313.650 2752.450 ;
        RECT 312.865 2752.140 313.450 2752.150 ;
        RECT 312.865 2752.135 313.195 2752.140 ;
        RECT 312.865 2728.660 313.195 2728.665 ;
        RECT 312.865 2728.650 313.450 2728.660 ;
        RECT 312.640 2728.350 313.450 2728.650 ;
        RECT 312.865 2728.340 313.450 2728.350 ;
        RECT 312.865 2728.335 313.195 2728.340 ;
        RECT 312.865 2558.660 313.195 2558.665 ;
        RECT 312.865 2558.650 313.450 2558.660 ;
        RECT 312.640 2558.350 313.450 2558.650 ;
        RECT 312.865 2558.340 313.450 2558.350 ;
        RECT 312.865 2558.335 313.195 2558.340 ;
        RECT 312.865 2517.860 313.195 2517.865 ;
        RECT 312.865 2517.850 313.450 2517.860 ;
        RECT 312.865 2517.550 313.650 2517.850 ;
        RECT 312.865 2517.540 313.450 2517.550 ;
        RECT 312.865 2517.535 313.195 2517.540 ;
        RECT 313.070 2511.420 313.450 2511.740 ;
        RECT 313.110 2511.060 313.410 2511.420 ;
        RECT 313.070 2510.740 313.450 2511.060 ;
        RECT 312.865 2481.140 313.195 2481.145 ;
        RECT 312.865 2481.130 313.450 2481.140 ;
        RECT 312.865 2480.830 313.650 2481.130 ;
        RECT 312.865 2480.820 313.450 2480.830 ;
        RECT 312.865 2480.815 313.195 2480.820 ;
        RECT 312.865 2456.660 313.195 2456.665 ;
        RECT 312.865 2456.650 313.450 2456.660 ;
        RECT 312.640 2456.350 313.450 2456.650 ;
        RECT 312.865 2456.340 313.450 2456.350 ;
        RECT 312.865 2456.335 313.195 2456.340 ;
        RECT 312.405 2225.450 312.735 2225.465 ;
        RECT 313.070 2225.450 313.450 2225.460 ;
        RECT 312.405 2225.150 313.450 2225.450 ;
        RECT 312.405 2225.135 312.735 2225.150 ;
        RECT 313.070 2225.140 313.450 2225.150 ;
        RECT 312.405 2201.650 312.735 2201.665 ;
        RECT 313.070 2201.650 313.450 2201.660 ;
        RECT 312.405 2201.350 313.450 2201.650 ;
        RECT 312.405 2201.335 312.735 2201.350 ;
        RECT 313.070 2201.340 313.450 2201.350 ;
        RECT 312.865 2150.660 313.195 2150.665 ;
        RECT 312.865 2150.650 313.450 2150.660 ;
        RECT 312.640 2150.350 313.450 2150.650 ;
        RECT 312.865 2150.340 313.450 2150.350 ;
        RECT 312.865 2150.335 313.195 2150.340 ;
        RECT 312.865 2113.260 313.195 2113.265 ;
        RECT 312.865 2113.250 313.450 2113.260 ;
        RECT 312.640 2112.950 313.450 2113.250 ;
        RECT 312.865 2112.940 313.450 2112.950 ;
        RECT 312.865 2112.935 313.195 2112.940 ;
        RECT 312.150 1840.570 312.530 1840.580 ;
        RECT 313.070 1840.570 313.450 1840.580 ;
        RECT 312.150 1840.270 313.450 1840.570 ;
        RECT 312.150 1840.260 312.530 1840.270 ;
        RECT 313.070 1840.260 313.450 1840.270 ;
        RECT 312.865 1038.860 313.195 1038.865 ;
        RECT 312.865 1038.850 313.450 1038.860 ;
        RECT 312.640 1038.550 313.450 1038.850 ;
        RECT 312.865 1038.540 313.450 1038.550 ;
        RECT 312.865 1038.535 313.195 1038.540 ;
        RECT 312.150 1000.770 312.530 1000.780 ;
        RECT 312.865 1000.770 313.195 1000.785 ;
        RECT 312.150 1000.470 313.195 1000.770 ;
        RECT 312.150 1000.460 312.530 1000.470 ;
        RECT 312.865 1000.455 313.195 1000.470 ;
        RECT 314.910 233.420 315.290 233.740 ;
        RECT 314.950 232.380 315.250 233.420 ;
        RECT 314.910 232.060 315.290 232.380 ;
        RECT 314.910 192.620 315.290 192.940 ;
        RECT 314.950 192.265 315.250 192.620 ;
        RECT 314.950 191.950 315.495 192.265 ;
        RECT 315.165 191.935 315.495 191.950 ;
        RECT 315.165 155.530 315.495 155.545 ;
        RECT 1261.845 155.530 1262.175 155.545 ;
        RECT 315.165 155.230 1262.175 155.530 ;
        RECT 315.165 155.215 315.495 155.230 ;
        RECT 1261.845 155.215 1262.175 155.230 ;
      LAYER via3 ;
        RECT 313.100 2759.620 313.420 2759.940 ;
        RECT 313.100 2752.140 313.420 2752.460 ;
        RECT 313.100 2728.340 313.420 2728.660 ;
        RECT 313.100 2558.340 313.420 2558.660 ;
        RECT 313.100 2517.540 313.420 2517.860 ;
        RECT 313.100 2511.420 313.420 2511.740 ;
        RECT 313.100 2510.740 313.420 2511.060 ;
        RECT 313.100 2480.820 313.420 2481.140 ;
        RECT 313.100 2456.340 313.420 2456.660 ;
        RECT 313.100 2225.140 313.420 2225.460 ;
        RECT 313.100 2201.340 313.420 2201.660 ;
        RECT 313.100 2150.340 313.420 2150.660 ;
        RECT 313.100 2112.940 313.420 2113.260 ;
        RECT 312.180 1840.260 312.500 1840.580 ;
        RECT 313.100 1840.260 313.420 1840.580 ;
        RECT 313.100 1038.540 313.420 1038.860 ;
        RECT 312.180 1000.460 312.500 1000.780 ;
        RECT 314.940 233.420 315.260 233.740 ;
        RECT 314.940 232.060 315.260 232.380 ;
        RECT 314.940 192.620 315.260 192.940 ;
      LAYER met4 ;
        RECT 313.095 2759.615 313.425 2759.945 ;
        RECT 313.110 2752.465 313.410 2759.615 ;
        RECT 313.095 2752.135 313.425 2752.465 ;
        RECT 313.095 2728.650 313.425 2728.665 ;
        RECT 313.095 2728.350 314.330 2728.650 ;
        RECT 313.095 2728.335 313.425 2728.350 ;
        RECT 314.030 2725.250 314.330 2728.350 ;
        RECT 314.030 2724.950 315.250 2725.250 ;
        RECT 314.950 2691.250 315.250 2724.950 ;
        RECT 314.950 2690.950 317.090 2691.250 ;
        RECT 316.790 2667.450 317.090 2690.950 ;
        RECT 314.950 2667.150 317.090 2667.450 ;
        RECT 314.950 2649.770 315.250 2667.150 ;
        RECT 314.030 2649.470 315.250 2649.770 ;
        RECT 314.030 2643.650 314.330 2649.470 ;
        RECT 314.030 2643.350 315.250 2643.650 ;
        RECT 314.950 2585.850 315.250 2643.350 ;
        RECT 313.110 2585.550 315.250 2585.850 ;
        RECT 313.110 2568.850 313.410 2585.550 ;
        RECT 313.110 2568.550 315.250 2568.850 ;
        RECT 313.095 2558.650 313.425 2558.665 ;
        RECT 314.950 2558.650 315.250 2568.550 ;
        RECT 313.095 2558.350 315.250 2558.650 ;
        RECT 313.095 2558.335 313.425 2558.350 ;
        RECT 313.095 2517.535 313.425 2517.865 ;
        RECT 313.110 2511.745 313.410 2517.535 ;
        RECT 313.095 2511.415 313.425 2511.745 ;
        RECT 313.095 2510.735 313.425 2511.065 ;
        RECT 313.110 2481.145 313.410 2510.735 ;
        RECT 313.095 2480.815 313.425 2481.145 ;
        RECT 313.095 2456.650 313.425 2456.665 ;
        RECT 313.095 2456.350 316.170 2456.650 ;
        RECT 313.095 2456.335 313.425 2456.350 ;
        RECT 315.870 2429.450 316.170 2456.350 ;
        RECT 314.030 2429.150 316.170 2429.450 ;
        RECT 314.030 2422.650 314.330 2429.150 ;
        RECT 314.030 2422.350 315.250 2422.650 ;
        RECT 313.095 2225.450 313.425 2225.465 ;
        RECT 314.950 2225.450 315.250 2422.350 ;
        RECT 313.095 2225.150 315.250 2225.450 ;
        RECT 313.095 2225.135 313.425 2225.150 ;
        RECT 313.095 2201.650 313.425 2201.665 ;
        RECT 313.095 2201.350 315.250 2201.650 ;
        RECT 313.095 2201.335 313.425 2201.350 ;
        RECT 313.095 2150.650 313.425 2150.665 ;
        RECT 314.950 2150.650 315.250 2201.350 ;
        RECT 313.095 2150.350 315.250 2150.650 ;
        RECT 313.095 2150.335 313.425 2150.350 ;
        RECT 313.095 2113.250 313.425 2113.265 ;
        RECT 313.095 2112.950 315.250 2113.250 ;
        RECT 313.095 2112.935 313.425 2112.950 ;
        RECT 314.950 1929.650 315.250 2112.950 ;
        RECT 312.190 1929.350 315.250 1929.650 ;
        RECT 312.190 1885.450 312.490 1929.350 ;
        RECT 312.190 1885.150 315.250 1885.450 ;
        RECT 314.950 1848.050 315.250 1885.150 ;
        RECT 312.190 1847.750 315.250 1848.050 ;
        RECT 312.190 1840.585 312.490 1847.750 ;
        RECT 312.175 1840.255 312.505 1840.585 ;
        RECT 313.095 1840.255 313.425 1840.585 ;
        RECT 313.110 1837.850 313.410 1840.255 ;
        RECT 313.110 1837.550 315.250 1837.850 ;
        RECT 314.950 1416.250 315.250 1837.550 ;
        RECT 314.030 1415.950 315.250 1416.250 ;
        RECT 314.030 1409.450 314.330 1415.950 ;
        RECT 314.030 1409.150 315.250 1409.450 ;
        RECT 313.095 1038.850 313.425 1038.865 ;
        RECT 314.950 1038.850 315.250 1409.150 ;
        RECT 313.095 1038.550 315.250 1038.850 ;
        RECT 313.095 1038.535 313.425 1038.550 ;
        RECT 312.175 1000.455 312.505 1000.785 ;
        RECT 312.190 977.650 312.490 1000.455 ;
        RECT 312.190 977.350 315.250 977.650 ;
        RECT 314.950 923.250 315.250 977.350 ;
        RECT 313.110 922.950 315.250 923.250 ;
        RECT 313.110 917.810 313.410 922.950 ;
        RECT 313.110 917.510 315.250 917.810 ;
        RECT 314.950 848.450 315.250 917.510 ;
        RECT 314.030 848.150 315.250 848.450 ;
        RECT 314.030 794.050 314.330 848.150 ;
        RECT 314.030 793.750 316.170 794.050 ;
        RECT 315.870 780.450 316.170 793.750 ;
        RECT 314.950 780.150 316.170 780.450 ;
        RECT 314.950 702.250 315.250 780.150 ;
        RECT 314.030 701.950 315.250 702.250 ;
        RECT 314.030 695.450 314.330 701.950 ;
        RECT 314.030 695.150 315.250 695.450 ;
        RECT 314.950 562.850 315.250 695.150 ;
        RECT 314.030 562.550 315.250 562.850 ;
        RECT 314.030 556.050 314.330 562.550 ;
        RECT 314.030 555.750 315.250 556.050 ;
        RECT 314.950 508.450 315.250 555.750 ;
        RECT 314.950 508.150 317.090 508.450 ;
        RECT 316.790 484.650 317.090 508.150 ;
        RECT 314.950 484.350 317.090 484.650 ;
        RECT 314.950 369.050 315.250 484.350 ;
        RECT 312.190 368.750 315.250 369.050 ;
        RECT 312.190 348.650 312.490 368.750 ;
        RECT 312.190 348.350 315.250 348.650 ;
        RECT 314.950 233.745 315.250 348.350 ;
        RECT 314.935 233.415 315.265 233.745 ;
        RECT 314.935 232.055 315.265 232.385 ;
        RECT 314.950 192.945 315.250 232.055 ;
        RECT 314.935 192.615 315.265 192.945 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.070 20.640 1311.390 20.700 ;
        RECT 1317.510 20.640 1317.830 20.700 ;
        RECT 1311.070 20.500 1317.830 20.640 ;
        RECT 1311.070 20.440 1311.390 20.500 ;
        RECT 1317.510 20.440 1317.830 20.500 ;
      LAYER via ;
        RECT 1311.100 20.440 1311.360 20.700 ;
        RECT 1317.540 20.440 1317.800 20.700 ;
      LAYER met2 ;
        RECT 1317.530 204.835 1317.810 205.205 ;
        RECT 1317.600 20.730 1317.740 204.835 ;
        RECT 1311.100 20.410 1311.360 20.730 ;
        RECT 1317.540 20.410 1317.800 20.730 ;
        RECT 1311.160 2.400 1311.300 20.410 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
      LAYER via2 ;
        RECT 1317.530 204.880 1317.810 205.160 ;
      LAYER met3 ;
        RECT 2606.000 2833.370 2610.000 2833.760 ;
        RECT 2624.110 2833.370 2624.490 2833.380 ;
        RECT 2606.000 2833.160 2624.490 2833.370 ;
        RECT 2609.580 2833.070 2624.490 2833.160 ;
        RECT 2624.110 2833.060 2624.490 2833.070 ;
        RECT 1317.505 205.170 1317.835 205.185 ;
        RECT 2624.110 205.170 2624.490 205.180 ;
        RECT 1317.505 204.870 2624.490 205.170 ;
        RECT 1317.505 204.855 1317.835 204.870 ;
        RECT 2624.110 204.860 2624.490 204.870 ;
      LAYER via3 ;
        RECT 2624.140 2833.060 2624.460 2833.380 ;
        RECT 2624.140 204.860 2624.460 205.180 ;
      LAYER met4 ;
        RECT 2624.135 2833.055 2624.465 2833.385 ;
        RECT 2624.150 205.185 2624.450 2833.055 ;
        RECT 2624.135 204.855 2624.465 205.185 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2511.820 2615.490 2511.880 ;
        RECT 2679.110 2511.820 2679.430 2511.880 ;
        RECT 2615.170 2511.680 2679.430 2511.820 ;
        RECT 2615.170 2511.620 2615.490 2511.680 ;
        RECT 2679.110 2511.620 2679.430 2511.680 ;
        RECT 1331.310 238.240 1331.630 238.300 ;
        RECT 2679.110 238.240 2679.430 238.300 ;
        RECT 1331.310 238.100 2679.430 238.240 ;
        RECT 1331.310 238.040 1331.630 238.100 ;
        RECT 2679.110 238.040 2679.430 238.100 ;
        RECT 1329.010 20.640 1329.330 20.700 ;
        RECT 1331.310 20.640 1331.630 20.700 ;
        RECT 1329.010 20.500 1331.630 20.640 ;
        RECT 1329.010 20.440 1329.330 20.500 ;
        RECT 1331.310 20.440 1331.630 20.500 ;
      LAYER via ;
        RECT 2615.200 2511.620 2615.460 2511.880 ;
        RECT 2679.140 2511.620 2679.400 2511.880 ;
        RECT 1331.340 238.040 1331.600 238.300 ;
        RECT 2679.140 238.040 2679.400 238.300 ;
        RECT 1329.040 20.440 1329.300 20.700 ;
        RECT 1331.340 20.440 1331.600 20.700 ;
      LAYER met2 ;
        RECT 2615.190 2514.795 2615.470 2515.165 ;
        RECT 2615.260 2511.910 2615.400 2514.795 ;
        RECT 2615.200 2511.590 2615.460 2511.910 ;
        RECT 2679.140 2511.590 2679.400 2511.910 ;
        RECT 2679.200 238.330 2679.340 2511.590 ;
        RECT 1331.340 238.010 1331.600 238.330 ;
        RECT 2679.140 238.010 2679.400 238.330 ;
        RECT 1331.400 20.730 1331.540 238.010 ;
        RECT 1329.040 20.410 1329.300 20.730 ;
        RECT 1331.340 20.410 1331.600 20.730 ;
        RECT 1329.100 2.400 1329.240 20.410 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2514.840 2615.470 2515.120 ;
      LAYER met3 ;
        RECT 2606.000 2515.130 2610.000 2515.520 ;
        RECT 2615.165 2515.130 2615.495 2515.145 ;
        RECT 2606.000 2514.920 2615.495 2515.130 ;
        RECT 2609.580 2514.830 2615.495 2514.920 ;
        RECT 2615.165 2514.815 2615.495 2514.830 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 512.510 244.020 512.830 244.080 ;
        RECT 517.110 244.020 517.430 244.080 ;
        RECT 512.510 243.880 517.430 244.020 ;
        RECT 512.510 243.820 512.830 243.880 ;
        RECT 517.110 243.820 517.430 243.880 ;
        RECT 517.110 25.400 517.430 25.460 ;
        RECT 686.390 25.400 686.710 25.460 ;
        RECT 517.110 25.260 686.710 25.400 ;
        RECT 517.110 25.200 517.430 25.260 ;
        RECT 686.390 25.200 686.710 25.260 ;
      LAYER via ;
        RECT 512.540 243.820 512.800 244.080 ;
        RECT 517.140 243.820 517.400 244.080 ;
        RECT 517.140 25.200 517.400 25.460 ;
        RECT 686.420 25.200 686.680 25.460 ;
      LAYER met2 ;
        RECT 512.490 260.000 512.770 264.000 ;
        RECT 512.600 244.110 512.740 260.000 ;
        RECT 512.540 243.790 512.800 244.110 ;
        RECT 517.140 243.790 517.400 244.110 ;
        RECT 517.200 25.490 517.340 243.790 ;
        RECT 517.140 25.170 517.400 25.490 ;
        RECT 686.420 25.170 686.680 25.490 ;
        RECT 686.480 2.400 686.620 25.170 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 304.130 129.100 304.450 129.160 ;
        RECT 1345.570 129.100 1345.890 129.160 ;
        RECT 304.130 128.960 1345.890 129.100 ;
        RECT 304.130 128.900 304.450 128.960 ;
        RECT 1345.570 128.900 1345.890 128.960 ;
        RECT 1345.570 14.180 1345.890 14.240 ;
        RECT 1345.570 14.040 1346.720 14.180 ;
        RECT 1345.570 13.980 1345.890 14.040 ;
        RECT 1346.580 13.900 1346.720 14.040 ;
        RECT 1346.490 13.640 1346.810 13.900 ;
      LAYER via ;
        RECT 304.160 128.900 304.420 129.160 ;
        RECT 1345.600 128.900 1345.860 129.160 ;
        RECT 1345.600 13.980 1345.860 14.240 ;
        RECT 1346.520 13.640 1346.780 13.900 ;
      LAYER met2 ;
        RECT 304.150 2461.755 304.430 2462.125 ;
        RECT 304.220 129.190 304.360 2461.755 ;
        RECT 304.160 128.870 304.420 129.190 ;
        RECT 1345.600 128.870 1345.860 129.190 ;
        RECT 1345.660 14.270 1345.800 128.870 ;
        RECT 1345.600 13.950 1345.860 14.270 ;
        RECT 1346.520 13.610 1346.780 13.930 ;
        RECT 1346.580 2.400 1346.720 13.610 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
      LAYER via2 ;
        RECT 304.150 2461.800 304.430 2462.080 ;
      LAYER met3 ;
        RECT 304.125 2462.090 304.455 2462.105 ;
        RECT 310.000 2462.090 314.000 2462.480 ;
        RECT 304.125 2461.880 314.000 2462.090 ;
        RECT 304.125 2461.790 310.500 2461.880 ;
        RECT 304.125 2461.775 304.455 2461.790 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1364.505 48.365 1364.675 137.955 ;
      LAYER mcon ;
        RECT 1364.505 137.785 1364.675 137.955 ;
      LAYER met1 ;
        RECT 1620.190 3284.640 1620.510 3284.700 ;
        RECT 2611.950 3284.640 2612.270 3284.700 ;
        RECT 1620.190 3284.500 2612.270 3284.640 ;
        RECT 1620.190 3284.440 1620.510 3284.500 ;
        RECT 2611.950 3284.440 2612.270 3284.500 ;
        RECT 2611.950 666.980 2612.270 667.040 ;
        RECT 2615.170 666.980 2615.490 667.040 ;
        RECT 2611.950 666.840 2615.490 666.980 ;
        RECT 2611.950 666.780 2612.270 666.840 ;
        RECT 2615.170 666.780 2615.490 666.840 ;
        RECT 2614.250 635.020 2614.570 635.080 ;
        RECT 2615.170 635.020 2615.490 635.080 ;
        RECT 2614.250 634.880 2615.490 635.020 ;
        RECT 2614.250 634.820 2614.570 634.880 ;
        RECT 2615.170 634.820 2615.490 634.880 ;
        RECT 1365.810 186.560 1366.130 186.620 ;
        RECT 1374.550 186.560 1374.870 186.620 ;
        RECT 1365.810 186.420 1374.870 186.560 ;
        RECT 1365.810 186.360 1366.130 186.420 ;
        RECT 1374.550 186.360 1374.870 186.420 ;
        RECT 1364.445 137.940 1364.735 137.985 ;
        RECT 1365.810 137.940 1366.130 138.000 ;
        RECT 1364.445 137.800 1366.130 137.940 ;
        RECT 1364.445 137.755 1364.735 137.800 ;
        RECT 1365.810 137.740 1366.130 137.800 ;
        RECT 1364.430 48.520 1364.750 48.580 ;
        RECT 1364.235 48.380 1364.750 48.520 ;
        RECT 1364.430 48.320 1364.750 48.380 ;
      LAYER via ;
        RECT 1620.220 3284.440 1620.480 3284.700 ;
        RECT 2611.980 3284.440 2612.240 3284.700 ;
        RECT 2611.980 666.780 2612.240 667.040 ;
        RECT 2615.200 666.780 2615.460 667.040 ;
        RECT 2614.280 634.820 2614.540 635.080 ;
        RECT 2615.200 634.820 2615.460 635.080 ;
        RECT 1365.840 186.360 1366.100 186.620 ;
        RECT 1374.580 186.360 1374.840 186.620 ;
        RECT 1365.840 137.740 1366.100 138.000 ;
        RECT 1364.460 48.320 1364.720 48.580 ;
      LAYER met2 ;
        RECT 1620.220 3284.410 1620.480 3284.730 ;
        RECT 2611.980 3284.410 2612.240 3284.730 ;
        RECT 1620.280 3260.000 1620.420 3284.410 ;
        RECT 1620.170 3256.000 1620.450 3260.000 ;
        RECT 2612.040 667.070 2612.180 3284.410 ;
        RECT 2611.980 666.750 2612.240 667.070 ;
        RECT 2615.200 666.750 2615.460 667.070 ;
        RECT 2615.260 635.110 2615.400 666.750 ;
        RECT 2614.280 634.790 2614.540 635.110 ;
        RECT 2615.200 634.790 2615.460 635.110 ;
        RECT 2614.340 490.125 2614.480 634.790 ;
        RECT 2614.270 489.755 2614.550 490.125 ;
        RECT 2614.270 358.515 2614.550 358.885 ;
        RECT 2614.340 280.005 2614.480 358.515 ;
        RECT 2614.270 279.635 2614.550 280.005 ;
        RECT 2608.750 267.395 2609.030 267.765 ;
        RECT 2608.820 231.725 2608.960 267.395 ;
        RECT 1374.570 231.355 1374.850 231.725 ;
        RECT 2608.750 231.355 2609.030 231.725 ;
        RECT 1374.640 186.650 1374.780 231.355 ;
        RECT 1365.840 186.330 1366.100 186.650 ;
        RECT 1374.580 186.330 1374.840 186.650 ;
        RECT 1365.900 138.030 1366.040 186.330 ;
        RECT 1365.840 137.710 1366.100 138.030 ;
        RECT 1364.460 48.290 1364.720 48.610 ;
        RECT 1364.520 2.400 1364.660 48.290 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
      LAYER via2 ;
        RECT 2614.270 489.800 2614.550 490.080 ;
        RECT 2614.270 358.560 2614.550 358.840 ;
        RECT 2614.270 279.680 2614.550 279.960 ;
        RECT 2608.750 267.440 2609.030 267.720 ;
        RECT 1374.570 231.400 1374.850 231.680 ;
        RECT 2608.750 231.400 2609.030 231.680 ;
      LAYER met3 ;
        RECT 2614.245 490.090 2614.575 490.105 ;
        RECT 2619.510 490.090 2619.890 490.100 ;
        RECT 2614.245 489.790 2619.890 490.090 ;
        RECT 2614.245 489.775 2614.575 489.790 ;
        RECT 2619.510 489.780 2619.890 489.790 ;
        RECT 2614.245 358.850 2614.575 358.865 ;
        RECT 2619.510 358.850 2619.890 358.860 ;
        RECT 2614.245 358.550 2619.890 358.850 ;
        RECT 2614.245 358.535 2614.575 358.550 ;
        RECT 2619.510 358.540 2619.890 358.550 ;
        RECT 2606.630 279.970 2607.010 279.980 ;
        RECT 2614.245 279.970 2614.575 279.985 ;
        RECT 2606.630 279.670 2614.575 279.970 ;
        RECT 2606.630 279.660 2607.010 279.670 ;
        RECT 2614.245 279.655 2614.575 279.670 ;
        RECT 2606.630 267.730 2607.010 267.740 ;
        RECT 2608.725 267.730 2609.055 267.745 ;
        RECT 2606.630 267.430 2609.055 267.730 ;
        RECT 2606.630 267.420 2607.010 267.430 ;
        RECT 2608.725 267.415 2609.055 267.430 ;
        RECT 1374.545 231.690 1374.875 231.705 ;
        RECT 2608.725 231.690 2609.055 231.705 ;
        RECT 1374.545 231.390 2609.055 231.690 ;
        RECT 1374.545 231.375 1374.875 231.390 ;
        RECT 2608.725 231.375 2609.055 231.390 ;
      LAYER via3 ;
        RECT 2619.540 489.780 2619.860 490.100 ;
        RECT 2619.540 358.540 2619.860 358.860 ;
        RECT 2606.660 279.660 2606.980 279.980 ;
        RECT 2606.660 267.420 2606.980 267.740 ;
      LAYER met4 ;
        RECT 2619.535 489.775 2619.865 490.105 ;
        RECT 2619.550 358.865 2619.850 489.775 ;
        RECT 2619.535 358.535 2619.865 358.865 ;
        RECT 2606.655 279.655 2606.985 279.985 ;
        RECT 2606.670 267.745 2606.970 279.655 ;
        RECT 2606.655 267.415 2606.985 267.745 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 277.910 386.480 278.230 386.540 ;
        RECT 296.770 386.480 297.090 386.540 ;
        RECT 277.910 386.340 297.090 386.480 ;
        RECT 277.910 386.280 278.230 386.340 ;
        RECT 296.770 386.280 297.090 386.340 ;
        RECT 277.910 33.560 278.230 33.620 ;
        RECT 1382.370 33.560 1382.690 33.620 ;
        RECT 277.910 33.420 1382.690 33.560 ;
        RECT 277.910 33.360 278.230 33.420 ;
        RECT 1382.370 33.360 1382.690 33.420 ;
      LAYER via ;
        RECT 277.940 386.280 278.200 386.540 ;
        RECT 296.800 386.280 297.060 386.540 ;
        RECT 277.940 33.360 278.200 33.620 ;
        RECT 1382.400 33.360 1382.660 33.620 ;
      LAYER met2 ;
        RECT 296.790 390.475 297.070 390.845 ;
        RECT 296.860 386.570 297.000 390.475 ;
        RECT 277.940 386.250 278.200 386.570 ;
        RECT 296.800 386.250 297.060 386.570 ;
        RECT 278.000 33.650 278.140 386.250 ;
        RECT 277.940 33.330 278.200 33.650 ;
        RECT 1382.400 33.330 1382.660 33.650 ;
        RECT 1382.460 2.400 1382.600 33.330 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
      LAYER via2 ;
        RECT 296.790 390.520 297.070 390.800 ;
      LAYER met3 ;
        RECT 296.765 390.810 297.095 390.825 ;
        RECT 310.000 390.810 314.000 391.200 ;
        RECT 296.765 390.600 314.000 390.810 ;
        RECT 296.765 390.510 310.500 390.600 ;
        RECT 296.765 390.495 297.095 390.510 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 245.710 2712.080 246.030 2712.140 ;
        RECT 296.770 2712.080 297.090 2712.140 ;
        RECT 245.710 2711.940 297.090 2712.080 ;
        RECT 245.710 2711.880 246.030 2711.940 ;
        RECT 296.770 2711.880 297.090 2711.940 ;
        RECT 245.710 47.840 246.030 47.900 ;
        RECT 1399.850 47.840 1400.170 47.900 ;
        RECT 245.710 47.700 1400.170 47.840 ;
        RECT 245.710 47.640 246.030 47.700 ;
        RECT 1399.850 47.640 1400.170 47.700 ;
      LAYER via ;
        RECT 245.740 2711.880 246.000 2712.140 ;
        RECT 296.800 2711.880 297.060 2712.140 ;
        RECT 245.740 47.640 246.000 47.900 ;
        RECT 1399.880 47.640 1400.140 47.900 ;
      LAYER met2 ;
        RECT 296.790 2714.715 297.070 2715.085 ;
        RECT 296.860 2712.170 297.000 2714.715 ;
        RECT 245.740 2711.850 246.000 2712.170 ;
        RECT 296.800 2711.850 297.060 2712.170 ;
        RECT 245.800 47.930 245.940 2711.850 ;
        RECT 245.740 47.610 246.000 47.930 ;
        RECT 1399.880 47.610 1400.140 47.930 ;
        RECT 1399.940 16.050 1400.080 47.610 ;
        RECT 1399.940 15.910 1400.540 16.050 ;
        RECT 1400.400 2.400 1400.540 15.910 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
      LAYER via2 ;
        RECT 296.790 2714.760 297.070 2715.040 ;
      LAYER met3 ;
        RECT 296.765 2715.050 297.095 2715.065 ;
        RECT 310.000 2715.050 314.000 2715.440 ;
        RECT 296.765 2714.840 314.000 2715.050 ;
        RECT 296.765 2714.750 310.500 2714.840 ;
        RECT 296.765 2714.735 297.095 2714.750 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 198.120 1421.330 198.180 ;
        RECT 2625.290 198.120 2625.610 198.180 ;
        RECT 1421.010 197.980 2625.610 198.120 ;
        RECT 1421.010 197.920 1421.330 197.980 ;
        RECT 2625.290 197.920 2625.610 197.980 ;
        RECT 1418.250 20.640 1418.570 20.700 ;
        RECT 1421.010 20.640 1421.330 20.700 ;
        RECT 1418.250 20.500 1421.330 20.640 ;
        RECT 1418.250 20.440 1418.570 20.500 ;
        RECT 1421.010 20.440 1421.330 20.500 ;
      LAYER via ;
        RECT 1421.040 197.920 1421.300 198.180 ;
        RECT 2625.320 197.920 2625.580 198.180 ;
        RECT 1418.280 20.440 1418.540 20.700 ;
        RECT 1421.040 20.440 1421.300 20.700 ;
      LAYER met2 ;
        RECT 2625.310 1078.635 2625.590 1079.005 ;
        RECT 2625.380 198.210 2625.520 1078.635 ;
        RECT 1421.040 197.890 1421.300 198.210 ;
        RECT 2625.320 197.890 2625.580 198.210 ;
        RECT 1421.100 20.730 1421.240 197.890 ;
        RECT 1418.280 20.410 1418.540 20.730 ;
        RECT 1421.040 20.410 1421.300 20.730 ;
        RECT 1418.340 2.400 1418.480 20.410 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
      LAYER via2 ;
        RECT 2625.310 1078.680 2625.590 1078.960 ;
      LAYER met3 ;
        RECT 2606.000 1078.970 2610.000 1079.360 ;
        RECT 2625.285 1078.970 2625.615 1078.985 ;
        RECT 2606.000 1078.760 2625.615 1078.970 ;
        RECT 2609.580 1078.670 2625.615 1078.760 ;
        RECT 2625.285 1078.655 2625.615 1078.670 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1648.710 3284.980 1649.030 3285.040 ;
        RECT 2632.190 3284.980 2632.510 3285.040 ;
        RECT 1648.710 3284.840 2632.510 3284.980 ;
        RECT 1648.710 3284.780 1649.030 3284.840 ;
        RECT 2632.190 3284.780 2632.510 3284.840 ;
        RECT 2632.190 338.200 2632.510 338.260 ;
        RECT 2643.230 338.200 2643.550 338.260 ;
        RECT 2632.190 338.060 2643.550 338.200 ;
        RECT 2632.190 338.000 2632.510 338.060 ;
        RECT 2643.230 338.000 2643.550 338.060 ;
        RECT 2632.190 275.980 2632.510 276.040 ;
        RECT 2643.230 275.980 2643.550 276.040 ;
        RECT 2632.190 275.840 2643.550 275.980 ;
        RECT 2632.190 275.780 2632.510 275.840 ;
        RECT 2643.230 275.780 2643.550 275.840 ;
        RECT 1441.710 218.180 1442.030 218.240 ;
        RECT 2632.190 218.180 2632.510 218.240 ;
        RECT 1441.710 218.040 2632.510 218.180 ;
        RECT 1441.710 217.980 1442.030 218.040 ;
        RECT 2632.190 217.980 2632.510 218.040 ;
        RECT 1435.730 16.560 1436.050 16.620 ;
        RECT 1441.710 16.560 1442.030 16.620 ;
        RECT 1435.730 16.420 1442.030 16.560 ;
        RECT 1435.730 16.360 1436.050 16.420 ;
        RECT 1441.710 16.360 1442.030 16.420 ;
      LAYER via ;
        RECT 1648.740 3284.780 1649.000 3285.040 ;
        RECT 2632.220 3284.780 2632.480 3285.040 ;
        RECT 2632.220 338.000 2632.480 338.260 ;
        RECT 2643.260 338.000 2643.520 338.260 ;
        RECT 2632.220 275.780 2632.480 276.040 ;
        RECT 2643.260 275.780 2643.520 276.040 ;
        RECT 1441.740 217.980 1442.000 218.240 ;
        RECT 2632.220 217.980 2632.480 218.240 ;
        RECT 1435.760 16.360 1436.020 16.620 ;
        RECT 1441.740 16.360 1442.000 16.620 ;
      LAYER met2 ;
        RECT 1648.740 3284.750 1649.000 3285.070 ;
        RECT 2632.220 3284.750 2632.480 3285.070 ;
        RECT 1648.800 3260.000 1648.940 3284.750 ;
        RECT 1648.690 3256.000 1648.970 3260.000 ;
        RECT 2632.280 338.290 2632.420 3284.750 ;
        RECT 2632.220 337.970 2632.480 338.290 ;
        RECT 2643.260 337.970 2643.520 338.290 ;
        RECT 2643.320 276.070 2643.460 337.970 ;
        RECT 2632.220 275.750 2632.480 276.070 ;
        RECT 2643.260 275.750 2643.520 276.070 ;
        RECT 2632.280 218.270 2632.420 275.750 ;
        RECT 1441.740 217.950 1442.000 218.270 ;
        RECT 2632.220 217.950 2632.480 218.270 ;
        RECT 1441.800 16.650 1441.940 217.950 ;
        RECT 1435.760 16.330 1436.020 16.650 ;
        RECT 1441.740 16.330 1442.000 16.650 ;
        RECT 1435.820 2.400 1435.960 16.330 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.690 45.715 1453.970 46.085 ;
        RECT 1453.760 2.400 1453.900 45.715 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
      LAYER via2 ;
        RECT 1453.690 45.760 1453.970 46.040 ;
      LAYER met3 ;
        RECT 310.000 2927.000 314.000 2927.600 ;
        RECT 252.350 2925.850 252.730 2925.860 ;
        RECT 310.350 2925.850 310.650 2927.000 ;
        RECT 252.350 2925.550 310.650 2925.850 ;
        RECT 252.350 2925.540 252.730 2925.550 ;
        RECT 252.350 46.050 252.730 46.060 ;
        RECT 1453.665 46.050 1453.995 46.065 ;
        RECT 252.350 45.750 1453.995 46.050 ;
        RECT 252.350 45.740 252.730 45.750 ;
        RECT 1453.665 45.735 1453.995 45.750 ;
      LAYER via3 ;
        RECT 252.380 2925.540 252.700 2925.860 ;
        RECT 252.380 45.740 252.700 46.060 ;
      LAYER met4 ;
        RECT 252.375 2925.535 252.705 2925.865 ;
        RECT 252.390 46.065 252.690 2925.535 ;
        RECT 252.375 45.735 252.705 46.065 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1098.550 244.020 1098.870 244.080 ;
        RECT 1103.610 244.020 1103.930 244.080 ;
        RECT 1098.550 243.880 1103.930 244.020 ;
        RECT 1098.550 243.820 1098.870 243.880 ;
        RECT 1103.610 243.820 1103.930 243.880 ;
        RECT 1103.610 26.080 1103.930 26.140 ;
        RECT 1471.610 26.080 1471.930 26.140 ;
        RECT 1103.610 25.940 1471.930 26.080 ;
        RECT 1103.610 25.880 1103.930 25.940 ;
        RECT 1471.610 25.880 1471.930 25.940 ;
      LAYER via ;
        RECT 1098.580 243.820 1098.840 244.080 ;
        RECT 1103.640 243.820 1103.900 244.080 ;
        RECT 1103.640 25.880 1103.900 26.140 ;
        RECT 1471.640 25.880 1471.900 26.140 ;
      LAYER met2 ;
        RECT 1098.530 260.000 1098.810 264.000 ;
        RECT 1098.640 244.110 1098.780 260.000 ;
        RECT 1098.580 243.790 1098.840 244.110 ;
        RECT 1103.640 243.790 1103.900 244.110 ;
        RECT 1103.700 26.170 1103.840 243.790 ;
        RECT 1103.640 25.850 1103.900 26.170 ;
        RECT 1471.640 25.850 1471.900 26.170 ;
        RECT 1471.700 2.400 1471.840 25.850 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 25.400 1490.330 25.460 ;
        RECT 2325.370 25.400 2325.690 25.460 ;
        RECT 1490.010 25.260 2325.690 25.400 ;
        RECT 1490.010 25.200 1490.330 25.260 ;
        RECT 2325.370 25.200 2325.690 25.260 ;
      LAYER via ;
        RECT 1490.040 25.200 1490.300 25.460 ;
        RECT 2325.400 25.200 2325.660 25.460 ;
      LAYER met2 ;
        RECT 2328.570 260.170 2328.850 264.000 ;
        RECT 2325.460 260.030 2328.850 260.170 ;
        RECT 2325.460 25.490 2325.600 260.030 ;
        RECT 2328.570 260.000 2328.850 260.030 ;
        RECT 1490.040 25.170 1490.300 25.490 ;
        RECT 2325.400 25.170 2325.660 25.490 ;
        RECT 1490.100 12.650 1490.240 25.170 ;
        RECT 1489.640 12.510 1490.240 12.650 ;
        RECT 1489.640 2.400 1489.780 12.510 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1849.270 3266.620 1849.590 3266.680 ;
        RECT 2632.650 3266.620 2632.970 3266.680 ;
        RECT 1849.270 3266.480 2632.970 3266.620 ;
        RECT 1849.270 3266.420 1849.590 3266.480 ;
        RECT 2632.650 3266.420 2632.970 3266.480 ;
        RECT 2632.650 383.420 2632.970 383.480 ;
        RECT 2642.770 383.420 2643.090 383.480 ;
        RECT 2632.650 383.280 2643.090 383.420 ;
        RECT 2632.650 383.220 2632.970 383.280 ;
        RECT 2642.770 383.220 2643.090 383.280 ;
        RECT 1507.030 20.640 1507.350 20.700 ;
        RECT 1510.710 20.640 1511.030 20.700 ;
        RECT 1507.030 20.500 1511.030 20.640 ;
        RECT 1507.030 20.440 1507.350 20.500 ;
        RECT 1510.710 20.440 1511.030 20.500 ;
      LAYER via ;
        RECT 1849.300 3266.420 1849.560 3266.680 ;
        RECT 2632.680 3266.420 2632.940 3266.680 ;
        RECT 2632.680 383.220 2632.940 383.480 ;
        RECT 2642.800 383.220 2643.060 383.480 ;
        RECT 1507.060 20.440 1507.320 20.700 ;
        RECT 1510.740 20.440 1511.000 20.700 ;
      LAYER met2 ;
        RECT 1849.300 3266.390 1849.560 3266.710 ;
        RECT 2632.680 3266.390 2632.940 3266.710 ;
        RECT 1849.360 3260.000 1849.500 3266.390 ;
        RECT 1849.250 3256.000 1849.530 3260.000 ;
        RECT 2632.740 383.510 2632.880 3266.390 ;
        RECT 2632.680 383.190 2632.940 383.510 ;
        RECT 2642.800 383.190 2643.060 383.510 ;
        RECT 2642.860 351.405 2643.000 383.190 ;
        RECT 2642.790 351.035 2643.070 351.405 ;
        RECT 1510.730 232.715 1511.010 233.085 ;
        RECT 1510.800 20.730 1510.940 232.715 ;
        RECT 1507.060 20.410 1507.320 20.730 ;
        RECT 1510.740 20.410 1511.000 20.730 ;
        RECT 1507.120 2.400 1507.260 20.410 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
      LAYER via2 ;
        RECT 2642.790 351.080 2643.070 351.360 ;
        RECT 1510.730 232.760 1511.010 233.040 ;
      LAYER met3 ;
        RECT 2619.510 351.370 2619.890 351.380 ;
        RECT 2642.765 351.370 2643.095 351.385 ;
        RECT 2619.510 351.070 2643.095 351.370 ;
        RECT 2619.510 351.060 2619.890 351.070 ;
        RECT 2642.765 351.055 2643.095 351.070 ;
        RECT 1510.705 233.050 1511.035 233.065 ;
        RECT 2619.510 233.050 2619.890 233.060 ;
        RECT 1510.705 232.750 2619.890 233.050 ;
        RECT 1510.705 232.735 1511.035 232.750 ;
        RECT 2619.510 232.740 2619.890 232.750 ;
      LAYER via3 ;
        RECT 2619.540 351.060 2619.860 351.380 ;
        RECT 2619.540 232.740 2619.860 233.060 ;
      LAYER met4 ;
        RECT 2619.535 351.055 2619.865 351.385 ;
        RECT 2619.550 233.065 2619.850 351.055 ;
        RECT 2619.535 232.735 2619.865 233.065 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 312.870 241.980 313.190 242.040 ;
        RECT 321.150 241.980 321.470 242.040 ;
        RECT 312.870 241.840 321.470 241.980 ;
        RECT 312.870 241.780 313.190 241.840 ;
        RECT 321.150 241.780 321.470 241.840 ;
        RECT 321.150 148.140 321.470 148.200 ;
        RECT 704.330 148.140 704.650 148.200 ;
        RECT 321.150 148.000 704.650 148.140 ;
        RECT 321.150 147.940 321.470 148.000 ;
        RECT 704.330 147.940 704.650 148.000 ;
      LAYER via ;
        RECT 312.900 241.780 313.160 242.040 ;
        RECT 321.180 241.780 321.440 242.040 ;
        RECT 321.180 147.940 321.440 148.200 ;
        RECT 704.360 147.940 704.620 148.200 ;
      LAYER met2 ;
        RECT 312.850 260.000 313.130 264.000 ;
        RECT 312.960 242.070 313.100 260.000 ;
        RECT 312.900 241.750 313.160 242.070 ;
        RECT 321.180 241.750 321.440 242.070 ;
        RECT 321.240 148.230 321.380 241.750 ;
        RECT 321.180 147.910 321.440 148.230 ;
        RECT 704.360 147.910 704.620 148.230 ;
        RECT 704.420 2.400 704.560 147.910 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2574.040 2615.490 2574.100 ;
        RECT 2678.650 2574.040 2678.970 2574.100 ;
        RECT 2615.170 2573.900 2678.970 2574.040 ;
        RECT 2615.170 2573.840 2615.490 2573.900 ;
        RECT 2678.650 2573.840 2678.970 2573.900 ;
        RECT 1531.410 238.580 1531.730 238.640 ;
        RECT 2678.650 238.580 2678.970 238.640 ;
        RECT 1531.410 238.440 2678.970 238.580 ;
        RECT 1531.410 238.380 1531.730 238.440 ;
        RECT 2678.650 238.380 2678.970 238.440 ;
        RECT 1524.970 16.220 1525.290 16.280 ;
        RECT 1531.410 16.220 1531.730 16.280 ;
        RECT 1524.970 16.080 1531.730 16.220 ;
        RECT 1524.970 16.020 1525.290 16.080 ;
        RECT 1531.410 16.020 1531.730 16.080 ;
      LAYER via ;
        RECT 2615.200 2573.840 2615.460 2574.100 ;
        RECT 2678.680 2573.840 2678.940 2574.100 ;
        RECT 1531.440 238.380 1531.700 238.640 ;
        RECT 2678.680 238.380 2678.940 238.640 ;
        RECT 1525.000 16.020 1525.260 16.280 ;
        RECT 1531.440 16.020 1531.700 16.280 ;
      LAYER met2 ;
        RECT 2615.190 2578.715 2615.470 2579.085 ;
        RECT 2615.260 2574.130 2615.400 2578.715 ;
        RECT 2615.200 2573.810 2615.460 2574.130 ;
        RECT 2678.680 2573.810 2678.940 2574.130 ;
        RECT 2678.740 238.670 2678.880 2573.810 ;
        RECT 1531.440 238.350 1531.700 238.670 ;
        RECT 2678.680 238.350 2678.940 238.670 ;
        RECT 1531.500 16.310 1531.640 238.350 ;
        RECT 1525.000 15.990 1525.260 16.310 ;
        RECT 1531.440 15.990 1531.700 16.310 ;
        RECT 1525.060 2.400 1525.200 15.990 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2578.760 2615.470 2579.040 ;
      LAYER met3 ;
        RECT 2606.000 2579.050 2610.000 2579.440 ;
        RECT 2615.165 2579.050 2615.495 2579.065 ;
        RECT 2606.000 2578.840 2615.495 2579.050 ;
        RECT 2609.580 2578.750 2615.495 2578.840 ;
        RECT 2615.165 2578.735 2615.495 2578.750 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1539.305 48.365 1539.475 96.475 ;
      LAYER mcon ;
        RECT 1539.305 96.305 1539.475 96.475 ;
      LAYER met1 ;
        RECT 312.410 121.620 312.730 121.680 ;
        RECT 1539.690 121.620 1540.010 121.680 ;
        RECT 312.410 121.480 1540.010 121.620 ;
        RECT 312.410 121.420 312.730 121.480 ;
        RECT 1539.690 121.420 1540.010 121.480 ;
        RECT 1539.230 96.460 1539.550 96.520 ;
        RECT 1539.035 96.320 1539.550 96.460 ;
        RECT 1539.230 96.260 1539.550 96.320 ;
        RECT 1539.230 48.520 1539.550 48.580 ;
        RECT 1539.035 48.380 1539.550 48.520 ;
        RECT 1539.230 48.320 1539.550 48.380 ;
        RECT 1539.230 14.180 1539.550 14.240 ;
        RECT 1539.230 14.040 1543.140 14.180 ;
        RECT 1539.230 13.980 1539.550 14.040 ;
        RECT 1543.000 13.900 1543.140 14.040 ;
        RECT 1542.910 13.640 1543.230 13.900 ;
      LAYER via ;
        RECT 312.440 121.420 312.700 121.680 ;
        RECT 1539.720 121.420 1539.980 121.680 ;
        RECT 1539.260 96.260 1539.520 96.520 ;
        RECT 1539.260 48.320 1539.520 48.580 ;
        RECT 1539.260 13.980 1539.520 14.240 ;
        RECT 1542.940 13.640 1543.200 13.900 ;
      LAYER met2 ;
        RECT 312.430 1190.155 312.710 1190.525 ;
        RECT 312.500 121.710 312.640 1190.155 ;
        RECT 312.440 121.390 312.700 121.710 ;
        RECT 1539.720 121.390 1539.980 121.710 ;
        RECT 1539.780 96.970 1539.920 121.390 ;
        RECT 1539.320 96.830 1539.920 96.970 ;
        RECT 1539.320 96.550 1539.460 96.830 ;
        RECT 1539.260 96.230 1539.520 96.550 ;
        RECT 1539.260 48.290 1539.520 48.610 ;
        RECT 1539.320 14.270 1539.460 48.290 ;
        RECT 1539.260 13.950 1539.520 14.270 ;
        RECT 1542.940 13.610 1543.200 13.930 ;
        RECT 1543.000 2.400 1543.140 13.610 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
      LAYER via2 ;
        RECT 312.430 1190.200 312.710 1190.480 ;
      LAYER met3 ;
        RECT 310.000 1193.000 314.000 1193.600 ;
        RECT 312.190 1190.505 312.490 1193.000 ;
        RECT 312.190 1190.190 312.735 1190.505 ;
        RECT 312.405 1190.175 312.735 1190.190 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 807.445 24.225 808.535 24.395 ;
      LAYER mcon ;
        RECT 808.365 24.225 808.535 24.395 ;
      LAYER met1 ;
        RECT 455.470 241.640 455.790 241.700 ;
        RECT 461.910 241.640 462.230 241.700 ;
        RECT 455.470 241.500 462.230 241.640 ;
        RECT 455.470 241.440 455.790 241.500 ;
        RECT 461.910 241.440 462.230 241.500 ;
        RECT 461.910 24.380 462.230 24.440 ;
        RECT 807.385 24.380 807.675 24.425 ;
        RECT 461.910 24.240 807.675 24.380 ;
        RECT 461.910 24.180 462.230 24.240 ;
        RECT 807.385 24.195 807.675 24.240 ;
        RECT 808.305 24.380 808.595 24.425 ;
        RECT 1560.850 24.380 1561.170 24.440 ;
        RECT 808.305 24.240 1561.170 24.380 ;
        RECT 808.305 24.195 808.595 24.240 ;
        RECT 1560.850 24.180 1561.170 24.240 ;
      LAYER via ;
        RECT 455.500 241.440 455.760 241.700 ;
        RECT 461.940 241.440 462.200 241.700 ;
        RECT 461.940 24.180 462.200 24.440 ;
        RECT 1560.880 24.180 1561.140 24.440 ;
      LAYER met2 ;
        RECT 455.450 260.000 455.730 264.000 ;
        RECT 455.560 241.730 455.700 260.000 ;
        RECT 455.500 241.410 455.760 241.730 ;
        RECT 461.940 241.410 462.200 241.730 ;
        RECT 462.000 24.470 462.140 241.410 ;
        RECT 461.940 24.150 462.200 24.470 ;
        RECT 1560.880 24.150 1561.140 24.470 ;
        RECT 1560.940 2.400 1561.080 24.150 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1918.520 2615.490 1918.580 ;
        RECT 2658.410 1918.520 2658.730 1918.580 ;
        RECT 2615.170 1918.380 2658.730 1918.520 ;
        RECT 2615.170 1918.320 2615.490 1918.380 ;
        RECT 2658.410 1918.320 2658.730 1918.380 ;
        RECT 1579.710 238.920 1580.030 238.980 ;
        RECT 2658.410 238.920 2658.730 238.980 ;
        RECT 1579.710 238.780 2658.730 238.920 ;
        RECT 1579.710 238.720 1580.030 238.780 ;
        RECT 2658.410 238.720 2658.730 238.780 ;
        RECT 1579.710 62.460 1580.030 62.520 ;
        RECT 1578.880 62.320 1580.030 62.460 ;
        RECT 1578.880 62.180 1579.020 62.320 ;
        RECT 1579.710 62.260 1580.030 62.320 ;
        RECT 1578.790 61.920 1579.110 62.180 ;
      LAYER via ;
        RECT 2615.200 1918.320 2615.460 1918.580 ;
        RECT 2658.440 1918.320 2658.700 1918.580 ;
        RECT 1579.740 238.720 1580.000 238.980 ;
        RECT 2658.440 238.720 2658.700 238.980 ;
        RECT 1579.740 62.260 1580.000 62.520 ;
        RECT 1578.820 61.920 1579.080 62.180 ;
      LAYER met2 ;
        RECT 2615.190 1923.195 2615.470 1923.565 ;
        RECT 2615.260 1918.610 2615.400 1923.195 ;
        RECT 2615.200 1918.290 2615.460 1918.610 ;
        RECT 2658.440 1918.290 2658.700 1918.610 ;
        RECT 2658.500 239.010 2658.640 1918.290 ;
        RECT 1579.740 238.690 1580.000 239.010 ;
        RECT 2658.440 238.690 2658.700 239.010 ;
        RECT 1579.800 62.550 1579.940 238.690 ;
        RECT 1579.740 62.230 1580.000 62.550 ;
        RECT 1578.820 61.890 1579.080 62.210 ;
        RECT 1578.880 2.400 1579.020 61.890 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1923.240 2615.470 1923.520 ;
      LAYER met3 ;
        RECT 2606.000 1923.530 2610.000 1923.920 ;
        RECT 2615.165 1923.530 2615.495 1923.545 ;
        RECT 2606.000 1923.320 2615.495 1923.530 ;
        RECT 2609.580 1923.230 2615.495 1923.320 ;
        RECT 2615.165 1923.215 2615.495 1923.230 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1920.110 3266.960 1920.430 3267.020 ;
        RECT 2643.230 3266.960 2643.550 3267.020 ;
        RECT 1920.110 3266.820 2643.550 3266.960 ;
        RECT 1920.110 3266.760 1920.430 3266.820 ;
        RECT 2643.230 3266.760 2643.550 3266.820 ;
        RECT 1596.270 20.640 1596.590 20.700 ;
        RECT 1600.410 20.640 1600.730 20.700 ;
        RECT 1596.270 20.500 1600.730 20.640 ;
        RECT 1596.270 20.440 1596.590 20.500 ;
        RECT 1600.410 20.440 1600.730 20.500 ;
      LAYER via ;
        RECT 1920.140 3266.760 1920.400 3267.020 ;
        RECT 2643.260 3266.760 2643.520 3267.020 ;
        RECT 1596.300 20.440 1596.560 20.700 ;
        RECT 1600.440 20.440 1600.700 20.700 ;
      LAYER met2 ;
        RECT 1920.140 3266.730 1920.400 3267.050 ;
        RECT 2643.260 3266.730 2643.520 3267.050 ;
        RECT 1920.200 3260.000 1920.340 3266.730 ;
        RECT 1920.090 3256.000 1920.370 3260.000 ;
        RECT 2643.320 400.365 2643.460 3266.730 ;
        RECT 2643.250 399.995 2643.530 400.365 ;
        RECT 1600.430 233.395 1600.710 233.765 ;
        RECT 1600.500 20.730 1600.640 233.395 ;
        RECT 1596.300 20.410 1596.560 20.730 ;
        RECT 1600.440 20.410 1600.700 20.730 ;
        RECT 1596.360 2.400 1596.500 20.410 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
      LAYER via2 ;
        RECT 2643.250 400.040 2643.530 400.320 ;
        RECT 1600.430 233.440 1600.710 233.720 ;
      LAYER met3 ;
        RECT 2612.150 400.330 2612.530 400.340 ;
        RECT 2643.225 400.330 2643.555 400.345 ;
        RECT 2612.150 400.030 2643.555 400.330 ;
        RECT 2612.150 400.020 2612.530 400.030 ;
        RECT 2643.225 400.015 2643.555 400.030 ;
        RECT 1600.405 233.730 1600.735 233.745 ;
        RECT 2592.830 233.730 2593.210 233.740 ;
        RECT 1600.405 233.430 2593.210 233.730 ;
        RECT 1600.405 233.415 1600.735 233.430 ;
        RECT 2592.830 233.420 2593.210 233.430 ;
      LAYER via3 ;
        RECT 2612.180 400.020 2612.500 400.340 ;
        RECT 2592.860 233.420 2593.180 233.740 ;
      LAYER met4 ;
        RECT 2612.175 400.015 2612.505 400.345 ;
        RECT 2612.190 379.690 2612.490 400.015 ;
        RECT 2592.430 378.510 2593.610 379.690 ;
        RECT 2611.750 378.510 2612.930 379.690 ;
        RECT 2592.870 233.745 2593.170 378.510 ;
        RECT 2592.855 233.415 2593.185 233.745 ;
      LAYER met5 ;
        RECT 2592.220 378.300 2613.140 379.900 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 218.520 1614.530 218.580 ;
        RECT 2705.330 218.520 2705.650 218.580 ;
        RECT 1614.210 218.380 2705.650 218.520 ;
        RECT 1614.210 218.320 1614.530 218.380 ;
        RECT 2705.330 218.320 2705.650 218.380 ;
      LAYER via ;
        RECT 1614.240 218.320 1614.500 218.580 ;
        RECT 2705.360 218.320 2705.620 218.580 ;
      LAYER met2 ;
        RECT 2450.050 3264.155 2450.330 3264.525 ;
        RECT 2705.350 3264.155 2705.630 3264.525 ;
        RECT 2450.120 3260.000 2450.260 3264.155 ;
        RECT 2450.010 3256.000 2450.290 3260.000 ;
        RECT 2705.420 218.610 2705.560 3264.155 ;
        RECT 1614.240 218.290 1614.500 218.610 ;
        RECT 2705.360 218.290 2705.620 218.610 ;
        RECT 1614.300 2.400 1614.440 218.290 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
      LAYER via2 ;
        RECT 2450.050 3264.200 2450.330 3264.480 ;
        RECT 2705.350 3264.200 2705.630 3264.480 ;
      LAYER met3 ;
        RECT 2450.025 3264.490 2450.355 3264.505 ;
        RECT 2705.325 3264.490 2705.655 3264.505 ;
        RECT 2450.025 3264.190 2705.655 3264.490 ;
        RECT 2450.025 3264.175 2450.355 3264.190 ;
        RECT 2705.325 3264.175 2705.655 3264.190 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 3022.500 2615.490 3022.560 ;
        RECT 2678.190 3022.500 2678.510 3022.560 ;
        RECT 2615.170 3022.360 2678.510 3022.500 ;
        RECT 2615.170 3022.300 2615.490 3022.360 ;
        RECT 2678.190 3022.300 2678.510 3022.360 ;
        RECT 1634.910 239.260 1635.230 239.320 ;
        RECT 2678.190 239.260 2678.510 239.320 ;
        RECT 1634.910 239.120 2678.510 239.260 ;
        RECT 1634.910 239.060 1635.230 239.120 ;
        RECT 2678.190 239.060 2678.510 239.120 ;
        RECT 1632.150 20.640 1632.470 20.700 ;
        RECT 1634.910 20.640 1635.230 20.700 ;
        RECT 1632.150 20.500 1635.230 20.640 ;
        RECT 1632.150 20.440 1632.470 20.500 ;
        RECT 1634.910 20.440 1635.230 20.500 ;
      LAYER via ;
        RECT 2615.200 3022.300 2615.460 3022.560 ;
        RECT 2678.220 3022.300 2678.480 3022.560 ;
        RECT 1634.940 239.060 1635.200 239.320 ;
        RECT 2678.220 239.060 2678.480 239.320 ;
        RECT 1632.180 20.440 1632.440 20.700 ;
        RECT 1634.940 20.440 1635.200 20.700 ;
      LAYER met2 ;
        RECT 2615.190 3023.435 2615.470 3023.805 ;
        RECT 2615.260 3022.590 2615.400 3023.435 ;
        RECT 2615.200 3022.270 2615.460 3022.590 ;
        RECT 2678.220 3022.270 2678.480 3022.590 ;
        RECT 2678.280 239.350 2678.420 3022.270 ;
        RECT 1634.940 239.030 1635.200 239.350 ;
        RECT 2678.220 239.030 2678.480 239.350 ;
        RECT 1635.000 20.730 1635.140 239.030 ;
        RECT 1632.180 20.410 1632.440 20.730 ;
        RECT 1634.940 20.410 1635.200 20.730 ;
        RECT 1632.240 2.400 1632.380 20.410 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
      LAYER via2 ;
        RECT 2615.190 3023.480 2615.470 3023.760 ;
      LAYER met3 ;
        RECT 2606.000 3023.770 2610.000 3024.160 ;
        RECT 2615.165 3023.770 2615.495 3023.785 ;
        RECT 2606.000 3023.560 2615.495 3023.770 ;
        RECT 2609.580 3023.470 2615.495 3023.560 ;
        RECT 2615.165 3023.455 2615.495 3023.470 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 3105.120 2615.490 3105.180 ;
        RECT 2691.990 3105.120 2692.310 3105.180 ;
        RECT 2615.170 3104.980 2692.310 3105.120 ;
        RECT 2615.170 3104.920 2615.490 3104.980 ;
        RECT 2691.990 3104.920 2692.310 3104.980 ;
        RECT 1655.610 234.160 1655.930 234.220 ;
        RECT 2691.990 234.160 2692.310 234.220 ;
        RECT 1655.610 234.020 2692.310 234.160 ;
        RECT 1655.610 233.960 1655.930 234.020 ;
        RECT 2691.990 233.960 2692.310 234.020 ;
        RECT 1650.090 20.640 1650.410 20.700 ;
        RECT 1655.610 20.640 1655.930 20.700 ;
        RECT 1650.090 20.500 1655.930 20.640 ;
        RECT 1650.090 20.440 1650.410 20.500 ;
        RECT 1655.610 20.440 1655.930 20.500 ;
      LAYER via ;
        RECT 2615.200 3104.920 2615.460 3105.180 ;
        RECT 2692.020 3104.920 2692.280 3105.180 ;
        RECT 1655.640 233.960 1655.900 234.220 ;
        RECT 2692.020 233.960 2692.280 234.220 ;
        RECT 1650.120 20.440 1650.380 20.700 ;
        RECT 1655.640 20.440 1655.900 20.700 ;
      LAYER met2 ;
        RECT 2615.190 3107.755 2615.470 3108.125 ;
        RECT 2615.260 3105.210 2615.400 3107.755 ;
        RECT 2615.200 3104.890 2615.460 3105.210 ;
        RECT 2692.020 3104.890 2692.280 3105.210 ;
        RECT 2692.080 234.250 2692.220 3104.890 ;
        RECT 1655.640 233.930 1655.900 234.250 ;
        RECT 2692.020 233.930 2692.280 234.250 ;
        RECT 1655.700 20.730 1655.840 233.930 ;
        RECT 1650.120 20.410 1650.380 20.730 ;
        RECT 1655.640 20.410 1655.900 20.730 ;
        RECT 1650.180 2.400 1650.320 20.410 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
      LAYER via2 ;
        RECT 2615.190 3107.800 2615.470 3108.080 ;
      LAYER met3 ;
        RECT 2606.000 3108.090 2610.000 3108.480 ;
        RECT 2615.165 3108.090 2615.495 3108.105 ;
        RECT 2606.000 3107.880 2615.495 3108.090 ;
        RECT 2609.580 3107.790 2615.495 3107.880 ;
        RECT 2615.165 3107.775 2615.495 3107.790 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1669.485 41.565 1669.655 89.675 ;
      LAYER mcon ;
        RECT 1669.485 89.505 1669.655 89.675 ;
      LAYER met1 ;
        RECT 1669.410 134.880 1669.730 134.940 ;
        RECT 2484.070 134.880 2484.390 134.940 ;
        RECT 1669.410 134.740 2484.390 134.880 ;
        RECT 1669.410 134.680 1669.730 134.740 ;
        RECT 2484.070 134.680 2484.390 134.740 ;
        RECT 1669.410 89.660 1669.730 89.720 ;
        RECT 1669.215 89.520 1669.730 89.660 ;
        RECT 1669.410 89.460 1669.730 89.520 ;
        RECT 1669.410 41.720 1669.730 41.780 ;
        RECT 1669.215 41.580 1669.730 41.720 ;
        RECT 1669.410 41.520 1669.730 41.580 ;
      LAYER via ;
        RECT 1669.440 134.680 1669.700 134.940 ;
        RECT 2484.100 134.680 2484.360 134.940 ;
        RECT 1669.440 89.460 1669.700 89.720 ;
        RECT 1669.440 41.520 1669.700 41.780 ;
      LAYER met2 ;
        RECT 2485.890 260.170 2486.170 264.000 ;
        RECT 2484.160 260.030 2486.170 260.170 ;
        RECT 2484.160 134.970 2484.300 260.030 ;
        RECT 2485.890 260.000 2486.170 260.030 ;
        RECT 1669.440 134.650 1669.700 134.970 ;
        RECT 2484.100 134.650 2484.360 134.970 ;
        RECT 1669.500 89.750 1669.640 134.650 ;
        RECT 1669.440 89.430 1669.700 89.750 ;
        RECT 1669.440 41.490 1669.700 41.810 ;
        RECT 1669.500 14.690 1669.640 41.490 ;
        RECT 1668.580 14.550 1669.640 14.690 ;
        RECT 1668.580 10.610 1668.720 14.550 ;
        RECT 1668.120 10.470 1668.720 10.610 ;
        RECT 1668.120 2.400 1668.260 10.470 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 421.160 2615.490 421.220 ;
        RECT 2644.610 421.160 2644.930 421.220 ;
        RECT 2615.170 421.020 2644.930 421.160 ;
        RECT 2615.170 420.960 2615.490 421.020 ;
        RECT 2644.610 420.960 2644.930 421.020 ;
        RECT 1690.110 239.600 1690.430 239.660 ;
        RECT 2644.610 239.600 2644.930 239.660 ;
        RECT 1690.110 239.460 2644.930 239.600 ;
        RECT 1690.110 239.400 1690.430 239.460 ;
        RECT 2644.610 239.400 2644.930 239.460 ;
        RECT 1685.510 16.560 1685.830 16.620 ;
        RECT 1690.110 16.560 1690.430 16.620 ;
        RECT 1685.510 16.420 1690.430 16.560 ;
        RECT 1685.510 16.360 1685.830 16.420 ;
        RECT 1690.110 16.360 1690.430 16.420 ;
      LAYER via ;
        RECT 2615.200 420.960 2615.460 421.220 ;
        RECT 2644.640 420.960 2644.900 421.220 ;
        RECT 1690.140 239.400 1690.400 239.660 ;
        RECT 2644.640 239.400 2644.900 239.660 ;
        RECT 1685.540 16.360 1685.800 16.620 ;
        RECT 1690.140 16.360 1690.400 16.620 ;
      LAYER met2 ;
        RECT 2615.190 423.115 2615.470 423.485 ;
        RECT 2615.260 421.250 2615.400 423.115 ;
        RECT 2615.200 420.930 2615.460 421.250 ;
        RECT 2644.640 420.930 2644.900 421.250 ;
        RECT 2644.700 239.690 2644.840 420.930 ;
        RECT 1690.140 239.370 1690.400 239.690 ;
        RECT 2644.640 239.370 2644.900 239.690 ;
        RECT 1690.200 16.650 1690.340 239.370 ;
        RECT 1685.540 16.330 1685.800 16.650 ;
        RECT 1690.140 16.330 1690.400 16.650 ;
        RECT 1685.600 2.400 1685.740 16.330 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
      LAYER via2 ;
        RECT 2615.190 423.160 2615.470 423.440 ;
      LAYER met3 ;
        RECT 2606.000 423.450 2610.000 423.840 ;
        RECT 2615.165 423.450 2615.495 423.465 ;
        RECT 2606.000 423.240 2615.495 423.450 ;
        RECT 2609.580 423.150 2615.495 423.240 ;
        RECT 2615.165 423.135 2615.495 423.150 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 724.185 41.565 724.355 89.675 ;
      LAYER mcon ;
        RECT 724.185 89.505 724.355 89.675 ;
      LAYER met1 ;
        RECT 724.110 168.880 724.430 168.940 ;
        RECT 2125.730 168.880 2126.050 168.940 ;
        RECT 724.110 168.740 2126.050 168.880 ;
        RECT 724.110 168.680 724.430 168.740 ;
        RECT 2125.730 168.680 2126.050 168.740 ;
        RECT 723.650 96.800 723.970 96.860 ;
        RECT 724.110 96.800 724.430 96.860 ;
        RECT 723.650 96.660 724.430 96.800 ;
        RECT 723.650 96.600 723.970 96.660 ;
        RECT 724.110 96.600 724.430 96.660 ;
        RECT 724.110 89.660 724.430 89.720 ;
        RECT 723.915 89.520 724.430 89.660 ;
        RECT 724.110 89.460 724.430 89.520 ;
        RECT 724.110 41.720 724.430 41.780 ;
        RECT 723.915 41.580 724.430 41.720 ;
        RECT 724.110 41.520 724.430 41.580 ;
        RECT 724.110 14.180 724.430 14.240 ;
        RECT 722.360 14.040 724.430 14.180 ;
        RECT 722.360 13.900 722.500 14.040 ;
        RECT 724.110 13.980 724.430 14.040 ;
        RECT 722.270 13.640 722.590 13.900 ;
      LAYER via ;
        RECT 724.140 168.680 724.400 168.940 ;
        RECT 2125.760 168.680 2126.020 168.940 ;
        RECT 723.680 96.600 723.940 96.860 ;
        RECT 724.140 96.600 724.400 96.860 ;
        RECT 724.140 89.460 724.400 89.720 ;
        RECT 724.140 41.520 724.400 41.780 ;
        RECT 724.140 13.980 724.400 14.240 ;
        RECT 722.300 13.640 722.560 13.900 ;
      LAYER met2 ;
        RECT 2128.010 260.170 2128.290 264.000 ;
        RECT 2125.820 260.030 2128.290 260.170 ;
        RECT 2125.820 168.970 2125.960 260.030 ;
        RECT 2128.010 260.000 2128.290 260.030 ;
        RECT 724.140 168.650 724.400 168.970 ;
        RECT 2125.760 168.650 2126.020 168.970 ;
        RECT 724.200 98.330 724.340 168.650 ;
        RECT 723.740 98.190 724.340 98.330 ;
        RECT 723.740 96.890 723.880 98.190 ;
        RECT 723.680 96.570 723.940 96.890 ;
        RECT 724.140 96.570 724.400 96.890 ;
        RECT 724.200 89.750 724.340 96.570 ;
        RECT 724.140 89.430 724.400 89.750 ;
        RECT 724.140 41.490 724.400 41.810 ;
        RECT 724.200 14.270 724.340 41.490 ;
        RECT 724.140 13.950 724.400 14.270 ;
        RECT 722.300 13.610 722.560 13.930 ;
        RECT 722.360 2.400 722.500 13.610 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 266.410 1083.480 266.730 1083.540 ;
        RECT 296.770 1083.480 297.090 1083.540 ;
        RECT 266.410 1083.340 297.090 1083.480 ;
        RECT 266.410 1083.280 266.730 1083.340 ;
        RECT 296.770 1083.280 297.090 1083.340 ;
        RECT 266.410 47.500 266.730 47.560 ;
        RECT 1703.450 47.500 1703.770 47.560 ;
        RECT 266.410 47.360 1703.770 47.500 ;
        RECT 266.410 47.300 266.730 47.360 ;
        RECT 1703.450 47.300 1703.770 47.360 ;
      LAYER via ;
        RECT 266.440 1083.280 266.700 1083.540 ;
        RECT 296.800 1083.280 297.060 1083.540 ;
        RECT 266.440 47.300 266.700 47.560 ;
        RECT 1703.480 47.300 1703.740 47.560 ;
      LAYER met2 ;
        RECT 296.790 1088.155 297.070 1088.525 ;
        RECT 296.860 1083.570 297.000 1088.155 ;
        RECT 266.440 1083.250 266.700 1083.570 ;
        RECT 296.800 1083.250 297.060 1083.570 ;
        RECT 266.500 47.590 266.640 1083.250 ;
        RECT 266.440 47.270 266.700 47.590 ;
        RECT 1703.480 47.270 1703.740 47.590 ;
        RECT 1703.540 2.400 1703.680 47.270 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
      LAYER via2 ;
        RECT 296.790 1088.200 297.070 1088.480 ;
      LAYER met3 ;
        RECT 296.765 1088.490 297.095 1088.505 ;
        RECT 310.000 1088.490 314.000 1088.880 ;
        RECT 296.765 1088.280 314.000 1088.490 ;
        RECT 296.765 1088.190 310.500 1088.280 ;
        RECT 296.765 1088.175 297.095 1088.190 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.450 3256.220 1979.770 3256.480 ;
        RECT 1979.540 3254.040 1979.680 3256.220 ;
        RECT 2686.010 3254.040 2686.330 3254.100 ;
        RECT 1979.540 3253.900 2686.330 3254.040 ;
        RECT 2686.010 3253.840 2686.330 3253.900 ;
        RECT 2480.390 231.780 2480.710 231.840 ;
        RECT 2686.010 231.780 2686.330 231.840 ;
        RECT 2480.390 231.640 2686.330 231.780 ;
        RECT 2480.390 231.580 2480.710 231.640 ;
        RECT 2686.010 231.580 2686.330 231.640 ;
        RECT 1721.390 19.620 1721.710 19.680 ;
        RECT 2480.390 19.620 2480.710 19.680 ;
        RECT 1721.390 19.480 2480.710 19.620 ;
        RECT 1721.390 19.420 1721.710 19.480 ;
        RECT 2480.390 19.420 2480.710 19.480 ;
      LAYER via ;
        RECT 1979.480 3256.220 1979.740 3256.480 ;
        RECT 2686.040 3253.840 2686.300 3254.100 ;
        RECT 2480.420 231.580 2480.680 231.840 ;
        RECT 2686.040 231.580 2686.300 231.840 ;
        RECT 1721.420 19.420 1721.680 19.680 ;
        RECT 2480.420 19.420 2480.680 19.680 ;
      LAYER met2 ;
        RECT 1978.050 3256.930 1978.330 3260.000 ;
        RECT 1978.050 3256.790 1979.680 3256.930 ;
        RECT 1978.050 3256.000 1978.330 3256.790 ;
        RECT 1979.540 3256.510 1979.680 3256.790 ;
        RECT 1979.480 3256.190 1979.740 3256.510 ;
        RECT 2686.040 3253.810 2686.300 3254.130 ;
        RECT 2686.100 231.870 2686.240 3253.810 ;
        RECT 2480.420 231.550 2480.680 231.870 ;
        RECT 2686.040 231.550 2686.300 231.870 ;
        RECT 2480.480 19.710 2480.620 231.550 ;
        RECT 1721.420 19.390 1721.680 19.710 ;
        RECT 2480.420 19.390 2480.680 19.710 ;
        RECT 1721.480 2.400 1721.620 19.390 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 676.500 2615.490 676.560 ;
        RECT 2653.810 676.500 2654.130 676.560 ;
        RECT 2615.170 676.360 2654.130 676.500 ;
        RECT 2615.170 676.300 2615.490 676.360 ;
        RECT 2653.810 676.300 2654.130 676.360 ;
        RECT 1745.310 237.560 1745.630 237.620 ;
        RECT 2653.810 237.560 2654.130 237.620 ;
        RECT 1745.310 237.420 2654.130 237.560 ;
        RECT 1745.310 237.360 1745.630 237.420 ;
        RECT 2653.810 237.360 2654.130 237.420 ;
        RECT 1739.330 20.640 1739.650 20.700 ;
        RECT 1745.310 20.640 1745.630 20.700 ;
        RECT 1739.330 20.500 1745.630 20.640 ;
        RECT 1739.330 20.440 1739.650 20.500 ;
        RECT 1745.310 20.440 1745.630 20.500 ;
      LAYER via ;
        RECT 2615.200 676.300 2615.460 676.560 ;
        RECT 2653.840 676.300 2654.100 676.560 ;
        RECT 1745.340 237.360 1745.600 237.620 ;
        RECT 2653.840 237.360 2654.100 237.620 ;
        RECT 1739.360 20.440 1739.620 20.700 ;
        RECT 1745.340 20.440 1745.600 20.700 ;
      LAYER met2 ;
        RECT 2615.200 676.445 2615.460 676.590 ;
        RECT 2615.190 676.075 2615.470 676.445 ;
        RECT 2653.840 676.270 2654.100 676.590 ;
        RECT 2653.900 237.650 2654.040 676.270 ;
        RECT 1745.340 237.330 1745.600 237.650 ;
        RECT 2653.840 237.330 2654.100 237.650 ;
        RECT 1745.400 20.730 1745.540 237.330 ;
        RECT 1739.360 20.410 1739.620 20.730 ;
        RECT 1745.340 20.410 1745.600 20.730 ;
        RECT 1739.420 2.400 1739.560 20.410 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
      LAYER via2 ;
        RECT 2615.190 676.120 2615.470 676.400 ;
      LAYER met3 ;
        RECT 2606.000 676.410 2610.000 676.800 ;
        RECT 2615.165 676.410 2615.495 676.425 ;
        RECT 2606.000 676.200 2615.495 676.410 ;
        RECT 2609.580 676.110 2615.495 676.200 ;
        RECT 2615.165 676.095 2615.495 676.110 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 305.970 232.800 306.290 232.860 ;
        RECT 1752.670 232.800 1752.990 232.860 ;
        RECT 305.970 232.660 1752.990 232.800 ;
        RECT 305.970 232.600 306.290 232.660 ;
        RECT 1752.670 232.600 1752.990 232.660 ;
        RECT 1752.670 37.640 1752.990 37.700 ;
        RECT 1756.810 37.640 1757.130 37.700 ;
        RECT 1752.670 37.500 1757.130 37.640 ;
        RECT 1752.670 37.440 1752.990 37.500 ;
        RECT 1756.810 37.440 1757.130 37.500 ;
      LAYER via ;
        RECT 306.000 232.600 306.260 232.860 ;
        RECT 1752.700 232.600 1752.960 232.860 ;
        RECT 1752.700 37.440 1752.960 37.700 ;
        RECT 1756.840 37.440 1757.100 37.700 ;
      LAYER met2 ;
        RECT 305.990 1870.155 306.270 1870.525 ;
        RECT 306.060 232.890 306.200 1870.155 ;
        RECT 306.000 232.570 306.260 232.890 ;
        RECT 1752.700 232.570 1752.960 232.890 ;
        RECT 1752.760 37.730 1752.900 232.570 ;
        RECT 1752.700 37.410 1752.960 37.730 ;
        RECT 1756.840 37.410 1757.100 37.730 ;
        RECT 1756.900 2.400 1757.040 37.410 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
      LAYER via2 ;
        RECT 305.990 1870.200 306.270 1870.480 ;
      LAYER met3 ;
        RECT 305.965 1870.490 306.295 1870.505 ;
        RECT 310.000 1870.490 314.000 1870.880 ;
        RECT 305.965 1870.280 314.000 1870.490 ;
        RECT 305.965 1870.190 310.500 1870.280 ;
        RECT 305.965 1870.175 306.295 1870.190 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1906.310 3267.300 1906.630 3267.360 ;
        RECT 2608.730 3267.300 2609.050 3267.360 ;
        RECT 1906.310 3267.160 2609.050 3267.300 ;
        RECT 1906.310 3267.100 1906.630 3267.160 ;
        RECT 2608.730 3267.100 2609.050 3267.160 ;
        RECT 1779.810 253.880 1780.130 253.940 ;
        RECT 2633.110 253.880 2633.430 253.940 ;
        RECT 1779.810 253.740 2633.430 253.880 ;
        RECT 1779.810 253.680 1780.130 253.740 ;
        RECT 2633.110 253.680 2633.430 253.740 ;
        RECT 1774.750 15.200 1775.070 15.260 ;
        RECT 1779.810 15.200 1780.130 15.260 ;
        RECT 1774.750 15.060 1780.130 15.200 ;
        RECT 1774.750 15.000 1775.070 15.060 ;
        RECT 1779.810 15.000 1780.130 15.060 ;
      LAYER via ;
        RECT 1906.340 3267.100 1906.600 3267.360 ;
        RECT 2608.760 3267.100 2609.020 3267.360 ;
        RECT 1779.840 253.680 1780.100 253.940 ;
        RECT 2633.140 253.680 2633.400 253.940 ;
        RECT 1774.780 15.000 1775.040 15.260 ;
        RECT 1779.840 15.000 1780.100 15.260 ;
      LAYER met2 ;
        RECT 1906.340 3267.070 1906.600 3267.390 ;
        RECT 2608.760 3267.070 2609.020 3267.390 ;
        RECT 1906.400 3260.000 1906.540 3267.070 ;
        RECT 1906.290 3256.000 1906.570 3260.000 ;
        RECT 2608.820 497.605 2608.960 3267.070 ;
        RECT 2608.750 497.235 2609.030 497.605 ;
        RECT 2607.830 433.995 2608.110 434.365 ;
        RECT 2607.900 386.765 2608.040 433.995 ;
        RECT 2607.830 386.395 2608.110 386.765 ;
        RECT 2633.130 385.035 2633.410 385.405 ;
        RECT 2633.200 253.970 2633.340 385.035 ;
        RECT 1779.840 253.650 1780.100 253.970 ;
        RECT 2633.140 253.650 2633.400 253.970 ;
        RECT 1779.900 15.290 1780.040 253.650 ;
        RECT 1774.780 14.970 1775.040 15.290 ;
        RECT 1779.840 14.970 1780.100 15.290 ;
        RECT 1774.840 2.400 1774.980 14.970 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
      LAYER via2 ;
        RECT 2608.750 497.280 2609.030 497.560 ;
        RECT 2607.830 434.040 2608.110 434.320 ;
        RECT 2607.830 386.440 2608.110 386.720 ;
        RECT 2633.130 385.080 2633.410 385.360 ;
      LAYER met3 ;
        RECT 2607.550 497.570 2607.930 497.580 ;
        RECT 2608.725 497.570 2609.055 497.585 ;
        RECT 2607.550 497.270 2609.055 497.570 ;
        RECT 2607.550 497.260 2607.930 497.270 ;
        RECT 2608.725 497.255 2609.055 497.270 ;
        RECT 2607.805 434.340 2608.135 434.345 ;
        RECT 2607.550 434.330 2608.135 434.340 ;
        RECT 2607.350 434.030 2608.135 434.330 ;
        RECT 2607.550 434.020 2608.135 434.030 ;
        RECT 2607.805 434.015 2608.135 434.020 ;
        RECT 2606.630 386.730 2607.010 386.740 ;
        RECT 2607.805 386.730 2608.135 386.745 ;
        RECT 2606.630 386.430 2608.135 386.730 ;
        RECT 2606.630 386.420 2607.010 386.430 ;
        RECT 2607.805 386.415 2608.135 386.430 ;
        RECT 2606.630 385.370 2607.010 385.380 ;
        RECT 2633.105 385.370 2633.435 385.385 ;
        RECT 2606.630 385.070 2633.435 385.370 ;
        RECT 2606.630 385.060 2607.010 385.070 ;
        RECT 2633.105 385.055 2633.435 385.070 ;
      LAYER via3 ;
        RECT 2607.580 497.260 2607.900 497.580 ;
        RECT 2607.580 434.020 2607.900 434.340 ;
        RECT 2606.660 386.420 2606.980 386.740 ;
        RECT 2606.660 385.060 2606.980 385.380 ;
      LAYER met4 ;
        RECT 2607.575 497.255 2607.905 497.585 ;
        RECT 2607.590 434.345 2607.890 497.255 ;
        RECT 2607.575 434.015 2607.905 434.345 ;
        RECT 2606.655 386.415 2606.985 386.745 ;
        RECT 2606.670 385.385 2606.970 386.415 ;
        RECT 2606.655 385.055 2606.985 385.385 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 300.450 212.060 300.770 212.120 ;
        RECT 1787.170 212.060 1787.490 212.120 ;
        RECT 300.450 211.920 1787.490 212.060 ;
        RECT 300.450 211.860 300.770 211.920 ;
        RECT 1787.170 211.860 1787.490 211.920 ;
        RECT 1787.170 62.120 1787.490 62.180 ;
        RECT 1792.690 62.120 1793.010 62.180 ;
        RECT 1787.170 61.980 1793.010 62.120 ;
        RECT 1787.170 61.920 1787.490 61.980 ;
        RECT 1792.690 61.920 1793.010 61.980 ;
      LAYER via ;
        RECT 300.480 211.860 300.740 212.120 ;
        RECT 1787.200 211.860 1787.460 212.120 ;
        RECT 1787.200 61.920 1787.460 62.180 ;
        RECT 1792.720 61.920 1792.980 62.180 ;
      LAYER met2 ;
        RECT 300.470 559.115 300.750 559.485 ;
        RECT 300.540 212.150 300.680 559.115 ;
        RECT 300.480 211.830 300.740 212.150 ;
        RECT 1787.200 211.830 1787.460 212.150 ;
        RECT 1787.260 62.210 1787.400 211.830 ;
        RECT 1787.200 61.890 1787.460 62.210 ;
        RECT 1792.720 61.890 1792.980 62.210 ;
        RECT 1792.780 2.400 1792.920 61.890 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
      LAYER via2 ;
        RECT 300.470 559.160 300.750 559.440 ;
      LAYER met3 ;
        RECT 300.445 559.450 300.775 559.465 ;
        RECT 310.000 559.450 314.000 559.840 ;
        RECT 300.445 559.240 314.000 559.450 ;
        RECT 300.445 559.150 310.500 559.240 ;
        RECT 300.445 559.135 300.775 559.150 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1871.425 24.225 1871.595 26.095 ;
      LAYER mcon ;
        RECT 1871.425 25.925 1871.595 26.095 ;
      LAYER met1 ;
        RECT 1871.365 26.080 1871.655 26.125 ;
        RECT 1925.170 26.080 1925.490 26.140 ;
        RECT 1871.365 25.940 1925.490 26.080 ;
        RECT 1871.365 25.895 1871.655 25.940 ;
        RECT 1925.170 25.880 1925.490 25.940 ;
        RECT 1810.630 24.380 1810.950 24.440 ;
        RECT 1871.365 24.380 1871.655 24.425 ;
        RECT 1810.630 24.240 1871.655 24.380 ;
        RECT 1810.630 24.180 1810.950 24.240 ;
        RECT 1871.365 24.195 1871.655 24.240 ;
      LAYER via ;
        RECT 1925.200 25.880 1925.460 26.140 ;
        RECT 1810.660 24.180 1810.920 24.440 ;
      LAYER met2 ;
        RECT 1928.370 260.170 1928.650 264.000 ;
        RECT 1925.260 260.030 1928.650 260.170 ;
        RECT 1925.260 26.170 1925.400 260.030 ;
        RECT 1928.370 260.000 1928.650 260.030 ;
        RECT 1925.200 25.850 1925.460 26.170 ;
        RECT 1810.660 24.150 1810.920 24.470 ;
        RECT 1810.720 2.400 1810.860 24.150 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1642.440 2615.490 1642.500 ;
        RECT 2686.930 1642.440 2687.250 1642.500 ;
        RECT 2615.170 1642.300 2687.250 1642.440 ;
        RECT 2615.170 1642.240 2615.490 1642.300 ;
        RECT 2686.930 1642.240 2687.250 1642.300 ;
        RECT 1835.010 232.800 1835.330 232.860 ;
        RECT 2686.930 232.800 2687.250 232.860 ;
        RECT 1835.010 232.660 2687.250 232.800 ;
        RECT 1835.010 232.600 1835.330 232.660 ;
        RECT 2686.930 232.600 2687.250 232.660 ;
        RECT 1828.570 14.860 1828.890 14.920 ;
        RECT 1835.010 14.860 1835.330 14.920 ;
        RECT 1828.570 14.720 1835.330 14.860 ;
        RECT 1828.570 14.660 1828.890 14.720 ;
        RECT 1835.010 14.660 1835.330 14.720 ;
      LAYER via ;
        RECT 2615.200 1642.240 2615.460 1642.500 ;
        RECT 2686.960 1642.240 2687.220 1642.500 ;
        RECT 1835.040 232.600 1835.300 232.860 ;
        RECT 2686.960 232.600 2687.220 232.860 ;
        RECT 1828.600 14.660 1828.860 14.920 ;
        RECT 1835.040 14.660 1835.300 14.920 ;
      LAYER met2 ;
        RECT 2615.190 1648.475 2615.470 1648.845 ;
        RECT 2615.260 1642.530 2615.400 1648.475 ;
        RECT 2615.200 1642.210 2615.460 1642.530 ;
        RECT 2686.960 1642.210 2687.220 1642.530 ;
        RECT 2687.020 232.890 2687.160 1642.210 ;
        RECT 1835.040 232.570 1835.300 232.890 ;
        RECT 2686.960 232.570 2687.220 232.890 ;
        RECT 1835.100 14.950 1835.240 232.570 ;
        RECT 1828.600 14.630 1828.860 14.950 ;
        RECT 1835.040 14.630 1835.300 14.950 ;
        RECT 1828.660 2.400 1828.800 14.630 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1648.520 2615.470 1648.800 ;
      LAYER met3 ;
        RECT 2606.000 1648.810 2610.000 1649.200 ;
        RECT 2615.165 1648.810 2615.495 1648.825 ;
        RECT 2606.000 1648.600 2615.495 1648.810 ;
        RECT 2609.580 1648.510 2615.495 1648.600 ;
        RECT 2615.165 1648.495 2615.495 1648.510 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 314.785 258.145 314.955 265.455 ;
      LAYER mcon ;
        RECT 314.785 265.285 314.955 265.455 ;
      LAYER met1 ;
        RECT 311.950 676.500 312.270 676.560 ;
        RECT 312.870 676.500 313.190 676.560 ;
        RECT 311.950 676.360 313.190 676.500 ;
        RECT 311.950 676.300 312.270 676.360 ;
        RECT 312.870 676.300 313.190 676.360 ;
        RECT 312.870 265.440 313.190 265.500 ;
        RECT 314.725 265.440 315.015 265.485 ;
        RECT 312.870 265.300 315.015 265.440 ;
        RECT 312.870 265.240 313.190 265.300 ;
        RECT 314.725 265.255 315.015 265.300 ;
        RECT 314.710 258.300 315.030 258.360 ;
        RECT 314.515 258.160 315.030 258.300 ;
        RECT 314.710 258.100 315.030 258.160 ;
        RECT 1842.370 62.120 1842.690 62.180 ;
        RECT 1846.050 62.120 1846.370 62.180 ;
        RECT 1842.370 61.980 1846.370 62.120 ;
        RECT 1842.370 61.920 1842.690 61.980 ;
        RECT 1846.050 61.920 1846.370 61.980 ;
      LAYER via ;
        RECT 311.980 676.300 312.240 676.560 ;
        RECT 312.900 676.300 313.160 676.560 ;
        RECT 312.900 265.240 313.160 265.500 ;
        RECT 314.740 258.100 315.000 258.360 ;
        RECT 1842.400 61.920 1842.660 62.180 ;
        RECT 1846.080 61.920 1846.340 62.180 ;
      LAYER met2 ;
        RECT 312.890 2775.915 313.170 2776.285 ;
        RECT 312.960 2766.085 313.100 2775.915 ;
        RECT 312.890 2765.715 313.170 2766.085 ;
        RECT 311.510 2413.475 311.790 2413.845 ;
        RECT 311.580 2367.605 311.720 2413.475 ;
        RECT 311.510 2367.235 311.790 2367.605 ;
        RECT 312.430 2272.715 312.710 2273.085 ;
        RECT 312.500 2270.365 312.640 2272.715 ;
        RECT 312.430 2269.995 312.710 2270.365 ;
        RECT 312.890 2259.795 313.170 2260.165 ;
        RECT 312.960 2224.805 313.100 2259.795 ;
        RECT 312.890 2224.435 313.170 2224.805 ;
        RECT 312.430 2129.915 312.710 2130.285 ;
        RECT 312.500 2109.885 312.640 2129.915 ;
        RECT 312.430 2109.515 312.710 2109.885 ;
        RECT 312.430 2044.915 312.710 2045.285 ;
        RECT 312.500 1980.685 312.640 2044.915 ;
        RECT 312.430 1980.315 312.710 1980.685 ;
        RECT 312.890 1946.315 313.170 1946.685 ;
        RECT 312.960 1895.685 313.100 1946.315 ;
        RECT 312.890 1895.315 313.170 1895.685 ;
        RECT 312.890 1840.915 313.170 1841.285 ;
        RECT 312.960 1835.845 313.100 1840.915 ;
        RECT 312.890 1835.475 313.170 1835.845 ;
        RECT 312.430 1810.995 312.710 1811.365 ;
        RECT 312.500 1733.165 312.640 1810.995 ;
        RECT 312.430 1732.795 312.710 1733.165 ;
        RECT 312.430 1682.475 312.710 1682.845 ;
        RECT 312.500 1611.445 312.640 1682.475 ;
        RECT 312.430 1611.075 312.710 1611.445 ;
        RECT 312.890 1497.515 313.170 1497.885 ;
        RECT 312.960 1491.085 313.100 1497.515 ;
        RECT 312.890 1490.715 313.170 1491.085 ;
        RECT 312.890 1483.235 313.170 1483.605 ;
        RECT 312.960 1446.885 313.100 1483.235 ;
        RECT 312.890 1446.515 313.170 1446.885 ;
        RECT 311.970 765.155 312.250 765.525 ;
        RECT 312.040 717.925 312.180 765.155 ;
        RECT 311.970 717.555 312.250 717.925 ;
        RECT 311.970 716.195 312.250 716.565 ;
        RECT 312.040 676.590 312.180 716.195 ;
        RECT 311.980 676.270 312.240 676.590 ;
        RECT 312.900 676.270 313.160 676.590 ;
        RECT 312.960 621.365 313.100 676.270 ;
        RECT 312.890 620.995 313.170 621.365 ;
        RECT 312.890 619.635 313.170 620.005 ;
        RECT 312.960 552.685 313.100 619.635 ;
        RECT 312.890 552.315 313.170 552.685 ;
        RECT 312.890 514.915 313.170 515.285 ;
        RECT 312.960 484.005 313.100 514.915 ;
        RECT 312.890 483.635 313.170 484.005 ;
        RECT 312.890 450.995 313.170 451.365 ;
        RECT 312.960 435.045 313.100 450.995 ;
        RECT 312.890 434.675 313.170 435.045 ;
        RECT 312.890 433.995 313.170 434.365 ;
        RECT 312.960 410.565 313.100 433.995 ;
        RECT 312.890 410.195 313.170 410.565 ;
        RECT 312.890 370.330 313.170 370.445 ;
        RECT 312.890 370.190 313.560 370.330 ;
        RECT 312.890 370.075 313.170 370.190 ;
        RECT 313.420 339.165 313.560 370.190 ;
        RECT 313.350 338.795 313.630 339.165 ;
        RECT 312.890 265.355 313.170 265.725 ;
        RECT 312.900 265.210 313.160 265.355 ;
        RECT 314.740 258.070 315.000 258.390 ;
        RECT 314.800 257.565 314.940 258.070 ;
        RECT 314.730 257.195 315.010 257.565 ;
        RECT 1842.390 92.635 1842.670 93.005 ;
        RECT 1842.460 62.210 1842.600 92.635 ;
        RECT 1842.400 61.890 1842.660 62.210 ;
        RECT 1846.080 61.890 1846.340 62.210 ;
        RECT 1846.140 2.400 1846.280 61.890 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
      LAYER via2 ;
        RECT 312.890 2775.960 313.170 2776.240 ;
        RECT 312.890 2765.760 313.170 2766.040 ;
        RECT 311.510 2413.520 311.790 2413.800 ;
        RECT 311.510 2367.280 311.790 2367.560 ;
        RECT 312.430 2272.760 312.710 2273.040 ;
        RECT 312.430 2270.040 312.710 2270.320 ;
        RECT 312.890 2259.840 313.170 2260.120 ;
        RECT 312.890 2224.480 313.170 2224.760 ;
        RECT 312.430 2129.960 312.710 2130.240 ;
        RECT 312.430 2109.560 312.710 2109.840 ;
        RECT 312.430 2044.960 312.710 2045.240 ;
        RECT 312.430 1980.360 312.710 1980.640 ;
        RECT 312.890 1946.360 313.170 1946.640 ;
        RECT 312.890 1895.360 313.170 1895.640 ;
        RECT 312.890 1840.960 313.170 1841.240 ;
        RECT 312.890 1835.520 313.170 1835.800 ;
        RECT 312.430 1811.040 312.710 1811.320 ;
        RECT 312.430 1732.840 312.710 1733.120 ;
        RECT 312.430 1682.520 312.710 1682.800 ;
        RECT 312.430 1611.120 312.710 1611.400 ;
        RECT 312.890 1497.560 313.170 1497.840 ;
        RECT 312.890 1490.760 313.170 1491.040 ;
        RECT 312.890 1483.280 313.170 1483.560 ;
        RECT 312.890 1446.560 313.170 1446.840 ;
        RECT 311.970 765.200 312.250 765.480 ;
        RECT 311.970 717.600 312.250 717.880 ;
        RECT 311.970 716.240 312.250 716.520 ;
        RECT 312.890 621.040 313.170 621.320 ;
        RECT 312.890 619.680 313.170 619.960 ;
        RECT 312.890 552.360 313.170 552.640 ;
        RECT 312.890 514.960 313.170 515.240 ;
        RECT 312.890 483.680 313.170 483.960 ;
        RECT 312.890 451.040 313.170 451.320 ;
        RECT 312.890 434.720 313.170 435.000 ;
        RECT 312.890 434.040 313.170 434.320 ;
        RECT 312.890 410.240 313.170 410.520 ;
        RECT 312.890 370.120 313.170 370.400 ;
        RECT 313.350 338.840 313.630 339.120 ;
        RECT 312.890 265.400 313.170 265.680 ;
        RECT 314.730 257.240 315.010 257.520 ;
        RECT 1842.390 92.680 1842.670 92.960 ;
      LAYER met3 ;
        RECT 310.000 2778.760 314.000 2779.360 ;
        RECT 313.110 2776.265 313.410 2778.760 ;
        RECT 312.865 2775.950 313.410 2776.265 ;
        RECT 312.865 2775.935 313.195 2775.950 ;
        RECT 312.865 2766.060 313.195 2766.065 ;
        RECT 312.865 2766.050 313.450 2766.060 ;
        RECT 312.865 2765.750 313.650 2766.050 ;
        RECT 312.865 2765.740 313.450 2765.750 ;
        RECT 312.865 2765.735 313.195 2765.740 ;
        RECT 310.310 2732.050 310.690 2732.060 ;
        RECT 313.070 2732.050 313.450 2732.060 ;
        RECT 310.310 2731.750 313.450 2732.050 ;
        RECT 310.310 2731.740 310.690 2731.750 ;
        RECT 313.070 2731.740 313.450 2731.750 ;
        RECT 310.310 2477.050 310.690 2477.060 ;
        RECT 313.070 2477.050 313.450 2477.060 ;
        RECT 310.310 2476.750 313.450 2477.050 ;
        RECT 310.310 2476.740 310.690 2476.750 ;
        RECT 313.070 2476.740 313.450 2476.750 ;
        RECT 310.310 2447.130 310.690 2447.140 ;
        RECT 310.310 2446.830 311.570 2447.130 ;
        RECT 310.310 2446.820 310.690 2446.830 ;
        RECT 311.270 2445.780 311.570 2446.830 ;
        RECT 311.230 2445.460 311.610 2445.780 ;
        RECT 311.230 2414.180 311.610 2414.500 ;
        RECT 311.270 2413.825 311.570 2414.180 ;
        RECT 311.270 2413.510 311.815 2413.825 ;
        RECT 311.485 2413.495 311.815 2413.510 ;
        RECT 311.485 2367.570 311.815 2367.585 ;
        RECT 313.070 2367.570 313.450 2367.580 ;
        RECT 311.485 2367.270 313.450 2367.570 ;
        RECT 311.485 2367.255 311.815 2367.270 ;
        RECT 313.070 2367.260 313.450 2367.270 ;
        RECT 313.070 2318.980 313.450 2319.300 ;
        RECT 313.110 2317.260 313.410 2318.980 ;
        RECT 313.070 2316.940 313.450 2317.260 ;
        RECT 312.405 2273.050 312.735 2273.065 ;
        RECT 313.070 2273.050 313.450 2273.060 ;
        RECT 312.405 2272.750 313.450 2273.050 ;
        RECT 312.405 2272.735 312.735 2272.750 ;
        RECT 313.070 2272.740 313.450 2272.750 ;
        RECT 312.405 2270.330 312.735 2270.345 ;
        RECT 313.070 2270.330 313.450 2270.340 ;
        RECT 312.405 2270.030 313.450 2270.330 ;
        RECT 312.405 2270.015 312.735 2270.030 ;
        RECT 313.070 2270.020 313.450 2270.030 ;
        RECT 312.865 2260.140 313.195 2260.145 ;
        RECT 312.865 2260.130 313.450 2260.140 ;
        RECT 312.865 2259.830 313.650 2260.130 ;
        RECT 312.865 2259.820 313.450 2259.830 ;
        RECT 312.865 2259.815 313.195 2259.820 ;
        RECT 312.865 2224.780 313.195 2224.785 ;
        RECT 312.865 2224.770 313.450 2224.780 ;
        RECT 312.640 2224.470 313.450 2224.770 ;
        RECT 312.865 2224.460 313.450 2224.470 ;
        RECT 312.865 2224.455 313.195 2224.460 ;
        RECT 312.405 2130.250 312.735 2130.265 ;
        RECT 313.070 2130.250 313.450 2130.260 ;
        RECT 312.405 2129.950 313.450 2130.250 ;
        RECT 312.405 2129.935 312.735 2129.950 ;
        RECT 313.070 2129.940 313.450 2129.950 ;
        RECT 312.405 2109.850 312.735 2109.865 ;
        RECT 313.070 2109.850 313.450 2109.860 ;
        RECT 312.405 2109.550 313.450 2109.850 ;
        RECT 312.405 2109.535 312.735 2109.550 ;
        RECT 313.070 2109.540 313.450 2109.550 ;
        RECT 312.405 2045.250 312.735 2045.265 ;
        RECT 313.070 2045.250 313.450 2045.260 ;
        RECT 312.405 2044.950 313.450 2045.250 ;
        RECT 312.405 2044.935 312.735 2044.950 ;
        RECT 313.070 2044.940 313.450 2044.950 ;
        RECT 312.405 1980.650 312.735 1980.665 ;
        RECT 313.070 1980.650 313.450 1980.660 ;
        RECT 312.405 1980.350 313.450 1980.650 ;
        RECT 312.405 1980.335 312.735 1980.350 ;
        RECT 313.070 1980.340 313.450 1980.350 ;
        RECT 312.865 1946.660 313.195 1946.665 ;
        RECT 312.865 1946.650 313.450 1946.660 ;
        RECT 312.640 1946.350 313.450 1946.650 ;
        RECT 312.865 1946.340 313.450 1946.350 ;
        RECT 312.865 1946.335 313.195 1946.340 ;
        RECT 312.865 1895.660 313.195 1895.665 ;
        RECT 312.865 1895.650 313.450 1895.660 ;
        RECT 312.640 1895.350 313.450 1895.650 ;
        RECT 312.865 1895.340 313.450 1895.350 ;
        RECT 312.865 1895.335 313.195 1895.340 ;
        RECT 312.865 1841.260 313.195 1841.265 ;
        RECT 312.865 1841.250 313.450 1841.260 ;
        RECT 312.640 1840.950 313.450 1841.250 ;
        RECT 312.865 1840.940 313.450 1840.950 ;
        RECT 312.865 1840.935 313.195 1840.940 ;
        RECT 312.865 1835.820 313.195 1835.825 ;
        RECT 312.865 1835.810 313.450 1835.820 ;
        RECT 312.865 1835.510 313.650 1835.810 ;
        RECT 312.865 1835.500 313.450 1835.510 ;
        RECT 312.865 1835.495 313.195 1835.500 ;
        RECT 312.405 1811.330 312.735 1811.345 ;
        RECT 313.070 1811.330 313.450 1811.340 ;
        RECT 312.405 1811.030 313.450 1811.330 ;
        RECT 312.405 1811.015 312.735 1811.030 ;
        RECT 313.070 1811.020 313.450 1811.030 ;
        RECT 312.405 1733.130 312.735 1733.145 ;
        RECT 312.190 1732.815 312.735 1733.130 ;
        RECT 312.190 1732.460 312.490 1732.815 ;
        RECT 312.150 1732.140 312.530 1732.460 ;
        RECT 312.150 1683.180 312.530 1683.500 ;
        RECT 312.190 1682.825 312.490 1683.180 ;
        RECT 312.190 1682.510 312.735 1682.825 ;
        RECT 312.405 1682.495 312.735 1682.510 ;
        RECT 312.405 1611.410 312.735 1611.425 ;
        RECT 313.070 1611.410 313.450 1611.420 ;
        RECT 312.405 1611.110 313.450 1611.410 ;
        RECT 312.405 1611.095 312.735 1611.110 ;
        RECT 313.070 1611.100 313.450 1611.110 ;
        RECT 312.865 1497.860 313.195 1497.865 ;
        RECT 312.865 1497.850 313.450 1497.860 ;
        RECT 312.640 1497.550 313.450 1497.850 ;
        RECT 312.865 1497.540 313.450 1497.550 ;
        RECT 312.865 1497.535 313.195 1497.540 ;
        RECT 312.150 1491.050 312.530 1491.060 ;
        RECT 312.865 1491.050 313.195 1491.065 ;
        RECT 312.150 1490.750 313.195 1491.050 ;
        RECT 312.150 1490.740 312.530 1490.750 ;
        RECT 312.865 1490.735 313.195 1490.750 ;
        RECT 312.150 1483.570 312.530 1483.580 ;
        RECT 312.865 1483.570 313.195 1483.585 ;
        RECT 312.150 1483.270 313.195 1483.570 ;
        RECT 312.150 1483.260 312.530 1483.270 ;
        RECT 312.865 1483.255 313.195 1483.270 ;
        RECT 312.865 1446.860 313.195 1446.865 ;
        RECT 312.865 1446.850 313.450 1446.860 ;
        RECT 312.640 1446.550 313.450 1446.850 ;
        RECT 312.865 1446.540 313.450 1446.550 ;
        RECT 312.865 1446.535 313.195 1446.540 ;
        RECT 311.230 1435.290 311.610 1435.300 ;
        RECT 313.070 1435.290 313.450 1435.300 ;
        RECT 311.230 1434.990 313.450 1435.290 ;
        RECT 311.230 1434.980 311.610 1434.990 ;
        RECT 313.070 1434.980 313.450 1434.990 ;
        RECT 313.070 1256.140 313.450 1256.460 ;
        RECT 313.110 1255.780 313.410 1256.140 ;
        RECT 313.070 1255.460 313.450 1255.780 ;
        RECT 311.230 1217.010 311.610 1217.020 ;
        RECT 313.070 1217.010 313.450 1217.020 ;
        RECT 311.230 1216.710 313.450 1217.010 ;
        RECT 311.230 1216.700 311.610 1216.710 ;
        RECT 313.070 1216.700 313.450 1216.710 ;
        RECT 310.310 1112.290 310.690 1112.300 ;
        RECT 310.310 1111.990 313.410 1112.290 ;
        RECT 310.310 1111.980 310.690 1111.990 ;
        RECT 313.110 1110.940 313.410 1111.990 ;
        RECT 313.070 1110.620 313.450 1110.940 ;
        RECT 311.945 765.490 312.275 765.505 ;
        RECT 313.070 765.490 313.450 765.500 ;
        RECT 311.945 765.190 313.450 765.490 ;
        RECT 311.945 765.175 312.275 765.190 ;
        RECT 313.070 765.180 313.450 765.190 ;
        RECT 311.945 717.900 312.275 717.905 ;
        RECT 311.945 717.890 312.530 717.900 ;
        RECT 311.945 717.590 312.730 717.890 ;
        RECT 311.945 717.580 312.530 717.590 ;
        RECT 311.945 717.575 312.275 717.580 ;
        RECT 312.150 716.900 312.530 717.220 ;
        RECT 312.190 716.545 312.490 716.900 ;
        RECT 311.945 716.230 312.490 716.545 ;
        RECT 311.945 716.215 312.275 716.230 ;
        RECT 312.865 621.330 313.195 621.345 ;
        RECT 312.865 621.015 313.410 621.330 ;
        RECT 313.110 619.985 313.410 621.015 ;
        RECT 312.865 619.670 313.410 619.985 ;
        RECT 312.865 619.655 313.195 619.670 ;
        RECT 312.865 552.660 313.195 552.665 ;
        RECT 312.865 552.650 313.450 552.660 ;
        RECT 312.640 552.350 313.450 552.650 ;
        RECT 312.865 552.340 313.450 552.350 ;
        RECT 312.865 552.335 313.195 552.340 ;
        RECT 312.865 515.260 313.195 515.265 ;
        RECT 312.865 515.250 313.450 515.260 ;
        RECT 312.640 514.950 313.450 515.250 ;
        RECT 312.865 514.940 313.450 514.950 ;
        RECT 312.865 514.935 313.195 514.940 ;
        RECT 312.865 483.980 313.195 483.985 ;
        RECT 312.865 483.970 313.450 483.980 ;
        RECT 312.865 483.670 313.650 483.970 ;
        RECT 312.865 483.660 313.450 483.670 ;
        RECT 312.865 483.655 313.195 483.660 ;
        RECT 312.865 451.340 313.195 451.345 ;
        RECT 312.865 451.330 313.450 451.340 ;
        RECT 312.640 451.030 313.450 451.330 ;
        RECT 312.865 451.020 313.450 451.030 ;
        RECT 312.865 451.015 313.195 451.020 ;
        RECT 312.865 435.010 313.195 435.025 ;
        RECT 312.865 434.695 313.410 435.010 ;
        RECT 313.110 434.345 313.410 434.695 ;
        RECT 312.865 434.030 313.410 434.345 ;
        RECT 312.865 434.015 313.195 434.030 ;
        RECT 312.865 410.530 313.195 410.545 ;
        RECT 312.865 410.215 313.410 410.530 ;
        RECT 313.110 409.180 313.410 410.215 ;
        RECT 313.070 408.860 313.450 409.180 ;
        RECT 312.865 370.420 313.195 370.425 ;
        RECT 312.865 370.410 313.450 370.420 ;
        RECT 312.640 370.110 313.450 370.410 ;
        RECT 312.865 370.100 313.450 370.110 ;
        RECT 312.865 370.095 313.195 370.100 ;
        RECT 313.325 339.130 313.655 339.145 ;
        RECT 313.110 338.815 313.655 339.130 ;
        RECT 313.110 338.460 313.410 338.815 ;
        RECT 313.070 338.140 313.450 338.460 ;
        RECT 312.150 265.690 312.530 265.700 ;
        RECT 312.865 265.690 313.195 265.705 ;
        RECT 312.150 265.390 313.195 265.690 ;
        RECT 312.150 265.380 312.530 265.390 ;
        RECT 312.865 265.375 313.195 265.390 ;
        RECT 314.705 257.530 315.035 257.545 ;
        RECT 316.750 257.530 317.130 257.540 ;
        RECT 314.705 257.230 317.130 257.530 ;
        RECT 314.705 257.215 315.035 257.230 ;
        RECT 316.750 257.220 317.130 257.230 ;
        RECT 313.990 217.410 314.370 217.420 ;
        RECT 316.750 217.410 317.130 217.420 ;
        RECT 313.990 217.110 317.130 217.410 ;
        RECT 313.990 217.100 314.370 217.110 ;
        RECT 316.750 217.100 317.130 217.110 ;
        RECT 313.990 158.930 314.370 158.940 ;
        RECT 316.750 158.930 317.130 158.940 ;
        RECT 313.990 158.630 317.130 158.930 ;
        RECT 313.990 158.620 314.370 158.630 ;
        RECT 316.750 158.620 317.130 158.630 ;
        RECT 314.910 92.970 315.290 92.980 ;
        RECT 1842.365 92.970 1842.695 92.985 ;
        RECT 314.910 92.670 1842.695 92.970 ;
        RECT 314.910 92.660 315.290 92.670 ;
        RECT 1842.365 92.655 1842.695 92.670 ;
      LAYER via3 ;
        RECT 313.100 2765.740 313.420 2766.060 ;
        RECT 310.340 2731.740 310.660 2732.060 ;
        RECT 313.100 2731.740 313.420 2732.060 ;
        RECT 310.340 2476.740 310.660 2477.060 ;
        RECT 313.100 2476.740 313.420 2477.060 ;
        RECT 310.340 2446.820 310.660 2447.140 ;
        RECT 311.260 2445.460 311.580 2445.780 ;
        RECT 311.260 2414.180 311.580 2414.500 ;
        RECT 313.100 2367.260 313.420 2367.580 ;
        RECT 313.100 2318.980 313.420 2319.300 ;
        RECT 313.100 2316.940 313.420 2317.260 ;
        RECT 313.100 2272.740 313.420 2273.060 ;
        RECT 313.100 2270.020 313.420 2270.340 ;
        RECT 313.100 2259.820 313.420 2260.140 ;
        RECT 313.100 2224.460 313.420 2224.780 ;
        RECT 313.100 2129.940 313.420 2130.260 ;
        RECT 313.100 2109.540 313.420 2109.860 ;
        RECT 313.100 2044.940 313.420 2045.260 ;
        RECT 313.100 1980.340 313.420 1980.660 ;
        RECT 313.100 1946.340 313.420 1946.660 ;
        RECT 313.100 1895.340 313.420 1895.660 ;
        RECT 313.100 1840.940 313.420 1841.260 ;
        RECT 313.100 1835.500 313.420 1835.820 ;
        RECT 313.100 1811.020 313.420 1811.340 ;
        RECT 312.180 1732.140 312.500 1732.460 ;
        RECT 312.180 1683.180 312.500 1683.500 ;
        RECT 313.100 1611.100 313.420 1611.420 ;
        RECT 313.100 1497.540 313.420 1497.860 ;
        RECT 312.180 1490.740 312.500 1491.060 ;
        RECT 312.180 1483.260 312.500 1483.580 ;
        RECT 313.100 1446.540 313.420 1446.860 ;
        RECT 311.260 1434.980 311.580 1435.300 ;
        RECT 313.100 1434.980 313.420 1435.300 ;
        RECT 313.100 1256.140 313.420 1256.460 ;
        RECT 313.100 1255.460 313.420 1255.780 ;
        RECT 311.260 1216.700 311.580 1217.020 ;
        RECT 313.100 1216.700 313.420 1217.020 ;
        RECT 310.340 1111.980 310.660 1112.300 ;
        RECT 313.100 1110.620 313.420 1110.940 ;
        RECT 313.100 765.180 313.420 765.500 ;
        RECT 312.180 717.580 312.500 717.900 ;
        RECT 312.180 716.900 312.500 717.220 ;
        RECT 313.100 552.340 313.420 552.660 ;
        RECT 313.100 514.940 313.420 515.260 ;
        RECT 313.100 483.660 313.420 483.980 ;
        RECT 313.100 451.020 313.420 451.340 ;
        RECT 313.100 408.860 313.420 409.180 ;
        RECT 313.100 370.100 313.420 370.420 ;
        RECT 313.100 338.140 313.420 338.460 ;
        RECT 312.180 265.380 312.500 265.700 ;
        RECT 316.780 257.220 317.100 257.540 ;
        RECT 314.020 217.100 314.340 217.420 ;
        RECT 316.780 217.100 317.100 217.420 ;
        RECT 314.020 158.620 314.340 158.940 ;
        RECT 316.780 158.620 317.100 158.940 ;
        RECT 314.940 92.660 315.260 92.980 ;
      LAYER met4 ;
        RECT 313.095 2766.050 313.425 2766.065 ;
        RECT 313.095 2765.750 314.330 2766.050 ;
        RECT 313.095 2765.735 313.425 2765.750 ;
        RECT 310.335 2731.735 310.665 2732.065 ;
        RECT 313.095 2732.050 313.425 2732.065 ;
        RECT 314.030 2732.050 314.330 2765.750 ;
        RECT 313.095 2731.750 314.330 2732.050 ;
        RECT 313.095 2731.735 313.425 2731.750 ;
        RECT 310.350 2647.490 310.650 2731.735 ;
        RECT 309.910 2646.310 311.090 2647.490 ;
        RECT 315.430 2646.310 316.610 2647.490 ;
        RECT 315.870 2582.450 316.170 2646.310 ;
        RECT 314.030 2582.150 316.170 2582.450 ;
        RECT 314.030 2572.250 314.330 2582.150 ;
        RECT 314.030 2571.950 316.170 2572.250 ;
        RECT 315.870 2531.450 316.170 2571.950 ;
        RECT 315.870 2531.150 317.090 2531.450 ;
        RECT 310.335 2476.735 310.665 2477.065 ;
        RECT 313.095 2477.050 313.425 2477.065 ;
        RECT 316.790 2477.050 317.090 2531.150 ;
        RECT 313.095 2476.750 317.090 2477.050 ;
        RECT 313.095 2476.735 313.425 2476.750 ;
        RECT 310.350 2447.145 310.650 2476.735 ;
        RECT 310.335 2446.815 310.665 2447.145 ;
        RECT 311.255 2445.455 311.585 2445.785 ;
        RECT 311.270 2414.505 311.570 2445.455 ;
        RECT 311.255 2414.175 311.585 2414.505 ;
        RECT 313.095 2367.255 313.425 2367.585 ;
        RECT 313.110 2319.305 313.410 2367.255 ;
        RECT 313.095 2318.975 313.425 2319.305 ;
        RECT 313.095 2317.250 313.425 2317.265 ;
        RECT 313.095 2316.950 314.330 2317.250 ;
        RECT 313.095 2316.935 313.425 2316.950 ;
        RECT 313.095 2273.050 313.425 2273.065 ;
        RECT 314.030 2273.050 314.330 2316.950 ;
        RECT 313.095 2272.750 314.330 2273.050 ;
        RECT 313.095 2272.735 313.425 2272.750 ;
        RECT 313.095 2270.015 313.425 2270.345 ;
        RECT 313.110 2260.145 313.410 2270.015 ;
        RECT 313.095 2259.815 313.425 2260.145 ;
        RECT 313.095 2224.455 313.425 2224.785 ;
        RECT 313.110 2208.450 313.410 2224.455 ;
        RECT 313.110 2208.150 316.170 2208.450 ;
        RECT 315.870 2147.250 316.170 2208.150 ;
        RECT 314.030 2146.950 316.170 2147.250 ;
        RECT 313.095 2130.250 313.425 2130.265 ;
        RECT 314.030 2130.250 314.330 2146.950 ;
        RECT 313.095 2129.950 314.330 2130.250 ;
        RECT 313.095 2129.935 313.425 2129.950 ;
        RECT 313.095 2109.850 313.425 2109.865 ;
        RECT 313.095 2109.550 314.330 2109.850 ;
        RECT 313.095 2109.535 313.425 2109.550 ;
        RECT 313.095 2045.250 313.425 2045.265 ;
        RECT 314.030 2045.250 314.330 2109.550 ;
        RECT 313.095 2044.950 314.330 2045.250 ;
        RECT 313.095 2044.935 313.425 2044.950 ;
        RECT 313.095 1980.650 313.425 1980.665 ;
        RECT 313.095 1980.350 314.330 1980.650 ;
        RECT 313.095 1980.335 313.425 1980.350 ;
        RECT 313.095 1946.650 313.425 1946.665 ;
        RECT 314.030 1946.650 314.330 1980.350 ;
        RECT 313.095 1946.350 314.330 1946.650 ;
        RECT 313.095 1946.335 313.425 1946.350 ;
        RECT 313.095 1895.650 313.425 1895.665 ;
        RECT 313.095 1895.350 316.170 1895.650 ;
        RECT 313.095 1895.335 313.425 1895.350 ;
        RECT 313.095 1841.250 313.425 1841.265 ;
        RECT 315.870 1841.250 316.170 1895.350 ;
        RECT 313.095 1840.950 316.170 1841.250 ;
        RECT 313.095 1840.935 313.425 1840.950 ;
        RECT 313.095 1835.495 313.425 1835.825 ;
        RECT 313.110 1811.345 313.410 1835.495 ;
        RECT 313.095 1811.015 313.425 1811.345 ;
        RECT 312.175 1732.135 312.505 1732.465 ;
        RECT 312.190 1683.505 312.490 1732.135 ;
        RECT 312.175 1683.175 312.505 1683.505 ;
        RECT 313.095 1611.095 313.425 1611.425 ;
        RECT 313.110 1497.865 313.410 1611.095 ;
        RECT 313.095 1497.535 313.425 1497.865 ;
        RECT 312.175 1490.735 312.505 1491.065 ;
        RECT 312.190 1483.585 312.490 1490.735 ;
        RECT 312.175 1483.255 312.505 1483.585 ;
        RECT 313.095 1446.535 313.425 1446.865 ;
        RECT 313.110 1435.305 313.410 1446.535 ;
        RECT 311.255 1434.975 311.585 1435.305 ;
        RECT 313.095 1434.975 313.425 1435.305 ;
        RECT 311.270 1402.650 311.570 1434.975 ;
        RECT 311.270 1402.350 314.330 1402.650 ;
        RECT 314.030 1310.850 314.330 1402.350 ;
        RECT 313.110 1310.550 314.330 1310.850 ;
        RECT 313.110 1256.465 313.410 1310.550 ;
        RECT 313.095 1256.135 313.425 1256.465 ;
        RECT 313.095 1255.455 313.425 1255.785 ;
        RECT 313.110 1217.025 313.410 1255.455 ;
        RECT 311.255 1216.695 311.585 1217.025 ;
        RECT 313.095 1216.695 313.425 1217.025 ;
        RECT 311.270 1178.250 311.570 1216.695 ;
        RECT 310.350 1177.950 311.570 1178.250 ;
        RECT 310.350 1112.305 310.650 1177.950 ;
        RECT 310.335 1111.975 310.665 1112.305 ;
        RECT 313.095 1110.615 313.425 1110.945 ;
        RECT 313.110 1089.850 313.410 1110.615 ;
        RECT 312.190 1089.550 313.410 1089.850 ;
        RECT 312.190 1035.450 312.490 1089.550 ;
        RECT 312.190 1035.150 316.170 1035.450 ;
        RECT 315.870 801.290 316.170 1035.150 ;
        RECT 311.750 800.110 312.930 801.290 ;
        RECT 315.430 800.110 316.610 801.290 ;
        RECT 312.190 797.450 312.490 800.110 ;
        RECT 312.190 797.150 313.180 797.450 ;
        RECT 312.880 796.770 313.180 797.150 ;
        RECT 312.880 796.470 313.410 796.770 ;
        RECT 313.110 765.505 313.410 796.470 ;
        RECT 313.095 765.175 313.425 765.505 ;
        RECT 312.175 717.575 312.505 717.905 ;
        RECT 312.190 717.225 312.490 717.575 ;
        RECT 312.175 716.895 312.505 717.225 ;
        RECT 313.095 552.650 313.425 552.665 ;
        RECT 313.095 552.350 314.330 552.650 ;
        RECT 313.095 552.335 313.425 552.350 ;
        RECT 313.095 515.250 313.425 515.265 ;
        RECT 314.030 515.250 314.330 552.350 ;
        RECT 313.095 514.950 314.330 515.250 ;
        RECT 313.095 514.935 313.425 514.950 ;
        RECT 313.095 483.655 313.425 483.985 ;
        RECT 313.110 451.345 313.410 483.655 ;
        RECT 313.095 451.015 313.425 451.345 ;
        RECT 313.095 408.855 313.425 409.185 ;
        RECT 313.110 406.450 313.410 408.855 ;
        RECT 313.110 406.150 314.330 406.450 ;
        RECT 314.030 379.250 314.330 406.150 ;
        RECT 313.110 378.950 314.330 379.250 ;
        RECT 313.110 370.425 313.410 378.950 ;
        RECT 313.095 370.095 313.425 370.425 ;
        RECT 313.095 338.135 313.425 338.465 ;
        RECT 313.110 304.450 313.410 338.135 ;
        RECT 312.190 304.150 313.410 304.450 ;
        RECT 312.190 265.705 312.490 304.150 ;
        RECT 312.175 265.375 312.505 265.705 ;
        RECT 316.775 257.215 317.105 257.545 ;
        RECT 316.790 217.425 317.090 257.215 ;
        RECT 314.015 217.095 314.345 217.425 ;
        RECT 316.775 217.095 317.105 217.425 ;
        RECT 314.030 158.945 314.330 217.095 ;
        RECT 314.015 158.615 314.345 158.945 ;
        RECT 316.775 158.615 317.105 158.945 ;
        RECT 316.790 134.450 317.090 158.615 ;
        RECT 314.950 134.150 317.090 134.450 ;
        RECT 314.950 92.985 315.250 134.150 ;
        RECT 314.935 92.655 315.265 92.985 ;
      LAYER met5 ;
        RECT 309.700 2646.100 316.820 2647.700 ;
        RECT 311.540 799.900 316.820 801.500 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1863.145 48.365 1863.315 96.475 ;
      LAYER mcon ;
        RECT 1863.145 96.305 1863.315 96.475 ;
      LAYER met1 ;
        RECT 1863.070 96.460 1863.390 96.520 ;
        RECT 1862.875 96.320 1863.390 96.460 ;
        RECT 1863.070 96.260 1863.390 96.320 ;
        RECT 1863.085 48.520 1863.375 48.565 ;
        RECT 1863.990 48.520 1864.310 48.580 ;
        RECT 1863.085 48.380 1864.310 48.520 ;
        RECT 1863.085 48.335 1863.375 48.380 ;
        RECT 1863.990 48.320 1864.310 48.380 ;
      LAYER via ;
        RECT 1863.100 96.260 1863.360 96.520 ;
        RECT 1864.020 48.320 1864.280 48.580 ;
      LAYER met2 ;
        RECT 1863.090 183.075 1863.370 183.445 ;
        RECT 1863.160 96.550 1863.300 183.075 ;
        RECT 1863.100 96.230 1863.360 96.550 ;
        RECT 1864.020 48.290 1864.280 48.610 ;
        RECT 1864.080 2.400 1864.220 48.290 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
      LAYER via2 ;
        RECT 1863.090 183.120 1863.370 183.400 ;
      LAYER met3 ;
        RECT 298.350 2271.690 298.730 2271.700 ;
        RECT 310.000 2271.690 314.000 2272.080 ;
        RECT 298.350 2271.480 314.000 2271.690 ;
        RECT 298.350 2271.390 310.500 2271.480 ;
        RECT 298.350 2271.380 298.730 2271.390 ;
        RECT 298.350 183.410 298.730 183.420 ;
        RECT 1863.065 183.410 1863.395 183.425 ;
        RECT 298.350 183.110 1863.395 183.410 ;
        RECT 298.350 183.100 298.730 183.110 ;
        RECT 1863.065 183.095 1863.395 183.110 ;
      LAYER via3 ;
        RECT 298.380 2271.380 298.700 2271.700 ;
        RECT 298.380 183.100 298.700 183.420 ;
      LAYER met4 ;
        RECT 298.375 2271.375 298.705 2271.705 ;
        RECT 298.390 183.425 298.690 2271.375 ;
        RECT 298.375 183.095 298.705 183.425 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 740.210 20.640 740.530 20.700 ;
        RECT 744.810 20.640 745.130 20.700 ;
        RECT 740.210 20.500 745.130 20.640 ;
        RECT 740.210 20.440 740.530 20.500 ;
        RECT 744.810 20.440 745.130 20.500 ;
      LAYER via ;
        RECT 740.240 20.440 740.500 20.700 ;
        RECT 744.840 20.440 745.100 20.700 ;
      LAYER met2 ;
        RECT 744.830 237.475 745.110 237.845 ;
        RECT 744.900 20.730 745.040 237.475 ;
        RECT 740.240 20.410 740.500 20.730 ;
        RECT 744.840 20.410 745.100 20.730 ;
        RECT 740.300 2.400 740.440 20.410 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 744.830 237.520 745.110 237.800 ;
      LAYER met3 ;
        RECT 2606.000 3212.600 2610.000 3213.200 ;
        RECT 2609.430 3210.090 2609.730 3212.600 ;
        RECT 2609.430 3209.790 2610.650 3210.090 ;
        RECT 2610.350 3208.730 2610.650 3209.790 ;
        RECT 2671.950 3208.730 2672.330 3208.740 ;
        RECT 2610.350 3208.430 2672.330 3208.730 ;
        RECT 2671.950 3208.420 2672.330 3208.430 ;
        RECT 744.805 237.810 745.135 237.825 ;
        RECT 2671.950 237.810 2672.330 237.820 ;
        RECT 744.805 237.510 2672.330 237.810 ;
        RECT 744.805 237.495 745.135 237.510 ;
        RECT 2671.950 237.500 2672.330 237.510 ;
      LAYER via3 ;
        RECT 2671.980 3208.420 2672.300 3208.740 ;
        RECT 2671.980 237.500 2672.300 237.820 ;
      LAYER met4 ;
        RECT 2671.975 3208.415 2672.305 3208.745 ;
        RECT 2671.990 237.825 2672.290 3208.415 ;
        RECT 2671.975 237.495 2672.305 237.825 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.910 3278.860 1635.230 3278.920 ;
        RECT 2663.470 3278.860 2663.790 3278.920 ;
        RECT 1634.910 3278.720 2663.790 3278.860 ;
        RECT 1634.910 3278.660 1635.230 3278.720 ;
        RECT 2663.470 3278.660 2663.790 3278.720 ;
        RECT 1881.930 34.240 1882.250 34.300 ;
        RECT 2663.470 34.240 2663.790 34.300 ;
        RECT 1881.930 34.100 2663.790 34.240 ;
        RECT 1881.930 34.040 1882.250 34.100 ;
        RECT 2663.470 34.040 2663.790 34.100 ;
      LAYER via ;
        RECT 1634.940 3278.660 1635.200 3278.920 ;
        RECT 2663.500 3278.660 2663.760 3278.920 ;
        RECT 1881.960 34.040 1882.220 34.300 ;
        RECT 2663.500 34.040 2663.760 34.300 ;
      LAYER met2 ;
        RECT 1634.940 3278.630 1635.200 3278.950 ;
        RECT 2663.500 3278.630 2663.760 3278.950 ;
        RECT 1635.000 3260.000 1635.140 3278.630 ;
        RECT 1634.890 3256.000 1635.170 3260.000 ;
        RECT 2663.560 34.330 2663.700 3278.630 ;
        RECT 1881.960 34.010 1882.220 34.330 ;
        RECT 2663.500 34.010 2663.760 34.330 ;
        RECT 1882.020 2.400 1882.160 34.010 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1899.870 25.060 1900.190 25.120 ;
        RECT 2339.170 25.060 2339.490 25.120 ;
        RECT 1899.870 24.920 2339.490 25.060 ;
        RECT 1899.870 24.860 1900.190 24.920 ;
        RECT 2339.170 24.860 2339.490 24.920 ;
      LAYER via ;
        RECT 1899.900 24.860 1900.160 25.120 ;
        RECT 2339.200 24.860 2339.460 25.120 ;
      LAYER met2 ;
        RECT 2343.290 260.170 2343.570 264.000 ;
        RECT 2339.260 260.030 2343.570 260.170 ;
        RECT 2339.260 25.150 2339.400 260.030 ;
        RECT 2343.290 260.000 2343.570 260.030 ;
        RECT 1899.900 24.830 1900.160 25.150 ;
        RECT 2339.200 24.830 2339.460 25.150 ;
        RECT 1899.960 2.400 1900.100 24.830 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 306.430 141.680 306.750 141.740 ;
        RECT 1911.370 141.680 1911.690 141.740 ;
        RECT 306.430 141.540 1911.690 141.680 ;
        RECT 306.430 141.480 306.750 141.540 ;
        RECT 1911.370 141.480 1911.690 141.540 ;
        RECT 1911.370 37.640 1911.690 37.700 ;
        RECT 1917.810 37.640 1918.130 37.700 ;
        RECT 1911.370 37.500 1918.130 37.640 ;
        RECT 1911.370 37.440 1911.690 37.500 ;
        RECT 1917.810 37.440 1918.130 37.500 ;
      LAYER via ;
        RECT 306.460 141.480 306.720 141.740 ;
        RECT 1911.400 141.480 1911.660 141.740 ;
        RECT 1911.400 37.440 1911.660 37.700 ;
        RECT 1917.840 37.440 1918.100 37.700 ;
      LAYER met2 ;
        RECT 306.450 1467.595 306.730 1467.965 ;
        RECT 306.520 141.770 306.660 1467.595 ;
        RECT 306.460 141.450 306.720 141.770 ;
        RECT 1911.400 141.450 1911.660 141.770 ;
        RECT 1911.460 37.730 1911.600 141.450 ;
        RECT 1911.400 37.410 1911.660 37.730 ;
        RECT 1917.840 37.410 1918.100 37.730 ;
        RECT 1917.900 2.400 1918.040 37.410 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
      LAYER via2 ;
        RECT 306.450 1467.640 306.730 1467.920 ;
      LAYER met3 ;
        RECT 306.425 1467.930 306.755 1467.945 ;
        RECT 310.000 1467.930 314.000 1468.320 ;
        RECT 306.425 1467.720 314.000 1467.930 ;
        RECT 306.425 1467.630 310.500 1467.720 ;
        RECT 306.425 1467.615 306.755 1467.630 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.490 203.900 311.810 203.960 ;
        RECT 1932.070 203.900 1932.390 203.960 ;
        RECT 311.490 203.760 1932.390 203.900 ;
        RECT 311.490 203.700 311.810 203.760 ;
        RECT 1932.070 203.700 1932.390 203.760 ;
        RECT 1932.070 62.260 1932.390 62.520 ;
        RECT 1932.160 61.780 1932.300 62.260 ;
        RECT 1935.290 61.780 1935.610 61.840 ;
        RECT 1932.160 61.640 1935.610 61.780 ;
        RECT 1935.290 61.580 1935.610 61.640 ;
      LAYER via ;
        RECT 311.520 203.700 311.780 203.960 ;
        RECT 1932.100 203.700 1932.360 203.960 ;
        RECT 1932.100 62.260 1932.360 62.520 ;
        RECT 1935.320 61.580 1935.580 61.840 ;
      LAYER met2 ;
        RECT 311.050 3035.675 311.330 3036.045 ;
        RECT 311.120 3008.165 311.260 3035.675 ;
        RECT 311.050 3007.795 311.330 3008.165 ;
        RECT 312.890 2667.795 313.170 2668.165 ;
        RECT 312.960 2649.805 313.100 2667.795 ;
        RECT 312.890 2649.435 313.170 2649.805 ;
        RECT 311.510 2600.475 311.790 2600.845 ;
        RECT 311.580 2553.245 311.720 2600.475 ;
        RECT 311.510 2552.875 311.790 2553.245 ;
        RECT 311.970 2365.875 312.250 2366.245 ;
        RECT 312.040 2318.645 312.180 2365.875 ;
        RECT 311.970 2318.275 312.250 2318.645 ;
        RECT 311.510 1978.955 311.790 1979.325 ;
        RECT 311.580 1932.405 311.720 1978.955 ;
        RECT 311.510 1932.035 311.790 1932.405 ;
        RECT 311.510 1834.795 311.790 1835.165 ;
        RECT 311.580 1739.285 311.720 1834.795 ;
        RECT 311.510 1738.915 311.790 1739.285 ;
        RECT 311.050 1690.635 311.330 1691.005 ;
        RECT 311.120 1684.885 311.260 1690.635 ;
        RECT 311.050 1684.515 311.330 1684.885 ;
        RECT 311.050 1683.155 311.330 1683.525 ;
        RECT 311.120 1640.685 311.260 1683.155 ;
        RECT 311.050 1640.315 311.330 1640.685 ;
        RECT 311.510 1555.995 311.790 1556.365 ;
        RECT 311.580 1491.085 311.720 1555.995 ;
        RECT 311.510 1490.715 311.790 1491.085 ;
        RECT 311.050 1483.235 311.330 1483.605 ;
        RECT 311.120 1436.685 311.260 1483.235 ;
        RECT 311.050 1436.315 311.330 1436.685 ;
        RECT 310.130 1434.955 310.410 1435.325 ;
        RECT 310.200 1380.245 310.340 1434.955 ;
        RECT 310.130 1379.875 310.410 1380.245 ;
        RECT 311.510 1355.395 311.790 1355.765 ;
        RECT 311.580 1307.485 311.720 1355.395 ;
        RECT 311.510 1307.115 311.790 1307.485 ;
        RECT 310.590 1282.635 310.870 1283.005 ;
        RECT 310.660 1153.125 310.800 1282.635 ;
        RECT 310.590 1152.755 310.870 1153.125 ;
        RECT 311.510 1054.155 311.790 1054.525 ;
        RECT 311.580 1007.605 311.720 1054.155 ;
        RECT 311.510 1007.235 311.790 1007.605 ;
        RECT 311.050 820.235 311.330 820.605 ;
        RECT 311.120 796.805 311.260 820.235 ;
        RECT 311.050 796.435 311.330 796.805 ;
        RECT 310.590 716.875 310.870 717.245 ;
        RECT 310.660 669.645 310.800 716.875 ;
        RECT 310.590 669.275 310.870 669.645 ;
        RECT 311.510 268.755 311.790 269.125 ;
        RECT 311.580 203.990 311.720 268.755 ;
        RECT 311.520 203.670 311.780 203.990 ;
        RECT 1932.100 203.670 1932.360 203.990 ;
        RECT 1932.160 62.550 1932.300 203.670 ;
        RECT 1932.100 62.230 1932.360 62.550 ;
        RECT 1935.320 61.550 1935.580 61.870 ;
        RECT 1935.380 2.400 1935.520 61.550 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
      LAYER via2 ;
        RECT 311.050 3035.720 311.330 3036.000 ;
        RECT 311.050 3007.840 311.330 3008.120 ;
        RECT 312.890 2667.840 313.170 2668.120 ;
        RECT 312.890 2649.480 313.170 2649.760 ;
        RECT 311.510 2600.520 311.790 2600.800 ;
        RECT 311.510 2552.920 311.790 2553.200 ;
        RECT 311.970 2365.920 312.250 2366.200 ;
        RECT 311.970 2318.320 312.250 2318.600 ;
        RECT 311.510 1979.000 311.790 1979.280 ;
        RECT 311.510 1932.080 311.790 1932.360 ;
        RECT 311.510 1834.840 311.790 1835.120 ;
        RECT 311.510 1738.960 311.790 1739.240 ;
        RECT 311.050 1690.680 311.330 1690.960 ;
        RECT 311.050 1684.560 311.330 1684.840 ;
        RECT 311.050 1683.200 311.330 1683.480 ;
        RECT 311.050 1640.360 311.330 1640.640 ;
        RECT 311.510 1556.040 311.790 1556.320 ;
        RECT 311.510 1490.760 311.790 1491.040 ;
        RECT 311.050 1483.280 311.330 1483.560 ;
        RECT 311.050 1436.360 311.330 1436.640 ;
        RECT 310.130 1435.000 310.410 1435.280 ;
        RECT 310.130 1379.920 310.410 1380.200 ;
        RECT 311.510 1355.440 311.790 1355.720 ;
        RECT 311.510 1307.160 311.790 1307.440 ;
        RECT 310.590 1282.680 310.870 1282.960 ;
        RECT 310.590 1152.800 310.870 1153.080 ;
        RECT 311.510 1054.200 311.790 1054.480 ;
        RECT 311.510 1007.280 311.790 1007.560 ;
        RECT 311.050 820.280 311.330 820.560 ;
        RECT 311.050 796.480 311.330 796.760 ;
        RECT 310.590 716.920 310.870 717.200 ;
        RECT 310.590 669.320 310.870 669.600 ;
        RECT 311.510 268.800 311.790 269.080 ;
      LAYER met3 ;
        RECT 310.000 3201.720 314.000 3202.320 ;
        RECT 310.310 3201.250 310.690 3201.260 ;
        RECT 312.190 3201.250 312.490 3201.720 ;
        RECT 310.310 3200.950 312.490 3201.250 ;
        RECT 310.310 3200.940 310.690 3200.950 ;
        RECT 310.310 3154.020 310.690 3154.340 ;
        RECT 310.350 3152.970 310.650 3154.020 ;
        RECT 311.230 3152.970 311.610 3152.980 ;
        RECT 310.350 3152.670 311.610 3152.970 ;
        RECT 311.230 3152.660 311.610 3152.670 ;
        RECT 313.070 3057.770 313.450 3057.780 ;
        RECT 312.190 3057.470 313.450 3057.770 ;
        RECT 312.190 3056.420 312.490 3057.470 ;
        RECT 313.070 3057.460 313.450 3057.470 ;
        RECT 312.150 3056.100 312.530 3056.420 ;
        RECT 311.025 3036.010 311.355 3036.025 ;
        RECT 312.150 3036.010 312.530 3036.020 ;
        RECT 311.025 3035.710 312.530 3036.010 ;
        RECT 311.025 3035.695 311.355 3035.710 ;
        RECT 312.150 3035.700 312.530 3035.710 ;
        RECT 310.310 3008.130 310.690 3008.140 ;
        RECT 311.025 3008.130 311.355 3008.145 ;
        RECT 310.310 3007.830 311.355 3008.130 ;
        RECT 310.310 3007.820 310.690 3007.830 ;
        RECT 311.025 3007.815 311.355 3007.830 ;
        RECT 311.230 2718.820 311.610 2719.140 ;
        RECT 311.270 2717.770 311.570 2718.820 ;
        RECT 312.150 2717.770 312.530 2717.780 ;
        RECT 311.270 2717.470 312.530 2717.770 ;
        RECT 312.150 2717.460 312.530 2717.470 ;
        RECT 312.150 2668.130 312.530 2668.140 ;
        RECT 312.865 2668.130 313.195 2668.145 ;
        RECT 312.150 2667.830 313.195 2668.130 ;
        RECT 312.150 2667.820 312.530 2667.830 ;
        RECT 312.865 2667.815 313.195 2667.830 ;
        RECT 312.865 2649.780 313.195 2649.785 ;
        RECT 312.865 2649.770 313.450 2649.780 ;
        RECT 312.640 2649.470 313.450 2649.770 ;
        RECT 312.865 2649.460 313.450 2649.470 ;
        RECT 312.865 2649.455 313.195 2649.460 ;
        RECT 312.150 2601.490 312.530 2601.500 ;
        RECT 313.070 2601.490 313.450 2601.500 ;
        RECT 312.150 2601.190 313.450 2601.490 ;
        RECT 312.150 2601.180 312.530 2601.190 ;
        RECT 313.070 2601.180 313.450 2601.190 ;
        RECT 311.485 2600.810 311.815 2600.825 ;
        RECT 312.150 2600.810 312.530 2600.820 ;
        RECT 311.485 2600.510 312.530 2600.810 ;
        RECT 311.485 2600.495 311.815 2600.510 ;
        RECT 312.150 2600.500 312.530 2600.510 ;
        RECT 311.485 2553.220 311.815 2553.225 ;
        RECT 311.230 2553.210 311.815 2553.220 ;
        RECT 311.030 2552.910 311.815 2553.210 ;
        RECT 311.230 2552.900 311.815 2552.910 ;
        RECT 311.485 2552.895 311.815 2552.900 ;
        RECT 311.230 2511.730 311.610 2511.740 ;
        RECT 312.150 2511.730 312.530 2511.740 ;
        RECT 311.230 2511.430 312.530 2511.730 ;
        RECT 311.230 2511.420 311.610 2511.430 ;
        RECT 312.150 2511.420 312.530 2511.430 ;
        RECT 309.390 2390.690 309.770 2390.700 ;
        RECT 312.150 2390.690 312.530 2390.700 ;
        RECT 309.390 2390.390 312.530 2390.690 ;
        RECT 309.390 2390.380 309.770 2390.390 ;
        RECT 312.150 2390.380 312.530 2390.390 ;
        RECT 311.945 2366.220 312.275 2366.225 ;
        RECT 311.945 2366.210 312.530 2366.220 ;
        RECT 311.720 2365.910 312.530 2366.210 ;
        RECT 311.945 2365.900 312.530 2365.910 ;
        RECT 311.945 2365.895 312.275 2365.900 ;
        RECT 309.390 2318.610 309.770 2318.620 ;
        RECT 311.945 2318.610 312.275 2318.625 ;
        RECT 309.390 2318.310 312.275 2318.610 ;
        RECT 309.390 2318.300 309.770 2318.310 ;
        RECT 311.945 2318.295 312.275 2318.310 ;
        RECT 312.150 2029.610 312.530 2029.620 ;
        RECT 310.350 2029.310 312.530 2029.610 ;
        RECT 310.350 2028.940 310.650 2029.310 ;
        RECT 312.150 2029.300 312.530 2029.310 ;
        RECT 310.310 2028.620 310.690 2028.940 ;
        RECT 309.390 1980.650 309.770 1980.660 ;
        RECT 309.390 1980.350 311.570 1980.650 ;
        RECT 309.390 1980.340 309.770 1980.350 ;
        RECT 311.270 1979.305 311.570 1980.350 ;
        RECT 311.270 1978.990 311.815 1979.305 ;
        RECT 311.485 1978.975 311.815 1978.990 ;
        RECT 311.485 1932.380 311.815 1932.385 ;
        RECT 311.230 1932.370 311.815 1932.380 ;
        RECT 311.230 1932.070 312.040 1932.370 ;
        RECT 311.230 1932.060 311.815 1932.070 ;
        RECT 311.485 1932.055 311.815 1932.060 ;
        RECT 310.310 1884.090 310.690 1884.100 ;
        RECT 310.310 1883.790 312.490 1884.090 ;
        RECT 310.310 1883.780 310.690 1883.790 ;
        RECT 311.230 1882.050 311.610 1882.060 ;
        RECT 312.190 1882.050 312.490 1883.790 ;
        RECT 311.230 1881.750 312.490 1882.050 ;
        RECT 311.230 1881.740 311.610 1881.750 ;
        RECT 311.485 1835.130 311.815 1835.145 ;
        RECT 312.150 1835.130 312.530 1835.140 ;
        RECT 311.485 1834.830 312.530 1835.130 ;
        RECT 311.485 1834.815 311.815 1834.830 ;
        RECT 312.150 1834.820 312.530 1834.830 ;
        RECT 311.485 1739.260 311.815 1739.265 ;
        RECT 311.230 1739.250 311.815 1739.260 ;
        RECT 311.230 1738.950 312.040 1739.250 ;
        RECT 311.230 1738.940 311.815 1738.950 ;
        RECT 311.485 1738.935 311.815 1738.940 ;
        RECT 311.025 1690.980 311.355 1690.985 ;
        RECT 311.025 1690.970 311.610 1690.980 ;
        RECT 310.800 1690.670 311.610 1690.970 ;
        RECT 311.025 1690.660 311.610 1690.670 ;
        RECT 311.025 1690.655 311.355 1690.660 ;
        RECT 311.025 1684.860 311.355 1684.865 ;
        RECT 311.025 1684.850 311.610 1684.860 ;
        RECT 311.025 1684.550 311.810 1684.850 ;
        RECT 311.025 1684.540 311.610 1684.550 ;
        RECT 311.025 1684.535 311.355 1684.540 ;
        RECT 311.025 1683.500 311.355 1683.505 ;
        RECT 311.025 1683.490 311.610 1683.500 ;
        RECT 310.800 1683.190 311.610 1683.490 ;
        RECT 311.025 1683.180 311.610 1683.190 ;
        RECT 311.025 1683.175 311.355 1683.180 ;
        RECT 310.310 1640.650 310.690 1640.660 ;
        RECT 311.025 1640.650 311.355 1640.665 ;
        RECT 310.310 1640.350 311.355 1640.650 ;
        RECT 310.310 1640.340 310.690 1640.350 ;
        RECT 311.025 1640.335 311.355 1640.350 ;
        RECT 310.310 1594.100 310.690 1594.420 ;
        RECT 310.350 1593.050 310.650 1594.100 ;
        RECT 311.230 1593.050 311.610 1593.060 ;
        RECT 310.350 1592.750 311.610 1593.050 ;
        RECT 311.230 1592.740 311.610 1592.750 ;
        RECT 311.485 1556.340 311.815 1556.345 ;
        RECT 311.230 1556.330 311.815 1556.340 ;
        RECT 311.030 1556.030 311.815 1556.330 ;
        RECT 311.230 1556.020 311.815 1556.030 ;
        RECT 311.485 1556.015 311.815 1556.020 ;
        RECT 311.485 1491.060 311.815 1491.065 ;
        RECT 311.230 1491.050 311.815 1491.060 ;
        RECT 311.030 1490.750 311.815 1491.050 ;
        RECT 311.230 1490.740 311.815 1490.750 ;
        RECT 311.485 1490.735 311.815 1490.740 ;
        RECT 311.025 1483.580 311.355 1483.585 ;
        RECT 311.025 1483.570 311.610 1483.580 ;
        RECT 310.800 1483.270 311.610 1483.570 ;
        RECT 311.025 1483.260 311.610 1483.270 ;
        RECT 311.025 1483.255 311.355 1483.260 ;
        RECT 311.025 1436.650 311.355 1436.665 ;
        RECT 309.430 1436.350 311.355 1436.650 ;
        RECT 309.430 1435.980 309.730 1436.350 ;
        RECT 311.025 1436.335 311.355 1436.350 ;
        RECT 309.390 1435.660 309.770 1435.980 ;
        RECT 309.390 1435.290 309.770 1435.300 ;
        RECT 310.105 1435.290 310.435 1435.305 ;
        RECT 309.390 1434.990 310.435 1435.290 ;
        RECT 309.390 1434.980 309.770 1434.990 ;
        RECT 310.105 1434.975 310.435 1434.990 ;
        RECT 310.105 1380.210 310.435 1380.225 ;
        RECT 311.230 1380.210 311.610 1380.220 ;
        RECT 310.105 1379.910 311.610 1380.210 ;
        RECT 310.105 1379.895 310.435 1379.910 ;
        RECT 311.230 1379.900 311.610 1379.910 ;
        RECT 311.485 1355.740 311.815 1355.745 ;
        RECT 311.230 1355.730 311.815 1355.740 ;
        RECT 311.030 1355.430 311.815 1355.730 ;
        RECT 311.230 1355.420 311.815 1355.430 ;
        RECT 311.485 1355.415 311.815 1355.420 ;
        RECT 311.485 1307.460 311.815 1307.465 ;
        RECT 311.230 1307.450 311.815 1307.460 ;
        RECT 311.030 1307.150 311.815 1307.450 ;
        RECT 311.230 1307.140 311.815 1307.150 ;
        RECT 311.485 1307.135 311.815 1307.140 ;
        RECT 310.565 1282.970 310.895 1282.985 ;
        RECT 311.230 1282.970 311.610 1282.980 ;
        RECT 310.565 1282.670 311.610 1282.970 ;
        RECT 310.565 1282.655 310.895 1282.670 ;
        RECT 311.230 1282.660 311.610 1282.670 ;
        RECT 310.565 1153.090 310.895 1153.105 ;
        RECT 311.230 1153.090 311.610 1153.100 ;
        RECT 310.565 1152.790 311.610 1153.090 ;
        RECT 310.565 1152.775 310.895 1152.790 ;
        RECT 311.230 1152.780 311.610 1152.790 ;
        RECT 311.230 1111.300 311.610 1111.620 ;
        RECT 311.270 1110.250 311.570 1111.300 ;
        RECT 312.150 1110.250 312.530 1110.260 ;
        RECT 311.270 1109.950 312.530 1110.250 ;
        RECT 312.150 1109.940 312.530 1109.950 ;
        RECT 311.230 1054.860 311.610 1055.180 ;
        RECT 311.270 1054.505 311.570 1054.860 ;
        RECT 311.270 1054.190 311.815 1054.505 ;
        RECT 311.485 1054.175 311.815 1054.190 ;
        RECT 311.485 1007.570 311.815 1007.585 ;
        RECT 312.150 1007.570 312.530 1007.580 ;
        RECT 311.485 1007.270 312.530 1007.570 ;
        RECT 311.485 1007.255 311.815 1007.270 ;
        RECT 312.150 1007.260 312.530 1007.270 ;
        RECT 312.150 1006.580 312.530 1006.900 ;
        RECT 311.230 1006.210 311.610 1006.220 ;
        RECT 312.190 1006.210 312.490 1006.580 ;
        RECT 311.230 1005.910 312.490 1006.210 ;
        RECT 311.230 1005.900 311.610 1005.910 ;
        RECT 311.230 917.500 311.610 917.820 ;
        RECT 311.270 917.130 311.570 917.500 ;
        RECT 312.150 917.130 312.530 917.140 ;
        RECT 311.270 916.830 312.530 917.130 ;
        RECT 312.150 916.820 312.530 916.830 ;
        RECT 312.150 821.250 312.530 821.260 ;
        RECT 311.270 820.950 312.530 821.250 ;
        RECT 311.270 820.585 311.570 820.950 ;
        RECT 312.150 820.940 312.530 820.950 ;
        RECT 311.025 820.270 311.570 820.585 ;
        RECT 311.025 820.255 311.355 820.270 ;
        RECT 310.310 796.770 310.690 796.780 ;
        RECT 311.025 796.770 311.355 796.785 ;
        RECT 310.310 796.470 311.355 796.770 ;
        RECT 310.310 796.460 310.690 796.470 ;
        RECT 311.025 796.455 311.355 796.470 ;
        RECT 310.310 726.050 310.690 726.060 ;
        RECT 310.310 725.750 311.570 726.050 ;
        RECT 310.310 725.740 310.690 725.750 ;
        RECT 311.270 724.870 311.570 725.750 ;
        RECT 311.230 724.550 311.610 724.870 ;
        RECT 310.565 717.210 310.895 717.225 ;
        RECT 311.230 717.210 311.610 717.220 ;
        RECT 310.565 716.910 311.610 717.210 ;
        RECT 310.565 716.895 310.895 716.910 ;
        RECT 311.230 716.900 311.610 716.910 ;
        RECT 309.390 669.610 309.770 669.620 ;
        RECT 310.565 669.610 310.895 669.625 ;
        RECT 309.390 669.310 310.895 669.610 ;
        RECT 309.390 669.300 309.770 669.310 ;
        RECT 310.565 669.295 310.895 669.310 ;
        RECT 309.390 628.130 309.770 628.140 ;
        RECT 311.230 628.130 311.610 628.140 ;
        RECT 309.390 627.830 311.610 628.130 ;
        RECT 309.390 627.820 309.770 627.830 ;
        RECT 311.230 627.820 311.610 627.830 ;
        RECT 311.230 580.220 311.610 580.540 ;
        RECT 311.270 579.180 311.570 580.220 ;
        RECT 311.230 578.860 311.610 579.180 ;
        RECT 310.310 383.330 310.690 383.340 ;
        RECT 313.070 383.330 313.450 383.340 ;
        RECT 310.310 383.030 313.450 383.330 ;
        RECT 310.310 383.020 310.690 383.030 ;
        RECT 313.070 383.020 313.450 383.030 ;
        RECT 310.310 269.090 310.690 269.100 ;
        RECT 311.485 269.090 311.815 269.105 ;
        RECT 310.310 268.790 311.815 269.090 ;
        RECT 310.310 268.780 310.690 268.790 ;
        RECT 311.485 268.775 311.815 268.790 ;
      LAYER via3 ;
        RECT 310.340 3200.940 310.660 3201.260 ;
        RECT 310.340 3154.020 310.660 3154.340 ;
        RECT 311.260 3152.660 311.580 3152.980 ;
        RECT 313.100 3057.460 313.420 3057.780 ;
        RECT 312.180 3056.100 312.500 3056.420 ;
        RECT 312.180 3035.700 312.500 3036.020 ;
        RECT 310.340 3007.820 310.660 3008.140 ;
        RECT 311.260 2718.820 311.580 2719.140 ;
        RECT 312.180 2717.460 312.500 2717.780 ;
        RECT 312.180 2667.820 312.500 2668.140 ;
        RECT 313.100 2649.460 313.420 2649.780 ;
        RECT 312.180 2601.180 312.500 2601.500 ;
        RECT 313.100 2601.180 313.420 2601.500 ;
        RECT 312.180 2600.500 312.500 2600.820 ;
        RECT 311.260 2552.900 311.580 2553.220 ;
        RECT 311.260 2511.420 311.580 2511.740 ;
        RECT 312.180 2511.420 312.500 2511.740 ;
        RECT 309.420 2390.380 309.740 2390.700 ;
        RECT 312.180 2390.380 312.500 2390.700 ;
        RECT 312.180 2365.900 312.500 2366.220 ;
        RECT 309.420 2318.300 309.740 2318.620 ;
        RECT 312.180 2029.300 312.500 2029.620 ;
        RECT 310.340 2028.620 310.660 2028.940 ;
        RECT 309.420 1980.340 309.740 1980.660 ;
        RECT 311.260 1932.060 311.580 1932.380 ;
        RECT 310.340 1883.780 310.660 1884.100 ;
        RECT 311.260 1881.740 311.580 1882.060 ;
        RECT 312.180 1834.820 312.500 1835.140 ;
        RECT 311.260 1738.940 311.580 1739.260 ;
        RECT 311.260 1690.660 311.580 1690.980 ;
        RECT 311.260 1684.540 311.580 1684.860 ;
        RECT 311.260 1683.180 311.580 1683.500 ;
        RECT 310.340 1640.340 310.660 1640.660 ;
        RECT 310.340 1594.100 310.660 1594.420 ;
        RECT 311.260 1592.740 311.580 1593.060 ;
        RECT 311.260 1556.020 311.580 1556.340 ;
        RECT 311.260 1490.740 311.580 1491.060 ;
        RECT 311.260 1483.260 311.580 1483.580 ;
        RECT 309.420 1435.660 309.740 1435.980 ;
        RECT 309.420 1434.980 309.740 1435.300 ;
        RECT 311.260 1379.900 311.580 1380.220 ;
        RECT 311.260 1355.420 311.580 1355.740 ;
        RECT 311.260 1307.140 311.580 1307.460 ;
        RECT 311.260 1282.660 311.580 1282.980 ;
        RECT 311.260 1152.780 311.580 1153.100 ;
        RECT 311.260 1111.300 311.580 1111.620 ;
        RECT 312.180 1109.940 312.500 1110.260 ;
        RECT 311.260 1054.860 311.580 1055.180 ;
        RECT 312.180 1007.260 312.500 1007.580 ;
        RECT 312.180 1006.580 312.500 1006.900 ;
        RECT 311.260 1005.900 311.580 1006.220 ;
        RECT 311.260 917.500 311.580 917.820 ;
        RECT 312.180 916.820 312.500 917.140 ;
        RECT 312.180 820.940 312.500 821.260 ;
        RECT 310.340 796.460 310.660 796.780 ;
        RECT 310.340 725.740 310.660 726.060 ;
        RECT 311.260 724.550 311.580 724.870 ;
        RECT 311.260 716.900 311.580 717.220 ;
        RECT 309.420 669.300 309.740 669.620 ;
        RECT 309.420 627.820 309.740 628.140 ;
        RECT 311.260 627.820 311.580 628.140 ;
        RECT 311.260 580.220 311.580 580.540 ;
        RECT 311.260 578.860 311.580 579.180 ;
        RECT 310.340 383.020 310.660 383.340 ;
        RECT 313.100 383.020 313.420 383.340 ;
        RECT 310.340 268.780 310.660 269.100 ;
      LAYER met4 ;
        RECT 310.335 3200.935 310.665 3201.265 ;
        RECT 310.350 3154.345 310.650 3200.935 ;
        RECT 310.335 3154.015 310.665 3154.345 ;
        RECT 311.255 3152.655 311.585 3152.985 ;
        RECT 311.270 3106.050 311.570 3152.655 ;
        RECT 311.270 3105.750 313.410 3106.050 ;
        RECT 313.110 3057.785 313.410 3105.750 ;
        RECT 313.095 3057.455 313.425 3057.785 ;
        RECT 312.175 3056.095 312.505 3056.425 ;
        RECT 312.190 3036.025 312.490 3056.095 ;
        RECT 312.175 3035.695 312.505 3036.025 ;
        RECT 310.335 3007.815 310.665 3008.145 ;
        RECT 310.350 2959.850 310.650 3007.815 ;
        RECT 310.350 2959.550 311.570 2959.850 ;
        RECT 311.270 2912.250 311.570 2959.550 ;
        RECT 311.270 2911.950 313.410 2912.250 ;
        RECT 313.110 2908.850 313.410 2911.950 ;
        RECT 313.110 2908.550 314.330 2908.850 ;
        RECT 314.030 2861.250 314.330 2908.550 ;
        RECT 314.030 2860.950 316.170 2861.250 ;
        RECT 315.870 2806.850 316.170 2860.950 ;
        RECT 315.870 2806.550 317.090 2806.850 ;
        RECT 316.790 2779.650 317.090 2806.550 ;
        RECT 311.270 2779.350 317.090 2779.650 ;
        RECT 311.270 2719.145 311.570 2779.350 ;
        RECT 311.255 2718.815 311.585 2719.145 ;
        RECT 312.175 2717.455 312.505 2717.785 ;
        RECT 312.190 2668.145 312.490 2717.455 ;
        RECT 312.175 2667.815 312.505 2668.145 ;
        RECT 313.095 2649.455 313.425 2649.785 ;
        RECT 313.110 2601.505 313.410 2649.455 ;
        RECT 312.175 2601.175 312.505 2601.505 ;
        RECT 313.095 2601.175 313.425 2601.505 ;
        RECT 312.190 2600.825 312.490 2601.175 ;
        RECT 312.175 2600.495 312.505 2600.825 ;
        RECT 311.255 2552.895 311.585 2553.225 ;
        RECT 311.270 2534.850 311.570 2552.895 ;
        RECT 311.270 2534.550 312.490 2534.850 ;
        RECT 312.190 2511.745 312.490 2534.550 ;
        RECT 311.255 2511.415 311.585 2511.745 ;
        RECT 312.175 2511.415 312.505 2511.745 ;
        RECT 311.270 2446.450 311.570 2511.415 ;
        RECT 309.430 2446.150 311.570 2446.450 ;
        RECT 309.430 2390.705 309.730 2446.150 ;
        RECT 309.415 2390.375 309.745 2390.705 ;
        RECT 312.175 2390.375 312.505 2390.705 ;
        RECT 312.190 2366.225 312.490 2390.375 ;
        RECT 312.175 2365.895 312.505 2366.225 ;
        RECT 309.415 2318.295 309.745 2318.625 ;
        RECT 309.430 2279.850 309.730 2318.295 ;
        RECT 309.430 2279.550 310.650 2279.850 ;
        RECT 310.350 2235.650 310.650 2279.550 ;
        RECT 310.350 2235.350 312.490 2235.650 ;
        RECT 312.190 2029.625 312.490 2235.350 ;
        RECT 312.175 2029.295 312.505 2029.625 ;
        RECT 310.335 2028.615 310.665 2028.945 ;
        RECT 310.350 2004.450 310.650 2028.615 ;
        RECT 309.430 2004.150 310.650 2004.450 ;
        RECT 309.430 1980.665 309.730 2004.150 ;
        RECT 309.415 1980.335 309.745 1980.665 ;
        RECT 311.255 1932.055 311.585 1932.385 ;
        RECT 311.270 1909.250 311.570 1932.055 ;
        RECT 310.350 1908.950 311.570 1909.250 ;
        RECT 310.350 1884.105 310.650 1908.950 ;
        RECT 310.335 1883.775 310.665 1884.105 ;
        RECT 311.255 1881.735 311.585 1882.065 ;
        RECT 311.270 1837.850 311.570 1881.735 ;
        RECT 311.270 1837.550 312.490 1837.850 ;
        RECT 312.190 1835.145 312.490 1837.550 ;
        RECT 312.175 1834.815 312.505 1835.145 ;
        RECT 311.255 1738.935 311.585 1739.265 ;
        RECT 311.270 1690.985 311.570 1738.935 ;
        RECT 311.255 1690.655 311.585 1690.985 ;
        RECT 311.255 1684.535 311.585 1684.865 ;
        RECT 311.270 1683.505 311.570 1684.535 ;
        RECT 311.255 1683.175 311.585 1683.505 ;
        RECT 310.335 1640.335 310.665 1640.665 ;
        RECT 310.350 1594.425 310.650 1640.335 ;
        RECT 310.335 1594.095 310.665 1594.425 ;
        RECT 311.255 1592.735 311.585 1593.065 ;
        RECT 311.270 1556.345 311.570 1592.735 ;
        RECT 311.255 1556.015 311.585 1556.345 ;
        RECT 311.255 1490.735 311.585 1491.065 ;
        RECT 311.270 1483.585 311.570 1490.735 ;
        RECT 311.255 1483.255 311.585 1483.585 ;
        RECT 309.415 1435.655 309.745 1435.985 ;
        RECT 309.430 1435.305 309.730 1435.655 ;
        RECT 309.415 1434.975 309.745 1435.305 ;
        RECT 311.255 1379.895 311.585 1380.225 ;
        RECT 311.270 1355.745 311.570 1379.895 ;
        RECT 311.255 1355.415 311.585 1355.745 ;
        RECT 311.255 1307.135 311.585 1307.465 ;
        RECT 311.270 1282.985 311.570 1307.135 ;
        RECT 311.255 1282.655 311.585 1282.985 ;
        RECT 311.255 1152.775 311.585 1153.105 ;
        RECT 311.270 1111.625 311.570 1152.775 ;
        RECT 311.255 1111.295 311.585 1111.625 ;
        RECT 312.175 1109.935 312.505 1110.265 ;
        RECT 312.190 1093.250 312.490 1109.935 ;
        RECT 311.270 1092.950 312.490 1093.250 ;
        RECT 311.270 1055.185 311.570 1092.950 ;
        RECT 311.255 1054.855 311.585 1055.185 ;
        RECT 312.175 1007.255 312.505 1007.585 ;
        RECT 312.190 1006.905 312.490 1007.255 ;
        RECT 312.175 1006.575 312.505 1006.905 ;
        RECT 311.255 1005.895 311.585 1006.225 ;
        RECT 311.270 917.825 311.570 1005.895 ;
        RECT 311.255 917.495 311.585 917.825 ;
        RECT 312.175 916.815 312.505 917.145 ;
        RECT 312.190 821.265 312.490 916.815 ;
        RECT 312.175 820.935 312.505 821.265 ;
        RECT 310.335 796.455 310.665 796.785 ;
        RECT 310.350 726.065 310.650 796.455 ;
        RECT 310.335 725.735 310.665 726.065 ;
        RECT 311.255 724.545 311.585 724.875 ;
        RECT 311.270 717.225 311.570 724.545 ;
        RECT 311.255 716.895 311.585 717.225 ;
        RECT 309.415 669.295 309.745 669.625 ;
        RECT 309.430 628.145 309.730 669.295 ;
        RECT 309.415 627.815 309.745 628.145 ;
        RECT 311.255 627.815 311.585 628.145 ;
        RECT 311.270 580.545 311.570 627.815 ;
        RECT 311.255 580.215 311.585 580.545 ;
        RECT 311.255 578.855 311.585 579.185 ;
        RECT 311.270 573.050 311.570 578.855 ;
        RECT 311.270 572.750 312.490 573.050 ;
        RECT 312.190 396.250 312.490 572.750 ;
        RECT 312.190 395.950 313.410 396.250 ;
        RECT 313.110 383.345 313.410 395.950 ;
        RECT 310.335 383.015 310.665 383.345 ;
        RECT 313.095 383.015 313.425 383.345 ;
        RECT 310.350 362.250 310.650 383.015 ;
        RECT 310.350 361.950 311.570 362.250 ;
        RECT 311.270 314.650 311.570 361.950 ;
        RECT 310.350 314.350 311.570 314.650 ;
        RECT 310.350 269.105 310.650 314.350 ;
        RECT 310.335 268.775 310.665 269.105 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.170 3258.970 574.450 3259.085 ;
        RECT 575.970 3258.970 576.250 3260.000 ;
        RECT 574.170 3258.830 576.250 3258.970 ;
        RECT 574.170 3258.715 574.450 3258.830 ;
        RECT 575.970 3256.000 576.250 3258.830 ;
        RECT 1012.090 33.730 1012.370 33.845 ;
        RECT 1013.930 33.730 1014.210 33.845 ;
        RECT 1012.090 33.590 1014.210 33.730 ;
        RECT 1012.090 33.475 1012.370 33.590 ;
        RECT 1013.930 33.475 1014.210 33.590 ;
        RECT 1953.250 33.475 1953.530 33.845 ;
        RECT 1953.320 2.400 1953.460 33.475 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
      LAYER via2 ;
        RECT 574.170 3258.760 574.450 3259.040 ;
        RECT 1012.090 33.520 1012.370 33.800 ;
        RECT 1013.930 33.520 1014.210 33.800 ;
        RECT 1953.250 33.520 1953.530 33.800 ;
      LAYER met3 ;
        RECT 267.070 3259.050 267.450 3259.060 ;
        RECT 574.145 3259.050 574.475 3259.065 ;
        RECT 267.070 3258.750 574.475 3259.050 ;
        RECT 267.070 3258.740 267.450 3258.750 ;
        RECT 574.145 3258.735 574.475 3258.750 ;
        RECT 1706.910 34.190 1731.130 34.490 ;
        RECT 267.070 33.810 267.450 33.820 ;
        RECT 1012.065 33.810 1012.395 33.825 ;
        RECT 267.070 33.510 1012.395 33.810 ;
        RECT 267.070 33.500 267.450 33.510 ;
        RECT 1012.065 33.495 1012.395 33.510 ;
        RECT 1013.905 33.810 1014.235 33.825 ;
        RECT 1706.910 33.810 1707.210 34.190 ;
        RECT 1013.905 33.510 1707.210 33.810 ;
        RECT 1730.830 33.810 1731.130 34.190 ;
        RECT 1953.225 33.810 1953.555 33.825 ;
        RECT 1730.830 33.510 1953.555 33.810 ;
        RECT 1013.905 33.495 1014.235 33.510 ;
        RECT 1953.225 33.495 1953.555 33.510 ;
      LAYER via3 ;
        RECT 267.100 3258.740 267.420 3259.060 ;
        RECT 267.100 33.500 267.420 33.820 ;
      LAYER met4 ;
        RECT 267.095 3258.735 267.425 3259.065 ;
        RECT 267.110 33.825 267.410 3258.735 ;
        RECT 267.095 33.495 267.425 33.825 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1284.390 244.020 1284.710 244.080 ;
        RECT 1289.910 244.020 1290.230 244.080 ;
        RECT 1284.390 243.880 1290.230 244.020 ;
        RECT 1284.390 243.820 1284.710 243.880 ;
        RECT 1289.910 243.820 1290.230 243.880 ;
        RECT 1289.910 25.740 1290.230 25.800 ;
        RECT 1971.170 25.740 1971.490 25.800 ;
        RECT 1289.910 25.600 1971.490 25.740 ;
        RECT 1289.910 25.540 1290.230 25.600 ;
        RECT 1971.170 25.540 1971.490 25.600 ;
      LAYER via ;
        RECT 1284.420 243.820 1284.680 244.080 ;
        RECT 1289.940 243.820 1290.200 244.080 ;
        RECT 1289.940 25.540 1290.200 25.800 ;
        RECT 1971.200 25.540 1971.460 25.800 ;
      LAYER met2 ;
        RECT 1284.370 260.000 1284.650 264.000 ;
        RECT 1284.480 244.110 1284.620 260.000 ;
        RECT 1284.420 243.790 1284.680 244.110 ;
        RECT 1289.940 243.790 1290.200 244.110 ;
        RECT 1290.000 25.830 1290.140 243.790 ;
        RECT 1289.940 25.510 1290.200 25.830 ;
        RECT 1971.200 25.510 1971.460 25.830 ;
        RECT 1971.260 2.400 1971.400 25.510 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1476.860 2615.490 1476.920 ;
        RECT 2705.790 1476.860 2706.110 1476.920 ;
        RECT 2615.170 1476.720 2706.110 1476.860 ;
        RECT 2615.170 1476.660 2615.490 1476.720 ;
        RECT 2705.790 1476.660 2706.110 1476.720 ;
        RECT 1993.710 217.500 1994.030 217.560 ;
        RECT 2705.790 217.500 2706.110 217.560 ;
        RECT 1993.710 217.360 2706.110 217.500 ;
        RECT 1993.710 217.300 1994.030 217.360 ;
        RECT 2705.790 217.300 2706.110 217.360 ;
        RECT 1989.110 16.900 1989.430 16.960 ;
        RECT 1993.710 16.900 1994.030 16.960 ;
        RECT 1989.110 16.760 1994.030 16.900 ;
        RECT 1989.110 16.700 1989.430 16.760 ;
        RECT 1993.710 16.700 1994.030 16.760 ;
      LAYER via ;
        RECT 2615.200 1476.660 2615.460 1476.920 ;
        RECT 2705.820 1476.660 2706.080 1476.920 ;
        RECT 1993.740 217.300 1994.000 217.560 ;
        RECT 2705.820 217.300 2706.080 217.560 ;
        RECT 1989.140 16.700 1989.400 16.960 ;
        RECT 1993.740 16.700 1994.000 16.960 ;
      LAYER met2 ;
        RECT 2615.190 1479.835 2615.470 1480.205 ;
        RECT 2615.260 1476.950 2615.400 1479.835 ;
        RECT 2615.200 1476.630 2615.460 1476.950 ;
        RECT 2705.820 1476.630 2706.080 1476.950 ;
        RECT 2705.880 217.590 2706.020 1476.630 ;
        RECT 1993.740 217.270 1994.000 217.590 ;
        RECT 2705.820 217.270 2706.080 217.590 ;
        RECT 1993.800 16.990 1993.940 217.270 ;
        RECT 1989.140 16.670 1989.400 16.990 ;
        RECT 1993.740 16.670 1994.000 16.990 ;
        RECT 1989.200 2.400 1989.340 16.670 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1479.880 2615.470 1480.160 ;
      LAYER met3 ;
        RECT 2606.000 1480.170 2610.000 1480.560 ;
        RECT 2615.165 1480.170 2615.495 1480.185 ;
        RECT 2606.000 1479.960 2615.495 1480.170 ;
        RECT 2609.580 1479.870 2615.495 1479.960 ;
        RECT 2615.165 1479.855 2615.495 1479.870 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2007.585 145.265 2007.755 163.115 ;
        RECT 2007.125 48.365 2007.295 137.955 ;
      LAYER mcon ;
        RECT 2007.585 162.945 2007.755 163.115 ;
        RECT 2007.125 137.785 2007.295 137.955 ;
      LAYER met1 ;
        RECT 2007.525 163.100 2007.815 163.145 ;
        RECT 2610.110 163.100 2610.430 163.160 ;
        RECT 2007.525 162.960 2610.430 163.100 ;
        RECT 2007.525 162.915 2007.815 162.960 ;
        RECT 2610.110 162.900 2610.430 162.960 ;
        RECT 2007.510 145.420 2007.830 145.480 ;
        RECT 2007.315 145.280 2007.830 145.420 ;
        RECT 2007.510 145.220 2007.830 145.280 ;
        RECT 2007.065 137.940 2007.355 137.985 ;
        RECT 2007.510 137.940 2007.830 138.000 ;
        RECT 2007.065 137.800 2007.830 137.940 ;
        RECT 2007.065 137.755 2007.355 137.800 ;
        RECT 2007.510 137.740 2007.830 137.800 ;
        RECT 2007.050 48.520 2007.370 48.580 ;
        RECT 2006.855 48.380 2007.370 48.520 ;
        RECT 2007.050 48.320 2007.370 48.380 ;
      LAYER via ;
        RECT 2610.140 162.900 2610.400 163.160 ;
        RECT 2007.540 145.220 2007.800 145.480 ;
        RECT 2007.540 137.740 2007.800 138.000 ;
        RECT 2007.080 48.320 2007.340 48.580 ;
      LAYER met2 ;
        RECT 2610.130 821.595 2610.410 821.965 ;
        RECT 2610.200 163.190 2610.340 821.595 ;
        RECT 2610.140 162.870 2610.400 163.190 ;
        RECT 2007.540 145.190 2007.800 145.510 ;
        RECT 2007.600 138.030 2007.740 145.190 ;
        RECT 2007.540 137.710 2007.800 138.030 ;
        RECT 2007.080 48.290 2007.340 48.610 ;
        RECT 2007.140 23.530 2007.280 48.290 ;
        RECT 2006.680 23.390 2007.280 23.530 ;
        RECT 2006.680 2.400 2006.820 23.390 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
      LAYER via2 ;
        RECT 2610.130 821.640 2610.410 821.920 ;
      LAYER met3 ;
        RECT 2606.000 824.440 2610.000 825.040 ;
        RECT 2609.430 821.930 2609.730 824.440 ;
        RECT 2610.105 821.930 2610.435 821.945 ;
        RECT 2609.430 821.630 2610.435 821.930 ;
        RECT 2610.105 821.615 2610.435 821.630 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2021.845 144.925 2022.015 193.035 ;
        RECT 2021.845 48.365 2022.015 96.475 ;
      LAYER mcon ;
        RECT 2021.845 192.865 2022.015 193.035 ;
        RECT 2021.845 96.305 2022.015 96.475 ;
      LAYER met1 ;
        RECT 298.150 196.760 298.470 196.820 ;
        RECT 2021.770 196.760 2022.090 196.820 ;
        RECT 298.150 196.620 2022.090 196.760 ;
        RECT 298.150 196.560 298.470 196.620 ;
        RECT 2021.770 196.560 2022.090 196.620 ;
        RECT 2021.770 193.020 2022.090 193.080 ;
        RECT 2021.575 192.880 2022.090 193.020 ;
        RECT 2021.770 192.820 2022.090 192.880 ;
        RECT 2021.770 145.080 2022.090 145.140 ;
        RECT 2021.575 144.940 2022.090 145.080 ;
        RECT 2021.770 144.880 2022.090 144.940 ;
        RECT 2021.770 96.460 2022.090 96.520 ;
        RECT 2021.575 96.320 2022.090 96.460 ;
        RECT 2021.770 96.260 2022.090 96.320 ;
        RECT 2021.770 48.520 2022.090 48.580 ;
        RECT 2021.575 48.380 2022.090 48.520 ;
        RECT 2021.770 48.320 2022.090 48.380 ;
        RECT 2021.770 14.180 2022.090 14.240 ;
        RECT 2021.770 14.040 2024.760 14.180 ;
        RECT 2021.770 13.980 2022.090 14.040 ;
        RECT 2024.620 13.900 2024.760 14.040 ;
        RECT 2024.530 13.640 2024.850 13.900 ;
      LAYER via ;
        RECT 298.180 196.560 298.440 196.820 ;
        RECT 2021.800 196.560 2022.060 196.820 ;
        RECT 2021.800 192.820 2022.060 193.080 ;
        RECT 2021.800 144.880 2022.060 145.140 ;
        RECT 2021.800 96.260 2022.060 96.520 ;
        RECT 2021.800 48.320 2022.060 48.580 ;
        RECT 2021.800 13.980 2022.060 14.240 ;
        RECT 2024.560 13.640 2024.820 13.900 ;
      LAYER met2 ;
        RECT 298.170 1066.395 298.450 1066.765 ;
        RECT 298.240 196.850 298.380 1066.395 ;
        RECT 298.180 196.530 298.440 196.850 ;
        RECT 2021.800 196.530 2022.060 196.850 ;
        RECT 2021.860 193.110 2022.000 196.530 ;
        RECT 2021.800 192.790 2022.060 193.110 ;
        RECT 2021.800 144.850 2022.060 145.170 ;
        RECT 2021.860 96.550 2022.000 144.850 ;
        RECT 2021.800 96.230 2022.060 96.550 ;
        RECT 2021.800 48.290 2022.060 48.610 ;
        RECT 2021.860 14.270 2022.000 48.290 ;
        RECT 2021.800 13.950 2022.060 14.270 ;
        RECT 2024.560 13.610 2024.820 13.930 ;
        RECT 2024.620 2.400 2024.760 13.610 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
      LAYER via2 ;
        RECT 298.170 1066.440 298.450 1066.720 ;
      LAYER met3 ;
        RECT 298.145 1066.730 298.475 1066.745 ;
        RECT 310.000 1066.730 314.000 1067.120 ;
        RECT 298.145 1066.520 314.000 1066.730 ;
        RECT 298.145 1066.430 310.500 1066.520 ;
        RECT 298.145 1066.415 298.475 1066.430 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.930 24.380 2043.250 24.440 ;
        RECT 2553.070 24.380 2553.390 24.440 ;
        RECT 2042.930 24.240 2553.390 24.380 ;
        RECT 2042.930 24.180 2043.250 24.240 ;
        RECT 2553.070 24.180 2553.390 24.240 ;
      LAYER via ;
        RECT 2042.960 24.180 2043.220 24.440 ;
        RECT 2553.100 24.180 2553.360 24.440 ;
      LAYER met2 ;
        RECT 2557.650 260.170 2557.930 264.000 ;
        RECT 2553.160 260.030 2557.930 260.170 ;
        RECT 2553.160 24.470 2553.300 260.030 ;
        RECT 2557.650 260.000 2557.930 260.030 ;
        RECT 2042.960 24.150 2043.220 24.470 ;
        RECT 2553.100 24.150 2553.360 24.470 ;
        RECT 2043.020 12.650 2043.160 24.150 ;
        RECT 2042.560 12.510 2043.160 12.650 ;
        RECT 2042.560 2.400 2042.700 12.510 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.610 14.180 758.930 14.240 ;
        RECT 757.780 14.040 758.930 14.180 ;
        RECT 757.780 13.900 757.920 14.040 ;
        RECT 758.610 13.980 758.930 14.040 ;
        RECT 757.690 13.640 758.010 13.900 ;
      LAYER via ;
        RECT 758.640 13.980 758.900 14.240 ;
        RECT 757.720 13.640 757.980 13.900 ;
      LAYER met2 ;
        RECT 758.630 113.035 758.910 113.405 ;
        RECT 758.700 14.270 758.840 113.035 ;
        RECT 758.640 13.950 758.900 14.270 ;
        RECT 757.720 13.610 757.980 13.930 ;
        RECT 757.780 2.400 757.920 13.610 ;
        RECT 757.570 -4.800 758.130 2.400 ;
      LAYER via2 ;
        RECT 758.630 113.080 758.910 113.360 ;
      LAYER met3 ;
        RECT 2606.000 2177.850 2610.000 2178.240 ;
        RECT 2625.030 2177.850 2625.410 2177.860 ;
        RECT 2606.000 2177.640 2625.410 2177.850 ;
        RECT 2609.580 2177.550 2625.410 2177.640 ;
        RECT 2625.030 2177.540 2625.410 2177.550 ;
        RECT 758.605 113.370 758.935 113.385 ;
        RECT 2625.030 113.370 2625.410 113.380 ;
        RECT 758.605 113.070 2625.410 113.370 ;
        RECT 758.605 113.055 758.935 113.070 ;
        RECT 2625.030 113.060 2625.410 113.070 ;
      LAYER via3 ;
        RECT 2625.060 2177.540 2625.380 2177.860 ;
        RECT 2625.060 113.060 2625.380 113.380 ;
      LAYER met4 ;
        RECT 2625.055 2177.535 2625.385 2177.865 ;
        RECT 2625.070 113.385 2625.370 2177.535 ;
        RECT 2625.055 113.055 2625.385 113.385 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2259.665 24.565 2259.835 25.755 ;
      LAYER mcon ;
        RECT 2259.665 25.585 2259.835 25.755 ;
      LAYER met1 ;
        RECT 2259.605 25.740 2259.895 25.785 ;
        RECT 2311.570 25.740 2311.890 25.800 ;
        RECT 2259.605 25.600 2311.890 25.740 ;
        RECT 2259.605 25.555 2259.895 25.600 ;
        RECT 2311.570 25.540 2311.890 25.600 ;
        RECT 2060.410 24.720 2060.730 24.780 ;
        RECT 2259.605 24.720 2259.895 24.765 ;
        RECT 2060.410 24.580 2259.895 24.720 ;
        RECT 2060.410 24.520 2060.730 24.580 ;
        RECT 2259.605 24.535 2259.895 24.580 ;
      LAYER via ;
        RECT 2311.600 25.540 2311.860 25.800 ;
        RECT 2060.440 24.520 2060.700 24.780 ;
      LAYER met2 ;
        RECT 2314.770 260.170 2315.050 264.000 ;
        RECT 2311.660 260.030 2315.050 260.170 ;
        RECT 2311.660 25.830 2311.800 260.030 ;
        RECT 2314.770 260.000 2315.050 260.030 ;
        RECT 2311.600 25.510 2311.860 25.830 ;
        RECT 2060.440 24.490 2060.700 24.810 ;
        RECT 2060.500 2.400 2060.640 24.490 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2083.410 260.000 2083.730 260.060 ;
        RECT 2612.870 260.000 2613.190 260.060 ;
        RECT 2083.410 259.860 2613.190 260.000 ;
        RECT 2083.410 259.800 2083.730 259.860 ;
        RECT 2612.870 259.800 2613.190 259.860 ;
        RECT 2078.350 16.900 2078.670 16.960 ;
        RECT 2083.410 16.900 2083.730 16.960 ;
        RECT 2078.350 16.760 2083.730 16.900 ;
        RECT 2078.350 16.700 2078.670 16.760 ;
        RECT 2083.410 16.700 2083.730 16.760 ;
      LAYER via ;
        RECT 2083.440 259.800 2083.700 260.060 ;
        RECT 2612.900 259.800 2613.160 260.060 ;
        RECT 2078.380 16.700 2078.640 16.960 ;
        RECT 2083.440 16.700 2083.700 16.960 ;
      LAYER met2 ;
        RECT 2612.890 507.435 2613.170 507.805 ;
        RECT 2612.960 260.090 2613.100 507.435 ;
        RECT 2083.440 259.770 2083.700 260.090 ;
        RECT 2612.900 259.770 2613.160 260.090 ;
        RECT 2083.500 16.990 2083.640 259.770 ;
        RECT 2078.380 16.670 2078.640 16.990 ;
        RECT 2083.440 16.670 2083.700 16.990 ;
        RECT 2078.440 2.400 2078.580 16.670 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
      LAYER via2 ;
        RECT 2612.890 507.480 2613.170 507.760 ;
      LAYER met3 ;
        RECT 2606.000 507.770 2610.000 508.160 ;
        RECT 2612.865 507.770 2613.195 507.785 ;
        RECT 2606.000 507.560 2613.195 507.770 ;
        RECT 2609.580 507.470 2613.195 507.560 ;
        RECT 2612.865 507.455 2613.195 507.470 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2097.230 168.795 2097.510 169.165 ;
        RECT 2097.300 14.690 2097.440 168.795 ;
        RECT 2096.380 14.550 2097.440 14.690 ;
        RECT 2096.380 13.330 2096.520 14.550 ;
        RECT 2095.920 13.190 2096.520 13.330 ;
        RECT 2095.920 2.400 2096.060 13.190 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
      LAYER via2 ;
        RECT 2097.230 168.840 2097.510 169.120 ;
      LAYER met3 ;
        RECT 2606.000 3043.960 2610.000 3044.560 ;
        RECT 2609.430 3043.500 2609.730 3043.960 ;
        RECT 2609.390 3043.180 2609.770 3043.500 ;
        RECT 2097.205 169.130 2097.535 169.145 ;
        RECT 2609.390 169.130 2609.770 169.140 ;
        RECT 2097.205 168.830 2609.770 169.130 ;
        RECT 2097.205 168.815 2097.535 168.830 ;
        RECT 2609.390 168.820 2609.770 168.830 ;
      LAYER via3 ;
        RECT 2609.420 3043.180 2609.740 3043.500 ;
        RECT 2609.420 168.820 2609.740 169.140 ;
      LAYER met4 ;
        RECT 2609.415 3043.175 2609.745 3043.505 ;
        RECT 2609.430 169.145 2609.730 3043.175 ;
        RECT 2609.415 168.815 2609.745 169.145 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2113.770 30.160 2114.090 30.220 ;
        RECT 2693.830 30.160 2694.150 30.220 ;
        RECT 2113.770 30.020 2694.150 30.160 ;
        RECT 2113.770 29.960 2114.090 30.020 ;
        RECT 2693.830 29.960 2694.150 30.020 ;
      LAYER via ;
        RECT 2113.800 29.960 2114.060 30.220 ;
        RECT 2693.860 29.960 2694.120 30.220 ;
      LAYER met2 ;
        RECT 1233.810 3273.675 1234.090 3274.045 ;
        RECT 1233.880 3260.000 1234.020 3273.675 ;
        RECT 1233.770 3256.000 1234.050 3260.000 ;
        RECT 2606.910 3253.275 2607.190 3253.645 ;
        RECT 2606.980 3248.885 2607.120 3253.275 ;
        RECT 2606.910 3248.515 2607.190 3248.885 ;
        RECT 2606.910 3165.555 2607.190 3165.925 ;
        RECT 2606.980 3119.685 2607.120 3165.555 ;
        RECT 2606.910 3119.315 2607.190 3119.685 ;
        RECT 2606.910 3115.915 2607.190 3116.285 ;
        RECT 2606.980 3072.085 2607.120 3115.915 ;
        RECT 2606.910 3071.715 2607.190 3072.085 ;
        RECT 2606.910 2986.715 2607.190 2987.085 ;
        RECT 2606.980 2942.885 2607.120 2986.715 ;
        RECT 2606.910 2942.515 2607.190 2942.885 ;
        RECT 2607.370 2490.315 2607.650 2490.685 ;
        RECT 2607.440 2443.085 2607.580 2490.315 ;
        RECT 2607.370 2442.715 2607.650 2443.085 ;
        RECT 2606.910 2362.475 2607.190 2362.845 ;
        RECT 2606.980 2328.845 2607.120 2362.475 ;
        RECT 2606.910 2328.475 2607.190 2328.845 ;
        RECT 2606.910 2232.595 2607.190 2232.965 ;
        RECT 2606.980 2174.485 2607.120 2232.595 ;
        RECT 2606.910 2174.115 2607.190 2174.485 ;
        RECT 2607.830 1868.115 2608.110 1868.485 ;
        RECT 2607.900 1857.605 2608.040 1868.115 ;
        RECT 2607.830 1857.235 2608.110 1857.605 ;
        RECT 2693.850 1610.395 2694.130 1610.765 ;
        RECT 2693.920 30.250 2694.060 1610.395 ;
        RECT 2113.800 29.930 2114.060 30.250 ;
        RECT 2693.860 29.930 2694.120 30.250 ;
        RECT 2113.860 2.400 2114.000 29.930 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
      LAYER via2 ;
        RECT 1233.810 3273.720 1234.090 3274.000 ;
        RECT 2606.910 3253.320 2607.190 3253.600 ;
        RECT 2606.910 3248.560 2607.190 3248.840 ;
        RECT 2606.910 3165.600 2607.190 3165.880 ;
        RECT 2606.910 3119.360 2607.190 3119.640 ;
        RECT 2606.910 3115.960 2607.190 3116.240 ;
        RECT 2606.910 3071.760 2607.190 3072.040 ;
        RECT 2606.910 2986.760 2607.190 2987.040 ;
        RECT 2606.910 2942.560 2607.190 2942.840 ;
        RECT 2607.370 2490.360 2607.650 2490.640 ;
        RECT 2607.370 2442.760 2607.650 2443.040 ;
        RECT 2606.910 2362.520 2607.190 2362.800 ;
        RECT 2606.910 2328.520 2607.190 2328.800 ;
        RECT 2606.910 2232.640 2607.190 2232.920 ;
        RECT 2606.910 2174.160 2607.190 2174.440 ;
        RECT 2607.830 1868.160 2608.110 1868.440 ;
        RECT 2607.830 1857.280 2608.110 1857.560 ;
        RECT 2693.850 1610.440 2694.130 1610.720 ;
      LAYER met3 ;
        RECT 1233.785 3274.010 1234.115 3274.025 ;
        RECT 2605.710 3274.010 2606.090 3274.020 ;
        RECT 1233.785 3273.710 2606.090 3274.010 ;
        RECT 1233.785 3273.695 1234.115 3273.710 ;
        RECT 2605.710 3273.700 2606.090 3273.710 ;
        RECT 2605.710 3253.610 2606.090 3253.620 ;
        RECT 2606.885 3253.610 2607.215 3253.625 ;
        RECT 2605.710 3253.310 2607.215 3253.610 ;
        RECT 2605.710 3253.300 2606.090 3253.310 ;
        RECT 2606.885 3253.295 2607.215 3253.310 ;
        RECT 2604.790 3248.850 2605.170 3248.860 ;
        RECT 2606.885 3248.850 2607.215 3248.865 ;
        RECT 2604.790 3248.550 2607.215 3248.850 ;
        RECT 2604.790 3248.540 2605.170 3248.550 ;
        RECT 2606.885 3248.535 2607.215 3248.550 ;
        RECT 2606.630 3166.260 2607.010 3166.580 ;
        RECT 2606.670 3165.905 2606.970 3166.260 ;
        RECT 2606.670 3165.590 2607.215 3165.905 ;
        RECT 2606.885 3165.575 2607.215 3165.590 ;
        RECT 2606.885 3119.660 2607.215 3119.665 ;
        RECT 2606.630 3119.650 2607.215 3119.660 ;
        RECT 2606.430 3119.350 2607.215 3119.650 ;
        RECT 2606.630 3119.340 2607.215 3119.350 ;
        RECT 2606.885 3119.335 2607.215 3119.340 ;
        RECT 2606.885 3116.260 2607.215 3116.265 ;
        RECT 2606.630 3116.250 2607.215 3116.260 ;
        RECT 2606.430 3115.950 2607.215 3116.250 ;
        RECT 2606.630 3115.940 2607.215 3115.950 ;
        RECT 2606.885 3115.935 2607.215 3115.940 ;
        RECT 2606.885 3072.060 2607.215 3072.065 ;
        RECT 2606.630 3072.050 2607.215 3072.060 ;
        RECT 2606.630 3071.750 2607.440 3072.050 ;
        RECT 2606.630 3071.740 2607.215 3071.750 ;
        RECT 2606.885 3071.735 2607.215 3071.740 ;
        RECT 2606.885 2987.060 2607.215 2987.065 ;
        RECT 2606.630 2987.050 2607.215 2987.060 ;
        RECT 2606.630 2986.750 2607.440 2987.050 ;
        RECT 2606.630 2986.740 2607.215 2986.750 ;
        RECT 2606.885 2986.735 2607.215 2986.740 ;
        RECT 2606.885 2942.860 2607.215 2942.865 ;
        RECT 2606.630 2942.850 2607.215 2942.860 ;
        RECT 2606.430 2942.550 2607.215 2942.850 ;
        RECT 2606.630 2942.540 2607.215 2942.550 ;
        RECT 2606.885 2942.535 2607.215 2942.540 ;
        RECT 2606.630 2863.660 2607.010 2863.980 ;
        RECT 2606.670 2862.620 2606.970 2863.660 ;
        RECT 2606.630 2862.300 2607.010 2862.620 ;
        RECT 2606.630 2517.850 2607.010 2517.860 ;
        RECT 2607.550 2517.850 2607.930 2517.860 ;
        RECT 2606.630 2517.550 2607.930 2517.850 ;
        RECT 2606.630 2517.540 2607.010 2517.550 ;
        RECT 2607.550 2517.540 2607.930 2517.550 ;
        RECT 2606.630 2490.650 2607.010 2490.660 ;
        RECT 2607.345 2490.650 2607.675 2490.665 ;
        RECT 2606.630 2490.350 2607.675 2490.650 ;
        RECT 2606.630 2490.340 2607.010 2490.350 ;
        RECT 2607.345 2490.335 2607.675 2490.350 ;
        RECT 2606.630 2443.050 2607.010 2443.060 ;
        RECT 2607.345 2443.050 2607.675 2443.065 ;
        RECT 2606.630 2442.750 2607.675 2443.050 ;
        RECT 2606.630 2442.740 2607.010 2442.750 ;
        RECT 2607.345 2442.735 2607.675 2442.750 ;
        RECT 2606.885 2362.820 2607.215 2362.825 ;
        RECT 2606.630 2362.810 2607.215 2362.820 ;
        RECT 2606.430 2362.510 2607.215 2362.810 ;
        RECT 2606.630 2362.500 2607.215 2362.510 ;
        RECT 2606.885 2362.495 2607.215 2362.500 ;
        RECT 2606.885 2328.820 2607.215 2328.825 ;
        RECT 2606.630 2328.810 2607.215 2328.820 ;
        RECT 2606.630 2328.510 2607.440 2328.810 ;
        RECT 2606.630 2328.500 2607.215 2328.510 ;
        RECT 2606.885 2328.495 2607.215 2328.500 ;
        RECT 2606.885 2232.940 2607.215 2232.945 ;
        RECT 2606.630 2232.930 2607.215 2232.940 ;
        RECT 2606.430 2232.630 2607.215 2232.930 ;
        RECT 2606.630 2232.620 2607.215 2232.630 ;
        RECT 2606.885 2232.615 2607.215 2232.620 ;
        RECT 2606.885 2174.460 2607.215 2174.465 ;
        RECT 2606.630 2174.450 2607.215 2174.460 ;
        RECT 2606.430 2174.150 2607.215 2174.450 ;
        RECT 2606.630 2174.140 2607.215 2174.150 ;
        RECT 2606.885 2174.135 2607.215 2174.140 ;
        RECT 2606.630 1868.450 2607.010 1868.460 ;
        RECT 2607.805 1868.450 2608.135 1868.465 ;
        RECT 2606.630 1868.150 2608.135 1868.450 ;
        RECT 2606.630 1868.140 2607.010 1868.150 ;
        RECT 2607.805 1868.135 2608.135 1868.150 ;
        RECT 2606.630 1857.570 2607.010 1857.580 ;
        RECT 2607.805 1857.570 2608.135 1857.585 ;
        RECT 2606.630 1857.270 2608.135 1857.570 ;
        RECT 2606.630 1857.260 2607.010 1857.270 ;
        RECT 2607.805 1857.255 2608.135 1857.270 ;
        RECT 2606.630 1610.730 2607.010 1610.740 ;
        RECT 2693.825 1610.730 2694.155 1610.745 ;
        RECT 2606.630 1610.430 2694.155 1610.730 ;
        RECT 2606.630 1610.420 2607.010 1610.430 ;
        RECT 2693.825 1610.415 2694.155 1610.430 ;
      LAYER via3 ;
        RECT 2605.740 3273.700 2606.060 3274.020 ;
        RECT 2605.740 3253.300 2606.060 3253.620 ;
        RECT 2604.820 3248.540 2605.140 3248.860 ;
        RECT 2606.660 3166.260 2606.980 3166.580 ;
        RECT 2606.660 3119.340 2606.980 3119.660 ;
        RECT 2606.660 3115.940 2606.980 3116.260 ;
        RECT 2606.660 3071.740 2606.980 3072.060 ;
        RECT 2606.660 2986.740 2606.980 2987.060 ;
        RECT 2606.660 2942.540 2606.980 2942.860 ;
        RECT 2606.660 2863.660 2606.980 2863.980 ;
        RECT 2606.660 2862.300 2606.980 2862.620 ;
        RECT 2606.660 2517.540 2606.980 2517.860 ;
        RECT 2607.580 2517.540 2607.900 2517.860 ;
        RECT 2606.660 2490.340 2606.980 2490.660 ;
        RECT 2606.660 2442.740 2606.980 2443.060 ;
        RECT 2606.660 2362.500 2606.980 2362.820 ;
        RECT 2606.660 2328.500 2606.980 2328.820 ;
        RECT 2606.660 2232.620 2606.980 2232.940 ;
        RECT 2606.660 2174.140 2606.980 2174.460 ;
        RECT 2606.660 1868.140 2606.980 1868.460 ;
        RECT 2606.660 1857.260 2606.980 1857.580 ;
        RECT 2606.660 1610.420 2606.980 1610.740 ;
      LAYER met4 ;
        RECT 2605.735 3273.695 2606.065 3274.025 ;
        RECT 2605.750 3253.625 2606.050 3273.695 ;
        RECT 2605.735 3253.295 2606.065 3253.625 ;
        RECT 2604.815 3248.535 2605.145 3248.865 ;
        RECT 2604.830 3214.850 2605.130 3248.535 ;
        RECT 2604.830 3214.550 2606.050 3214.850 ;
        RECT 2605.750 3211.450 2606.050 3214.550 ;
        RECT 2605.750 3211.150 2606.970 3211.450 ;
        RECT 2606.670 3166.585 2606.970 3211.150 ;
        RECT 2606.655 3166.255 2606.985 3166.585 ;
        RECT 2606.655 3119.650 2606.985 3119.665 ;
        RECT 2604.830 3119.350 2606.985 3119.650 ;
        RECT 2604.830 3116.250 2605.130 3119.350 ;
        RECT 2606.655 3119.335 2606.985 3119.350 ;
        RECT 2606.655 3116.250 2606.985 3116.265 ;
        RECT 2604.830 3115.950 2606.985 3116.250 ;
        RECT 2606.655 3115.935 2606.985 3115.950 ;
        RECT 2606.655 3072.050 2606.985 3072.065 ;
        RECT 2605.750 3071.750 2606.985 3072.050 ;
        RECT 2605.750 3061.850 2606.050 3071.750 ;
        RECT 2606.655 3071.735 2606.985 3071.750 ;
        RECT 2604.830 3061.550 2606.050 3061.850 ;
        RECT 2604.830 3014.250 2605.130 3061.550 ;
        RECT 2604.830 3013.950 2606.050 3014.250 ;
        RECT 2605.750 2987.050 2606.050 3013.950 ;
        RECT 2606.655 2987.050 2606.985 2987.065 ;
        RECT 2605.750 2986.750 2606.985 2987.050 ;
        RECT 2606.655 2986.735 2606.985 2986.750 ;
        RECT 2606.655 2942.850 2606.985 2942.865 ;
        RECT 2604.830 2942.550 2606.985 2942.850 ;
        RECT 2604.830 2891.850 2605.130 2942.550 ;
        RECT 2606.655 2942.535 2606.985 2942.550 ;
        RECT 2604.830 2891.550 2606.050 2891.850 ;
        RECT 2605.750 2871.450 2606.050 2891.550 ;
        RECT 2605.750 2871.150 2606.970 2871.450 ;
        RECT 2606.670 2863.985 2606.970 2871.150 ;
        RECT 2606.655 2863.655 2606.985 2863.985 ;
        RECT 2606.655 2862.295 2606.985 2862.625 ;
        RECT 2606.670 2817.050 2606.970 2862.295 ;
        RECT 2604.830 2816.750 2606.970 2817.050 ;
        RECT 2604.830 2762.650 2605.130 2816.750 ;
        RECT 2603.910 2762.350 2605.130 2762.650 ;
        RECT 2603.910 2681.050 2604.210 2762.350 ;
        RECT 2603.910 2680.750 2605.130 2681.050 ;
        RECT 2604.830 2667.450 2605.130 2680.750 ;
        RECT 2603.910 2667.150 2605.130 2667.450 ;
        RECT 2603.910 2650.450 2604.210 2667.150 ;
        RECT 2603.910 2650.150 2606.050 2650.450 ;
        RECT 2605.750 2558.650 2606.050 2650.150 ;
        RECT 2605.750 2558.350 2607.890 2558.650 ;
        RECT 2607.590 2517.865 2607.890 2558.350 ;
        RECT 2606.655 2517.850 2606.985 2517.865 ;
        RECT 2605.750 2517.550 2606.985 2517.850 ;
        RECT 2605.750 2490.650 2606.050 2517.550 ;
        RECT 2606.655 2517.535 2606.985 2517.550 ;
        RECT 2607.575 2517.535 2607.905 2517.865 ;
        RECT 2606.655 2490.650 2606.985 2490.665 ;
        RECT 2605.750 2490.350 2606.985 2490.650 ;
        RECT 2606.655 2490.335 2606.985 2490.350 ;
        RECT 2606.655 2443.050 2606.985 2443.065 ;
        RECT 2604.830 2442.750 2606.985 2443.050 ;
        RECT 2604.830 2364.850 2605.130 2442.750 ;
        RECT 2606.655 2442.735 2606.985 2442.750 ;
        RECT 2604.830 2364.550 2606.970 2364.850 ;
        RECT 2606.670 2362.825 2606.970 2364.550 ;
        RECT 2606.655 2362.495 2606.985 2362.825 ;
        RECT 2606.655 2328.495 2606.985 2328.825 ;
        RECT 2606.670 2310.450 2606.970 2328.495 ;
        RECT 2604.830 2310.150 2606.970 2310.450 ;
        RECT 2604.830 2290.050 2605.130 2310.150 ;
        RECT 2604.830 2289.750 2607.890 2290.050 ;
        RECT 2607.590 2279.850 2607.890 2289.750 ;
        RECT 2604.830 2279.550 2607.890 2279.850 ;
        RECT 2604.830 2235.650 2605.130 2279.550 ;
        RECT 2604.830 2235.350 2606.970 2235.650 ;
        RECT 2606.670 2232.945 2606.970 2235.350 ;
        RECT 2606.655 2232.615 2606.985 2232.945 ;
        RECT 2606.655 2174.450 2606.985 2174.465 ;
        RECT 2604.830 2174.150 2606.985 2174.450 ;
        RECT 2604.830 1922.850 2605.130 2174.150 ;
        RECT 2606.655 2174.135 2606.985 2174.150 ;
        RECT 2604.830 1922.550 2606.050 1922.850 ;
        RECT 2605.750 1916.050 2606.050 1922.550 ;
        RECT 2604.830 1915.750 2606.050 1916.050 ;
        RECT 2604.830 1868.450 2605.130 1915.750 ;
        RECT 2606.655 1868.450 2606.985 1868.465 ;
        RECT 2604.830 1868.150 2606.985 1868.450 ;
        RECT 2606.655 1868.135 2606.985 1868.150 ;
        RECT 2606.655 1857.255 2606.985 1857.585 ;
        RECT 2606.670 1854.850 2606.970 1857.255 ;
        RECT 2604.830 1854.550 2606.970 1854.850 ;
        RECT 2604.830 1810.650 2605.130 1854.550 ;
        RECT 2604.830 1810.350 2606.970 1810.650 ;
        RECT 2606.670 1776.650 2606.970 1810.350 ;
        RECT 2604.830 1776.350 2606.970 1776.650 ;
        RECT 2604.830 1627.050 2605.130 1776.350 ;
        RECT 2604.830 1626.750 2606.050 1627.050 ;
        RECT 2605.750 1610.730 2606.050 1626.750 ;
        RECT 2606.655 1610.730 2606.985 1610.745 ;
        RECT 2605.750 1610.430 2606.985 1610.730 ;
        RECT 2606.655 1610.415 2606.985 1610.430 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 65.860 427.730 65.920 ;
        RECT 2125.730 65.860 2126.050 65.920 ;
        RECT 427.410 65.720 2126.050 65.860 ;
        RECT 427.410 65.660 427.730 65.720 ;
        RECT 2125.730 65.660 2126.050 65.720 ;
        RECT 2125.730 37.640 2126.050 37.700 ;
        RECT 2131.710 37.640 2132.030 37.700 ;
        RECT 2125.730 37.500 2132.030 37.640 ;
        RECT 2125.730 37.440 2126.050 37.500 ;
        RECT 2131.710 37.440 2132.030 37.500 ;
      LAYER via ;
        RECT 427.440 65.660 427.700 65.920 ;
        RECT 2125.760 65.660 2126.020 65.920 ;
        RECT 2125.760 37.440 2126.020 37.700 ;
        RECT 2131.740 37.440 2132.000 37.700 ;
      LAYER met2 ;
        RECT 426.930 260.170 427.210 264.000 ;
        RECT 426.930 260.030 427.640 260.170 ;
        RECT 426.930 260.000 427.210 260.030 ;
        RECT 427.500 65.950 427.640 260.030 ;
        RECT 427.440 65.630 427.700 65.950 ;
        RECT 2125.760 65.630 2126.020 65.950 ;
        RECT 2125.820 37.730 2125.960 65.630 ;
        RECT 2125.760 37.410 2126.020 37.730 ;
        RECT 2131.740 37.410 2132.000 37.730 ;
        RECT 2131.800 2.400 2131.940 37.410 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 155.960 1773.230 156.020 ;
        RECT 2145.970 155.960 2146.290 156.020 ;
        RECT 1772.910 155.820 2146.290 155.960 ;
        RECT 1772.910 155.760 1773.230 155.820 ;
        RECT 2145.970 155.760 2146.290 155.820 ;
        RECT 2145.970 62.120 2146.290 62.180 ;
        RECT 2149.650 62.120 2149.970 62.180 ;
        RECT 2145.970 61.980 2149.970 62.120 ;
        RECT 2145.970 61.920 2146.290 61.980 ;
        RECT 2149.650 61.920 2149.970 61.980 ;
      LAYER via ;
        RECT 1772.940 155.760 1773.200 156.020 ;
        RECT 2146.000 155.760 2146.260 156.020 ;
        RECT 2146.000 61.920 2146.260 62.180 ;
        RECT 2149.680 61.920 2149.940 62.180 ;
      LAYER met2 ;
        RECT 1771.050 260.170 1771.330 264.000 ;
        RECT 1771.050 260.030 1773.140 260.170 ;
        RECT 1771.050 260.000 1771.330 260.030 ;
        RECT 1773.000 156.050 1773.140 260.030 ;
        RECT 1772.940 155.730 1773.200 156.050 ;
        RECT 2146.000 155.730 2146.260 156.050 ;
        RECT 2146.060 62.210 2146.200 155.730 ;
        RECT 2146.000 61.890 2146.260 62.210 ;
        RECT 2149.680 61.890 2149.940 62.210 ;
        RECT 2149.740 2.400 2149.880 61.890 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2132.170 48.520 2132.490 48.580 ;
        RECT 2167.590 48.520 2167.910 48.580 ;
        RECT 2132.170 48.380 2167.910 48.520 ;
        RECT 2132.170 48.320 2132.490 48.380 ;
        RECT 2167.590 48.320 2167.910 48.380 ;
      LAYER via ;
        RECT 2132.200 48.320 2132.460 48.580 ;
        RECT 2167.620 48.320 2167.880 48.580 ;
      LAYER met2 ;
        RECT 2132.190 86.515 2132.470 86.885 ;
        RECT 2132.260 48.610 2132.400 86.515 ;
        RECT 2132.200 48.290 2132.460 48.610 ;
        RECT 2167.620 48.290 2167.880 48.610 ;
        RECT 2167.680 2.400 2167.820 48.290 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
      LAYER via2 ;
        RECT 2132.190 86.560 2132.470 86.840 ;
      LAYER met3 ;
        RECT 305.710 2588.570 306.090 2588.580 ;
        RECT 310.000 2588.570 314.000 2588.960 ;
        RECT 305.710 2588.360 314.000 2588.570 ;
        RECT 305.710 2588.270 310.500 2588.360 ;
        RECT 305.710 2588.260 306.090 2588.270 ;
        RECT 305.710 86.850 306.090 86.860 ;
        RECT 2132.165 86.850 2132.495 86.865 ;
        RECT 305.710 86.550 2132.495 86.850 ;
        RECT 305.710 86.540 306.090 86.550 ;
        RECT 2132.165 86.535 2132.495 86.550 ;
      LAYER via3 ;
        RECT 305.740 2588.260 306.060 2588.580 ;
        RECT 305.740 86.540 306.060 86.860 ;
      LAYER met4 ;
        RECT 305.735 2588.255 306.065 2588.585 ;
        RECT 305.750 86.865 306.050 2588.255 ;
        RECT 305.735 86.535 306.065 86.865 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 297.690 217.160 298.010 217.220 ;
        RECT 2180.470 217.160 2180.790 217.220 ;
        RECT 297.690 217.020 2180.790 217.160 ;
        RECT 297.690 216.960 298.010 217.020 ;
        RECT 2180.470 216.960 2180.790 217.020 ;
        RECT 2180.470 62.120 2180.790 62.180 ;
        RECT 2185.070 62.120 2185.390 62.180 ;
        RECT 2180.470 61.980 2185.390 62.120 ;
        RECT 2180.470 61.920 2180.790 61.980 ;
        RECT 2185.070 61.920 2185.390 61.980 ;
      LAYER via ;
        RECT 297.720 216.960 297.980 217.220 ;
        RECT 2180.500 216.960 2180.760 217.220 ;
        RECT 2180.500 61.920 2180.760 62.180 ;
        RECT 2185.100 61.920 2185.360 62.180 ;
      LAYER met2 ;
        RECT 297.710 1003.835 297.990 1004.205 ;
        RECT 297.780 217.250 297.920 1003.835 ;
        RECT 297.720 216.930 297.980 217.250 ;
        RECT 2180.500 216.930 2180.760 217.250 ;
        RECT 2180.560 62.210 2180.700 216.930 ;
        RECT 2180.500 61.890 2180.760 62.210 ;
        RECT 2185.100 61.890 2185.360 62.210 ;
        RECT 2185.160 2.400 2185.300 61.890 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
      LAYER via2 ;
        RECT 297.710 1003.880 297.990 1004.160 ;
      LAYER met3 ;
        RECT 297.685 1004.170 298.015 1004.185 ;
        RECT 310.000 1004.170 314.000 1004.560 ;
        RECT 297.685 1003.960 314.000 1004.170 ;
        RECT 297.685 1003.870 310.500 1003.960 ;
        RECT 297.685 1003.855 298.015 1003.870 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2283.970 26.420 2284.290 26.480 ;
        RECT 2259.220 26.280 2284.290 26.420 ;
        RECT 2203.010 25.740 2203.330 25.800 ;
        RECT 2259.220 25.740 2259.360 26.280 ;
        RECT 2283.970 26.220 2284.290 26.280 ;
        RECT 2203.010 25.600 2259.360 25.740 ;
        RECT 2203.010 25.540 2203.330 25.600 ;
      LAYER via ;
        RECT 2203.040 25.540 2203.300 25.800 ;
        RECT 2284.000 26.220 2284.260 26.480 ;
      LAYER met2 ;
        RECT 2285.330 260.170 2285.610 264.000 ;
        RECT 2284.060 260.030 2285.610 260.170 ;
        RECT 2284.060 26.510 2284.200 260.030 ;
        RECT 2285.330 260.000 2285.610 260.030 ;
        RECT 2284.000 26.190 2284.260 26.510 ;
        RECT 2203.040 25.510 2203.300 25.830 ;
        RECT 2203.100 2.400 2203.240 25.510 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2583.430 3261.180 2583.750 3261.240 ;
        RECT 2663.930 3261.180 2664.250 3261.240 ;
        RECT 2583.430 3261.040 2664.250 3261.180 ;
        RECT 2583.430 3260.980 2583.750 3261.040 ;
        RECT 2663.930 3260.980 2664.250 3261.040 ;
      LAYER via ;
        RECT 2583.460 3260.980 2583.720 3261.240 ;
        RECT 2663.960 3260.980 2664.220 3261.240 ;
      LAYER met2 ;
        RECT 704.810 3270.955 705.090 3271.325 ;
        RECT 2583.450 3270.955 2583.730 3271.325 ;
        RECT 704.880 3260.000 705.020 3270.955 ;
        RECT 2583.520 3261.270 2583.660 3270.955 ;
        RECT 2583.460 3260.950 2583.720 3261.270 ;
        RECT 2663.960 3260.950 2664.220 3261.270 ;
        RECT 704.770 3256.000 705.050 3260.000 ;
        RECT 2664.020 18.205 2664.160 3260.950 ;
        RECT 2220.970 17.835 2221.250 18.205 ;
        RECT 2663.950 17.835 2664.230 18.205 ;
        RECT 2221.040 2.400 2221.180 17.835 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
      LAYER via2 ;
        RECT 704.810 3271.000 705.090 3271.280 ;
        RECT 2583.450 3271.000 2583.730 3271.280 ;
        RECT 2220.970 17.880 2221.250 18.160 ;
        RECT 2663.950 17.880 2664.230 18.160 ;
      LAYER met3 ;
        RECT 704.785 3271.290 705.115 3271.305 ;
        RECT 2583.425 3271.290 2583.755 3271.305 ;
        RECT 704.785 3270.990 2583.755 3271.290 ;
        RECT 704.785 3270.975 705.115 3270.990 ;
        RECT 2583.425 3270.975 2583.755 3270.990 ;
        RECT 2220.945 18.170 2221.275 18.185 ;
        RECT 2663.925 18.170 2664.255 18.185 ;
        RECT 2220.945 17.870 2664.255 18.170 ;
        RECT 2220.945 17.855 2221.275 17.870 ;
        RECT 2663.925 17.855 2664.255 17.870 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 100.200 779.630 100.260 ;
        RECT 2608.270 100.200 2608.590 100.260 ;
        RECT 779.310 100.060 2608.590 100.200 ;
        RECT 779.310 100.000 779.630 100.060 ;
        RECT 2608.270 100.000 2608.590 100.060 ;
        RECT 775.630 20.640 775.950 20.700 ;
        RECT 779.310 20.640 779.630 20.700 ;
        RECT 775.630 20.500 779.630 20.640 ;
        RECT 775.630 20.440 775.950 20.500 ;
        RECT 779.310 20.440 779.630 20.500 ;
      LAYER via ;
        RECT 779.340 100.000 779.600 100.260 ;
        RECT 2608.300 100.000 2608.560 100.260 ;
        RECT 775.660 20.440 775.920 20.700 ;
        RECT 779.340 20.440 779.600 20.700 ;
      LAYER met2 ;
        RECT 2608.290 378.915 2608.570 379.285 ;
        RECT 2608.360 100.290 2608.500 378.915 ;
        RECT 779.340 99.970 779.600 100.290 ;
        RECT 2608.300 99.970 2608.560 100.290 ;
        RECT 779.400 20.730 779.540 99.970 ;
        RECT 775.660 20.410 775.920 20.730 ;
        RECT 779.340 20.410 779.600 20.730 ;
        RECT 775.720 2.400 775.860 20.410 ;
        RECT 775.510 -4.800 776.070 2.400 ;
      LAYER via2 ;
        RECT 2608.290 378.960 2608.570 379.240 ;
      LAYER met3 ;
        RECT 2606.000 381.080 2610.000 381.680 ;
        RECT 2608.265 379.250 2608.595 379.265 ;
        RECT 2609.430 379.250 2609.730 381.080 ;
        RECT 2608.265 378.950 2609.730 379.250 ;
        RECT 2608.265 378.935 2608.595 378.950 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1020.810 3257.780 1021.130 3257.840 ;
        RECT 2645.990 3257.780 2646.310 3257.840 ;
        RECT 1020.810 3257.640 2646.310 3257.780 ;
        RECT 1020.810 3257.580 1021.130 3257.640 ;
        RECT 2645.990 3257.580 2646.310 3257.640 ;
        RECT 2645.990 297.400 2646.310 297.460 ;
        RECT 2657.490 297.400 2657.810 297.460 ;
        RECT 2645.990 297.260 2657.810 297.400 ;
        RECT 2645.990 297.200 2646.310 297.260 ;
        RECT 2657.490 297.200 2657.810 297.260 ;
      LAYER via ;
        RECT 1020.840 3257.580 1021.100 3257.840 ;
        RECT 2646.020 3257.580 2646.280 3257.840 ;
        RECT 2646.020 297.200 2646.280 297.460 ;
        RECT 2657.520 297.200 2657.780 297.460 ;
      LAYER met2 ;
        RECT 1019.410 3257.610 1019.690 3260.000 ;
        RECT 1020.840 3257.610 1021.100 3257.870 ;
        RECT 1019.410 3257.550 1021.100 3257.610 ;
        RECT 2646.020 3257.550 2646.280 3257.870 ;
        RECT 1019.410 3257.470 1021.040 3257.550 ;
        RECT 1019.410 3256.000 1019.690 3257.470 ;
        RECT 2646.080 297.490 2646.220 3257.550 ;
        RECT 2646.020 297.170 2646.280 297.490 ;
        RECT 2657.520 297.170 2657.780 297.490 ;
        RECT 2657.580 18.885 2657.720 297.170 ;
        RECT 2238.910 18.515 2239.190 18.885 ;
        RECT 2657.510 18.515 2657.790 18.885 ;
        RECT 2238.980 2.400 2239.120 18.515 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
      LAYER via2 ;
        RECT 2238.910 18.560 2239.190 18.840 ;
        RECT 2657.510 18.560 2657.790 18.840 ;
      LAYER met3 ;
        RECT 2238.885 18.850 2239.215 18.865 ;
        RECT 2657.485 18.850 2657.815 18.865 ;
        RECT 2238.885 18.550 2657.815 18.850 ;
        RECT 2238.885 18.535 2239.215 18.550 ;
        RECT 2657.485 18.535 2657.815 18.550 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2318.545 15.725 2318.715 16.915 ;
        RECT 2342.465 16.745 2342.635 17.935 ;
        RECT 2387.085 15.385 2387.255 17.935 ;
        RECT 2452.865 15.385 2453.035 17.935 ;
        RECT 2501.165 15.385 2501.335 17.935 ;
        RECT 2549.465 15.385 2549.635 17.935 ;
      LAYER mcon ;
        RECT 2342.465 17.765 2342.635 17.935 ;
        RECT 2318.545 16.745 2318.715 16.915 ;
        RECT 2387.085 17.765 2387.255 17.935 ;
        RECT 2452.865 17.765 2453.035 17.935 ;
        RECT 2501.165 17.765 2501.335 17.935 ;
        RECT 2549.465 17.765 2549.635 17.935 ;
      LAYER met1 ;
        RECT 2206.230 3274.440 2206.550 3274.500 ;
        RECT 2553.070 3274.440 2553.390 3274.500 ;
        RECT 2206.230 3274.300 2553.390 3274.440 ;
        RECT 2206.230 3274.240 2206.550 3274.300 ;
        RECT 2553.070 3274.240 2553.390 3274.300 ;
        RECT 2553.070 3261.520 2553.390 3261.580 ;
        RECT 2618.390 3261.520 2618.710 3261.580 ;
        RECT 2553.070 3261.380 2618.710 3261.520 ;
        RECT 2553.070 3261.320 2553.390 3261.380 ;
        RECT 2618.390 3261.320 2618.710 3261.380 ;
        RECT 2618.390 669.360 2618.710 669.420 ;
        RECT 2640.010 669.360 2640.330 669.420 ;
        RECT 2618.390 669.220 2640.330 669.360 ;
        RECT 2618.390 669.160 2618.710 669.220 ;
        RECT 2640.010 669.160 2640.330 669.220 ;
        RECT 2342.405 17.920 2342.695 17.965 ;
        RECT 2387.025 17.920 2387.315 17.965 ;
        RECT 2342.405 17.780 2387.315 17.920 ;
        RECT 2342.405 17.735 2342.695 17.780 ;
        RECT 2387.025 17.735 2387.315 17.780 ;
        RECT 2452.805 17.920 2453.095 17.965 ;
        RECT 2501.105 17.920 2501.395 17.965 ;
        RECT 2452.805 17.780 2501.395 17.920 ;
        RECT 2452.805 17.735 2453.095 17.780 ;
        RECT 2501.105 17.735 2501.395 17.780 ;
        RECT 2549.405 17.920 2549.695 17.965 ;
        RECT 2549.405 17.780 2580.900 17.920 ;
        RECT 2549.405 17.735 2549.695 17.780 ;
        RECT 2580.760 17.580 2580.900 17.780 ;
        RECT 2640.010 17.580 2640.330 17.640 ;
        RECT 2580.760 17.440 2640.330 17.580 ;
        RECT 2640.010 17.380 2640.330 17.440 ;
        RECT 2318.485 16.900 2318.775 16.945 ;
        RECT 2342.405 16.900 2342.695 16.945 ;
        RECT 2318.485 16.760 2342.695 16.900 ;
        RECT 2318.485 16.715 2318.775 16.760 ;
        RECT 2342.405 16.715 2342.695 16.760 ;
        RECT 2256.370 15.880 2256.690 15.940 ;
        RECT 2318.485 15.880 2318.775 15.925 ;
        RECT 2256.370 15.740 2318.775 15.880 ;
        RECT 2256.370 15.680 2256.690 15.740 ;
        RECT 2318.485 15.695 2318.775 15.740 ;
        RECT 2387.025 15.540 2387.315 15.585 ;
        RECT 2452.805 15.540 2453.095 15.585 ;
        RECT 2387.025 15.400 2453.095 15.540 ;
        RECT 2387.025 15.355 2387.315 15.400 ;
        RECT 2452.805 15.355 2453.095 15.400 ;
        RECT 2501.105 15.540 2501.395 15.585 ;
        RECT 2549.405 15.540 2549.695 15.585 ;
        RECT 2501.105 15.400 2549.695 15.540 ;
        RECT 2501.105 15.355 2501.395 15.400 ;
        RECT 2549.405 15.355 2549.695 15.400 ;
      LAYER via ;
        RECT 2206.260 3274.240 2206.520 3274.500 ;
        RECT 2553.100 3274.240 2553.360 3274.500 ;
        RECT 2553.100 3261.320 2553.360 3261.580 ;
        RECT 2618.420 3261.320 2618.680 3261.580 ;
        RECT 2618.420 669.160 2618.680 669.420 ;
        RECT 2640.040 669.160 2640.300 669.420 ;
        RECT 2640.040 17.380 2640.300 17.640 ;
        RECT 2256.400 15.680 2256.660 15.940 ;
      LAYER met2 ;
        RECT 2206.260 3274.210 2206.520 3274.530 ;
        RECT 2553.100 3274.210 2553.360 3274.530 ;
        RECT 2206.320 3260.000 2206.460 3274.210 ;
        RECT 2553.160 3261.610 2553.300 3274.210 ;
        RECT 2553.100 3261.290 2553.360 3261.610 ;
        RECT 2618.420 3261.290 2618.680 3261.610 ;
        RECT 2206.210 3256.000 2206.490 3260.000 ;
        RECT 2618.480 669.450 2618.620 3261.290 ;
        RECT 2618.420 669.130 2618.680 669.450 ;
        RECT 2640.040 669.130 2640.300 669.450 ;
        RECT 2640.100 17.670 2640.240 669.130 ;
        RECT 2640.040 17.350 2640.300 17.670 ;
        RECT 2256.400 15.650 2256.660 15.970 ;
        RECT 2256.460 2.400 2256.600 15.650 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2270.170 62.120 2270.490 62.180 ;
        RECT 2274.310 62.120 2274.630 62.180 ;
        RECT 2270.170 61.980 2274.630 62.120 ;
        RECT 2270.170 61.920 2270.490 61.980 ;
        RECT 2274.310 61.920 2274.630 61.980 ;
      LAYER via ;
        RECT 2270.200 61.920 2270.460 62.180 ;
        RECT 2274.340 61.920 2274.600 62.180 ;
      LAYER met2 ;
        RECT 2270.190 223.875 2270.470 224.245 ;
        RECT 2270.260 62.210 2270.400 223.875 ;
        RECT 2270.200 61.890 2270.460 62.210 ;
        RECT 2274.340 61.890 2274.600 62.210 ;
        RECT 2274.400 2.400 2274.540 61.890 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
      LAYER via2 ;
        RECT 2270.190 223.920 2270.470 224.200 ;
      LAYER met3 ;
        RECT 300.190 918.490 300.570 918.500 ;
        RECT 310.000 918.490 314.000 918.880 ;
        RECT 300.190 918.280 314.000 918.490 ;
        RECT 300.190 918.190 310.500 918.280 ;
        RECT 300.190 918.180 300.570 918.190 ;
        RECT 300.190 224.210 300.570 224.220 ;
        RECT 2270.165 224.210 2270.495 224.225 ;
        RECT 300.190 223.910 2270.495 224.210 ;
        RECT 300.190 223.900 300.570 223.910 ;
        RECT 2270.165 223.895 2270.495 223.910 ;
      LAYER via3 ;
        RECT 300.220 918.180 300.540 918.500 ;
        RECT 300.220 223.900 300.540 224.220 ;
      LAYER met4 ;
        RECT 300.215 918.175 300.545 918.505 ;
        RECT 300.230 224.225 300.530 918.175 ;
        RECT 300.215 223.895 300.545 224.225 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2290.890 134.115 2291.170 134.485 ;
        RECT 2290.960 3.130 2291.100 134.115 ;
        RECT 2290.960 2.990 2292.020 3.130 ;
        RECT 2291.880 2.960 2292.020 2.990 ;
        RECT 2291.880 2.820 2292.480 2.960 ;
        RECT 2292.340 2.400 2292.480 2.820 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
      LAYER via2 ;
        RECT 2290.890 134.160 2291.170 134.440 ;
      LAYER met3 ;
        RECT 306.630 1658.330 307.010 1658.340 ;
        RECT 310.000 1658.330 314.000 1658.720 ;
        RECT 306.630 1658.120 314.000 1658.330 ;
        RECT 306.630 1658.030 310.500 1658.120 ;
        RECT 306.630 1658.020 307.010 1658.030 ;
        RECT 306.630 134.450 307.010 134.460 ;
        RECT 2290.865 134.450 2291.195 134.465 ;
        RECT 306.630 134.150 2291.195 134.450 ;
        RECT 306.630 134.140 307.010 134.150 ;
        RECT 2290.865 134.135 2291.195 134.150 ;
      LAYER via3 ;
        RECT 306.660 1658.020 306.980 1658.340 ;
        RECT 306.660 134.140 306.980 134.460 ;
      LAYER met4 ;
        RECT 306.655 1658.015 306.985 1658.345 ;
        RECT 306.670 134.465 306.970 1658.015 ;
        RECT 306.655 134.135 306.985 134.465 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1317.050 74.360 1317.370 74.420 ;
        RECT 2304.670 74.360 2304.990 74.420 ;
        RECT 1317.050 74.220 2304.990 74.360 ;
        RECT 1317.050 74.160 1317.370 74.220 ;
        RECT 2304.670 74.160 2304.990 74.220 ;
        RECT 2304.670 48.180 2304.990 48.240 ;
        RECT 2310.190 48.180 2310.510 48.240 ;
        RECT 2304.670 48.040 2310.510 48.180 ;
        RECT 2304.670 47.980 2304.990 48.040 ;
        RECT 2310.190 47.980 2310.510 48.040 ;
      LAYER via ;
        RECT 1317.080 74.160 1317.340 74.420 ;
        RECT 2304.700 74.160 2304.960 74.420 ;
        RECT 2304.700 47.980 2304.960 48.240 ;
        RECT 2310.220 47.980 2310.480 48.240 ;
      LAYER met2 ;
        RECT 1313.810 260.170 1314.090 264.000 ;
        RECT 1313.810 260.030 1317.280 260.170 ;
        RECT 1313.810 260.000 1314.090 260.030 ;
        RECT 1317.140 74.450 1317.280 260.030 ;
        RECT 1317.080 74.130 1317.340 74.450 ;
        RECT 2304.700 74.130 2304.960 74.450 ;
        RECT 2304.760 48.270 2304.900 74.130 ;
        RECT 2304.700 47.950 2304.960 48.270 ;
        RECT 2310.220 47.950 2310.480 48.270 ;
        RECT 2310.280 2.400 2310.420 47.950 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 257.210 828.620 257.530 828.880 ;
        RECT 257.300 828.200 257.440 828.620 ;
        RECT 257.210 827.940 257.530 828.200 ;
      LAYER via ;
        RECT 257.240 828.620 257.500 828.880 ;
        RECT 257.240 827.940 257.500 828.200 ;
      LAYER met2 ;
        RECT 257.230 3260.075 257.510 3260.445 ;
        RECT 560.370 3260.075 560.650 3260.445 ;
        RECT 257.300 828.910 257.440 3260.075 ;
        RECT 560.440 3259.650 560.580 3260.075 ;
        RECT 562.170 3259.650 562.450 3260.000 ;
        RECT 560.440 3259.510 562.450 3259.650 ;
        RECT 562.170 3256.000 562.450 3259.510 ;
        RECT 257.240 828.590 257.500 828.910 ;
        RECT 257.240 827.910 257.500 828.230 ;
        RECT 257.300 32.485 257.440 827.910 ;
        RECT 257.230 32.115 257.510 32.485 ;
        RECT 2328.150 32.115 2328.430 32.485 ;
        RECT 2328.220 2.400 2328.360 32.115 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
      LAYER via2 ;
        RECT 257.230 3260.120 257.510 3260.400 ;
        RECT 560.370 3260.120 560.650 3260.400 ;
        RECT 257.230 32.160 257.510 32.440 ;
        RECT 2328.150 32.160 2328.430 32.440 ;
      LAYER met3 ;
        RECT 257.205 3260.410 257.535 3260.425 ;
        RECT 560.345 3260.410 560.675 3260.425 ;
        RECT 257.205 3260.110 560.675 3260.410 ;
        RECT 257.205 3260.095 257.535 3260.110 ;
        RECT 560.345 3260.095 560.675 3260.110 ;
        RECT 257.205 32.450 257.535 32.465 ;
        RECT 2328.125 32.450 2328.455 32.465 ;
        RECT 257.205 32.150 2328.455 32.450 ;
        RECT 257.205 32.135 257.535 32.150 ;
        RECT 2328.125 32.135 2328.455 32.150 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1118.160 2615.490 1118.220 ;
        RECT 2659.330 1118.160 2659.650 1118.220 ;
        RECT 2615.170 1118.020 2659.650 1118.160 ;
        RECT 2615.170 1117.960 2615.490 1118.020 ;
        RECT 2659.330 1117.960 2659.650 1118.020 ;
        RECT 2345.150 16.900 2345.470 16.960 ;
        RECT 2559.970 16.900 2560.290 16.960 ;
        RECT 2345.150 16.760 2560.290 16.900 ;
        RECT 2345.150 16.700 2345.470 16.760 ;
        RECT 2559.970 16.700 2560.290 16.760 ;
        RECT 2561.350 16.900 2561.670 16.960 ;
        RECT 2659.330 16.900 2659.650 16.960 ;
        RECT 2561.350 16.760 2659.650 16.900 ;
        RECT 2561.350 16.700 2561.670 16.760 ;
        RECT 2659.330 16.700 2659.650 16.760 ;
      LAYER via ;
        RECT 2615.200 1117.960 2615.460 1118.220 ;
        RECT 2659.360 1117.960 2659.620 1118.220 ;
        RECT 2345.180 16.700 2345.440 16.960 ;
        RECT 2560.000 16.700 2560.260 16.960 ;
        RECT 2561.380 16.700 2561.640 16.960 ;
        RECT 2659.360 16.700 2659.620 16.960 ;
      LAYER met2 ;
        RECT 2615.190 1120.795 2615.470 1121.165 ;
        RECT 2615.260 1118.250 2615.400 1120.795 ;
        RECT 2615.200 1117.930 2615.460 1118.250 ;
        RECT 2659.360 1117.930 2659.620 1118.250 ;
        RECT 2659.420 16.990 2659.560 1117.930 ;
        RECT 2345.180 16.670 2345.440 16.990 ;
        RECT 2560.000 16.730 2560.260 16.990 ;
        RECT 2561.380 16.730 2561.640 16.990 ;
        RECT 2560.000 16.670 2561.640 16.730 ;
        RECT 2659.360 16.670 2659.620 16.990 ;
        RECT 2345.240 14.010 2345.380 16.670 ;
        RECT 2560.060 16.590 2561.580 16.670 ;
        RECT 2345.240 13.870 2345.840 14.010 ;
        RECT 2345.700 2.400 2345.840 13.870 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1120.840 2615.470 1121.120 ;
      LAYER met3 ;
        RECT 2606.000 1121.130 2610.000 1121.520 ;
        RECT 2615.165 1121.130 2615.495 1121.145 ;
        RECT 2606.000 1120.920 2615.495 1121.130 ;
        RECT 2609.580 1120.830 2615.495 1120.920 ;
        RECT 2615.165 1120.815 2615.495 1120.830 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 231.910 2373.780 232.230 2373.840 ;
        RECT 296.770 2373.780 297.090 2373.840 ;
        RECT 231.910 2373.640 297.090 2373.780 ;
        RECT 231.910 2373.580 232.230 2373.640 ;
        RECT 296.770 2373.580 297.090 2373.640 ;
        RECT 231.910 46.140 232.230 46.200 ;
        RECT 2363.550 46.140 2363.870 46.200 ;
        RECT 231.910 46.000 2363.870 46.140 ;
        RECT 231.910 45.940 232.230 46.000 ;
        RECT 2363.550 45.940 2363.870 46.000 ;
      LAYER via ;
        RECT 231.940 2373.580 232.200 2373.840 ;
        RECT 296.800 2373.580 297.060 2373.840 ;
        RECT 231.940 45.940 232.200 46.200 ;
        RECT 2363.580 45.940 2363.840 46.200 ;
      LAYER met2 ;
        RECT 296.790 2377.435 297.070 2377.805 ;
        RECT 296.860 2373.870 297.000 2377.435 ;
        RECT 231.940 2373.550 232.200 2373.870 ;
        RECT 296.800 2373.550 297.060 2373.870 ;
        RECT 232.000 46.230 232.140 2373.550 ;
        RECT 231.940 45.910 232.200 46.230 ;
        RECT 2363.580 45.910 2363.840 46.230 ;
        RECT 2363.640 2.400 2363.780 45.910 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 296.790 2377.480 297.070 2377.760 ;
      LAYER met3 ;
        RECT 296.765 2377.770 297.095 2377.785 ;
        RECT 310.000 2377.770 314.000 2378.160 ;
        RECT 296.765 2377.560 314.000 2377.770 ;
        RECT 296.765 2377.470 310.500 2377.560 ;
        RECT 296.765 2377.455 297.095 2377.470 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2057.190 244.020 2057.510 244.080 ;
        RECT 2062.710 244.020 2063.030 244.080 ;
        RECT 2057.190 243.880 2063.030 244.020 ;
        RECT 2057.190 243.820 2057.510 243.880 ;
        RECT 2062.710 243.820 2063.030 243.880 ;
        RECT 2062.710 24.040 2063.030 24.100 ;
        RECT 2381.490 24.040 2381.810 24.100 ;
        RECT 2062.710 23.900 2381.810 24.040 ;
        RECT 2062.710 23.840 2063.030 23.900 ;
        RECT 2381.490 23.840 2381.810 23.900 ;
      LAYER via ;
        RECT 2057.220 243.820 2057.480 244.080 ;
        RECT 2062.740 243.820 2063.000 244.080 ;
        RECT 2062.740 23.840 2063.000 24.100 ;
        RECT 2381.520 23.840 2381.780 24.100 ;
      LAYER met2 ;
        RECT 2057.170 260.000 2057.450 264.000 ;
        RECT 2057.280 244.110 2057.420 260.000 ;
        RECT 2057.220 243.790 2057.480 244.110 ;
        RECT 2062.740 243.790 2063.000 244.110 ;
        RECT 2062.800 24.130 2062.940 243.790 ;
        RECT 2062.740 23.810 2063.000 24.130 ;
        RECT 2381.520 23.810 2381.780 24.130 ;
        RECT 2381.580 2.400 2381.720 23.810 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2400.885 241.485 2401.055 261.035 ;
        RECT 2400.885 144.925 2401.055 193.035 ;
        RECT 2400.885 48.365 2401.055 96.475 ;
      LAYER mcon ;
        RECT 2400.885 260.865 2401.055 261.035 ;
        RECT 2400.885 192.865 2401.055 193.035 ;
        RECT 2400.885 96.305 2401.055 96.475 ;
      LAYER met1 ;
        RECT 2615.170 2235.740 2615.490 2235.800 ;
        RECT 2679.570 2235.740 2679.890 2235.800 ;
        RECT 2615.170 2235.600 2679.890 2235.740 ;
        RECT 2615.170 2235.540 2615.490 2235.600 ;
        RECT 2679.570 2235.540 2679.890 2235.600 ;
        RECT 2400.825 261.020 2401.115 261.065 ;
        RECT 2679.570 261.020 2679.890 261.080 ;
        RECT 2400.825 260.880 2679.890 261.020 ;
        RECT 2400.825 260.835 2401.115 260.880 ;
        RECT 2679.570 260.820 2679.890 260.880 ;
        RECT 2400.810 241.640 2401.130 241.700 ;
        RECT 2400.615 241.500 2401.130 241.640 ;
        RECT 2400.810 241.440 2401.130 241.500 ;
        RECT 2400.810 193.020 2401.130 193.080 ;
        RECT 2400.615 192.880 2401.130 193.020 ;
        RECT 2400.810 192.820 2401.130 192.880 ;
        RECT 2400.810 145.080 2401.130 145.140 ;
        RECT 2400.615 144.940 2401.130 145.080 ;
        RECT 2400.810 144.880 2401.130 144.940 ;
        RECT 2400.810 96.460 2401.130 96.520 ;
        RECT 2400.615 96.320 2401.130 96.460 ;
        RECT 2400.810 96.260 2401.130 96.320 ;
        RECT 2400.810 48.520 2401.130 48.580 ;
        RECT 2400.615 48.380 2401.130 48.520 ;
        RECT 2400.810 48.320 2401.130 48.380 ;
        RECT 2400.810 14.180 2401.130 14.240 ;
        RECT 2399.520 14.040 2401.130 14.180 ;
        RECT 2399.520 13.900 2399.660 14.040 ;
        RECT 2400.810 13.980 2401.130 14.040 ;
        RECT 2399.430 13.640 2399.750 13.900 ;
      LAYER via ;
        RECT 2615.200 2235.540 2615.460 2235.800 ;
        RECT 2679.600 2235.540 2679.860 2235.800 ;
        RECT 2679.600 260.820 2679.860 261.080 ;
        RECT 2400.840 241.440 2401.100 241.700 ;
        RECT 2400.840 192.820 2401.100 193.080 ;
        RECT 2400.840 144.880 2401.100 145.140 ;
        RECT 2400.840 96.260 2401.100 96.520 ;
        RECT 2400.840 48.320 2401.100 48.580 ;
        RECT 2400.840 13.980 2401.100 14.240 ;
        RECT 2399.460 13.640 2399.720 13.900 ;
      LAYER met2 ;
        RECT 2615.190 2240.075 2615.470 2240.445 ;
        RECT 2615.260 2235.830 2615.400 2240.075 ;
        RECT 2615.200 2235.510 2615.460 2235.830 ;
        RECT 2679.600 2235.510 2679.860 2235.830 ;
        RECT 2679.660 261.110 2679.800 2235.510 ;
        RECT 2679.600 260.790 2679.860 261.110 ;
        RECT 2400.840 241.410 2401.100 241.730 ;
        RECT 2400.900 193.110 2401.040 241.410 ;
        RECT 2400.840 192.790 2401.100 193.110 ;
        RECT 2400.840 144.850 2401.100 145.170 ;
        RECT 2400.900 96.550 2401.040 144.850 ;
        RECT 2400.840 96.230 2401.100 96.550 ;
        RECT 2400.840 48.290 2401.100 48.610 ;
        RECT 2400.900 14.270 2401.040 48.290 ;
        RECT 2400.840 13.950 2401.100 14.270 ;
        RECT 2399.460 13.610 2399.720 13.930 ;
        RECT 2399.520 2.400 2399.660 13.610 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2240.120 2615.470 2240.400 ;
      LAYER met3 ;
        RECT 2606.000 2240.410 2610.000 2240.800 ;
        RECT 2615.165 2240.410 2615.495 2240.425 ;
        RECT 2606.000 2240.200 2615.495 2240.410 ;
        RECT 2609.580 2240.110 2615.495 2240.200 ;
        RECT 2615.165 2240.095 2615.495 2240.110 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 252.150 1759.740 252.470 1759.800 ;
        RECT 296.770 1759.740 297.090 1759.800 ;
        RECT 252.150 1759.600 297.090 1759.740 ;
        RECT 252.150 1759.540 252.470 1759.600 ;
        RECT 296.770 1759.540 297.090 1759.600 ;
        RECT 252.150 33.220 252.470 33.280 ;
        RECT 793.570 33.220 793.890 33.280 ;
        RECT 252.150 33.080 793.890 33.220 ;
        RECT 252.150 33.020 252.470 33.080 ;
        RECT 793.570 33.020 793.890 33.080 ;
      LAYER via ;
        RECT 252.180 1759.540 252.440 1759.800 ;
        RECT 296.800 1759.540 297.060 1759.800 ;
        RECT 252.180 33.020 252.440 33.280 ;
        RECT 793.600 33.020 793.860 33.280 ;
      LAYER met2 ;
        RECT 296.790 1764.075 297.070 1764.445 ;
        RECT 296.860 1759.830 297.000 1764.075 ;
        RECT 252.180 1759.510 252.440 1759.830 ;
        RECT 296.800 1759.510 297.060 1759.830 ;
        RECT 252.240 33.310 252.380 1759.510 ;
        RECT 252.180 32.990 252.440 33.310 ;
        RECT 793.600 32.990 793.860 33.310 ;
        RECT 793.660 2.400 793.800 32.990 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 296.790 1764.120 297.070 1764.400 ;
      LAYER met3 ;
        RECT 296.765 1764.410 297.095 1764.425 ;
        RECT 310.000 1764.410 314.000 1764.800 ;
        RECT 296.765 1764.200 314.000 1764.410 ;
        RECT 296.765 1764.110 310.500 1764.200 ;
        RECT 296.765 1764.095 297.095 1764.110 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 25.060 639.330 25.120 ;
        RECT 1511.170 25.060 1511.490 25.120 ;
        RECT 639.010 24.920 1511.490 25.060 ;
        RECT 639.010 24.860 639.330 24.920 ;
        RECT 1511.170 24.860 1511.490 24.920 ;
      LAYER via ;
        RECT 639.040 24.860 639.300 25.120 ;
        RECT 1511.200 24.860 1511.460 25.120 ;
      LAYER met2 ;
        RECT 1513.450 260.170 1513.730 264.000 ;
        RECT 1511.260 260.030 1513.730 260.170 ;
        RECT 1511.260 25.150 1511.400 260.030 ;
        RECT 1513.450 260.000 1513.730 260.030 ;
        RECT 639.040 24.830 639.300 25.150 ;
        RECT 1511.200 24.830 1511.460 25.150 ;
        RECT 639.100 2.400 639.240 24.830 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2590.790 241.640 2591.110 241.700 ;
        RECT 2599.990 241.640 2600.310 241.700 ;
        RECT 2590.790 241.500 2600.310 241.640 ;
        RECT 2590.790 241.440 2591.110 241.500 ;
        RECT 2599.990 241.440 2600.310 241.500 ;
        RECT 2428.410 135.560 2428.730 135.620 ;
        RECT 2590.790 135.560 2591.110 135.620 ;
        RECT 2428.410 135.420 2591.110 135.560 ;
        RECT 2428.410 135.360 2428.730 135.420 ;
        RECT 2590.790 135.360 2591.110 135.420 ;
        RECT 2422.890 17.920 2423.210 17.980 ;
        RECT 2428.410 17.920 2428.730 17.980 ;
        RECT 2422.890 17.780 2428.730 17.920 ;
        RECT 2422.890 17.720 2423.210 17.780 ;
        RECT 2428.410 17.720 2428.730 17.780 ;
      LAYER via ;
        RECT 2590.820 241.440 2591.080 241.700 ;
        RECT 2600.020 241.440 2600.280 241.700 ;
        RECT 2428.440 135.360 2428.700 135.620 ;
        RECT 2590.820 135.360 2591.080 135.620 ;
        RECT 2422.920 17.720 2423.180 17.980 ;
        RECT 2428.440 17.720 2428.700 17.980 ;
      LAYER met2 ;
        RECT 2599.970 260.000 2600.250 264.000 ;
        RECT 2600.080 241.730 2600.220 260.000 ;
        RECT 2590.820 241.410 2591.080 241.730 ;
        RECT 2600.020 241.410 2600.280 241.730 ;
        RECT 2590.880 135.650 2591.020 241.410 ;
        RECT 2428.440 135.330 2428.700 135.650 ;
        RECT 2590.820 135.330 2591.080 135.650 ;
        RECT 2428.500 18.010 2428.640 135.330 ;
        RECT 2422.920 17.690 2423.180 18.010 ;
        RECT 2428.440 17.690 2428.700 18.010 ;
        RECT 2422.980 2.400 2423.120 17.690 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2439.985 89.845 2440.155 137.955 ;
        RECT 2440.905 2.805 2441.075 48.195 ;
      LAYER mcon ;
        RECT 2439.985 137.785 2440.155 137.955 ;
        RECT 2440.905 48.025 2441.075 48.195 ;
      LAYER met1 ;
        RECT 2442.210 258.300 2442.530 258.360 ;
        RECT 2611.030 258.300 2611.350 258.360 ;
        RECT 2442.210 258.160 2611.350 258.300 ;
        RECT 2442.210 258.100 2442.530 258.160 ;
        RECT 2611.030 258.100 2611.350 258.160 ;
        RECT 2442.210 186.560 2442.530 186.620 ;
        RECT 2443.130 186.560 2443.450 186.620 ;
        RECT 2442.210 186.420 2443.450 186.560 ;
        RECT 2442.210 186.360 2442.530 186.420 ;
        RECT 2443.130 186.360 2443.450 186.420 ;
        RECT 2439.925 137.940 2440.215 137.985 ;
        RECT 2442.210 137.940 2442.530 138.000 ;
        RECT 2439.925 137.800 2442.530 137.940 ;
        RECT 2439.925 137.755 2440.215 137.800 ;
        RECT 2442.210 137.740 2442.530 137.800 ;
        RECT 2439.910 90.000 2440.230 90.060 ;
        RECT 2439.715 89.860 2440.230 90.000 ;
        RECT 2439.910 89.800 2440.230 89.860 ;
        RECT 2440.830 48.180 2441.150 48.240 ;
        RECT 2440.635 48.040 2441.150 48.180 ;
        RECT 2440.830 47.980 2441.150 48.040 ;
        RECT 2440.830 2.960 2441.150 3.020 ;
        RECT 2440.635 2.820 2441.150 2.960 ;
        RECT 2440.830 2.760 2441.150 2.820 ;
      LAYER via ;
        RECT 2442.240 258.100 2442.500 258.360 ;
        RECT 2611.060 258.100 2611.320 258.360 ;
        RECT 2442.240 186.360 2442.500 186.620 ;
        RECT 2443.160 186.360 2443.420 186.620 ;
        RECT 2442.240 137.740 2442.500 138.000 ;
        RECT 2439.940 89.800 2440.200 90.060 ;
        RECT 2440.860 47.980 2441.120 48.240 ;
        RECT 2440.860 2.760 2441.120 3.020 ;
      LAYER met2 ;
        RECT 2611.050 633.915 2611.330 634.285 ;
        RECT 2611.120 258.390 2611.260 633.915 ;
        RECT 2442.240 258.070 2442.500 258.390 ;
        RECT 2611.060 258.070 2611.320 258.390 ;
        RECT 2442.300 234.445 2442.440 258.070 ;
        RECT 2442.230 234.075 2442.510 234.445 ;
        RECT 2443.150 234.075 2443.430 234.445 ;
        RECT 2443.220 186.650 2443.360 234.075 ;
        RECT 2442.240 186.330 2442.500 186.650 ;
        RECT 2443.160 186.330 2443.420 186.650 ;
        RECT 2442.300 138.030 2442.440 186.330 ;
        RECT 2442.240 137.710 2442.500 138.030 ;
        RECT 2439.940 89.770 2440.200 90.090 ;
        RECT 2440.000 48.805 2440.140 89.770 ;
        RECT 2439.930 48.435 2440.210 48.805 ;
        RECT 2440.850 48.435 2441.130 48.805 ;
        RECT 2440.920 48.270 2441.060 48.435 ;
        RECT 2440.860 47.950 2441.120 48.270 ;
        RECT 2440.860 2.730 2441.120 3.050 ;
        RECT 2440.920 2.400 2441.060 2.730 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
      LAYER via2 ;
        RECT 2611.050 633.960 2611.330 634.240 ;
        RECT 2442.230 234.120 2442.510 234.400 ;
        RECT 2443.150 234.120 2443.430 234.400 ;
        RECT 2439.930 48.480 2440.210 48.760 ;
        RECT 2440.850 48.480 2441.130 48.760 ;
      LAYER met3 ;
        RECT 2606.000 634.250 2610.000 634.640 ;
        RECT 2611.025 634.250 2611.355 634.265 ;
        RECT 2606.000 634.040 2611.355 634.250 ;
        RECT 2609.580 633.950 2611.355 634.040 ;
        RECT 2611.025 633.935 2611.355 633.950 ;
        RECT 2442.205 234.410 2442.535 234.425 ;
        RECT 2443.125 234.410 2443.455 234.425 ;
        RECT 2442.205 234.110 2443.455 234.410 ;
        RECT 2442.205 234.095 2442.535 234.110 ;
        RECT 2443.125 234.095 2443.455 234.110 ;
        RECT 2439.905 48.770 2440.235 48.785 ;
        RECT 2440.825 48.770 2441.155 48.785 ;
        RECT 2439.905 48.470 2441.155 48.770 ;
        RECT 2439.905 48.455 2440.235 48.470 ;
        RECT 2440.825 48.455 2441.155 48.470 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.050 162.080 627.370 162.140 ;
        RECT 2456.930 162.080 2457.250 162.140 ;
        RECT 627.050 161.940 2457.250 162.080 ;
        RECT 627.050 161.880 627.370 161.940 ;
        RECT 2456.930 161.880 2457.250 161.940 ;
        RECT 2456.930 14.180 2457.250 14.240 ;
        RECT 2456.930 14.040 2459.000 14.180 ;
        RECT 2456.930 13.980 2457.250 14.040 ;
        RECT 2458.860 13.900 2459.000 14.040 ;
        RECT 2458.770 13.640 2459.090 13.900 ;
      LAYER via ;
        RECT 627.080 161.880 627.340 162.140 ;
        RECT 2456.960 161.880 2457.220 162.140 ;
        RECT 2456.960 13.980 2457.220 14.240 ;
        RECT 2458.800 13.640 2459.060 13.900 ;
      LAYER met2 ;
        RECT 626.570 260.170 626.850 264.000 ;
        RECT 626.570 260.030 627.280 260.170 ;
        RECT 626.570 260.000 626.850 260.030 ;
        RECT 627.140 162.170 627.280 260.030 ;
        RECT 627.080 161.850 627.340 162.170 ;
        RECT 2456.960 161.850 2457.220 162.170 ;
        RECT 2457.020 14.270 2457.160 161.850 ;
        RECT 2456.960 13.950 2457.220 14.270 ;
        RECT 2458.800 13.610 2459.060 13.930 ;
        RECT 2458.860 2.400 2459.000 13.610 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 441.210 127.740 441.530 127.800 ;
        RECT 2470.270 127.740 2470.590 127.800 ;
        RECT 441.210 127.600 2470.590 127.740 ;
        RECT 441.210 127.540 441.530 127.600 ;
        RECT 2470.270 127.540 2470.590 127.600 ;
        RECT 2470.270 37.640 2470.590 37.700 ;
        RECT 2476.710 37.640 2477.030 37.700 ;
        RECT 2470.270 37.500 2477.030 37.640 ;
        RECT 2470.270 37.440 2470.590 37.500 ;
        RECT 2476.710 37.440 2477.030 37.500 ;
      LAYER via ;
        RECT 441.240 127.540 441.500 127.800 ;
        RECT 2470.300 127.540 2470.560 127.800 ;
        RECT 2470.300 37.440 2470.560 37.700 ;
        RECT 2476.740 37.440 2477.000 37.700 ;
      LAYER met2 ;
        RECT 440.730 260.170 441.010 264.000 ;
        RECT 440.730 260.030 441.440 260.170 ;
        RECT 440.730 260.000 441.010 260.030 ;
        RECT 441.300 127.830 441.440 260.030 ;
        RECT 441.240 127.510 441.500 127.830 ;
        RECT 2470.300 127.510 2470.560 127.830 ;
        RECT 2470.360 37.730 2470.500 127.510 ;
        RECT 2470.300 37.410 2470.560 37.730 ;
        RECT 2476.740 37.410 2477.000 37.730 ;
        RECT 2476.800 2.400 2476.940 37.410 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1856.300 2615.490 1856.360 ;
        RECT 2666.230 1856.300 2666.550 1856.360 ;
        RECT 2615.170 1856.160 2666.550 1856.300 ;
        RECT 2615.170 1856.100 2615.490 1856.160 ;
        RECT 2666.230 1856.100 2666.550 1856.160 ;
        RECT 2497.410 244.360 2497.730 244.420 ;
        RECT 2666.230 244.360 2666.550 244.420 ;
        RECT 2497.410 244.220 2666.550 244.360 ;
        RECT 2497.410 244.160 2497.730 244.220 ;
        RECT 2666.230 244.160 2666.550 244.220 ;
        RECT 2494.650 20.640 2494.970 20.700 ;
        RECT 2497.410 20.640 2497.730 20.700 ;
        RECT 2494.650 20.500 2497.730 20.640 ;
        RECT 2494.650 20.440 2494.970 20.500 ;
        RECT 2497.410 20.440 2497.730 20.500 ;
      LAYER via ;
        RECT 2615.200 1856.100 2615.460 1856.360 ;
        RECT 2666.260 1856.100 2666.520 1856.360 ;
        RECT 2497.440 244.160 2497.700 244.420 ;
        RECT 2666.260 244.160 2666.520 244.420 ;
        RECT 2494.680 20.440 2494.940 20.700 ;
        RECT 2497.440 20.440 2497.700 20.700 ;
      LAYER met2 ;
        RECT 2615.190 1860.635 2615.470 1861.005 ;
        RECT 2615.260 1856.390 2615.400 1860.635 ;
        RECT 2615.200 1856.070 2615.460 1856.390 ;
        RECT 2666.260 1856.070 2666.520 1856.390 ;
        RECT 2666.320 244.450 2666.460 1856.070 ;
        RECT 2497.440 244.130 2497.700 244.450 ;
        RECT 2666.260 244.130 2666.520 244.450 ;
        RECT 2497.500 20.730 2497.640 244.130 ;
        RECT 2494.680 20.410 2494.940 20.730 ;
        RECT 2497.440 20.410 2497.700 20.730 ;
        RECT 2494.740 2.400 2494.880 20.410 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1860.680 2615.470 1860.960 ;
      LAYER met3 ;
        RECT 2606.000 1860.970 2610.000 1861.360 ;
        RECT 2615.165 1860.970 2615.495 1860.985 ;
        RECT 2606.000 1860.760 2615.495 1860.970 ;
        RECT 2609.580 1860.670 2615.495 1860.760 ;
        RECT 2615.165 1860.655 2615.495 1860.670 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2512.205 48.365 2512.375 96.475 ;
      LAYER mcon ;
        RECT 2512.205 96.305 2512.375 96.475 ;
      LAYER met1 ;
        RECT 311.950 113.800 312.270 113.860 ;
        RECT 2511.670 113.800 2511.990 113.860 ;
        RECT 311.950 113.660 2511.990 113.800 ;
        RECT 311.950 113.600 312.270 113.660 ;
        RECT 2511.670 113.600 2511.990 113.660 ;
        RECT 2511.670 96.460 2511.990 96.520 ;
        RECT 2512.145 96.460 2512.435 96.505 ;
        RECT 2511.670 96.320 2512.435 96.460 ;
        RECT 2511.670 96.260 2511.990 96.320 ;
        RECT 2512.145 96.275 2512.435 96.320 ;
        RECT 2511.670 48.520 2511.990 48.580 ;
        RECT 2512.145 48.520 2512.435 48.565 ;
        RECT 2511.670 48.380 2512.435 48.520 ;
        RECT 2511.670 48.320 2511.990 48.380 ;
        RECT 2512.145 48.335 2512.435 48.380 ;
        RECT 2511.670 14.180 2511.990 14.240 ;
        RECT 2511.670 14.040 2512.360 14.180 ;
        RECT 2511.670 13.980 2511.990 14.040 ;
        RECT 2512.220 13.900 2512.360 14.040 ;
        RECT 2512.130 13.640 2512.450 13.900 ;
      LAYER via ;
        RECT 311.980 113.600 312.240 113.860 ;
        RECT 2511.700 113.600 2511.960 113.860 ;
        RECT 2511.700 96.260 2511.960 96.520 ;
        RECT 2511.700 48.320 2511.960 48.580 ;
        RECT 2511.700 13.980 2511.960 14.240 ;
        RECT 2512.160 13.640 2512.420 13.900 ;
      LAYER met2 ;
        RECT 311.970 662.475 312.250 662.845 ;
        RECT 312.040 113.890 312.180 662.475 ;
        RECT 311.980 113.570 312.240 113.890 ;
        RECT 2511.700 113.570 2511.960 113.890 ;
        RECT 2511.760 96.550 2511.900 113.570 ;
        RECT 2511.700 96.230 2511.960 96.550 ;
        RECT 2511.700 48.290 2511.960 48.610 ;
        RECT 2511.760 14.270 2511.900 48.290 ;
        RECT 2511.700 13.950 2511.960 14.270 ;
        RECT 2512.160 13.610 2512.420 13.930 ;
        RECT 2512.220 2.400 2512.360 13.610 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
      LAYER via2 ;
        RECT 311.970 662.520 312.250 662.800 ;
      LAYER met3 ;
        RECT 310.000 665.320 314.000 665.920 ;
        RECT 312.190 662.825 312.490 665.320 ;
        RECT 311.945 662.510 312.490 662.825 ;
        RECT 311.945 662.495 312.275 662.510 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1113.270 244.020 1113.590 244.080 ;
        RECT 1117.410 244.020 1117.730 244.080 ;
        RECT 1113.270 243.880 1117.730 244.020 ;
        RECT 1113.270 243.820 1113.590 243.880 ;
        RECT 1117.410 243.820 1117.730 243.880 ;
        RECT 1117.410 94.080 1117.730 94.140 ;
        RECT 2525.930 94.080 2526.250 94.140 ;
        RECT 1117.410 93.940 2526.250 94.080 ;
        RECT 1117.410 93.880 1117.730 93.940 ;
        RECT 2525.930 93.880 2526.250 93.940 ;
        RECT 2525.930 14.180 2526.250 14.240 ;
        RECT 2525.930 14.040 2530.300 14.180 ;
        RECT 2525.930 13.980 2526.250 14.040 ;
        RECT 2530.160 13.900 2530.300 14.040 ;
        RECT 2530.070 13.640 2530.390 13.900 ;
      LAYER via ;
        RECT 1113.300 243.820 1113.560 244.080 ;
        RECT 1117.440 243.820 1117.700 244.080 ;
        RECT 1117.440 93.880 1117.700 94.140 ;
        RECT 2525.960 93.880 2526.220 94.140 ;
        RECT 2525.960 13.980 2526.220 14.240 ;
        RECT 2530.100 13.640 2530.360 13.900 ;
      LAYER met2 ;
        RECT 1113.250 260.000 1113.530 264.000 ;
        RECT 1113.360 244.110 1113.500 260.000 ;
        RECT 1113.300 243.790 1113.560 244.110 ;
        RECT 1117.440 243.790 1117.700 244.110 ;
        RECT 1117.500 94.170 1117.640 243.790 ;
        RECT 1117.440 93.850 1117.700 94.170 ;
        RECT 2525.960 93.850 2526.220 94.170 ;
        RECT 2526.020 14.270 2526.160 93.850 ;
        RECT 2525.960 13.950 2526.220 14.270 ;
        RECT 2530.100 13.610 2530.360 13.930 ;
        RECT 2530.160 2.400 2530.300 13.610 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 225.470 2608.380 225.790 2608.440 ;
        RECT 296.770 2608.380 297.090 2608.440 ;
        RECT 225.470 2608.240 297.090 2608.380 ;
        RECT 225.470 2608.180 225.790 2608.240 ;
        RECT 296.770 2608.180 297.090 2608.240 ;
      LAYER via ;
        RECT 225.500 2608.180 225.760 2608.440 ;
        RECT 296.800 2608.180 297.060 2608.440 ;
      LAYER met2 ;
        RECT 296.790 2609.995 297.070 2610.365 ;
        RECT 296.860 2608.470 297.000 2609.995 ;
        RECT 225.500 2608.150 225.760 2608.470 ;
        RECT 296.800 2608.150 297.060 2608.470 ;
        RECT 225.560 45.405 225.700 2608.150 ;
        RECT 225.490 45.035 225.770 45.405 ;
        RECT 2548.030 45.035 2548.310 45.405 ;
        RECT 2548.100 2.400 2548.240 45.035 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
      LAYER via2 ;
        RECT 296.790 2610.040 297.070 2610.320 ;
        RECT 225.490 45.080 225.770 45.360 ;
        RECT 2548.030 45.080 2548.310 45.360 ;
      LAYER met3 ;
        RECT 296.765 2610.330 297.095 2610.345 ;
        RECT 310.000 2610.330 314.000 2610.720 ;
        RECT 296.765 2610.120 314.000 2610.330 ;
        RECT 296.765 2610.030 310.500 2610.120 ;
        RECT 296.765 2610.015 297.095 2610.030 ;
        RECT 225.465 45.370 225.795 45.385 ;
        RECT 2548.005 45.370 2548.335 45.385 ;
        RECT 225.465 45.070 2548.335 45.370 ;
        RECT 225.465 45.055 225.795 45.070 ;
        RECT 2548.005 45.055 2548.335 45.070 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 225.010 2525.760 225.330 2525.820 ;
        RECT 296.770 2525.760 297.090 2525.820 ;
        RECT 225.010 2525.620 297.090 2525.760 ;
        RECT 225.010 2525.560 225.330 2525.620 ;
        RECT 296.770 2525.560 297.090 2525.620 ;
      LAYER via ;
        RECT 225.040 2525.560 225.300 2525.820 ;
        RECT 296.800 2525.560 297.060 2525.820 ;
      LAYER met2 ;
        RECT 225.040 2525.530 225.300 2525.850 ;
        RECT 296.790 2525.675 297.070 2526.045 ;
        RECT 296.800 2525.530 297.060 2525.675 ;
        RECT 225.100 44.725 225.240 2525.530 ;
        RECT 225.030 44.355 225.310 44.725 ;
        RECT 2565.970 44.355 2566.250 44.725 ;
        RECT 2566.040 2.400 2566.180 44.355 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
      LAYER via2 ;
        RECT 296.790 2525.720 297.070 2526.000 ;
        RECT 225.030 44.400 225.310 44.680 ;
        RECT 2565.970 44.400 2566.250 44.680 ;
      LAYER met3 ;
        RECT 296.765 2526.010 297.095 2526.025 ;
        RECT 310.000 2526.010 314.000 2526.400 ;
        RECT 296.765 2525.800 314.000 2526.010 ;
        RECT 296.765 2525.710 310.500 2525.800 ;
        RECT 296.765 2525.695 297.095 2525.710 ;
        RECT 225.005 44.690 225.335 44.705 ;
        RECT 2565.945 44.690 2566.275 44.705 ;
        RECT 225.005 44.390 2566.275 44.690 ;
        RECT 225.005 44.375 225.335 44.390 ;
        RECT 2565.945 44.375 2566.275 44.390 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2580.690 140.915 2580.970 141.285 ;
        RECT 2580.760 3.130 2580.900 140.915 ;
        RECT 2580.760 2.990 2583.660 3.130 ;
        RECT 2583.520 2.960 2583.660 2.990 ;
        RECT 2583.520 2.820 2584.120 2.960 ;
        RECT 2583.980 2.400 2584.120 2.820 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
      LAYER via2 ;
        RECT 2580.690 140.960 2580.970 141.240 ;
      LAYER met3 ;
        RECT 290.990 2440.330 291.370 2440.340 ;
        RECT 310.000 2440.330 314.000 2440.720 ;
        RECT 290.990 2440.120 314.000 2440.330 ;
        RECT 290.990 2440.030 310.500 2440.120 ;
        RECT 290.990 2440.020 291.370 2440.030 ;
        RECT 290.990 141.250 291.370 141.260 ;
        RECT 2580.665 141.250 2580.995 141.265 ;
        RECT 290.990 140.950 2580.995 141.250 ;
        RECT 290.990 140.940 291.370 140.950 ;
        RECT 2580.665 140.935 2580.995 140.950 ;
      LAYER via3 ;
        RECT 291.020 2440.020 291.340 2440.340 ;
        RECT 291.020 140.940 291.340 141.260 ;
      LAYER met4 ;
        RECT 291.015 2440.015 291.345 2440.345 ;
        RECT 291.030 141.265 291.330 2440.015 ;
        RECT 291.015 140.935 291.345 141.265 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 20.640 817.810 20.700 ;
        RECT 820.710 20.640 821.030 20.700 ;
        RECT 817.490 20.500 821.030 20.640 ;
        RECT 817.490 20.440 817.810 20.500 ;
        RECT 820.710 20.440 821.030 20.500 ;
      LAYER via ;
        RECT 817.520 20.440 817.780 20.700 ;
        RECT 820.740 20.440 821.000 20.700 ;
      LAYER met2 ;
        RECT 2378.250 3257.610 2378.530 3260.000 ;
        RECT 2379.670 3257.610 2379.950 3257.725 ;
        RECT 2378.250 3257.470 2379.950 3257.610 ;
        RECT 2378.250 3256.000 2378.530 3257.470 ;
        RECT 2379.670 3257.355 2379.950 3257.470 ;
        RECT 820.730 259.235 821.010 259.605 ;
        RECT 820.800 20.730 820.940 259.235 ;
        RECT 817.520 20.410 817.780 20.730 ;
        RECT 820.740 20.410 821.000 20.730 ;
        RECT 817.580 2.400 817.720 20.410 ;
        RECT 817.370 -4.800 817.930 2.400 ;
      LAYER via2 ;
        RECT 2379.670 3257.400 2379.950 3257.680 ;
        RECT 820.730 259.280 821.010 259.560 ;
      LAYER met3 ;
        RECT 2379.645 3257.690 2379.975 3257.705 ;
        RECT 2656.310 3257.690 2656.690 3257.700 ;
        RECT 2379.645 3257.390 2656.690 3257.690 ;
        RECT 2379.645 3257.375 2379.975 3257.390 ;
        RECT 2656.310 3257.380 2656.690 3257.390 ;
        RECT 2656.310 1641.330 2656.690 1641.340 ;
        RECT 2659.070 1641.330 2659.450 1641.340 ;
        RECT 2656.310 1641.030 2659.450 1641.330 ;
        RECT 2656.310 1641.020 2656.690 1641.030 ;
        RECT 2659.070 1641.020 2659.450 1641.030 ;
        RECT 2656.310 1595.770 2656.690 1595.780 ;
        RECT 2659.070 1595.770 2659.450 1595.780 ;
        RECT 2656.310 1595.470 2659.450 1595.770 ;
        RECT 2656.310 1595.460 2656.690 1595.470 ;
        RECT 2659.070 1595.460 2659.450 1595.470 ;
        RECT 820.705 259.570 821.035 259.585 ;
        RECT 2656.310 259.570 2656.690 259.580 ;
        RECT 820.705 259.270 2656.690 259.570 ;
        RECT 820.705 259.255 821.035 259.270 ;
        RECT 2656.310 259.260 2656.690 259.270 ;
      LAYER via3 ;
        RECT 2656.340 3257.380 2656.660 3257.700 ;
        RECT 2656.340 1641.020 2656.660 1641.340 ;
        RECT 2659.100 1641.020 2659.420 1641.340 ;
        RECT 2656.340 1595.460 2656.660 1595.780 ;
        RECT 2659.100 1595.460 2659.420 1595.780 ;
        RECT 2656.340 259.260 2656.660 259.580 ;
      LAYER met4 ;
        RECT 2656.335 3257.375 2656.665 3257.705 ;
        RECT 2656.350 1641.345 2656.650 3257.375 ;
        RECT 2656.335 1641.015 2656.665 1641.345 ;
        RECT 2659.095 1641.015 2659.425 1641.345 ;
        RECT 2659.110 1595.785 2659.410 1641.015 ;
        RECT 2656.335 1595.455 2656.665 1595.785 ;
        RECT 2659.095 1595.455 2659.425 1595.785 ;
        RECT 2656.350 259.585 2656.650 1595.455 ;
        RECT 2656.335 259.255 2656.665 259.585 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1613.290 86.600 1613.610 86.660 ;
        RECT 2601.370 86.600 2601.690 86.660 ;
        RECT 1613.290 86.460 2601.690 86.600 ;
        RECT 1613.290 86.400 1613.610 86.460 ;
        RECT 2601.370 86.400 2601.690 86.460 ;
      LAYER via ;
        RECT 1613.320 86.400 1613.580 86.660 ;
        RECT 2601.400 86.400 2601.660 86.660 ;
      LAYER met2 ;
        RECT 1613.730 260.170 1614.010 264.000 ;
        RECT 1613.380 260.030 1614.010 260.170 ;
        RECT 1613.380 86.690 1613.520 260.030 ;
        RECT 1613.730 260.000 1614.010 260.030 ;
        RECT 1613.320 86.370 1613.580 86.690 ;
        RECT 2601.400 86.370 2601.660 86.690 ;
        RECT 2601.460 2.400 2601.600 86.370 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2.960 2615.490 3.020 ;
        RECT 2619.310 2.960 2619.630 3.020 ;
        RECT 2615.170 2.820 2619.630 2.960 ;
        RECT 2615.170 2.760 2615.490 2.820 ;
        RECT 2619.310 2.760 2619.630 2.820 ;
      LAYER via ;
        RECT 2615.200 2.760 2615.460 3.020 ;
        RECT 2619.340 2.760 2619.600 3.020 ;
      LAYER met2 ;
        RECT 2615.190 72.235 2615.470 72.605 ;
        RECT 2615.260 3.050 2615.400 72.235 ;
        RECT 2615.200 2.730 2615.460 3.050 ;
        RECT 2619.340 2.730 2619.600 3.050 ;
        RECT 2619.400 2.400 2619.540 2.730 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
      LAYER via2 ;
        RECT 2615.190 72.280 2615.470 72.560 ;
      LAYER met3 ;
        RECT 295.590 3011.530 295.970 3011.540 ;
        RECT 310.000 3011.530 314.000 3011.920 ;
        RECT 295.590 3011.320 314.000 3011.530 ;
        RECT 295.590 3011.230 310.500 3011.320 ;
        RECT 295.590 3011.220 295.970 3011.230 ;
        RECT 295.590 72.570 295.970 72.580 ;
        RECT 2615.165 72.570 2615.495 72.585 ;
        RECT 295.590 72.270 2615.495 72.570 ;
        RECT 295.590 72.260 295.970 72.270 ;
        RECT 2615.165 72.255 2615.495 72.270 ;
      LAYER via3 ;
        RECT 295.620 3011.220 295.940 3011.540 ;
        RECT 295.620 72.260 295.940 72.580 ;
      LAYER met4 ;
        RECT 295.615 3011.215 295.945 3011.545 ;
        RECT 295.630 72.585 295.930 3011.215 ;
        RECT 295.615 72.255 295.945 72.585 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1827.650 121.280 1827.970 121.340 ;
        RECT 2636.790 121.280 2637.110 121.340 ;
        RECT 1827.650 121.140 2637.110 121.280 ;
        RECT 1827.650 121.080 1827.970 121.140 ;
        RECT 2636.790 121.080 2637.110 121.140 ;
      LAYER via ;
        RECT 1827.680 121.080 1827.940 121.340 ;
        RECT 2636.820 121.080 2637.080 121.340 ;
      LAYER met2 ;
        RECT 1828.090 260.170 1828.370 264.000 ;
        RECT 1827.740 260.030 1828.370 260.170 ;
        RECT 1827.740 121.370 1827.880 260.030 ;
        RECT 1828.090 260.000 1828.370 260.030 ;
        RECT 1827.680 121.050 1827.940 121.370 ;
        RECT 2636.820 121.050 2637.080 121.370 ;
        RECT 2636.880 3.130 2637.020 121.050 ;
        RECT 2636.880 2.990 2637.480 3.130 ;
        RECT 2637.340 2.400 2637.480 2.990 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.930 189.620 295.250 189.680 ;
        RECT 2651.050 189.620 2651.370 189.680 ;
        RECT 294.930 189.480 2651.370 189.620 ;
        RECT 294.930 189.420 295.250 189.480 ;
        RECT 2651.050 189.420 2651.370 189.480 ;
        RECT 2650.590 2.960 2650.910 3.020 ;
        RECT 2655.190 2.960 2655.510 3.020 ;
        RECT 2650.590 2.820 2655.510 2.960 ;
        RECT 2650.590 2.760 2650.910 2.820 ;
        RECT 2655.190 2.760 2655.510 2.820 ;
      LAYER via ;
        RECT 294.960 189.420 295.220 189.680 ;
        RECT 2651.080 189.420 2651.340 189.680 ;
        RECT 2650.620 2.760 2650.880 3.020 ;
        RECT 2655.220 2.760 2655.480 3.020 ;
      LAYER met2 ;
        RECT 294.950 1890.555 295.230 1890.925 ;
        RECT 295.020 189.710 295.160 1890.555 ;
        RECT 294.960 189.390 295.220 189.710 ;
        RECT 2651.080 189.390 2651.340 189.710 ;
        RECT 2651.140 14.690 2651.280 189.390 ;
        RECT 2650.680 14.550 2651.280 14.690 ;
        RECT 2650.680 3.050 2650.820 14.550 ;
        RECT 2650.620 2.730 2650.880 3.050 ;
        RECT 2655.220 2.730 2655.480 3.050 ;
        RECT 2655.280 2.400 2655.420 2.730 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
      LAYER via2 ;
        RECT 294.950 1890.600 295.230 1890.880 ;
      LAYER met3 ;
        RECT 294.925 1890.890 295.255 1890.905 ;
        RECT 310.000 1890.890 314.000 1891.280 ;
        RECT 294.925 1890.680 314.000 1890.890 ;
        RECT 294.925 1890.590 310.500 1890.680 ;
        RECT 294.925 1890.575 295.255 1890.590 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2263.270 3260.500 2263.590 3260.560 ;
        RECT 2670.370 3260.500 2670.690 3260.560 ;
        RECT 2263.270 3260.360 2670.690 3260.500 ;
        RECT 2263.270 3260.300 2263.590 3260.360 ;
        RECT 2670.370 3260.300 2670.690 3260.360 ;
      LAYER via ;
        RECT 2263.300 3260.300 2263.560 3260.560 ;
        RECT 2670.400 3260.300 2670.660 3260.560 ;
      LAYER met2 ;
        RECT 2263.300 3260.270 2263.560 3260.590 ;
        RECT 2670.400 3260.270 2670.660 3260.590 ;
        RECT 2263.360 3260.000 2263.500 3260.270 ;
        RECT 2263.250 3256.000 2263.530 3260.000 ;
        RECT 2670.460 20.130 2670.600 3260.270 ;
        RECT 2670.460 19.990 2672.900 20.130 ;
        RECT 2672.760 2.400 2672.900 19.990 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2688.845 3091.365 2689.015 3139.475 ;
        RECT 2688.845 2994.805 2689.015 3042.915 ;
        RECT 2688.845 2898.245 2689.015 2946.355 ;
        RECT 2690.685 2.805 2690.855 14.195 ;
      LAYER mcon ;
        RECT 2688.845 3139.305 2689.015 3139.475 ;
        RECT 2688.845 3042.745 2689.015 3042.915 ;
        RECT 2688.845 2946.185 2689.015 2946.355 ;
        RECT 2690.685 14.025 2690.855 14.195 ;
      LAYER met1 ;
        RECT 2688.310 3188.220 2688.630 3188.480 ;
        RECT 2615.170 3188.080 2615.490 3188.140 ;
        RECT 2688.400 3188.080 2688.540 3188.220 ;
        RECT 2615.170 3187.940 2688.540 3188.080 ;
        RECT 2615.170 3187.880 2615.490 3187.940 ;
        RECT 2688.770 3139.460 2689.090 3139.520 ;
        RECT 2688.575 3139.320 2689.090 3139.460 ;
        RECT 2688.770 3139.260 2689.090 3139.320 ;
        RECT 2688.770 3091.520 2689.090 3091.580 ;
        RECT 2688.575 3091.380 2689.090 3091.520 ;
        RECT 2688.770 3091.320 2689.090 3091.380 ;
        RECT 2688.770 3042.900 2689.090 3042.960 ;
        RECT 2688.575 3042.760 2689.090 3042.900 ;
        RECT 2688.770 3042.700 2689.090 3042.760 ;
        RECT 2688.770 2994.960 2689.090 2995.020 ;
        RECT 2688.575 2994.820 2689.090 2994.960 ;
        RECT 2688.770 2994.760 2689.090 2994.820 ;
        RECT 2688.770 2946.340 2689.090 2946.400 ;
        RECT 2688.575 2946.200 2689.090 2946.340 ;
        RECT 2688.770 2946.140 2689.090 2946.200 ;
        RECT 2688.770 2898.400 2689.090 2898.460 ;
        RECT 2688.575 2898.260 2689.090 2898.400 ;
        RECT 2688.770 2898.200 2689.090 2898.260 ;
        RECT 2688.770 2801.500 2689.090 2801.560 ;
        RECT 2689.690 2801.500 2690.010 2801.560 ;
        RECT 2688.770 2801.360 2690.010 2801.500 ;
        RECT 2688.770 2801.300 2689.090 2801.360 ;
        RECT 2689.690 2801.300 2690.010 2801.360 ;
        RECT 2688.770 2704.940 2689.090 2705.000 ;
        RECT 2689.690 2704.940 2690.010 2705.000 ;
        RECT 2688.770 2704.800 2690.010 2704.940 ;
        RECT 2688.770 2704.740 2689.090 2704.800 ;
        RECT 2689.690 2704.740 2690.010 2704.800 ;
        RECT 2688.770 2608.380 2689.090 2608.440 ;
        RECT 2689.690 2608.380 2690.010 2608.440 ;
        RECT 2688.770 2608.240 2690.010 2608.380 ;
        RECT 2688.770 2608.180 2689.090 2608.240 ;
        RECT 2689.690 2608.180 2690.010 2608.240 ;
        RECT 2688.770 2511.820 2689.090 2511.880 ;
        RECT 2689.690 2511.820 2690.010 2511.880 ;
        RECT 2688.770 2511.680 2690.010 2511.820 ;
        RECT 2688.770 2511.620 2689.090 2511.680 ;
        RECT 2689.690 2511.620 2690.010 2511.680 ;
        RECT 2688.770 2463.200 2689.090 2463.260 ;
        RECT 2689.690 2463.200 2690.010 2463.260 ;
        RECT 2688.770 2463.060 2690.010 2463.200 ;
        RECT 2688.770 2463.000 2689.090 2463.060 ;
        RECT 2689.690 2463.000 2690.010 2463.060 ;
        RECT 2688.770 14.180 2689.090 14.240 ;
        RECT 2690.625 14.180 2690.915 14.225 ;
        RECT 2688.770 14.040 2690.915 14.180 ;
        RECT 2688.770 13.980 2689.090 14.040 ;
        RECT 2690.625 13.995 2690.915 14.040 ;
        RECT 2690.610 2.960 2690.930 3.020 ;
        RECT 2690.415 2.820 2690.930 2.960 ;
        RECT 2690.610 2.760 2690.930 2.820 ;
      LAYER via ;
        RECT 2688.340 3188.220 2688.600 3188.480 ;
        RECT 2615.200 3187.880 2615.460 3188.140 ;
        RECT 2688.800 3139.260 2689.060 3139.520 ;
        RECT 2688.800 3091.320 2689.060 3091.580 ;
        RECT 2688.800 3042.700 2689.060 3042.960 ;
        RECT 2688.800 2994.760 2689.060 2995.020 ;
        RECT 2688.800 2946.140 2689.060 2946.400 ;
        RECT 2688.800 2898.200 2689.060 2898.460 ;
        RECT 2688.800 2801.300 2689.060 2801.560 ;
        RECT 2689.720 2801.300 2689.980 2801.560 ;
        RECT 2688.800 2704.740 2689.060 2705.000 ;
        RECT 2689.720 2704.740 2689.980 2705.000 ;
        RECT 2688.800 2608.180 2689.060 2608.440 ;
        RECT 2689.720 2608.180 2689.980 2608.440 ;
        RECT 2688.800 2511.620 2689.060 2511.880 ;
        RECT 2689.720 2511.620 2689.980 2511.880 ;
        RECT 2688.800 2463.000 2689.060 2463.260 ;
        RECT 2689.720 2463.000 2689.980 2463.260 ;
        RECT 2688.800 13.980 2689.060 14.240 ;
        RECT 2690.640 2.760 2690.900 3.020 ;
      LAYER met2 ;
        RECT 2615.190 3192.075 2615.470 3192.445 ;
        RECT 2615.260 3188.170 2615.400 3192.075 ;
        RECT 2688.340 3188.250 2688.600 3188.510 ;
        RECT 2688.340 3188.190 2689.000 3188.250 ;
        RECT 2615.200 3187.850 2615.460 3188.170 ;
        RECT 2688.400 3188.110 2689.000 3188.190 ;
        RECT 2688.860 3139.550 2689.000 3188.110 ;
        RECT 2688.800 3139.230 2689.060 3139.550 ;
        RECT 2688.800 3091.290 2689.060 3091.610 ;
        RECT 2688.860 3042.990 2689.000 3091.290 ;
        RECT 2688.800 3042.670 2689.060 3042.990 ;
        RECT 2688.800 2994.730 2689.060 2995.050 ;
        RECT 2688.860 2946.430 2689.000 2994.730 ;
        RECT 2688.800 2946.110 2689.060 2946.430 ;
        RECT 2688.800 2898.170 2689.060 2898.490 ;
        RECT 2688.860 2849.725 2689.000 2898.170 ;
        RECT 2688.790 2849.355 2689.070 2849.725 ;
        RECT 2689.710 2849.355 2689.990 2849.725 ;
        RECT 2689.780 2801.590 2689.920 2849.355 ;
        RECT 2688.800 2801.270 2689.060 2801.590 ;
        RECT 2689.720 2801.270 2689.980 2801.590 ;
        RECT 2688.860 2753.165 2689.000 2801.270 ;
        RECT 2688.790 2752.795 2689.070 2753.165 ;
        RECT 2689.710 2752.795 2689.990 2753.165 ;
        RECT 2689.780 2705.030 2689.920 2752.795 ;
        RECT 2688.800 2704.710 2689.060 2705.030 ;
        RECT 2689.720 2704.710 2689.980 2705.030 ;
        RECT 2688.860 2656.605 2689.000 2704.710 ;
        RECT 2688.790 2656.235 2689.070 2656.605 ;
        RECT 2689.710 2656.235 2689.990 2656.605 ;
        RECT 2689.780 2608.470 2689.920 2656.235 ;
        RECT 2688.800 2608.150 2689.060 2608.470 ;
        RECT 2689.720 2608.150 2689.980 2608.470 ;
        RECT 2688.860 2560.045 2689.000 2608.150 ;
        RECT 2688.790 2559.675 2689.070 2560.045 ;
        RECT 2689.710 2559.675 2689.990 2560.045 ;
        RECT 2689.780 2511.910 2689.920 2559.675 ;
        RECT 2688.800 2511.590 2689.060 2511.910 ;
        RECT 2689.720 2511.590 2689.980 2511.910 ;
        RECT 2688.860 2463.290 2689.000 2511.590 ;
        RECT 2688.800 2462.970 2689.060 2463.290 ;
        RECT 2689.720 2462.970 2689.980 2463.290 ;
        RECT 2689.780 2415.205 2689.920 2462.970 ;
        RECT 2688.790 2414.835 2689.070 2415.205 ;
        RECT 2689.710 2414.835 2689.990 2415.205 ;
        RECT 2688.860 14.270 2689.000 2414.835 ;
        RECT 2688.800 13.950 2689.060 14.270 ;
        RECT 2690.640 2.730 2690.900 3.050 ;
        RECT 2690.700 2.400 2690.840 2.730 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
      LAYER via2 ;
        RECT 2615.190 3192.120 2615.470 3192.400 ;
        RECT 2688.790 2849.400 2689.070 2849.680 ;
        RECT 2689.710 2849.400 2689.990 2849.680 ;
        RECT 2688.790 2752.840 2689.070 2753.120 ;
        RECT 2689.710 2752.840 2689.990 2753.120 ;
        RECT 2688.790 2656.280 2689.070 2656.560 ;
        RECT 2689.710 2656.280 2689.990 2656.560 ;
        RECT 2688.790 2559.720 2689.070 2560.000 ;
        RECT 2689.710 2559.720 2689.990 2560.000 ;
        RECT 2688.790 2414.880 2689.070 2415.160 ;
        RECT 2689.710 2414.880 2689.990 2415.160 ;
      LAYER met3 ;
        RECT 2606.000 3192.410 2610.000 3192.800 ;
        RECT 2615.165 3192.410 2615.495 3192.425 ;
        RECT 2606.000 3192.200 2615.495 3192.410 ;
        RECT 2609.580 3192.110 2615.495 3192.200 ;
        RECT 2615.165 3192.095 2615.495 3192.110 ;
        RECT 2688.765 2849.690 2689.095 2849.705 ;
        RECT 2689.685 2849.690 2690.015 2849.705 ;
        RECT 2688.765 2849.390 2690.015 2849.690 ;
        RECT 2688.765 2849.375 2689.095 2849.390 ;
        RECT 2689.685 2849.375 2690.015 2849.390 ;
        RECT 2688.765 2753.130 2689.095 2753.145 ;
        RECT 2689.685 2753.130 2690.015 2753.145 ;
        RECT 2688.765 2752.830 2690.015 2753.130 ;
        RECT 2688.765 2752.815 2689.095 2752.830 ;
        RECT 2689.685 2752.815 2690.015 2752.830 ;
        RECT 2688.765 2656.570 2689.095 2656.585 ;
        RECT 2689.685 2656.570 2690.015 2656.585 ;
        RECT 2688.765 2656.270 2690.015 2656.570 ;
        RECT 2688.765 2656.255 2689.095 2656.270 ;
        RECT 2689.685 2656.255 2690.015 2656.270 ;
        RECT 2688.765 2560.010 2689.095 2560.025 ;
        RECT 2689.685 2560.010 2690.015 2560.025 ;
        RECT 2688.765 2559.710 2690.015 2560.010 ;
        RECT 2688.765 2559.695 2689.095 2559.710 ;
        RECT 2689.685 2559.695 2690.015 2559.710 ;
        RECT 2688.765 2415.170 2689.095 2415.185 ;
        RECT 2689.685 2415.170 2690.015 2415.185 ;
        RECT 2688.765 2414.870 2690.015 2415.170 ;
        RECT 2688.765 2414.855 2689.095 2414.870 ;
        RECT 2689.685 2414.855 2690.015 2414.870 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2042.470 243.340 2042.790 243.400 ;
        RECT 2048.910 243.340 2049.230 243.400 ;
        RECT 2042.470 243.200 2049.230 243.340 ;
        RECT 2042.470 243.140 2042.790 243.200 ;
        RECT 2048.910 243.140 2049.230 243.200 ;
        RECT 2048.910 79.800 2049.230 79.860 ;
        RECT 2704.870 79.800 2705.190 79.860 ;
        RECT 2048.910 79.660 2705.190 79.800 ;
        RECT 2048.910 79.600 2049.230 79.660 ;
        RECT 2704.870 79.600 2705.190 79.660 ;
      LAYER via ;
        RECT 2042.500 243.140 2042.760 243.400 ;
        RECT 2048.940 243.140 2049.200 243.400 ;
        RECT 2048.940 79.600 2049.200 79.860 ;
        RECT 2704.900 79.600 2705.160 79.860 ;
      LAYER met2 ;
        RECT 2042.450 260.000 2042.730 264.000 ;
        RECT 2042.560 243.430 2042.700 260.000 ;
        RECT 2042.500 243.110 2042.760 243.430 ;
        RECT 2048.940 243.110 2049.200 243.430 ;
        RECT 2049.000 79.890 2049.140 243.110 ;
        RECT 2048.940 79.570 2049.200 79.890 ;
        RECT 2704.900 79.570 2705.160 79.890 ;
        RECT 2704.960 18.090 2705.100 79.570 ;
        RECT 2704.960 17.950 2708.780 18.090 ;
        RECT 2708.640 2.400 2708.780 17.950 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1497.600 2615.490 1497.660 ;
        RECT 2725.570 1497.600 2725.890 1497.660 ;
        RECT 2615.170 1497.460 2725.890 1497.600 ;
        RECT 2615.170 1497.400 2615.490 1497.460 ;
        RECT 2725.570 1497.400 2725.890 1497.460 ;
        RECT 2725.110 48.520 2725.430 48.580 ;
        RECT 2726.490 48.520 2726.810 48.580 ;
        RECT 2725.110 48.380 2726.810 48.520 ;
        RECT 2725.110 48.320 2725.430 48.380 ;
        RECT 2726.490 48.320 2726.810 48.380 ;
      LAYER via ;
        RECT 2615.200 1497.400 2615.460 1497.660 ;
        RECT 2725.600 1497.400 2725.860 1497.660 ;
        RECT 2725.140 48.320 2725.400 48.580 ;
        RECT 2726.520 48.320 2726.780 48.580 ;
      LAYER met2 ;
        RECT 2615.190 1500.235 2615.470 1500.605 ;
        RECT 2615.260 1497.690 2615.400 1500.235 ;
        RECT 2615.200 1497.370 2615.460 1497.690 ;
        RECT 2725.600 1497.370 2725.860 1497.690 ;
        RECT 2725.660 72.490 2725.800 1497.370 ;
        RECT 2725.200 72.350 2725.800 72.490 ;
        RECT 2725.200 48.610 2725.340 72.350 ;
        RECT 2725.140 48.290 2725.400 48.610 ;
        RECT 2726.520 48.290 2726.780 48.610 ;
        RECT 2726.580 2.400 2726.720 48.290 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1500.280 2615.470 1500.560 ;
      LAYER met3 ;
        RECT 2606.000 1500.570 2610.000 1500.960 ;
        RECT 2615.165 1500.570 2615.495 1500.585 ;
        RECT 2606.000 1500.360 2615.495 1500.570 ;
        RECT 2609.580 1500.270 2615.495 1500.360 ;
        RECT 2615.165 1500.255 2615.495 1500.270 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1835.560 2615.490 1835.620 ;
        RECT 2701.190 1835.560 2701.510 1835.620 ;
        RECT 2615.170 1835.420 2701.510 1835.560 ;
        RECT 2615.170 1835.360 2615.490 1835.420 ;
        RECT 2701.190 1835.360 2701.510 1835.420 ;
        RECT 2701.190 18.260 2701.510 18.320 ;
        RECT 2744.430 18.260 2744.750 18.320 ;
        RECT 2701.190 18.120 2744.750 18.260 ;
        RECT 2701.190 18.060 2701.510 18.120 ;
        RECT 2744.430 18.060 2744.750 18.120 ;
      LAYER via ;
        RECT 2615.200 1835.360 2615.460 1835.620 ;
        RECT 2701.220 1835.360 2701.480 1835.620 ;
        RECT 2701.220 18.060 2701.480 18.320 ;
        RECT 2744.460 18.060 2744.720 18.320 ;
      LAYER met2 ;
        RECT 2615.190 1838.875 2615.470 1839.245 ;
        RECT 2615.260 1835.650 2615.400 1838.875 ;
        RECT 2615.200 1835.330 2615.460 1835.650 ;
        RECT 2701.220 1835.330 2701.480 1835.650 ;
        RECT 2701.280 18.350 2701.420 1835.330 ;
        RECT 2701.220 18.030 2701.480 18.350 ;
        RECT 2744.460 18.030 2744.720 18.350 ;
        RECT 2744.520 2.400 2744.660 18.030 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1838.920 2615.470 1839.200 ;
      LAYER met3 ;
        RECT 2606.000 1839.210 2610.000 1839.600 ;
        RECT 2615.165 1839.210 2615.495 1839.225 ;
        RECT 2606.000 1839.000 2615.495 1839.210 ;
        RECT 2609.580 1838.910 2615.495 1839.000 ;
        RECT 2615.165 1838.895 2615.495 1838.910 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 304.590 231.100 304.910 231.160 ;
        RECT 2760.070 231.100 2760.390 231.160 ;
        RECT 304.590 230.960 2760.390 231.100 ;
        RECT 304.590 230.900 304.910 230.960 ;
        RECT 2760.070 230.900 2760.390 230.960 ;
        RECT 2759.610 48.520 2759.930 48.580 ;
        RECT 2761.910 48.520 2762.230 48.580 ;
        RECT 2759.610 48.380 2762.230 48.520 ;
        RECT 2759.610 48.320 2759.930 48.380 ;
        RECT 2761.910 48.320 2762.230 48.380 ;
      LAYER via ;
        RECT 304.620 230.900 304.880 231.160 ;
        RECT 2760.100 230.900 2760.360 231.160 ;
        RECT 2759.640 48.320 2759.900 48.580 ;
        RECT 2761.940 48.320 2762.200 48.580 ;
      LAYER met2 ;
        RECT 304.610 474.795 304.890 475.165 ;
        RECT 304.680 231.190 304.820 474.795 ;
        RECT 304.620 230.870 304.880 231.190 ;
        RECT 2760.100 230.870 2760.360 231.190 ;
        RECT 2760.160 72.490 2760.300 230.870 ;
        RECT 2759.700 72.350 2760.300 72.490 ;
        RECT 2759.700 48.610 2759.840 72.350 ;
        RECT 2759.640 48.290 2759.900 48.610 ;
        RECT 2761.940 48.290 2762.200 48.610 ;
        RECT 2762.000 2.400 2762.140 48.290 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
      LAYER via2 ;
        RECT 304.610 474.840 304.890 475.120 ;
      LAYER met3 ;
        RECT 304.585 475.130 304.915 475.145 ;
        RECT 310.000 475.130 314.000 475.520 ;
        RECT 304.585 474.920 314.000 475.130 ;
        RECT 304.585 474.830 310.500 474.920 ;
        RECT 304.585 474.815 304.915 474.830 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 835.045 48.365 835.215 96.475 ;
      LAYER mcon ;
        RECT 835.045 96.305 835.215 96.475 ;
      LAYER met1 ;
        RECT 296.310 252.860 296.630 252.920 ;
        RECT 834.970 252.860 835.290 252.920 ;
        RECT 296.310 252.720 835.290 252.860 ;
        RECT 296.310 252.660 296.630 252.720 ;
        RECT 834.970 252.660 835.290 252.720 ;
        RECT 834.970 144.740 835.290 144.800 ;
        RECT 835.890 144.740 836.210 144.800 ;
        RECT 834.970 144.600 836.210 144.740 ;
        RECT 834.970 144.540 835.290 144.600 ;
        RECT 835.890 144.540 836.210 144.600 ;
        RECT 834.970 96.460 835.290 96.520 ;
        RECT 834.775 96.320 835.290 96.460 ;
        RECT 834.970 96.260 835.290 96.320 ;
        RECT 834.985 48.520 835.275 48.565 ;
        RECT 835.430 48.520 835.750 48.580 ;
        RECT 834.985 48.380 835.750 48.520 ;
        RECT 834.985 48.335 835.275 48.380 ;
        RECT 835.430 48.320 835.750 48.380 ;
      LAYER via ;
        RECT 296.340 252.660 296.600 252.920 ;
        RECT 835.000 252.660 835.260 252.920 ;
        RECT 835.000 144.540 835.260 144.800 ;
        RECT 835.920 144.540 836.180 144.800 ;
        RECT 835.000 96.260 835.260 96.520 ;
        RECT 835.460 48.320 835.720 48.580 ;
      LAYER met2 ;
        RECT 296.330 2080.955 296.610 2081.325 ;
        RECT 296.400 252.950 296.540 2080.955 ;
        RECT 296.340 252.630 296.600 252.950 ;
        RECT 835.000 252.630 835.260 252.950 ;
        RECT 835.060 241.130 835.200 252.630 ;
        RECT 834.600 240.990 835.200 241.130 ;
        RECT 834.600 194.325 834.740 240.990 ;
        RECT 834.530 193.955 834.810 194.325 ;
        RECT 834.990 193.275 835.270 193.645 ;
        RECT 835.060 144.830 835.200 193.275 ;
        RECT 835.000 144.510 835.260 144.830 ;
        RECT 835.920 144.510 836.180 144.830 ;
        RECT 835.980 97.085 836.120 144.510 ;
        RECT 834.990 96.715 835.270 97.085 ;
        RECT 835.910 96.715 836.190 97.085 ;
        RECT 835.060 96.550 835.200 96.715 ;
        RECT 835.000 96.230 835.260 96.550 ;
        RECT 835.460 48.290 835.720 48.610 ;
        RECT 835.520 2.400 835.660 48.290 ;
        RECT 835.310 -4.800 835.870 2.400 ;
      LAYER via2 ;
        RECT 296.330 2081.000 296.610 2081.280 ;
        RECT 834.530 194.000 834.810 194.280 ;
        RECT 834.990 193.320 835.270 193.600 ;
        RECT 834.990 96.760 835.270 97.040 ;
        RECT 835.910 96.760 836.190 97.040 ;
      LAYER met3 ;
        RECT 296.305 2081.290 296.635 2081.305 ;
        RECT 310.000 2081.290 314.000 2081.680 ;
        RECT 296.305 2081.080 314.000 2081.290 ;
        RECT 296.305 2080.990 310.500 2081.080 ;
        RECT 296.305 2080.975 296.635 2080.990 ;
        RECT 834.505 194.290 834.835 194.305 ;
        RECT 834.505 193.990 835.970 194.290 ;
        RECT 834.505 193.975 834.835 193.990 ;
        RECT 834.965 193.610 835.295 193.625 ;
        RECT 835.670 193.610 835.970 193.990 ;
        RECT 834.965 193.310 835.970 193.610 ;
        RECT 834.965 193.295 835.295 193.310 ;
        RECT 834.965 97.050 835.295 97.065 ;
        RECT 835.885 97.050 836.215 97.065 ;
        RECT 834.965 96.750 836.215 97.050 ;
        RECT 834.965 96.735 835.295 96.750 ;
        RECT 835.885 96.735 836.215 96.750 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1048.410 3257.100 1048.730 3257.160 ;
        RECT 2773.870 3257.100 2774.190 3257.160 ;
        RECT 1048.410 3256.960 2774.190 3257.100 ;
        RECT 1048.410 3256.900 1048.730 3256.960 ;
        RECT 2773.870 3256.900 2774.190 3256.960 ;
        RECT 2773.870 37.980 2774.190 38.040 ;
        RECT 2779.850 37.980 2780.170 38.040 ;
        RECT 2773.870 37.840 2780.170 37.980 ;
        RECT 2773.870 37.780 2774.190 37.840 ;
        RECT 2779.850 37.780 2780.170 37.840 ;
      LAYER via ;
        RECT 1048.440 3256.900 1048.700 3257.160 ;
        RECT 2773.900 3256.900 2774.160 3257.160 ;
        RECT 2773.900 37.780 2774.160 38.040 ;
        RECT 2779.880 37.780 2780.140 38.040 ;
      LAYER met2 ;
        RECT 1047.930 3256.930 1048.210 3260.000 ;
        RECT 1048.440 3256.930 1048.700 3257.190 ;
        RECT 1047.930 3256.870 1048.700 3256.930 ;
        RECT 2773.900 3256.870 2774.160 3257.190 ;
        RECT 1047.930 3256.790 1048.640 3256.870 ;
        RECT 1047.930 3256.000 1048.210 3256.790 ;
        RECT 2773.960 38.070 2774.100 3256.870 ;
        RECT 2773.900 37.750 2774.160 38.070 ;
        RECT 2779.880 37.750 2780.140 38.070 ;
        RECT 2779.940 2.400 2780.080 37.750 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 447.190 3260.500 447.510 3260.560 ;
        RECT 458.230 3260.500 458.550 3260.560 ;
        RECT 447.190 3260.360 458.550 3260.500 ;
        RECT 447.190 3260.300 447.510 3260.360 ;
        RECT 458.230 3260.300 458.550 3260.360 ;
        RECT 2794.570 62.120 2794.890 62.180 ;
        RECT 2797.790 62.120 2798.110 62.180 ;
        RECT 2794.570 61.980 2798.110 62.120 ;
        RECT 2794.570 61.920 2794.890 61.980 ;
        RECT 2797.790 61.920 2798.110 61.980 ;
      LAYER via ;
        RECT 447.220 3260.300 447.480 3260.560 ;
        RECT 458.260 3260.300 458.520 3260.560 ;
        RECT 2794.600 61.920 2794.860 62.180 ;
        RECT 2797.820 61.920 2798.080 62.180 ;
      LAYER met2 ;
        RECT 447.220 3260.270 447.480 3260.590 ;
        RECT 458.260 3260.270 458.520 3260.590 ;
        RECT 447.280 3260.000 447.420 3260.270 ;
        RECT 447.170 3256.000 447.450 3260.000 ;
        RECT 458.320 3259.765 458.460 3260.270 ;
        RECT 458.250 3259.395 458.530 3259.765 ;
        RECT 2794.590 3259.395 2794.870 3259.765 ;
        RECT 2794.660 62.210 2794.800 3259.395 ;
        RECT 2794.600 61.890 2794.860 62.210 ;
        RECT 2797.820 61.890 2798.080 62.210 ;
        RECT 2797.880 2.400 2798.020 61.890 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
      LAYER via2 ;
        RECT 458.250 3259.440 458.530 3259.720 ;
        RECT 2794.590 3259.440 2794.870 3259.720 ;
      LAYER met3 ;
        RECT 458.225 3259.730 458.555 3259.745 ;
        RECT 2794.565 3259.730 2794.895 3259.745 ;
        RECT 458.225 3259.430 2794.895 3259.730 ;
        RECT 458.225 3259.415 458.555 3259.430 ;
        RECT 2794.565 3259.415 2794.895 3259.430 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.750 210.275 2816.030 210.645 ;
        RECT 2815.820 2.400 2815.960 210.275 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
      LAYER via2 ;
        RECT 2815.750 210.320 2816.030 210.600 ;
      LAYER met3 ;
        RECT 301.110 982.410 301.490 982.420 ;
        RECT 310.000 982.410 314.000 982.800 ;
        RECT 301.110 982.200 314.000 982.410 ;
        RECT 301.110 982.110 310.500 982.200 ;
        RECT 301.110 982.100 301.490 982.110 ;
        RECT 301.110 210.610 301.490 210.620 ;
        RECT 2815.725 210.610 2816.055 210.625 ;
        RECT 301.110 210.310 2816.055 210.610 ;
        RECT 301.110 210.300 301.490 210.310 ;
        RECT 2815.725 210.295 2816.055 210.310 ;
      LAYER via3 ;
        RECT 301.140 982.100 301.460 982.420 ;
        RECT 301.140 210.300 301.460 210.620 ;
      LAYER met4 ;
        RECT 301.135 982.095 301.465 982.425 ;
        RECT 301.150 210.625 301.450 982.095 ;
        RECT 301.135 210.295 301.465 210.625 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1127.070 244.020 1127.390 244.080 ;
        RECT 1131.210 244.020 1131.530 244.080 ;
        RECT 1127.070 243.880 1131.530 244.020 ;
        RECT 1127.070 243.820 1127.390 243.880 ;
        RECT 1131.210 243.820 1131.530 243.880 ;
        RECT 1131.210 32.880 1131.530 32.940 ;
        RECT 2833.670 32.880 2833.990 32.940 ;
        RECT 1131.210 32.740 2833.990 32.880 ;
        RECT 1131.210 32.680 1131.530 32.740 ;
        RECT 2833.670 32.680 2833.990 32.740 ;
      LAYER via ;
        RECT 1127.100 243.820 1127.360 244.080 ;
        RECT 1131.240 243.820 1131.500 244.080 ;
        RECT 1131.240 32.680 1131.500 32.940 ;
        RECT 2833.700 32.680 2833.960 32.940 ;
      LAYER met2 ;
        RECT 1127.050 260.000 1127.330 264.000 ;
        RECT 1127.160 244.110 1127.300 260.000 ;
        RECT 1127.100 243.790 1127.360 244.110 ;
        RECT 1131.240 243.790 1131.500 244.110 ;
        RECT 1131.300 32.970 1131.440 243.790 ;
        RECT 1131.240 32.650 1131.500 32.970 ;
        RECT 2833.700 32.650 2833.960 32.970 ;
        RECT 2833.760 2.400 2833.900 32.650 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2850.305 3236.205 2850.475 3259.155 ;
        RECT 2849.845 3139.645 2850.015 3187.755 ;
        RECT 2849.845 3043.085 2850.015 3091.195 ;
        RECT 2849.845 2946.525 2850.015 2994.295 ;
        RECT 2849.845 2849.625 2850.015 2898.075 ;
        RECT 2849.845 2173.705 2850.015 2221.815 ;
        RECT 2849.845 2077.145 2850.015 2125.255 ;
        RECT 2850.305 1980.245 2850.475 2028.355 ;
        RECT 2850.305 1883.685 2850.475 1931.795 ;
        RECT 2849.845 1787.125 2850.015 1834.895 ;
        RECT 2849.845 1690.565 2850.015 1738.675 ;
        RECT 2849.845 1594.005 2850.015 1642.115 ;
        RECT 2849.845 1497.445 2850.015 1545.555 ;
        RECT 2849.845 1400.885 2850.015 1448.995 ;
        RECT 2849.845 1304.325 2850.015 1352.435 ;
        RECT 2849.845 1207.765 2850.015 1255.875 ;
        RECT 2849.845 531.505 2850.015 579.615 ;
        RECT 2849.845 434.945 2850.015 483.055 ;
        RECT 2849.845 338.045 2850.015 386.155 ;
        RECT 2850.305 241.485 2850.475 289.595 ;
        RECT 2850.305 144.925 2850.475 193.035 ;
        RECT 2849.845 48.365 2850.015 96.475 ;
      LAYER mcon ;
        RECT 2850.305 3258.985 2850.475 3259.155 ;
        RECT 2849.845 3187.585 2850.015 3187.755 ;
        RECT 2849.845 3091.025 2850.015 3091.195 ;
        RECT 2849.845 2994.125 2850.015 2994.295 ;
        RECT 2849.845 2897.905 2850.015 2898.075 ;
        RECT 2849.845 2221.645 2850.015 2221.815 ;
        RECT 2849.845 2125.085 2850.015 2125.255 ;
        RECT 2850.305 2028.185 2850.475 2028.355 ;
        RECT 2850.305 1931.625 2850.475 1931.795 ;
        RECT 2849.845 1834.725 2850.015 1834.895 ;
        RECT 2849.845 1738.505 2850.015 1738.675 ;
        RECT 2849.845 1641.945 2850.015 1642.115 ;
        RECT 2849.845 1545.385 2850.015 1545.555 ;
        RECT 2849.845 1448.825 2850.015 1448.995 ;
        RECT 2849.845 1352.265 2850.015 1352.435 ;
        RECT 2849.845 1255.705 2850.015 1255.875 ;
        RECT 2849.845 579.445 2850.015 579.615 ;
        RECT 2849.845 482.885 2850.015 483.055 ;
        RECT 2849.845 385.985 2850.015 386.155 ;
        RECT 2850.305 289.425 2850.475 289.595 ;
        RECT 2850.305 192.865 2850.475 193.035 ;
        RECT 2849.845 96.305 2850.015 96.475 ;
      LAYER met1 ;
        RECT 1793.610 3259.140 1793.930 3259.200 ;
        RECT 2850.245 3259.140 2850.535 3259.185 ;
        RECT 1793.610 3259.000 2850.535 3259.140 ;
        RECT 1793.610 3258.940 1793.930 3259.000 ;
        RECT 2850.245 3258.955 2850.535 3259.000 ;
        RECT 2849.770 3236.360 2850.090 3236.420 ;
        RECT 2850.245 3236.360 2850.535 3236.405 ;
        RECT 2849.770 3236.220 2850.535 3236.360 ;
        RECT 2849.770 3236.160 2850.090 3236.220 ;
        RECT 2850.245 3236.175 2850.535 3236.220 ;
        RECT 2849.770 3187.740 2850.090 3187.800 ;
        RECT 2849.770 3187.600 2850.285 3187.740 ;
        RECT 2849.770 3187.540 2850.090 3187.600 ;
        RECT 2849.770 3139.800 2850.090 3139.860 ;
        RECT 2849.770 3139.660 2850.285 3139.800 ;
        RECT 2849.770 3139.600 2850.090 3139.660 ;
        RECT 2849.770 3091.180 2850.090 3091.240 ;
        RECT 2849.770 3091.040 2850.285 3091.180 ;
        RECT 2849.770 3090.980 2850.090 3091.040 ;
        RECT 2849.770 3043.240 2850.090 3043.300 ;
        RECT 2849.770 3043.100 2850.285 3043.240 ;
        RECT 2849.770 3043.040 2850.090 3043.100 ;
        RECT 2849.770 2995.780 2850.090 2996.040 ;
        RECT 2849.860 2995.020 2850.000 2995.780 ;
        RECT 2849.770 2994.760 2850.090 2995.020 ;
        RECT 2849.770 2994.280 2850.090 2994.340 ;
        RECT 2849.770 2994.140 2850.285 2994.280 ;
        RECT 2849.770 2994.080 2850.090 2994.140 ;
        RECT 2849.770 2946.680 2850.090 2946.740 ;
        RECT 2849.770 2946.540 2850.285 2946.680 ;
        RECT 2849.770 2946.480 2850.090 2946.540 ;
        RECT 2849.770 2898.060 2850.090 2898.120 ;
        RECT 2849.770 2897.920 2850.285 2898.060 ;
        RECT 2849.770 2897.860 2850.090 2897.920 ;
        RECT 2849.770 2849.780 2850.090 2849.840 ;
        RECT 2849.770 2849.640 2850.285 2849.780 ;
        RECT 2849.770 2849.580 2850.090 2849.640 ;
        RECT 2849.770 2753.220 2850.090 2753.280 ;
        RECT 2850.690 2753.220 2851.010 2753.280 ;
        RECT 2849.770 2753.080 2851.010 2753.220 ;
        RECT 2849.770 2753.020 2850.090 2753.080 ;
        RECT 2850.690 2753.020 2851.010 2753.080 ;
        RECT 2849.770 2656.660 2850.090 2656.720 ;
        RECT 2850.690 2656.660 2851.010 2656.720 ;
        RECT 2849.770 2656.520 2851.010 2656.660 ;
        RECT 2849.770 2656.460 2850.090 2656.520 ;
        RECT 2850.690 2656.460 2851.010 2656.520 ;
        RECT 2849.770 2560.100 2850.090 2560.160 ;
        RECT 2850.690 2560.100 2851.010 2560.160 ;
        RECT 2849.770 2559.960 2851.010 2560.100 ;
        RECT 2849.770 2559.900 2850.090 2559.960 ;
        RECT 2850.690 2559.900 2851.010 2559.960 ;
        RECT 2849.770 2414.920 2850.090 2414.980 ;
        RECT 2850.690 2414.920 2851.010 2414.980 ;
        RECT 2849.770 2414.780 2851.010 2414.920 ;
        RECT 2849.770 2414.720 2850.090 2414.780 ;
        RECT 2850.690 2414.720 2851.010 2414.780 ;
        RECT 2849.770 2318.360 2850.090 2318.420 ;
        RECT 2850.690 2318.360 2851.010 2318.420 ;
        RECT 2849.770 2318.220 2851.010 2318.360 ;
        RECT 2849.770 2318.160 2850.090 2318.220 ;
        RECT 2850.690 2318.160 2851.010 2318.220 ;
        RECT 2849.770 2221.800 2850.090 2221.860 ;
        RECT 2849.770 2221.660 2850.285 2221.800 ;
        RECT 2849.770 2221.600 2850.090 2221.660 ;
        RECT 2849.770 2173.860 2850.090 2173.920 ;
        RECT 2849.770 2173.720 2850.285 2173.860 ;
        RECT 2849.770 2173.660 2850.090 2173.720 ;
        RECT 2849.770 2125.240 2850.090 2125.300 ;
        RECT 2849.770 2125.100 2850.285 2125.240 ;
        RECT 2849.770 2125.040 2850.090 2125.100 ;
        RECT 2849.770 2077.300 2850.090 2077.360 ;
        RECT 2849.770 2077.160 2850.285 2077.300 ;
        RECT 2849.770 2077.100 2850.090 2077.160 ;
        RECT 2849.770 2028.340 2850.090 2028.400 ;
        RECT 2850.245 2028.340 2850.535 2028.385 ;
        RECT 2849.770 2028.200 2850.535 2028.340 ;
        RECT 2849.770 2028.140 2850.090 2028.200 ;
        RECT 2850.245 2028.155 2850.535 2028.200 ;
        RECT 2849.770 1980.400 2850.090 1980.460 ;
        RECT 2850.245 1980.400 2850.535 1980.445 ;
        RECT 2849.770 1980.260 2850.535 1980.400 ;
        RECT 2849.770 1980.200 2850.090 1980.260 ;
        RECT 2850.245 1980.215 2850.535 1980.260 ;
        RECT 2849.770 1931.780 2850.090 1931.840 ;
        RECT 2850.245 1931.780 2850.535 1931.825 ;
        RECT 2849.770 1931.640 2850.535 1931.780 ;
        RECT 2849.770 1931.580 2850.090 1931.640 ;
        RECT 2850.245 1931.595 2850.535 1931.640 ;
        RECT 2849.770 1883.840 2850.090 1883.900 ;
        RECT 2850.245 1883.840 2850.535 1883.885 ;
        RECT 2849.770 1883.700 2850.535 1883.840 ;
        RECT 2849.770 1883.640 2850.090 1883.700 ;
        RECT 2850.245 1883.655 2850.535 1883.700 ;
        RECT 2849.770 1834.880 2850.090 1834.940 ;
        RECT 2849.770 1834.740 2850.285 1834.880 ;
        RECT 2849.770 1834.680 2850.090 1834.740 ;
        RECT 2849.770 1787.280 2850.090 1787.340 ;
        RECT 2849.770 1787.140 2850.285 1787.280 ;
        RECT 2849.770 1787.080 2850.090 1787.140 ;
        RECT 2849.770 1738.660 2850.090 1738.720 ;
        RECT 2849.770 1738.520 2850.285 1738.660 ;
        RECT 2849.770 1738.460 2850.090 1738.520 ;
        RECT 2849.770 1690.720 2850.090 1690.780 ;
        RECT 2849.770 1690.580 2850.285 1690.720 ;
        RECT 2849.770 1690.520 2850.090 1690.580 ;
        RECT 2849.770 1642.100 2850.090 1642.160 ;
        RECT 2849.770 1641.960 2850.285 1642.100 ;
        RECT 2849.770 1641.900 2850.090 1641.960 ;
        RECT 2849.770 1594.160 2850.090 1594.220 ;
        RECT 2849.770 1594.020 2850.285 1594.160 ;
        RECT 2849.770 1593.960 2850.090 1594.020 ;
        RECT 2849.770 1545.540 2850.090 1545.600 ;
        RECT 2849.770 1545.400 2850.285 1545.540 ;
        RECT 2849.770 1545.340 2850.090 1545.400 ;
        RECT 2849.770 1497.600 2850.090 1497.660 ;
        RECT 2849.770 1497.460 2850.285 1497.600 ;
        RECT 2849.770 1497.400 2850.090 1497.460 ;
        RECT 2849.770 1448.980 2850.090 1449.040 ;
        RECT 2849.770 1448.840 2850.285 1448.980 ;
        RECT 2849.770 1448.780 2850.090 1448.840 ;
        RECT 2849.770 1401.040 2850.090 1401.100 ;
        RECT 2849.770 1400.900 2850.285 1401.040 ;
        RECT 2849.770 1400.840 2850.090 1400.900 ;
        RECT 2849.770 1352.420 2850.090 1352.480 ;
        RECT 2849.770 1352.280 2850.285 1352.420 ;
        RECT 2849.770 1352.220 2850.090 1352.280 ;
        RECT 2849.770 1304.480 2850.090 1304.540 ;
        RECT 2849.770 1304.340 2850.285 1304.480 ;
        RECT 2849.770 1304.280 2850.090 1304.340 ;
        RECT 2849.770 1255.860 2850.090 1255.920 ;
        RECT 2849.770 1255.720 2850.285 1255.860 ;
        RECT 2849.770 1255.660 2850.090 1255.720 ;
        RECT 2849.770 1207.920 2850.090 1207.980 ;
        RECT 2849.770 1207.780 2850.285 1207.920 ;
        RECT 2849.770 1207.720 2850.090 1207.780 ;
        RECT 2849.770 1111.020 2850.090 1111.080 ;
        RECT 2850.690 1111.020 2851.010 1111.080 ;
        RECT 2849.770 1110.880 2851.010 1111.020 ;
        RECT 2849.770 1110.820 2850.090 1110.880 ;
        RECT 2850.690 1110.820 2851.010 1110.880 ;
        RECT 2849.770 1014.460 2850.090 1014.520 ;
        RECT 2850.690 1014.460 2851.010 1014.520 ;
        RECT 2849.770 1014.320 2851.010 1014.460 ;
        RECT 2849.770 1014.260 2850.090 1014.320 ;
        RECT 2850.690 1014.260 2851.010 1014.320 ;
        RECT 2849.770 917.900 2850.090 917.960 ;
        RECT 2850.690 917.900 2851.010 917.960 ;
        RECT 2849.770 917.760 2851.010 917.900 ;
        RECT 2849.770 917.700 2850.090 917.760 ;
        RECT 2850.690 917.700 2851.010 917.760 ;
        RECT 2849.770 772.720 2850.090 772.780 ;
        RECT 2850.690 772.720 2851.010 772.780 ;
        RECT 2849.770 772.580 2851.010 772.720 ;
        RECT 2849.770 772.520 2850.090 772.580 ;
        RECT 2850.690 772.520 2851.010 772.580 ;
        RECT 2849.770 676.160 2850.090 676.220 ;
        RECT 2850.690 676.160 2851.010 676.220 ;
        RECT 2849.770 676.020 2851.010 676.160 ;
        RECT 2849.770 675.960 2850.090 676.020 ;
        RECT 2850.690 675.960 2851.010 676.020 ;
        RECT 2849.770 579.600 2850.090 579.660 ;
        RECT 2849.770 579.460 2850.285 579.600 ;
        RECT 2849.770 579.400 2850.090 579.460 ;
        RECT 2849.770 531.660 2850.090 531.720 ;
        RECT 2849.770 531.520 2850.285 531.660 ;
        RECT 2849.770 531.460 2850.090 531.520 ;
        RECT 2849.770 483.040 2850.090 483.100 ;
        RECT 2849.770 482.900 2850.285 483.040 ;
        RECT 2849.770 482.840 2850.090 482.900 ;
        RECT 2849.770 435.100 2850.090 435.160 ;
        RECT 2849.770 434.960 2850.285 435.100 ;
        RECT 2849.770 434.900 2850.090 434.960 ;
        RECT 2849.770 386.140 2850.090 386.200 ;
        RECT 2849.770 386.000 2850.285 386.140 ;
        RECT 2849.770 385.940 2850.090 386.000 ;
        RECT 2849.770 338.200 2850.090 338.260 ;
        RECT 2849.770 338.060 2850.285 338.200 ;
        RECT 2849.770 338.000 2850.090 338.060 ;
        RECT 2849.770 289.580 2850.090 289.640 ;
        RECT 2850.245 289.580 2850.535 289.625 ;
        RECT 2849.770 289.440 2850.535 289.580 ;
        RECT 2849.770 289.380 2850.090 289.440 ;
        RECT 2850.245 289.395 2850.535 289.440 ;
        RECT 2849.770 241.640 2850.090 241.700 ;
        RECT 2850.245 241.640 2850.535 241.685 ;
        RECT 2849.770 241.500 2850.535 241.640 ;
        RECT 2849.770 241.440 2850.090 241.500 ;
        RECT 2850.245 241.455 2850.535 241.500 ;
        RECT 2849.770 193.020 2850.090 193.080 ;
        RECT 2850.245 193.020 2850.535 193.065 ;
        RECT 2849.770 192.880 2850.535 193.020 ;
        RECT 2849.770 192.820 2850.090 192.880 ;
        RECT 2850.245 192.835 2850.535 192.880 ;
        RECT 2849.770 145.080 2850.090 145.140 ;
        RECT 2850.245 145.080 2850.535 145.125 ;
        RECT 2849.770 144.940 2850.535 145.080 ;
        RECT 2849.770 144.880 2850.090 144.940 ;
        RECT 2850.245 144.895 2850.535 144.940 ;
        RECT 2849.770 96.460 2850.090 96.520 ;
        RECT 2849.770 96.320 2850.285 96.460 ;
        RECT 2849.770 96.260 2850.090 96.320 ;
        RECT 2849.785 48.520 2850.075 48.565 ;
        RECT 2851.150 48.520 2851.470 48.580 ;
        RECT 2849.785 48.380 2851.470 48.520 ;
        RECT 2849.785 48.335 2850.075 48.380 ;
        RECT 2851.150 48.320 2851.470 48.380 ;
      LAYER via ;
        RECT 1793.640 3258.940 1793.900 3259.200 ;
        RECT 2849.800 3236.160 2850.060 3236.420 ;
        RECT 2849.800 3187.540 2850.060 3187.800 ;
        RECT 2849.800 3139.600 2850.060 3139.860 ;
        RECT 2849.800 3090.980 2850.060 3091.240 ;
        RECT 2849.800 3043.040 2850.060 3043.300 ;
        RECT 2849.800 2995.780 2850.060 2996.040 ;
        RECT 2849.800 2994.760 2850.060 2995.020 ;
        RECT 2849.800 2994.080 2850.060 2994.340 ;
        RECT 2849.800 2946.480 2850.060 2946.740 ;
        RECT 2849.800 2897.860 2850.060 2898.120 ;
        RECT 2849.800 2849.580 2850.060 2849.840 ;
        RECT 2849.800 2753.020 2850.060 2753.280 ;
        RECT 2850.720 2753.020 2850.980 2753.280 ;
        RECT 2849.800 2656.460 2850.060 2656.720 ;
        RECT 2850.720 2656.460 2850.980 2656.720 ;
        RECT 2849.800 2559.900 2850.060 2560.160 ;
        RECT 2850.720 2559.900 2850.980 2560.160 ;
        RECT 2849.800 2414.720 2850.060 2414.980 ;
        RECT 2850.720 2414.720 2850.980 2414.980 ;
        RECT 2849.800 2318.160 2850.060 2318.420 ;
        RECT 2850.720 2318.160 2850.980 2318.420 ;
        RECT 2849.800 2221.600 2850.060 2221.860 ;
        RECT 2849.800 2173.660 2850.060 2173.920 ;
        RECT 2849.800 2125.040 2850.060 2125.300 ;
        RECT 2849.800 2077.100 2850.060 2077.360 ;
        RECT 2849.800 2028.140 2850.060 2028.400 ;
        RECT 2849.800 1980.200 2850.060 1980.460 ;
        RECT 2849.800 1931.580 2850.060 1931.840 ;
        RECT 2849.800 1883.640 2850.060 1883.900 ;
        RECT 2849.800 1834.680 2850.060 1834.940 ;
        RECT 2849.800 1787.080 2850.060 1787.340 ;
        RECT 2849.800 1738.460 2850.060 1738.720 ;
        RECT 2849.800 1690.520 2850.060 1690.780 ;
        RECT 2849.800 1641.900 2850.060 1642.160 ;
        RECT 2849.800 1593.960 2850.060 1594.220 ;
        RECT 2849.800 1545.340 2850.060 1545.600 ;
        RECT 2849.800 1497.400 2850.060 1497.660 ;
        RECT 2849.800 1448.780 2850.060 1449.040 ;
        RECT 2849.800 1400.840 2850.060 1401.100 ;
        RECT 2849.800 1352.220 2850.060 1352.480 ;
        RECT 2849.800 1304.280 2850.060 1304.540 ;
        RECT 2849.800 1255.660 2850.060 1255.920 ;
        RECT 2849.800 1207.720 2850.060 1207.980 ;
        RECT 2849.800 1110.820 2850.060 1111.080 ;
        RECT 2850.720 1110.820 2850.980 1111.080 ;
        RECT 2849.800 1014.260 2850.060 1014.520 ;
        RECT 2850.720 1014.260 2850.980 1014.520 ;
        RECT 2849.800 917.700 2850.060 917.960 ;
        RECT 2850.720 917.700 2850.980 917.960 ;
        RECT 2849.800 772.520 2850.060 772.780 ;
        RECT 2850.720 772.520 2850.980 772.780 ;
        RECT 2849.800 675.960 2850.060 676.220 ;
        RECT 2850.720 675.960 2850.980 676.220 ;
        RECT 2849.800 579.400 2850.060 579.660 ;
        RECT 2849.800 531.460 2850.060 531.720 ;
        RECT 2849.800 482.840 2850.060 483.100 ;
        RECT 2849.800 434.900 2850.060 435.160 ;
        RECT 2849.800 385.940 2850.060 386.200 ;
        RECT 2849.800 338.000 2850.060 338.260 ;
        RECT 2849.800 289.380 2850.060 289.640 ;
        RECT 2849.800 241.440 2850.060 241.700 ;
        RECT 2849.800 192.820 2850.060 193.080 ;
        RECT 2849.800 144.880 2850.060 145.140 ;
        RECT 2849.800 96.260 2850.060 96.520 ;
        RECT 2851.180 48.320 2851.440 48.580 ;
      LAYER met2 ;
        RECT 1792.210 3258.970 1792.490 3260.000 ;
        RECT 1793.640 3258.970 1793.900 3259.230 ;
        RECT 1792.210 3258.910 1793.900 3258.970 ;
        RECT 1792.210 3258.830 1793.840 3258.910 ;
        RECT 1792.210 3256.000 1792.490 3258.830 ;
        RECT 2849.800 3236.130 2850.060 3236.450 ;
        RECT 2849.860 3187.830 2850.000 3236.130 ;
        RECT 2849.800 3187.510 2850.060 3187.830 ;
        RECT 2849.800 3139.570 2850.060 3139.890 ;
        RECT 2849.860 3091.270 2850.000 3139.570 ;
        RECT 2849.800 3090.950 2850.060 3091.270 ;
        RECT 2849.800 3043.010 2850.060 3043.330 ;
        RECT 2849.860 2996.070 2850.000 3043.010 ;
        RECT 2849.800 2995.750 2850.060 2996.070 ;
        RECT 2849.800 2994.730 2850.060 2995.050 ;
        RECT 2849.860 2994.370 2850.000 2994.730 ;
        RECT 2849.800 2994.050 2850.060 2994.370 ;
        RECT 2849.800 2946.450 2850.060 2946.770 ;
        RECT 2849.860 2898.150 2850.000 2946.450 ;
        RECT 2849.800 2897.830 2850.060 2898.150 ;
        RECT 2849.800 2849.550 2850.060 2849.870 ;
        RECT 2849.860 2801.445 2850.000 2849.550 ;
        RECT 2849.790 2801.075 2850.070 2801.445 ;
        RECT 2850.710 2801.075 2850.990 2801.445 ;
        RECT 2850.780 2753.310 2850.920 2801.075 ;
        RECT 2849.800 2752.990 2850.060 2753.310 ;
        RECT 2850.720 2752.990 2850.980 2753.310 ;
        RECT 2849.860 2704.885 2850.000 2752.990 ;
        RECT 2849.790 2704.515 2850.070 2704.885 ;
        RECT 2850.710 2704.515 2850.990 2704.885 ;
        RECT 2850.780 2656.750 2850.920 2704.515 ;
        RECT 2849.800 2656.430 2850.060 2656.750 ;
        RECT 2850.720 2656.430 2850.980 2656.750 ;
        RECT 2849.860 2608.325 2850.000 2656.430 ;
        RECT 2849.790 2607.955 2850.070 2608.325 ;
        RECT 2850.710 2607.955 2850.990 2608.325 ;
        RECT 2850.780 2560.190 2850.920 2607.955 ;
        RECT 2849.800 2559.870 2850.060 2560.190 ;
        RECT 2850.720 2559.870 2850.980 2560.190 ;
        RECT 2849.860 2511.765 2850.000 2559.870 ;
        RECT 2849.790 2511.395 2850.070 2511.765 ;
        RECT 2850.710 2511.395 2850.990 2511.765 ;
        RECT 2850.780 2463.485 2850.920 2511.395 ;
        RECT 2849.790 2463.115 2850.070 2463.485 ;
        RECT 2850.710 2463.115 2850.990 2463.485 ;
        RECT 2849.860 2415.010 2850.000 2463.115 ;
        RECT 2849.800 2414.690 2850.060 2415.010 ;
        RECT 2850.720 2414.690 2850.980 2415.010 ;
        RECT 2850.780 2366.925 2850.920 2414.690 ;
        RECT 2849.790 2366.555 2850.070 2366.925 ;
        RECT 2850.710 2366.555 2850.990 2366.925 ;
        RECT 2849.860 2318.450 2850.000 2366.555 ;
        RECT 2849.800 2318.130 2850.060 2318.450 ;
        RECT 2850.720 2318.130 2850.980 2318.450 ;
        RECT 2850.780 2270.365 2850.920 2318.130 ;
        RECT 2849.790 2269.995 2850.070 2270.365 ;
        RECT 2850.710 2269.995 2850.990 2270.365 ;
        RECT 2849.860 2221.890 2850.000 2269.995 ;
        RECT 2849.800 2221.570 2850.060 2221.890 ;
        RECT 2849.800 2173.630 2850.060 2173.950 ;
        RECT 2849.860 2125.330 2850.000 2173.630 ;
        RECT 2849.800 2125.010 2850.060 2125.330 ;
        RECT 2849.800 2077.070 2850.060 2077.390 ;
        RECT 2849.860 2028.430 2850.000 2077.070 ;
        RECT 2849.800 2028.110 2850.060 2028.430 ;
        RECT 2849.800 1980.170 2850.060 1980.490 ;
        RECT 2849.860 1931.870 2850.000 1980.170 ;
        RECT 2849.800 1931.550 2850.060 1931.870 ;
        RECT 2849.800 1883.610 2850.060 1883.930 ;
        RECT 2849.860 1836.525 2850.000 1883.610 ;
        RECT 2849.790 1836.155 2850.070 1836.525 ;
        RECT 2849.790 1835.475 2850.070 1835.845 ;
        RECT 2849.860 1834.970 2850.000 1835.475 ;
        RECT 2849.800 1834.650 2850.060 1834.970 ;
        RECT 2849.800 1787.050 2850.060 1787.370 ;
        RECT 2849.860 1739.965 2850.000 1787.050 ;
        RECT 2849.790 1739.595 2850.070 1739.965 ;
        RECT 2849.790 1738.915 2850.070 1739.285 ;
        RECT 2849.860 1738.750 2850.000 1738.915 ;
        RECT 2849.800 1738.430 2850.060 1738.750 ;
        RECT 2849.800 1690.490 2850.060 1690.810 ;
        RECT 2849.860 1642.190 2850.000 1690.490 ;
        RECT 2849.800 1641.870 2850.060 1642.190 ;
        RECT 2849.800 1593.930 2850.060 1594.250 ;
        RECT 2849.860 1545.630 2850.000 1593.930 ;
        RECT 2849.800 1545.310 2850.060 1545.630 ;
        RECT 2849.800 1497.370 2850.060 1497.690 ;
        RECT 2849.860 1449.070 2850.000 1497.370 ;
        RECT 2849.800 1448.750 2850.060 1449.070 ;
        RECT 2849.800 1400.810 2850.060 1401.130 ;
        RECT 2849.860 1352.510 2850.000 1400.810 ;
        RECT 2849.800 1352.190 2850.060 1352.510 ;
        RECT 2849.800 1304.250 2850.060 1304.570 ;
        RECT 2849.860 1257.165 2850.000 1304.250 ;
        RECT 2849.790 1256.795 2850.070 1257.165 ;
        RECT 2849.790 1256.115 2850.070 1256.485 ;
        RECT 2849.860 1255.950 2850.000 1256.115 ;
        RECT 2849.800 1255.630 2850.060 1255.950 ;
        RECT 2849.800 1207.690 2850.060 1208.010 ;
        RECT 2849.860 1159.245 2850.000 1207.690 ;
        RECT 2849.790 1158.875 2850.070 1159.245 ;
        RECT 2850.710 1158.875 2850.990 1159.245 ;
        RECT 2850.780 1111.110 2850.920 1158.875 ;
        RECT 2849.800 1110.790 2850.060 1111.110 ;
        RECT 2850.720 1110.790 2850.980 1111.110 ;
        RECT 2849.860 1062.685 2850.000 1110.790 ;
        RECT 2849.790 1062.315 2850.070 1062.685 ;
        RECT 2850.710 1062.315 2850.990 1062.685 ;
        RECT 2850.780 1014.550 2850.920 1062.315 ;
        RECT 2849.800 1014.230 2850.060 1014.550 ;
        RECT 2850.720 1014.230 2850.980 1014.550 ;
        RECT 2849.860 966.125 2850.000 1014.230 ;
        RECT 2849.790 965.755 2850.070 966.125 ;
        RECT 2850.710 965.755 2850.990 966.125 ;
        RECT 2850.780 917.990 2850.920 965.755 ;
        RECT 2849.800 917.670 2850.060 917.990 ;
        RECT 2850.720 917.670 2850.980 917.990 ;
        RECT 2849.860 869.565 2850.000 917.670 ;
        RECT 2849.790 869.195 2850.070 869.565 ;
        RECT 2850.710 869.195 2850.990 869.565 ;
        RECT 2850.780 821.285 2850.920 869.195 ;
        RECT 2849.790 820.915 2850.070 821.285 ;
        RECT 2850.710 820.915 2850.990 821.285 ;
        RECT 2849.860 772.810 2850.000 820.915 ;
        RECT 2849.800 772.490 2850.060 772.810 ;
        RECT 2850.720 772.490 2850.980 772.810 ;
        RECT 2850.780 724.725 2850.920 772.490 ;
        RECT 2849.790 724.355 2850.070 724.725 ;
        RECT 2850.710 724.355 2850.990 724.725 ;
        RECT 2849.860 676.250 2850.000 724.355 ;
        RECT 2849.800 675.930 2850.060 676.250 ;
        RECT 2850.720 675.930 2850.980 676.250 ;
        RECT 2850.780 628.165 2850.920 675.930 ;
        RECT 2849.790 627.795 2850.070 628.165 ;
        RECT 2850.710 627.795 2850.990 628.165 ;
        RECT 2849.860 579.690 2850.000 627.795 ;
        RECT 2849.800 579.370 2850.060 579.690 ;
        RECT 2849.800 531.430 2850.060 531.750 ;
        RECT 2849.860 483.130 2850.000 531.430 ;
        RECT 2849.800 482.810 2850.060 483.130 ;
        RECT 2849.800 434.870 2850.060 435.190 ;
        RECT 2849.860 386.230 2850.000 434.870 ;
        RECT 2849.800 385.910 2850.060 386.230 ;
        RECT 2849.800 337.970 2850.060 338.290 ;
        RECT 2849.860 289.670 2850.000 337.970 ;
        RECT 2849.800 289.350 2850.060 289.670 ;
        RECT 2849.800 241.410 2850.060 241.730 ;
        RECT 2849.860 194.325 2850.000 241.410 ;
        RECT 2849.790 193.955 2850.070 194.325 ;
        RECT 2849.790 193.275 2850.070 193.645 ;
        RECT 2849.860 193.110 2850.000 193.275 ;
        RECT 2849.800 192.790 2850.060 193.110 ;
        RECT 2849.800 144.850 2850.060 145.170 ;
        RECT 2849.860 97.765 2850.000 144.850 ;
        RECT 2849.790 97.395 2850.070 97.765 ;
        RECT 2849.790 96.715 2850.070 97.085 ;
        RECT 2849.860 96.550 2850.000 96.715 ;
        RECT 2849.800 96.230 2850.060 96.550 ;
        RECT 2851.180 48.290 2851.440 48.610 ;
        RECT 2851.240 2.400 2851.380 48.290 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
      LAYER via2 ;
        RECT 2849.790 2801.120 2850.070 2801.400 ;
        RECT 2850.710 2801.120 2850.990 2801.400 ;
        RECT 2849.790 2704.560 2850.070 2704.840 ;
        RECT 2850.710 2704.560 2850.990 2704.840 ;
        RECT 2849.790 2608.000 2850.070 2608.280 ;
        RECT 2850.710 2608.000 2850.990 2608.280 ;
        RECT 2849.790 2511.440 2850.070 2511.720 ;
        RECT 2850.710 2511.440 2850.990 2511.720 ;
        RECT 2849.790 2463.160 2850.070 2463.440 ;
        RECT 2850.710 2463.160 2850.990 2463.440 ;
        RECT 2849.790 2366.600 2850.070 2366.880 ;
        RECT 2850.710 2366.600 2850.990 2366.880 ;
        RECT 2849.790 2270.040 2850.070 2270.320 ;
        RECT 2850.710 2270.040 2850.990 2270.320 ;
        RECT 2849.790 1836.200 2850.070 1836.480 ;
        RECT 2849.790 1835.520 2850.070 1835.800 ;
        RECT 2849.790 1739.640 2850.070 1739.920 ;
        RECT 2849.790 1738.960 2850.070 1739.240 ;
        RECT 2849.790 1256.840 2850.070 1257.120 ;
        RECT 2849.790 1256.160 2850.070 1256.440 ;
        RECT 2849.790 1158.920 2850.070 1159.200 ;
        RECT 2850.710 1158.920 2850.990 1159.200 ;
        RECT 2849.790 1062.360 2850.070 1062.640 ;
        RECT 2850.710 1062.360 2850.990 1062.640 ;
        RECT 2849.790 965.800 2850.070 966.080 ;
        RECT 2850.710 965.800 2850.990 966.080 ;
        RECT 2849.790 869.240 2850.070 869.520 ;
        RECT 2850.710 869.240 2850.990 869.520 ;
        RECT 2849.790 820.960 2850.070 821.240 ;
        RECT 2850.710 820.960 2850.990 821.240 ;
        RECT 2849.790 724.400 2850.070 724.680 ;
        RECT 2850.710 724.400 2850.990 724.680 ;
        RECT 2849.790 627.840 2850.070 628.120 ;
        RECT 2850.710 627.840 2850.990 628.120 ;
        RECT 2849.790 194.000 2850.070 194.280 ;
        RECT 2849.790 193.320 2850.070 193.600 ;
        RECT 2849.790 97.440 2850.070 97.720 ;
        RECT 2849.790 96.760 2850.070 97.040 ;
      LAYER met3 ;
        RECT 2849.765 2801.410 2850.095 2801.425 ;
        RECT 2850.685 2801.410 2851.015 2801.425 ;
        RECT 2849.765 2801.110 2851.015 2801.410 ;
        RECT 2849.765 2801.095 2850.095 2801.110 ;
        RECT 2850.685 2801.095 2851.015 2801.110 ;
        RECT 2849.765 2704.850 2850.095 2704.865 ;
        RECT 2850.685 2704.850 2851.015 2704.865 ;
        RECT 2849.765 2704.550 2851.015 2704.850 ;
        RECT 2849.765 2704.535 2850.095 2704.550 ;
        RECT 2850.685 2704.535 2851.015 2704.550 ;
        RECT 2849.765 2608.290 2850.095 2608.305 ;
        RECT 2850.685 2608.290 2851.015 2608.305 ;
        RECT 2849.765 2607.990 2851.015 2608.290 ;
        RECT 2849.765 2607.975 2850.095 2607.990 ;
        RECT 2850.685 2607.975 2851.015 2607.990 ;
        RECT 2849.765 2511.730 2850.095 2511.745 ;
        RECT 2850.685 2511.730 2851.015 2511.745 ;
        RECT 2849.765 2511.430 2851.015 2511.730 ;
        RECT 2849.765 2511.415 2850.095 2511.430 ;
        RECT 2850.685 2511.415 2851.015 2511.430 ;
        RECT 2849.765 2463.450 2850.095 2463.465 ;
        RECT 2850.685 2463.450 2851.015 2463.465 ;
        RECT 2849.765 2463.150 2851.015 2463.450 ;
        RECT 2849.765 2463.135 2850.095 2463.150 ;
        RECT 2850.685 2463.135 2851.015 2463.150 ;
        RECT 2849.765 2366.890 2850.095 2366.905 ;
        RECT 2850.685 2366.890 2851.015 2366.905 ;
        RECT 2849.765 2366.590 2851.015 2366.890 ;
        RECT 2849.765 2366.575 2850.095 2366.590 ;
        RECT 2850.685 2366.575 2851.015 2366.590 ;
        RECT 2849.765 2270.330 2850.095 2270.345 ;
        RECT 2850.685 2270.330 2851.015 2270.345 ;
        RECT 2849.765 2270.030 2851.015 2270.330 ;
        RECT 2849.765 2270.015 2850.095 2270.030 ;
        RECT 2850.685 2270.015 2851.015 2270.030 ;
        RECT 2849.765 1836.490 2850.095 1836.505 ;
        RECT 2849.550 1836.175 2850.095 1836.490 ;
        RECT 2849.550 1835.825 2849.850 1836.175 ;
        RECT 2849.550 1835.510 2850.095 1835.825 ;
        RECT 2849.765 1835.495 2850.095 1835.510 ;
        RECT 2849.765 1739.930 2850.095 1739.945 ;
        RECT 2849.550 1739.615 2850.095 1739.930 ;
        RECT 2849.550 1739.265 2849.850 1739.615 ;
        RECT 2849.550 1738.950 2850.095 1739.265 ;
        RECT 2849.765 1738.935 2850.095 1738.950 ;
        RECT 2849.765 1257.130 2850.095 1257.145 ;
        RECT 2849.550 1256.815 2850.095 1257.130 ;
        RECT 2849.550 1256.465 2849.850 1256.815 ;
        RECT 2849.550 1256.150 2850.095 1256.465 ;
        RECT 2849.765 1256.135 2850.095 1256.150 ;
        RECT 2849.765 1159.210 2850.095 1159.225 ;
        RECT 2850.685 1159.210 2851.015 1159.225 ;
        RECT 2849.765 1158.910 2851.015 1159.210 ;
        RECT 2849.765 1158.895 2850.095 1158.910 ;
        RECT 2850.685 1158.895 2851.015 1158.910 ;
        RECT 2849.765 1062.650 2850.095 1062.665 ;
        RECT 2850.685 1062.650 2851.015 1062.665 ;
        RECT 2849.765 1062.350 2851.015 1062.650 ;
        RECT 2849.765 1062.335 2850.095 1062.350 ;
        RECT 2850.685 1062.335 2851.015 1062.350 ;
        RECT 2849.765 966.090 2850.095 966.105 ;
        RECT 2850.685 966.090 2851.015 966.105 ;
        RECT 2849.765 965.790 2851.015 966.090 ;
        RECT 2849.765 965.775 2850.095 965.790 ;
        RECT 2850.685 965.775 2851.015 965.790 ;
        RECT 2849.765 869.530 2850.095 869.545 ;
        RECT 2850.685 869.530 2851.015 869.545 ;
        RECT 2849.765 869.230 2851.015 869.530 ;
        RECT 2849.765 869.215 2850.095 869.230 ;
        RECT 2850.685 869.215 2851.015 869.230 ;
        RECT 2849.765 821.250 2850.095 821.265 ;
        RECT 2850.685 821.250 2851.015 821.265 ;
        RECT 2849.765 820.950 2851.015 821.250 ;
        RECT 2849.765 820.935 2850.095 820.950 ;
        RECT 2850.685 820.935 2851.015 820.950 ;
        RECT 2849.765 724.690 2850.095 724.705 ;
        RECT 2850.685 724.690 2851.015 724.705 ;
        RECT 2849.765 724.390 2851.015 724.690 ;
        RECT 2849.765 724.375 2850.095 724.390 ;
        RECT 2850.685 724.375 2851.015 724.390 ;
        RECT 2849.765 628.130 2850.095 628.145 ;
        RECT 2850.685 628.130 2851.015 628.145 ;
        RECT 2849.765 627.830 2851.015 628.130 ;
        RECT 2849.765 627.815 2850.095 627.830 ;
        RECT 2850.685 627.815 2851.015 627.830 ;
        RECT 2849.765 194.290 2850.095 194.305 ;
        RECT 2849.550 193.975 2850.095 194.290 ;
        RECT 2849.550 193.625 2849.850 193.975 ;
        RECT 2849.550 193.310 2850.095 193.625 ;
        RECT 2849.765 193.295 2850.095 193.310 ;
        RECT 2849.765 97.730 2850.095 97.745 ;
        RECT 2849.550 97.415 2850.095 97.730 ;
        RECT 2849.550 97.065 2849.850 97.415 ;
        RECT 2849.550 96.750 2850.095 97.065 ;
        RECT 2849.765 96.735 2850.095 96.750 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1097.420 2615.490 1097.480 ;
        RECT 2863.570 1097.420 2863.890 1097.480 ;
        RECT 2615.170 1097.280 2863.890 1097.420 ;
        RECT 2615.170 1097.220 2615.490 1097.280 ;
        RECT 2863.570 1097.220 2863.890 1097.280 ;
      LAYER via ;
        RECT 2615.200 1097.220 2615.460 1097.480 ;
        RECT 2863.600 1097.220 2863.860 1097.480 ;
      LAYER met2 ;
        RECT 2615.190 1099.035 2615.470 1099.405 ;
        RECT 2615.260 1097.510 2615.400 1099.035 ;
        RECT 2615.200 1097.190 2615.460 1097.510 ;
        RECT 2863.600 1097.190 2863.860 1097.510 ;
        RECT 2863.660 19.450 2863.800 1097.190 ;
        RECT 2863.660 19.310 2869.320 19.450 ;
        RECT 2869.180 2.400 2869.320 19.310 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1099.080 2615.470 1099.360 ;
      LAYER met3 ;
        RECT 2606.000 1099.370 2610.000 1099.760 ;
        RECT 2615.165 1099.370 2615.495 1099.385 ;
        RECT 2606.000 1099.160 2615.495 1099.370 ;
        RECT 2609.580 1099.070 2615.495 1099.160 ;
        RECT 2615.165 1099.055 2615.495 1099.070 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1559.010 169.220 1559.330 169.280 ;
        RECT 2873.690 169.220 2874.010 169.280 ;
        RECT 1559.010 169.080 2874.010 169.220 ;
        RECT 1559.010 169.020 1559.330 169.080 ;
        RECT 2873.690 169.020 2874.010 169.080 ;
        RECT 2873.690 20.640 2874.010 20.700 ;
        RECT 2887.030 20.640 2887.350 20.700 ;
        RECT 2873.690 20.500 2887.350 20.640 ;
        RECT 2873.690 20.440 2874.010 20.500 ;
        RECT 2887.030 20.440 2887.350 20.500 ;
      LAYER via ;
        RECT 1559.040 169.020 1559.300 169.280 ;
        RECT 2873.720 169.020 2873.980 169.280 ;
        RECT 2873.720 20.440 2873.980 20.700 ;
        RECT 2887.060 20.440 2887.320 20.700 ;
      LAYER met2 ;
        RECT 1556.690 260.170 1556.970 264.000 ;
        RECT 1556.690 260.030 1559.240 260.170 ;
        RECT 1556.690 260.000 1556.970 260.030 ;
        RECT 1559.100 169.310 1559.240 260.030 ;
        RECT 1559.040 168.990 1559.300 169.310 ;
        RECT 2873.720 168.990 2873.980 169.310 ;
        RECT 2873.780 20.730 2873.920 168.990 ;
        RECT 2873.720 20.410 2873.980 20.730 ;
        RECT 2887.060 20.410 2887.320 20.730 ;
        RECT 2887.120 2.400 2887.260 20.410 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2442.670 247.760 2442.990 247.820 ;
        RECT 2708.550 247.760 2708.870 247.820 ;
        RECT 2442.670 247.620 2708.870 247.760 ;
        RECT 2442.670 247.560 2442.990 247.620 ;
        RECT 2708.550 247.560 2708.870 247.620 ;
        RECT 2708.550 18.940 2708.870 19.000 ;
        RECT 2708.550 18.800 2745.120 18.940 ;
        RECT 2708.550 18.740 2708.870 18.800 ;
        RECT 2744.980 17.920 2745.120 18.800 ;
        RECT 2904.970 17.920 2905.290 17.980 ;
        RECT 2744.980 17.780 2905.290 17.920 ;
        RECT 2904.970 17.720 2905.290 17.780 ;
      LAYER via ;
        RECT 2442.700 247.560 2442.960 247.820 ;
        RECT 2708.580 247.560 2708.840 247.820 ;
        RECT 2708.580 18.740 2708.840 19.000 ;
        RECT 2905.000 17.720 2905.260 17.980 ;
      LAYER met2 ;
        RECT 2442.650 260.000 2442.930 264.000 ;
        RECT 2442.760 247.850 2442.900 260.000 ;
        RECT 2442.700 247.530 2442.960 247.850 ;
        RECT 2708.580 247.530 2708.840 247.850 ;
        RECT 2708.640 19.030 2708.780 247.530 ;
        RECT 2708.580 18.710 2708.840 19.030 ;
        RECT 2905.000 17.690 2905.260 18.010 ;
        RECT 2905.060 2.400 2905.200 17.690 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 541.030 244.020 541.350 244.080 ;
        RECT 544.710 244.020 545.030 244.080 ;
        RECT 541.030 243.880 545.030 244.020 ;
        RECT 541.030 243.820 541.350 243.880 ;
        RECT 544.710 243.820 545.030 243.880 ;
        RECT 544.710 26.080 545.030 26.140 ;
        RECT 852.910 26.080 853.230 26.140 ;
        RECT 544.710 25.940 853.230 26.080 ;
        RECT 544.710 25.880 545.030 25.940 ;
        RECT 852.910 25.880 853.230 25.940 ;
      LAYER via ;
        RECT 541.060 243.820 541.320 244.080 ;
        RECT 544.740 243.820 545.000 244.080 ;
        RECT 544.740 25.880 545.000 26.140 ;
        RECT 852.940 25.880 853.200 26.140 ;
      LAYER met2 ;
        RECT 541.010 260.000 541.290 264.000 ;
        RECT 541.120 244.110 541.260 260.000 ;
        RECT 541.060 243.790 541.320 244.110 ;
        RECT 544.740 243.790 545.000 244.110 ;
        RECT 544.800 26.170 544.940 243.790 ;
        RECT 544.740 25.850 545.000 26.170 ;
        RECT 852.940 25.850 853.200 26.170 ;
        RECT 853.000 2.400 853.140 25.850 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 310.185 3181.125 310.355 3229.235 ;
        RECT 309.725 3043.425 309.895 3132.675 ;
        RECT 309.725 2939.385 309.895 2960.295 ;
        RECT 309.265 2891.105 309.435 2912.355 ;
        RECT 308.805 2408.305 308.975 2456.415 ;
        RECT 309.265 2070.005 309.435 2118.115 ;
        RECT 309.265 1193.825 309.435 1241.935 ;
        RECT 309.725 699.805 309.895 724.455 ;
        RECT 870.005 144.925 870.175 193.035 ;
        RECT 869.545 48.365 869.715 96.475 ;
      LAYER mcon ;
        RECT 310.185 3229.065 310.355 3229.235 ;
        RECT 309.725 3132.505 309.895 3132.675 ;
        RECT 309.725 2960.125 309.895 2960.295 ;
        RECT 309.265 2912.185 309.435 2912.355 ;
        RECT 308.805 2456.245 308.975 2456.415 ;
        RECT 309.265 2117.945 309.435 2118.115 ;
        RECT 309.265 1241.765 309.435 1241.935 ;
        RECT 309.725 724.285 309.895 724.455 ;
        RECT 870.005 192.865 870.175 193.035 ;
        RECT 869.545 96.305 869.715 96.475 ;
      LAYER met1 ;
        RECT 310.110 3229.220 310.430 3229.280 ;
        RECT 309.915 3229.080 310.430 3229.220 ;
        RECT 310.110 3229.020 310.430 3229.080 ;
        RECT 310.110 3181.280 310.430 3181.340 ;
        RECT 309.915 3181.140 310.430 3181.280 ;
        RECT 310.110 3181.080 310.430 3181.140 ;
        RECT 309.650 3140.140 309.970 3140.200 ;
        RECT 310.570 3140.140 310.890 3140.200 ;
        RECT 309.650 3140.000 310.890 3140.140 ;
        RECT 309.650 3139.940 309.970 3140.000 ;
        RECT 310.570 3139.940 310.890 3140.000 ;
        RECT 309.650 3132.660 309.970 3132.720 ;
        RECT 309.455 3132.520 309.970 3132.660 ;
        RECT 309.650 3132.460 309.970 3132.520 ;
        RECT 309.650 3043.580 309.970 3043.640 ;
        RECT 309.455 3043.440 309.970 3043.580 ;
        RECT 309.650 3043.380 309.970 3043.440 ;
        RECT 309.650 2960.280 309.970 2960.340 ;
        RECT 309.455 2960.140 309.970 2960.280 ;
        RECT 309.650 2960.080 309.970 2960.140 ;
        RECT 309.650 2939.540 309.970 2939.600 ;
        RECT 309.455 2939.400 309.970 2939.540 ;
        RECT 309.650 2939.340 309.970 2939.400 ;
        RECT 309.205 2912.340 309.495 2912.385 ;
        RECT 309.650 2912.340 309.970 2912.400 ;
        RECT 309.205 2912.200 309.970 2912.340 ;
        RECT 309.205 2912.155 309.495 2912.200 ;
        RECT 309.650 2912.140 309.970 2912.200 ;
        RECT 309.190 2891.260 309.510 2891.320 ;
        RECT 308.995 2891.120 309.510 2891.260 ;
        RECT 309.190 2891.060 309.510 2891.120 ;
        RECT 309.190 2815.100 309.510 2815.160 ;
        RECT 310.110 2815.100 310.430 2815.160 ;
        RECT 309.190 2814.960 310.430 2815.100 ;
        RECT 309.190 2814.900 309.510 2814.960 ;
        RECT 310.110 2814.900 310.430 2814.960 ;
        RECT 308.730 2746.420 309.050 2746.480 ;
        RECT 309.650 2746.420 309.970 2746.480 ;
        RECT 308.730 2746.280 309.970 2746.420 ;
        RECT 308.730 2746.220 309.050 2746.280 ;
        RECT 309.650 2746.220 309.970 2746.280 ;
        RECT 308.730 2697.800 309.050 2697.860 ;
        RECT 309.650 2697.800 309.970 2697.860 ;
        RECT 308.730 2697.660 309.970 2697.800 ;
        RECT 308.730 2697.600 309.050 2697.660 ;
        RECT 309.650 2697.600 309.970 2697.660 ;
        RECT 308.270 2649.520 308.590 2649.580 ;
        RECT 309.650 2649.520 309.970 2649.580 ;
        RECT 308.270 2649.380 309.970 2649.520 ;
        RECT 308.270 2649.320 308.590 2649.380 ;
        RECT 309.650 2649.320 309.970 2649.380 ;
        RECT 309.190 2560.100 309.510 2560.160 ;
        RECT 309.650 2560.100 309.970 2560.160 ;
        RECT 309.190 2559.960 309.970 2560.100 ;
        RECT 309.190 2559.900 309.510 2559.960 ;
        RECT 309.650 2559.900 309.970 2559.960 ;
        RECT 308.745 2456.400 309.035 2456.445 ;
        RECT 310.110 2456.400 310.430 2456.460 ;
        RECT 308.745 2456.260 310.430 2456.400 ;
        RECT 308.745 2456.215 309.035 2456.260 ;
        RECT 310.110 2456.200 310.430 2456.260 ;
        RECT 308.730 2408.460 309.050 2408.520 ;
        RECT 308.535 2408.320 309.050 2408.460 ;
        RECT 308.730 2408.260 309.050 2408.320 ;
        RECT 309.650 2366.440 309.970 2366.700 ;
        RECT 309.740 2366.300 309.880 2366.440 ;
        RECT 310.570 2366.300 310.890 2366.360 ;
        RECT 309.740 2366.160 310.890 2366.300 ;
        RECT 310.570 2366.100 310.890 2366.160 ;
        RECT 308.730 2235.400 309.050 2235.460 ;
        RECT 310.110 2235.400 310.430 2235.460 ;
        RECT 308.730 2235.260 310.430 2235.400 ;
        RECT 308.730 2235.200 309.050 2235.260 ;
        RECT 310.110 2235.200 310.430 2235.260 ;
        RECT 308.730 2221.800 309.050 2221.860 ;
        RECT 310.110 2221.800 310.430 2221.860 ;
        RECT 308.730 2221.660 310.430 2221.800 ;
        RECT 308.730 2221.600 309.050 2221.660 ;
        RECT 310.110 2221.600 310.430 2221.660 ;
        RECT 309.205 2118.100 309.495 2118.145 ;
        RECT 310.110 2118.100 310.430 2118.160 ;
        RECT 309.205 2117.960 310.430 2118.100 ;
        RECT 309.205 2117.915 309.495 2117.960 ;
        RECT 310.110 2117.900 310.430 2117.960 ;
        RECT 309.190 2070.160 309.510 2070.220 ;
        RECT 308.995 2070.020 309.510 2070.160 ;
        RECT 309.190 2069.960 309.510 2070.020 ;
        RECT 309.190 2046.020 309.510 2046.080 ;
        RECT 310.110 2046.020 310.430 2046.080 ;
        RECT 309.190 2045.880 310.430 2046.020 ;
        RECT 309.190 2045.820 309.510 2045.880 ;
        RECT 310.110 2045.820 310.430 2045.880 ;
        RECT 310.110 1801.220 310.430 1801.280 ;
        RECT 309.740 1801.080 310.430 1801.220 ;
        RECT 309.740 1800.940 309.880 1801.080 ;
        RECT 310.110 1801.020 310.430 1801.080 ;
        RECT 309.650 1800.680 309.970 1800.940 ;
        RECT 309.650 1786.740 309.970 1787.000 ;
        RECT 309.740 1786.600 309.880 1786.740 ;
        RECT 310.110 1786.600 310.430 1786.660 ;
        RECT 309.740 1786.460 310.430 1786.600 ;
        RECT 310.110 1786.400 310.430 1786.460 ;
        RECT 309.650 1594.160 309.970 1594.220 ;
        RECT 310.570 1594.160 310.890 1594.220 ;
        RECT 309.650 1594.020 310.890 1594.160 ;
        RECT 309.650 1593.960 309.970 1594.020 ;
        RECT 310.570 1593.960 310.890 1594.020 ;
        RECT 309.650 1545.880 309.970 1545.940 ;
        RECT 310.110 1545.880 310.430 1545.940 ;
        RECT 309.650 1545.740 310.430 1545.880 ;
        RECT 309.650 1545.680 309.970 1545.740 ;
        RECT 310.110 1545.680 310.430 1545.740 ;
        RECT 310.110 1490.800 310.430 1490.860 ;
        RECT 310.570 1490.800 310.890 1490.860 ;
        RECT 310.110 1490.660 310.890 1490.800 ;
        RECT 310.110 1490.600 310.430 1490.660 ;
        RECT 310.570 1490.600 310.890 1490.660 ;
        RECT 309.650 1401.040 309.970 1401.100 ;
        RECT 310.570 1401.040 310.890 1401.100 ;
        RECT 309.650 1400.900 310.890 1401.040 ;
        RECT 309.650 1400.840 309.970 1400.900 ;
        RECT 310.570 1400.840 310.890 1400.900 ;
        RECT 309.650 1352.760 309.970 1352.820 ;
        RECT 310.110 1352.760 310.430 1352.820 ;
        RECT 309.650 1352.620 310.430 1352.760 ;
        RECT 309.650 1352.560 309.970 1352.620 ;
        RECT 310.110 1352.560 310.430 1352.620 ;
        RECT 309.205 1241.920 309.495 1241.965 ;
        RECT 310.110 1241.920 310.430 1241.980 ;
        RECT 309.205 1241.780 310.430 1241.920 ;
        RECT 309.205 1241.735 309.495 1241.780 ;
        RECT 310.110 1241.720 310.430 1241.780 ;
        RECT 309.190 1193.980 309.510 1194.040 ;
        RECT 308.995 1193.840 309.510 1193.980 ;
        RECT 309.190 1193.780 309.510 1193.840 ;
        RECT 309.190 1128.360 309.510 1128.420 ;
        RECT 310.570 1128.360 310.890 1128.420 ;
        RECT 309.190 1128.220 310.890 1128.360 ;
        RECT 309.190 1128.160 309.510 1128.220 ;
        RECT 310.570 1128.160 310.890 1128.220 ;
        RECT 309.650 917.900 309.970 917.960 ;
        RECT 310.570 917.900 310.890 917.960 ;
        RECT 309.650 917.760 310.890 917.900 ;
        RECT 309.650 917.700 309.970 917.760 ;
        RECT 310.570 917.700 310.890 917.760 ;
        RECT 309.190 796.860 309.510 796.920 ;
        RECT 310.570 796.860 310.890 796.920 ;
        RECT 309.190 796.720 310.890 796.860 ;
        RECT 309.190 796.660 309.510 796.720 ;
        RECT 310.570 796.660 310.890 796.720 ;
        RECT 309.650 724.440 309.970 724.500 ;
        RECT 309.455 724.300 309.970 724.440 ;
        RECT 309.650 724.240 309.970 724.300 ;
        RECT 309.650 699.960 309.970 700.020 ;
        RECT 309.455 699.820 309.970 699.960 ;
        RECT 309.650 699.760 309.970 699.820 ;
        RECT 308.730 627.880 309.050 627.940 ;
        RECT 309.650 627.880 309.970 627.940 ;
        RECT 308.730 627.740 309.970 627.880 ;
        RECT 308.730 627.680 309.050 627.740 ;
        RECT 309.650 627.680 309.970 627.740 ;
        RECT 309.650 435.100 309.970 435.160 ;
        RECT 310.110 435.100 310.430 435.160 ;
        RECT 309.650 434.960 310.430 435.100 ;
        RECT 309.650 434.900 309.970 434.960 ;
        RECT 310.110 434.900 310.430 434.960 ;
        RECT 869.470 241.640 869.790 241.700 ;
        RECT 870.390 241.640 870.710 241.700 ;
        RECT 869.470 241.500 870.710 241.640 ;
        RECT 869.470 241.440 869.790 241.500 ;
        RECT 870.390 241.440 870.710 241.500 ;
        RECT 869.470 193.020 869.790 193.080 ;
        RECT 869.945 193.020 870.235 193.065 ;
        RECT 869.470 192.880 870.235 193.020 ;
        RECT 869.470 192.820 869.790 192.880 ;
        RECT 869.945 192.835 870.235 192.880 ;
        RECT 869.470 145.080 869.790 145.140 ;
        RECT 869.945 145.080 870.235 145.125 ;
        RECT 869.470 144.940 870.235 145.080 ;
        RECT 869.470 144.880 869.790 144.940 ;
        RECT 869.945 144.895 870.235 144.940 ;
        RECT 869.470 96.460 869.790 96.520 ;
        RECT 869.470 96.320 869.985 96.460 ;
        RECT 869.470 96.260 869.790 96.320 ;
        RECT 869.470 48.520 869.790 48.580 ;
        RECT 869.470 48.380 869.985 48.520 ;
        RECT 869.470 48.320 869.790 48.380 ;
      LAYER via ;
        RECT 310.140 3229.020 310.400 3229.280 ;
        RECT 310.140 3181.080 310.400 3181.340 ;
        RECT 309.680 3139.940 309.940 3140.200 ;
        RECT 310.600 3139.940 310.860 3140.200 ;
        RECT 309.680 3132.460 309.940 3132.720 ;
        RECT 309.680 3043.380 309.940 3043.640 ;
        RECT 309.680 2960.080 309.940 2960.340 ;
        RECT 309.680 2939.340 309.940 2939.600 ;
        RECT 309.680 2912.140 309.940 2912.400 ;
        RECT 309.220 2891.060 309.480 2891.320 ;
        RECT 309.220 2814.900 309.480 2815.160 ;
        RECT 310.140 2814.900 310.400 2815.160 ;
        RECT 308.760 2746.220 309.020 2746.480 ;
        RECT 309.680 2746.220 309.940 2746.480 ;
        RECT 308.760 2697.600 309.020 2697.860 ;
        RECT 309.680 2697.600 309.940 2697.860 ;
        RECT 308.300 2649.320 308.560 2649.580 ;
        RECT 309.680 2649.320 309.940 2649.580 ;
        RECT 309.220 2559.900 309.480 2560.160 ;
        RECT 309.680 2559.900 309.940 2560.160 ;
        RECT 310.140 2456.200 310.400 2456.460 ;
        RECT 308.760 2408.260 309.020 2408.520 ;
        RECT 309.680 2366.440 309.940 2366.700 ;
        RECT 310.600 2366.100 310.860 2366.360 ;
        RECT 308.760 2235.200 309.020 2235.460 ;
        RECT 310.140 2235.200 310.400 2235.460 ;
        RECT 308.760 2221.600 309.020 2221.860 ;
        RECT 310.140 2221.600 310.400 2221.860 ;
        RECT 310.140 2117.900 310.400 2118.160 ;
        RECT 309.220 2069.960 309.480 2070.220 ;
        RECT 309.220 2045.820 309.480 2046.080 ;
        RECT 310.140 2045.820 310.400 2046.080 ;
        RECT 310.140 1801.020 310.400 1801.280 ;
        RECT 309.680 1800.680 309.940 1800.940 ;
        RECT 309.680 1786.740 309.940 1787.000 ;
        RECT 310.140 1786.400 310.400 1786.660 ;
        RECT 309.680 1593.960 309.940 1594.220 ;
        RECT 310.600 1593.960 310.860 1594.220 ;
        RECT 309.680 1545.680 309.940 1545.940 ;
        RECT 310.140 1545.680 310.400 1545.940 ;
        RECT 310.140 1490.600 310.400 1490.860 ;
        RECT 310.600 1490.600 310.860 1490.860 ;
        RECT 309.680 1400.840 309.940 1401.100 ;
        RECT 310.600 1400.840 310.860 1401.100 ;
        RECT 309.680 1352.560 309.940 1352.820 ;
        RECT 310.140 1352.560 310.400 1352.820 ;
        RECT 310.140 1241.720 310.400 1241.980 ;
        RECT 309.220 1193.780 309.480 1194.040 ;
        RECT 309.220 1128.160 309.480 1128.420 ;
        RECT 310.600 1128.160 310.860 1128.420 ;
        RECT 309.680 917.700 309.940 917.960 ;
        RECT 310.600 917.700 310.860 917.960 ;
        RECT 309.220 796.660 309.480 796.920 ;
        RECT 310.600 796.660 310.860 796.920 ;
        RECT 309.680 724.240 309.940 724.500 ;
        RECT 309.680 699.760 309.940 700.020 ;
        RECT 308.760 627.680 309.020 627.940 ;
        RECT 309.680 627.680 309.940 627.940 ;
        RECT 309.680 434.900 309.940 435.160 ;
        RECT 310.140 434.900 310.400 435.160 ;
        RECT 869.500 241.440 869.760 241.700 ;
        RECT 870.420 241.440 870.680 241.700 ;
        RECT 869.500 192.820 869.760 193.080 ;
        RECT 869.500 144.880 869.760 145.140 ;
        RECT 869.500 96.260 869.760 96.520 ;
        RECT 869.500 48.320 869.760 48.580 ;
      LAYER met2 ;
        RECT 1518.550 3261.435 1518.830 3261.805 ;
        RECT 1518.620 3259.650 1518.760 3261.435 ;
        RECT 1519.890 3259.650 1520.170 3260.000 ;
        RECT 1518.620 3259.510 1520.170 3259.650 ;
        RECT 1519.890 3256.000 1520.170 3259.510 ;
        RECT 312.890 3251.915 313.170 3252.285 ;
        RECT 312.960 3237.325 313.100 3251.915 ;
        RECT 312.890 3236.955 313.170 3237.325 ;
        RECT 310.130 3236.275 310.410 3236.645 ;
        RECT 310.200 3229.310 310.340 3236.275 ;
        RECT 310.140 3228.990 310.400 3229.310 ;
        RECT 310.140 3181.050 310.400 3181.370 ;
        RECT 310.200 3154.250 310.340 3181.050 ;
        RECT 310.200 3154.110 310.800 3154.250 ;
        RECT 310.660 3140.230 310.800 3154.110 ;
        RECT 309.680 3139.910 309.940 3140.230 ;
        RECT 310.600 3139.910 310.860 3140.230 ;
        RECT 309.740 3132.750 309.880 3139.910 ;
        RECT 309.680 3132.430 309.940 3132.750 ;
        RECT 309.680 3043.350 309.940 3043.670 ;
        RECT 309.740 3012.130 309.880 3043.350 ;
        RECT 309.280 3011.990 309.880 3012.130 ;
        RECT 309.280 3008.050 309.420 3011.990 ;
        RECT 309.280 3007.910 309.880 3008.050 ;
        RECT 309.740 2960.370 309.880 3007.910 ;
        RECT 309.680 2960.050 309.940 2960.370 ;
        RECT 309.680 2939.310 309.940 2939.630 ;
        RECT 309.740 2912.430 309.880 2939.310 ;
        RECT 309.680 2912.110 309.940 2912.430 ;
        RECT 309.220 2891.030 309.480 2891.350 ;
        RECT 309.280 2815.190 309.420 2891.030 ;
        RECT 309.220 2814.870 309.480 2815.190 ;
        RECT 310.140 2814.870 310.400 2815.190 ;
        RECT 310.200 2794.530 310.340 2814.870 ;
        RECT 309.740 2794.390 310.340 2794.530 ;
        RECT 308.820 2746.510 308.960 2746.665 ;
        RECT 309.740 2746.510 309.880 2794.390 ;
        RECT 308.760 2746.250 309.020 2746.510 ;
        RECT 309.680 2746.250 309.940 2746.510 ;
        RECT 308.760 2746.190 309.940 2746.250 ;
        RECT 308.820 2746.110 309.880 2746.190 ;
        RECT 309.740 2697.890 309.880 2746.110 ;
        RECT 308.760 2697.570 309.020 2697.890 ;
        RECT 309.680 2697.570 309.940 2697.890 ;
        RECT 308.820 2649.805 308.960 2697.570 ;
        RECT 308.300 2649.290 308.560 2649.610 ;
        RECT 308.750 2649.435 309.030 2649.805 ;
        RECT 309.670 2649.435 309.950 2649.805 ;
        RECT 309.680 2649.290 309.940 2649.435 ;
        RECT 308.360 2601.525 308.500 2649.290 ;
        RECT 308.290 2601.155 308.570 2601.525 ;
        RECT 309.210 2601.155 309.490 2601.525 ;
        RECT 309.280 2560.190 309.420 2601.155 ;
        RECT 309.220 2559.870 309.480 2560.190 ;
        RECT 309.680 2559.870 309.940 2560.190 ;
        RECT 309.740 2536.810 309.880 2559.870 ;
        RECT 309.280 2536.670 309.880 2536.810 ;
        RECT 309.280 2535.450 309.420 2536.670 ;
        RECT 309.280 2535.310 310.340 2535.450 ;
        RECT 310.200 2456.490 310.340 2535.310 ;
        RECT 310.140 2456.170 310.400 2456.490 ;
        RECT 308.760 2408.230 309.020 2408.550 ;
        RECT 308.820 2366.925 308.960 2408.230 ;
        RECT 308.750 2366.555 309.030 2366.925 ;
        RECT 309.670 2366.555 309.950 2366.925 ;
        RECT 309.680 2366.410 309.940 2366.555 ;
        RECT 310.600 2366.070 310.860 2366.390 ;
        RECT 310.660 2332.130 310.800 2366.070 ;
        RECT 310.200 2331.990 310.800 2332.130 ;
        RECT 310.200 2294.050 310.340 2331.990 ;
        RECT 308.820 2293.910 310.340 2294.050 ;
        RECT 308.820 2235.490 308.960 2293.910 ;
        RECT 308.760 2235.170 309.020 2235.490 ;
        RECT 310.140 2235.170 310.400 2235.490 ;
        RECT 310.200 2221.890 310.340 2235.170 ;
        RECT 308.760 2221.570 309.020 2221.890 ;
        RECT 310.140 2221.570 310.400 2221.890 ;
        RECT 308.820 2173.805 308.960 2221.570 ;
        RECT 308.750 2173.435 309.030 2173.805 ;
        RECT 309.670 2173.435 309.950 2173.805 ;
        RECT 309.740 2149.210 309.880 2173.435 ;
        RECT 309.740 2149.070 310.800 2149.210 ;
        RECT 310.660 2126.205 310.800 2149.070 ;
        RECT 310.590 2125.835 310.870 2126.205 ;
        RECT 310.130 2125.155 310.410 2125.525 ;
        RECT 310.200 2118.190 310.340 2125.155 ;
        RECT 310.140 2117.870 310.400 2118.190 ;
        RECT 309.220 2069.930 309.480 2070.250 ;
        RECT 309.280 2046.110 309.420 2069.930 ;
        RECT 309.220 2045.790 309.480 2046.110 ;
        RECT 310.140 2045.790 310.400 2046.110 ;
        RECT 310.200 2004.370 310.340 2045.790 ;
        RECT 309.740 2004.230 310.340 2004.370 ;
        RECT 309.740 1956.090 309.880 2004.230 ;
        RECT 309.740 1955.950 310.340 1956.090 ;
        RECT 310.200 1897.610 310.340 1955.950 ;
        RECT 309.740 1897.470 310.340 1897.610 ;
        RECT 309.740 1859.530 309.880 1897.470 ;
        RECT 309.740 1859.390 310.340 1859.530 ;
        RECT 310.200 1801.310 310.340 1859.390 ;
        RECT 310.140 1800.990 310.400 1801.310 ;
        RECT 309.680 1800.650 309.940 1800.970 ;
        RECT 309.740 1787.030 309.880 1800.650 ;
        RECT 309.680 1786.710 309.940 1787.030 ;
        RECT 310.140 1786.370 310.400 1786.690 ;
        RECT 310.200 1643.405 310.340 1786.370 ;
        RECT 310.130 1643.035 310.410 1643.405 ;
        RECT 310.590 1641.675 310.870 1642.045 ;
        RECT 310.660 1594.250 310.800 1641.675 ;
        RECT 309.680 1593.930 309.940 1594.250 ;
        RECT 310.600 1593.930 310.860 1594.250 ;
        RECT 309.740 1545.970 309.880 1593.930 ;
        RECT 309.680 1545.650 309.940 1545.970 ;
        RECT 310.140 1545.650 310.400 1545.970 ;
        RECT 310.200 1490.890 310.340 1545.650 ;
        RECT 310.140 1490.570 310.400 1490.890 ;
        RECT 310.600 1490.570 310.860 1490.890 ;
        RECT 310.660 1401.130 310.800 1490.570 ;
        RECT 309.680 1400.810 309.940 1401.130 ;
        RECT 310.600 1400.810 310.860 1401.130 ;
        RECT 309.740 1352.850 309.880 1400.810 ;
        RECT 309.680 1352.530 309.940 1352.850 ;
        RECT 310.140 1352.530 310.400 1352.850 ;
        RECT 310.200 1242.010 310.340 1352.530 ;
        RECT 310.140 1241.690 310.400 1242.010 ;
        RECT 309.220 1193.750 309.480 1194.070 ;
        RECT 309.280 1158.450 309.420 1193.750 ;
        RECT 309.280 1158.310 309.880 1158.450 ;
        RECT 309.740 1157.090 309.880 1158.310 ;
        RECT 309.280 1156.950 309.880 1157.090 ;
        RECT 309.280 1128.450 309.420 1156.950 ;
        RECT 309.220 1128.130 309.480 1128.450 ;
        RECT 310.600 1128.130 310.860 1128.450 ;
        RECT 310.660 917.990 310.800 1128.130 ;
        RECT 309.680 917.845 309.940 917.990 ;
        RECT 310.600 917.845 310.860 917.990 ;
        RECT 309.670 917.475 309.950 917.845 ;
        RECT 310.590 917.475 310.870 917.845 ;
        RECT 310.660 869.620 310.800 917.475 ;
        RECT 310.200 869.480 310.800 869.620 ;
        RECT 310.200 845.650 310.340 869.480 ;
        RECT 309.280 845.510 310.340 845.650 ;
        RECT 309.280 796.950 309.420 845.510 ;
        RECT 309.220 796.630 309.480 796.950 ;
        RECT 310.600 796.630 310.860 796.950 ;
        RECT 310.660 724.725 310.800 796.630 ;
        RECT 309.670 724.355 309.950 724.725 ;
        RECT 310.590 724.355 310.870 724.725 ;
        RECT 309.680 724.210 309.940 724.355 ;
        RECT 309.680 699.730 309.940 700.050 ;
        RECT 309.740 676.330 309.880 699.730 ;
        RECT 309.740 676.190 310.340 676.330 ;
        RECT 310.200 628.050 310.340 676.190 ;
        RECT 309.740 627.970 310.340 628.050 ;
        RECT 308.760 627.650 309.020 627.970 ;
        RECT 309.680 627.910 310.340 627.970 ;
        RECT 309.680 627.650 309.940 627.910 ;
        RECT 308.820 579.885 308.960 627.650 ;
        RECT 308.750 579.515 309.030 579.885 ;
        RECT 310.130 579.515 310.410 579.885 ;
        RECT 310.200 531.490 310.340 579.515 ;
        RECT 309.740 531.350 310.340 531.490 ;
        RECT 309.740 507.010 309.880 531.350 ;
        RECT 309.740 506.870 310.340 507.010 ;
        RECT 310.200 496.130 310.340 506.870 ;
        RECT 309.740 495.990 310.340 496.130 ;
        RECT 309.740 483.325 309.880 495.990 ;
        RECT 309.670 482.955 309.950 483.325 ;
        RECT 309.670 482.275 309.950 482.645 ;
        RECT 309.740 435.190 309.880 482.275 ;
        RECT 309.680 434.870 309.940 435.190 ;
        RECT 310.140 434.870 310.400 435.190 ;
        RECT 310.200 410.450 310.340 434.870 ;
        RECT 309.740 410.310 310.340 410.450 ;
        RECT 309.740 365.685 309.880 410.310 ;
        RECT 309.670 365.315 309.950 365.685 ;
        RECT 870.410 244.955 870.690 245.325 ;
        RECT 870.480 241.730 870.620 244.955 ;
        RECT 869.500 241.410 869.760 241.730 ;
        RECT 870.420 241.410 870.680 241.730 ;
        RECT 869.560 193.110 869.700 241.410 ;
        RECT 869.500 192.790 869.760 193.110 ;
        RECT 869.500 144.850 869.760 145.170 ;
        RECT 869.560 96.550 869.700 144.850 ;
        RECT 869.500 96.230 869.760 96.550 ;
        RECT 869.500 48.290 869.760 48.610 ;
        RECT 869.560 14.180 869.700 48.290 ;
        RECT 869.560 14.040 870.160 14.180 ;
        RECT 870.020 13.330 870.160 14.040 ;
        RECT 870.020 13.190 871.080 13.330 ;
        RECT 870.940 2.400 871.080 13.190 ;
        RECT 870.730 -4.800 871.290 2.400 ;
      LAYER via2 ;
        RECT 1518.550 3261.480 1518.830 3261.760 ;
        RECT 312.890 3251.960 313.170 3252.240 ;
        RECT 312.890 3237.000 313.170 3237.280 ;
        RECT 310.130 3236.320 310.410 3236.600 ;
        RECT 308.750 2649.480 309.030 2649.760 ;
        RECT 309.670 2649.480 309.950 2649.760 ;
        RECT 308.290 2601.200 308.570 2601.480 ;
        RECT 309.210 2601.200 309.490 2601.480 ;
        RECT 308.750 2366.600 309.030 2366.880 ;
        RECT 309.670 2366.600 309.950 2366.880 ;
        RECT 308.750 2173.480 309.030 2173.760 ;
        RECT 309.670 2173.480 309.950 2173.760 ;
        RECT 310.590 2125.880 310.870 2126.160 ;
        RECT 310.130 2125.200 310.410 2125.480 ;
        RECT 310.130 1643.080 310.410 1643.360 ;
        RECT 310.590 1641.720 310.870 1642.000 ;
        RECT 309.670 917.520 309.950 917.800 ;
        RECT 310.590 917.520 310.870 917.800 ;
        RECT 309.670 724.400 309.950 724.680 ;
        RECT 310.590 724.400 310.870 724.680 ;
        RECT 308.750 579.560 309.030 579.840 ;
        RECT 310.130 579.560 310.410 579.840 ;
        RECT 309.670 483.000 309.950 483.280 ;
        RECT 309.670 482.320 309.950 482.600 ;
        RECT 309.670 365.360 309.950 365.640 ;
        RECT 870.410 245.000 870.690 245.280 ;
      LAYER met3 ;
        RECT 1518.525 3261.780 1518.855 3261.785 ;
        RECT 1518.270 3261.770 1518.855 3261.780 ;
        RECT 1518.070 3261.470 1518.855 3261.770 ;
        RECT 1518.270 3261.460 1518.855 3261.470 ;
        RECT 1518.525 3261.455 1518.855 3261.460 ;
        RECT 312.865 3252.250 313.195 3252.265 ;
        RECT 1518.270 3252.250 1518.650 3252.260 ;
        RECT 312.865 3251.950 1518.650 3252.250 ;
        RECT 312.865 3251.935 313.195 3251.950 ;
        RECT 1518.270 3251.940 1518.650 3251.950 ;
        RECT 312.865 3237.290 313.195 3237.305 ;
        RECT 310.120 3236.990 313.195 3237.290 ;
        RECT 310.120 3236.625 310.420 3236.990 ;
        RECT 312.865 3236.975 313.195 3236.990 ;
        RECT 310.105 3236.295 310.435 3236.625 ;
        RECT 308.725 2649.770 309.055 2649.785 ;
        RECT 309.645 2649.770 309.975 2649.785 ;
        RECT 308.725 2649.470 309.975 2649.770 ;
        RECT 308.725 2649.455 309.055 2649.470 ;
        RECT 309.645 2649.455 309.975 2649.470 ;
        RECT 308.265 2601.490 308.595 2601.505 ;
        RECT 309.185 2601.490 309.515 2601.505 ;
        RECT 308.265 2601.190 309.515 2601.490 ;
        RECT 308.265 2601.175 308.595 2601.190 ;
        RECT 309.185 2601.175 309.515 2601.190 ;
        RECT 308.725 2366.890 309.055 2366.905 ;
        RECT 309.645 2366.890 309.975 2366.905 ;
        RECT 308.725 2366.590 309.975 2366.890 ;
        RECT 308.725 2366.575 309.055 2366.590 ;
        RECT 309.645 2366.575 309.975 2366.590 ;
        RECT 308.725 2173.770 309.055 2173.785 ;
        RECT 309.645 2173.770 309.975 2173.785 ;
        RECT 308.725 2173.470 309.975 2173.770 ;
        RECT 308.725 2173.455 309.055 2173.470 ;
        RECT 309.645 2173.455 309.975 2173.470 ;
        RECT 310.565 2126.170 310.895 2126.185 ;
        RECT 310.350 2125.855 310.895 2126.170 ;
        RECT 310.350 2125.505 310.650 2125.855 ;
        RECT 310.105 2125.190 310.650 2125.505 ;
        RECT 310.105 2125.175 310.435 2125.190 ;
        RECT 310.105 1643.370 310.435 1643.385 ;
        RECT 310.105 1643.055 310.650 1643.370 ;
        RECT 310.350 1642.025 310.650 1643.055 ;
        RECT 310.350 1641.710 310.895 1642.025 ;
        RECT 310.565 1641.695 310.895 1641.710 ;
        RECT 309.645 917.810 309.975 917.825 ;
        RECT 310.565 917.810 310.895 917.825 ;
        RECT 309.645 917.510 310.895 917.810 ;
        RECT 309.645 917.495 309.975 917.510 ;
        RECT 310.565 917.495 310.895 917.510 ;
        RECT 309.645 724.690 309.975 724.705 ;
        RECT 310.565 724.690 310.895 724.705 ;
        RECT 309.645 724.390 310.895 724.690 ;
        RECT 309.645 724.375 309.975 724.390 ;
        RECT 310.565 724.375 310.895 724.390 ;
        RECT 308.725 579.850 309.055 579.865 ;
        RECT 310.105 579.850 310.435 579.865 ;
        RECT 308.725 579.550 310.435 579.850 ;
        RECT 308.725 579.535 309.055 579.550 ;
        RECT 310.105 579.535 310.435 579.550 ;
        RECT 309.645 483.290 309.975 483.305 ;
        RECT 309.645 482.990 310.650 483.290 ;
        RECT 309.645 482.975 309.975 482.990 ;
        RECT 309.645 482.610 309.975 482.625 ;
        RECT 310.350 482.610 310.650 482.990 ;
        RECT 309.645 482.310 310.650 482.610 ;
        RECT 309.645 482.295 309.975 482.310 ;
        RECT 309.645 365.650 309.975 365.665 ;
        RECT 313.070 365.650 313.450 365.660 ;
        RECT 309.645 365.350 313.450 365.650 ;
        RECT 309.645 365.335 309.975 365.350 ;
        RECT 313.070 365.340 313.450 365.350 ;
        RECT 315.830 245.290 316.210 245.300 ;
        RECT 870.385 245.290 870.715 245.305 ;
        RECT 315.830 244.990 870.715 245.290 ;
        RECT 315.830 244.980 316.210 244.990 ;
        RECT 870.385 244.975 870.715 244.990 ;
      LAYER via3 ;
        RECT 1518.300 3261.460 1518.620 3261.780 ;
        RECT 1518.300 3251.940 1518.620 3252.260 ;
        RECT 313.100 365.340 313.420 365.660 ;
        RECT 315.860 244.980 316.180 245.300 ;
      LAYER met4 ;
        RECT 1518.295 3261.455 1518.625 3261.785 ;
        RECT 1518.310 3252.265 1518.610 3261.455 ;
        RECT 1518.295 3251.935 1518.625 3252.265 ;
        RECT 313.095 365.650 313.425 365.665 ;
        RECT 313.095 365.350 314.330 365.650 ;
        RECT 313.095 365.335 313.425 365.350 ;
        RECT 314.030 355.450 314.330 365.350 ;
        RECT 314.030 355.150 316.170 355.450 ;
        RECT 315.870 245.305 316.170 355.150 ;
        RECT 315.855 244.975 316.185 245.305 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 309.265 252.025 309.435 289.595 ;
      LAYER mcon ;
        RECT 309.265 289.425 309.435 289.595 ;
      LAYER met1 ;
        RECT 309.190 289.580 309.510 289.640 ;
        RECT 308.995 289.440 309.510 289.580 ;
        RECT 309.190 289.380 309.510 289.440 ;
        RECT 309.205 252.180 309.495 252.225 ;
        RECT 883.730 252.180 884.050 252.240 ;
        RECT 309.205 252.040 884.050 252.180 ;
        RECT 309.205 251.995 309.495 252.040 ;
        RECT 883.730 251.980 884.050 252.040 ;
        RECT 883.730 20.640 884.050 20.700 ;
        RECT 888.790 20.640 889.110 20.700 ;
        RECT 883.730 20.500 889.110 20.640 ;
        RECT 883.730 20.440 884.050 20.500 ;
        RECT 888.790 20.440 889.110 20.500 ;
      LAYER via ;
        RECT 309.220 289.380 309.480 289.640 ;
        RECT 883.760 251.980 884.020 252.240 ;
        RECT 883.760 20.440 884.020 20.700 ;
        RECT 888.820 20.440 889.080 20.700 ;
      LAYER met2 ;
        RECT 1732.450 3261.435 1732.730 3261.805 ;
        RECT 1732.520 3259.650 1732.660 3261.435 ;
        RECT 1734.250 3259.650 1734.530 3260.000 ;
        RECT 1732.520 3259.510 1734.530 3259.650 ;
        RECT 1734.250 3256.000 1734.530 3259.510 ;
        RECT 309.210 372.115 309.490 372.485 ;
        RECT 309.280 289.670 309.420 372.115 ;
        RECT 309.220 289.350 309.480 289.670 ;
        RECT 883.760 251.950 884.020 252.270 ;
        RECT 883.820 20.730 883.960 251.950 ;
        RECT 883.760 20.410 884.020 20.730 ;
        RECT 888.820 20.410 889.080 20.730 ;
        RECT 888.880 2.400 889.020 20.410 ;
        RECT 888.670 -4.800 889.230 2.400 ;
      LAYER via2 ;
        RECT 1732.450 3261.480 1732.730 3261.760 ;
        RECT 309.210 372.160 309.490 372.440 ;
      LAYER met3 ;
        RECT 1730.790 3261.770 1731.170 3261.780 ;
        RECT 1732.425 3261.770 1732.755 3261.785 ;
        RECT 1730.790 3261.470 1732.755 3261.770 ;
        RECT 1730.790 3261.460 1731.170 3261.470 ;
        RECT 1732.425 3261.455 1732.755 3261.470 ;
        RECT 299.270 3251.570 299.650 3251.580 ;
        RECT 1730.790 3251.570 1731.170 3251.580 ;
        RECT 299.270 3251.270 1731.170 3251.570 ;
        RECT 299.270 3251.260 299.650 3251.270 ;
        RECT 1730.790 3251.260 1731.170 3251.270 ;
        RECT 299.270 555.370 299.650 555.380 ;
        RECT 311.230 555.370 311.610 555.380 ;
        RECT 299.270 555.070 311.610 555.370 ;
        RECT 299.270 555.060 299.650 555.070 ;
        RECT 311.230 555.060 311.610 555.070 ;
        RECT 309.185 372.450 309.515 372.465 ;
        RECT 311.230 372.450 311.610 372.460 ;
        RECT 309.185 372.150 311.610 372.450 ;
        RECT 309.185 372.135 309.515 372.150 ;
        RECT 311.230 372.140 311.610 372.150 ;
      LAYER via3 ;
        RECT 1730.820 3261.460 1731.140 3261.780 ;
        RECT 299.300 3251.260 299.620 3251.580 ;
        RECT 1730.820 3251.260 1731.140 3251.580 ;
        RECT 299.300 555.060 299.620 555.380 ;
        RECT 311.260 555.060 311.580 555.380 ;
        RECT 311.260 372.140 311.580 372.460 ;
      LAYER met4 ;
        RECT 1730.815 3261.455 1731.145 3261.785 ;
        RECT 1730.830 3251.585 1731.130 3261.455 ;
        RECT 299.295 3251.255 299.625 3251.585 ;
        RECT 1730.815 3251.255 1731.145 3251.585 ;
        RECT 299.310 555.385 299.610 3251.255 ;
        RECT 299.295 555.055 299.625 555.385 ;
        RECT 311.255 555.055 311.585 555.385 ;
        RECT 311.270 372.465 311.570 555.055 ;
        RECT 311.255 372.135 311.585 372.465 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 910.410 204.240 910.730 204.300 ;
        RECT 1297.270 204.240 1297.590 204.300 ;
        RECT 910.410 204.100 1297.590 204.240 ;
        RECT 910.410 204.040 910.730 204.100 ;
        RECT 1297.270 204.040 1297.590 204.100 ;
        RECT 906.730 20.640 907.050 20.700 ;
        RECT 910.410 20.640 910.730 20.700 ;
        RECT 906.730 20.500 910.730 20.640 ;
        RECT 906.730 20.440 907.050 20.500 ;
        RECT 910.410 20.440 910.730 20.500 ;
      LAYER via ;
        RECT 910.440 204.040 910.700 204.300 ;
        RECT 1297.300 204.040 1297.560 204.300 ;
        RECT 906.760 20.440 907.020 20.700 ;
        RECT 910.440 20.440 910.700 20.700 ;
      LAYER met2 ;
        RECT 1299.090 260.170 1299.370 264.000 ;
        RECT 1297.360 260.030 1299.370 260.170 ;
        RECT 1297.360 204.330 1297.500 260.030 ;
        RECT 1299.090 260.000 1299.370 260.030 ;
        RECT 910.440 204.010 910.700 204.330 ;
        RECT 1297.300 204.010 1297.560 204.330 ;
        RECT 910.500 20.730 910.640 204.010 ;
        RECT 906.760 20.410 907.020 20.730 ;
        RECT 910.440 20.410 910.700 20.730 ;
        RECT 906.820 2.400 906.960 20.410 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.630 310.660 2615.950 310.720 ;
        RECT 2642.770 310.660 2643.090 310.720 ;
        RECT 2615.630 310.520 2643.090 310.660 ;
        RECT 2615.630 310.460 2615.950 310.520 ;
        RECT 2642.770 310.460 2643.090 310.520 ;
        RECT 924.210 224.640 924.530 224.700 ;
        RECT 2642.770 224.640 2643.090 224.700 ;
        RECT 924.210 224.500 2643.090 224.640 ;
        RECT 924.210 224.440 924.530 224.500 ;
        RECT 2642.770 224.440 2643.090 224.500 ;
      LAYER via ;
        RECT 2615.660 310.460 2615.920 310.720 ;
        RECT 2642.800 310.460 2643.060 310.720 ;
        RECT 924.240 224.440 924.500 224.700 ;
        RECT 2642.800 224.440 2643.060 224.700 ;
      LAYER met2 ;
        RECT 2615.650 317.035 2615.930 317.405 ;
        RECT 2615.720 310.750 2615.860 317.035 ;
        RECT 2615.660 310.430 2615.920 310.750 ;
        RECT 2642.800 310.430 2643.060 310.750 ;
        RECT 2642.860 224.730 2643.000 310.430 ;
        RECT 924.240 224.410 924.500 224.730 ;
        RECT 2642.800 224.410 2643.060 224.730 ;
        RECT 924.300 2.400 924.440 224.410 ;
        RECT 924.090 -4.800 924.650 2.400 ;
      LAYER via2 ;
        RECT 2615.650 317.080 2615.930 317.360 ;
      LAYER met3 ;
        RECT 2606.000 317.370 2610.000 317.760 ;
        RECT 2615.625 317.370 2615.955 317.385 ;
        RECT 2606.000 317.160 2615.955 317.370 ;
        RECT 2609.580 317.070 2615.955 317.160 ;
        RECT 2615.625 317.055 2615.955 317.070 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 247.090 3278.520 247.410 3278.580 ;
        RECT 761.830 3278.520 762.150 3278.580 ;
        RECT 247.090 3278.380 762.150 3278.520 ;
        RECT 247.090 3278.320 247.410 3278.380 ;
        RECT 761.830 3278.320 762.150 3278.380 ;
        RECT 247.090 44.100 247.410 44.160 ;
        RECT 942.150 44.100 942.470 44.160 ;
        RECT 247.090 43.960 942.470 44.100 ;
        RECT 247.090 43.900 247.410 43.960 ;
        RECT 942.150 43.900 942.470 43.960 ;
      LAYER via ;
        RECT 247.120 3278.320 247.380 3278.580 ;
        RECT 761.860 3278.320 762.120 3278.580 ;
        RECT 247.120 43.900 247.380 44.160 ;
        RECT 942.180 43.900 942.440 44.160 ;
      LAYER met2 ;
        RECT 247.120 3278.290 247.380 3278.610 ;
        RECT 761.860 3278.290 762.120 3278.610 ;
        RECT 247.180 44.190 247.320 3278.290 ;
        RECT 761.920 3260.000 762.060 3278.290 ;
        RECT 761.810 3256.000 762.090 3260.000 ;
        RECT 247.120 43.870 247.380 44.190 ;
        RECT 942.180 43.870 942.440 44.190 ;
        RECT 942.240 2.400 942.380 43.870 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 33.220 960.410 33.280 ;
        RECT 2139.070 33.220 2139.390 33.280 ;
        RECT 960.090 33.080 2139.390 33.220 ;
        RECT 960.090 33.020 960.410 33.080 ;
        RECT 2139.070 33.020 2139.390 33.080 ;
      LAYER via ;
        RECT 960.120 33.020 960.380 33.280 ;
        RECT 2139.100 33.020 2139.360 33.280 ;
      LAYER met2 ;
        RECT 2142.730 260.170 2143.010 264.000 ;
        RECT 2139.160 260.030 2143.010 260.170 ;
        RECT 2139.160 33.310 2139.300 260.030 ;
        RECT 2142.730 260.000 2143.010 260.030 ;
        RECT 960.120 32.990 960.380 33.310 ;
        RECT 2139.100 32.990 2139.360 33.310 ;
        RECT 960.180 2.400 960.320 32.990 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 979.485 144.925 979.655 193.035 ;
        RECT 979.485 48.365 979.655 96.475 ;
      LAYER mcon ;
        RECT 979.485 192.865 979.655 193.035 ;
        RECT 979.485 96.305 979.655 96.475 ;
      LAYER met1 ;
        RECT 2615.170 2615.180 2615.490 2615.240 ;
        RECT 2692.450 2615.180 2692.770 2615.240 ;
        RECT 2615.170 2615.040 2692.770 2615.180 ;
        RECT 2615.170 2614.980 2615.490 2615.040 ;
        RECT 2692.450 2614.980 2692.770 2615.040 ;
        RECT 978.950 224.980 979.270 225.040 ;
        RECT 2692.450 224.980 2692.770 225.040 ;
        RECT 978.950 224.840 2692.770 224.980 ;
        RECT 978.950 224.780 979.270 224.840 ;
        RECT 2692.450 224.780 2692.770 224.840 ;
        RECT 979.410 193.020 979.730 193.080 ;
        RECT 979.215 192.880 979.730 193.020 ;
        RECT 979.410 192.820 979.730 192.880 ;
        RECT 979.410 145.080 979.730 145.140 ;
        RECT 979.215 144.940 979.730 145.080 ;
        RECT 979.410 144.880 979.730 144.940 ;
        RECT 979.410 96.460 979.730 96.520 ;
        RECT 979.215 96.320 979.730 96.460 ;
        RECT 979.410 96.260 979.730 96.320 ;
        RECT 979.410 48.520 979.730 48.580 ;
        RECT 979.215 48.380 979.730 48.520 ;
        RECT 979.410 48.320 979.730 48.380 ;
      LAYER via ;
        RECT 2615.200 2614.980 2615.460 2615.240 ;
        RECT 2692.480 2614.980 2692.740 2615.240 ;
        RECT 978.980 224.780 979.240 225.040 ;
        RECT 2692.480 224.780 2692.740 225.040 ;
        RECT 979.440 192.820 979.700 193.080 ;
        RECT 979.440 144.880 979.700 145.140 ;
        RECT 979.440 96.260 979.700 96.520 ;
        RECT 979.440 48.320 979.700 48.580 ;
      LAYER met2 ;
        RECT 2615.190 2620.875 2615.470 2621.245 ;
        RECT 2615.260 2615.270 2615.400 2620.875 ;
        RECT 2615.200 2614.950 2615.460 2615.270 ;
        RECT 2692.480 2614.950 2692.740 2615.270 ;
        RECT 2692.540 225.070 2692.680 2614.950 ;
        RECT 978.980 224.750 979.240 225.070 ;
        RECT 2692.480 224.750 2692.740 225.070 ;
        RECT 979.040 193.530 979.180 224.750 ;
        RECT 979.040 193.390 979.640 193.530 ;
        RECT 979.500 193.110 979.640 193.390 ;
        RECT 979.440 192.790 979.700 193.110 ;
        RECT 979.440 144.850 979.700 145.170 ;
        RECT 979.500 96.550 979.640 144.850 ;
        RECT 979.440 96.230 979.700 96.550 ;
        RECT 979.440 48.290 979.700 48.610 ;
        RECT 979.500 14.010 979.640 48.290 ;
        RECT 979.040 13.870 979.640 14.010 ;
        RECT 979.040 12.650 979.180 13.870 ;
        RECT 978.120 12.510 979.180 12.650 ;
        RECT 978.120 2.400 978.260 12.510 ;
        RECT 977.910 -4.800 978.470 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2620.920 2615.470 2621.200 ;
      LAYER met3 ;
        RECT 2606.000 2621.210 2610.000 2621.600 ;
        RECT 2615.165 2621.210 2615.495 2621.225 ;
        RECT 2606.000 2621.000 2615.495 2621.210 ;
        RECT 2609.580 2620.910 2615.495 2621.000 ;
        RECT 2615.165 2620.895 2615.495 2620.910 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 655.645 145.265 655.815 193.035 ;
        RECT 655.645 57.205 655.815 96.475 ;
      LAYER mcon ;
        RECT 655.645 192.865 655.815 193.035 ;
        RECT 655.645 96.305 655.815 96.475 ;
      LAYER met1 ;
        RECT 303.210 3259.820 303.530 3259.880 ;
        RECT 1332.230 3259.820 1332.550 3259.880 ;
        RECT 303.210 3259.680 1332.550 3259.820 ;
        RECT 303.210 3259.620 303.530 3259.680 ;
        RECT 1332.230 3259.620 1332.550 3259.680 ;
        RECT 303.210 600.680 303.530 600.740 ;
        RECT 304.590 600.680 304.910 600.740 ;
        RECT 303.210 600.540 304.910 600.680 ;
        RECT 303.210 600.480 303.530 600.540 ;
        RECT 304.590 600.480 304.910 600.540 ;
        RECT 282.510 475.900 282.830 475.960 ;
        RECT 304.590 475.900 304.910 475.960 ;
        RECT 282.510 475.760 304.910 475.900 ;
        RECT 282.510 475.700 282.830 475.760 ;
        RECT 304.590 475.700 304.910 475.760 ;
        RECT 282.510 379.680 282.830 379.740 ;
        RECT 286.190 379.680 286.510 379.740 ;
        RECT 282.510 379.540 286.510 379.680 ;
        RECT 282.510 379.480 282.830 379.540 ;
        RECT 286.190 379.480 286.510 379.540 ;
        RECT 655.570 193.020 655.890 193.080 ;
        RECT 655.375 192.880 655.890 193.020 ;
        RECT 655.570 192.820 655.890 192.880 ;
        RECT 655.570 145.420 655.890 145.480 ;
        RECT 655.375 145.280 655.890 145.420 ;
        RECT 655.570 145.220 655.890 145.280 ;
        RECT 655.570 144.740 655.890 144.800 ;
        RECT 656.490 144.740 656.810 144.800 ;
        RECT 655.570 144.600 656.810 144.740 ;
        RECT 655.570 144.540 655.890 144.600 ;
        RECT 656.490 144.540 656.810 144.600 ;
        RECT 655.570 96.460 655.890 96.520 ;
        RECT 655.375 96.320 655.890 96.460 ;
        RECT 655.570 96.260 655.890 96.320 ;
        RECT 655.585 57.360 655.875 57.405 ;
        RECT 656.950 57.360 657.270 57.420 ;
        RECT 655.585 57.220 657.270 57.360 ;
        RECT 655.585 57.175 655.875 57.220 ;
        RECT 656.950 57.160 657.270 57.220 ;
      LAYER via ;
        RECT 303.240 3259.620 303.500 3259.880 ;
        RECT 1332.260 3259.620 1332.520 3259.880 ;
        RECT 303.240 600.480 303.500 600.740 ;
        RECT 304.620 600.480 304.880 600.740 ;
        RECT 282.540 475.700 282.800 475.960 ;
        RECT 304.620 475.700 304.880 475.960 ;
        RECT 282.540 379.480 282.800 379.740 ;
        RECT 286.220 379.480 286.480 379.740 ;
        RECT 655.600 192.820 655.860 193.080 ;
        RECT 655.600 145.220 655.860 145.480 ;
        RECT 655.600 144.540 655.860 144.800 ;
        RECT 656.520 144.540 656.780 144.800 ;
        RECT 655.600 96.260 655.860 96.520 ;
        RECT 656.980 57.160 657.240 57.420 ;
      LAYER met2 ;
        RECT 303.240 3259.590 303.500 3259.910 ;
        RECT 1332.260 3259.650 1332.520 3259.910 ;
        RECT 1334.050 3259.650 1334.330 3260.000 ;
        RECT 1332.260 3259.590 1334.330 3259.650 ;
        RECT 303.300 600.770 303.440 3259.590 ;
        RECT 1332.320 3259.510 1334.330 3259.590 ;
        RECT 1334.050 3256.000 1334.330 3259.510 ;
        RECT 303.240 600.450 303.500 600.770 ;
        RECT 304.620 600.450 304.880 600.770 ;
        RECT 304.680 475.990 304.820 600.450 ;
        RECT 282.540 475.670 282.800 475.990 ;
        RECT 304.620 475.670 304.880 475.990 ;
        RECT 282.600 379.770 282.740 475.670 ;
        RECT 282.540 379.450 282.800 379.770 ;
        RECT 286.220 379.450 286.480 379.770 ;
        RECT 286.280 263.005 286.420 379.450 ;
        RECT 286.210 262.635 286.490 263.005 ;
        RECT 654.210 262.890 654.490 263.005 ;
        RECT 654.210 262.750 655.800 262.890 ;
        RECT 654.210 262.635 654.490 262.750 ;
        RECT 655.660 241.130 655.800 262.750 ;
        RECT 655.200 240.990 655.800 241.130 ;
        RECT 655.200 194.325 655.340 240.990 ;
        RECT 655.130 193.955 655.410 194.325 ;
        RECT 655.590 193.275 655.870 193.645 ;
        RECT 655.660 193.110 655.800 193.275 ;
        RECT 655.600 192.790 655.860 193.110 ;
        RECT 655.600 145.190 655.860 145.510 ;
        RECT 655.660 144.830 655.800 145.190 ;
        RECT 655.600 144.510 655.860 144.830 ;
        RECT 656.520 144.510 656.780 144.830 ;
        RECT 656.580 97.085 656.720 144.510 ;
        RECT 655.590 96.715 655.870 97.085 ;
        RECT 656.510 96.715 656.790 97.085 ;
        RECT 655.660 96.550 655.800 96.715 ;
        RECT 655.600 96.230 655.860 96.550 ;
        RECT 656.980 57.130 657.240 57.450 ;
        RECT 657.040 2.400 657.180 57.130 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 286.210 262.680 286.490 262.960 ;
        RECT 654.210 262.680 654.490 262.960 ;
        RECT 655.130 194.000 655.410 194.280 ;
        RECT 655.590 193.320 655.870 193.600 ;
        RECT 655.590 96.760 655.870 97.040 ;
        RECT 656.510 96.760 656.790 97.040 ;
      LAYER met3 ;
        RECT 286.185 262.970 286.515 262.985 ;
        RECT 654.185 262.970 654.515 262.985 ;
        RECT 286.185 262.670 654.515 262.970 ;
        RECT 286.185 262.655 286.515 262.670 ;
        RECT 654.185 262.655 654.515 262.670 ;
        RECT 655.105 194.290 655.435 194.305 ;
        RECT 655.105 193.990 656.570 194.290 ;
        RECT 655.105 193.975 655.435 193.990 ;
        RECT 655.565 193.610 655.895 193.625 ;
        RECT 656.270 193.610 656.570 193.990 ;
        RECT 655.565 193.310 656.570 193.610 ;
        RECT 655.565 193.295 655.895 193.310 ;
        RECT 655.565 97.050 655.895 97.065 ;
        RECT 656.485 97.050 656.815 97.065 ;
        RECT 655.565 96.750 656.815 97.050 ;
        RECT 655.565 96.735 655.895 96.750 ;
        RECT 656.485 96.735 656.815 96.750 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2870.520 2615.490 2870.580 ;
        RECT 2686.470 2870.520 2686.790 2870.580 ;
        RECT 2615.170 2870.380 2686.790 2870.520 ;
        RECT 2615.170 2870.320 2615.490 2870.380 ;
        RECT 2686.470 2870.320 2686.790 2870.380 ;
        RECT 1000.110 225.320 1000.430 225.380 ;
        RECT 2686.470 225.320 2686.790 225.380 ;
        RECT 1000.110 225.180 2686.790 225.320 ;
        RECT 1000.110 225.120 1000.430 225.180 ;
        RECT 2686.470 225.120 2686.790 225.180 ;
        RECT 995.970 15.880 996.290 15.940 ;
        RECT 1000.110 15.880 1000.430 15.940 ;
        RECT 995.970 15.740 1000.430 15.880 ;
        RECT 995.970 15.680 996.290 15.740 ;
        RECT 1000.110 15.680 1000.430 15.740 ;
      LAYER via ;
        RECT 2615.200 2870.320 2615.460 2870.580 ;
        RECT 2686.500 2870.320 2686.760 2870.580 ;
        RECT 1000.140 225.120 1000.400 225.380 ;
        RECT 2686.500 225.120 2686.760 225.380 ;
        RECT 996.000 15.680 996.260 15.940 ;
        RECT 1000.140 15.680 1000.400 15.940 ;
      LAYER met2 ;
        RECT 2615.190 2875.195 2615.470 2875.565 ;
        RECT 2615.260 2870.610 2615.400 2875.195 ;
        RECT 2615.200 2870.290 2615.460 2870.610 ;
        RECT 2686.500 2870.290 2686.760 2870.610 ;
        RECT 2686.560 225.410 2686.700 2870.290 ;
        RECT 1000.140 225.090 1000.400 225.410 ;
        RECT 2686.500 225.090 2686.760 225.410 ;
        RECT 1000.200 15.970 1000.340 225.090 ;
        RECT 996.000 15.650 996.260 15.970 ;
        RECT 1000.140 15.650 1000.400 15.970 ;
        RECT 996.060 2.400 996.200 15.650 ;
        RECT 995.850 -4.800 996.410 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2875.240 2615.470 2875.520 ;
      LAYER met3 ;
        RECT 2606.000 2875.530 2610.000 2875.920 ;
        RECT 2615.165 2875.530 2615.495 2875.545 ;
        RECT 2606.000 2875.320 2615.495 2875.530 ;
        RECT 2609.580 2875.230 2615.495 2875.320 ;
        RECT 2615.165 2875.215 2615.495 2875.230 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1013.525 23.885 1013.695 34.595 ;
      LAYER mcon ;
        RECT 1013.525 34.425 1013.695 34.595 ;
      LAYER met1 ;
        RECT 289.410 3267.640 289.730 3267.700 ;
        RECT 791.270 3267.640 791.590 3267.700 ;
        RECT 289.410 3267.500 791.590 3267.640 ;
        RECT 289.410 3267.440 289.730 3267.500 ;
        RECT 791.270 3267.440 791.590 3267.500 ;
        RECT 289.410 385.800 289.730 385.860 ;
        RECT 303.670 385.800 303.990 385.860 ;
        RECT 289.410 385.660 303.990 385.800 ;
        RECT 289.410 385.600 289.730 385.660 ;
        RECT 303.670 385.600 303.990 385.660 ;
        RECT 278.830 283.800 279.150 283.860 ;
        RECT 303.670 283.800 303.990 283.860 ;
        RECT 278.830 283.660 303.990 283.800 ;
        RECT 278.830 283.600 279.150 283.660 ;
        RECT 303.670 283.600 303.990 283.660 ;
        RECT 278.830 58.040 279.150 58.100 ;
        RECT 1013.450 58.040 1013.770 58.100 ;
        RECT 278.830 57.900 1013.770 58.040 ;
        RECT 278.830 57.840 279.150 57.900 ;
        RECT 1013.450 57.840 1013.770 57.900 ;
        RECT 1013.450 34.580 1013.770 34.640 ;
        RECT 1013.255 34.440 1013.770 34.580 ;
        RECT 1013.450 34.380 1013.770 34.440 ;
        RECT 1013.450 24.040 1013.770 24.100 ;
        RECT 1013.255 23.900 1013.770 24.040 ;
        RECT 1013.450 23.840 1013.770 23.900 ;
      LAYER via ;
        RECT 289.440 3267.440 289.700 3267.700 ;
        RECT 791.300 3267.440 791.560 3267.700 ;
        RECT 289.440 385.600 289.700 385.860 ;
        RECT 303.700 385.600 303.960 385.860 ;
        RECT 278.860 283.600 279.120 283.860 ;
        RECT 303.700 283.600 303.960 283.860 ;
        RECT 278.860 57.840 279.120 58.100 ;
        RECT 1013.480 57.840 1013.740 58.100 ;
        RECT 1013.480 34.380 1013.740 34.640 ;
        RECT 1013.480 23.840 1013.740 24.100 ;
      LAYER met2 ;
        RECT 289.440 3267.410 289.700 3267.730 ;
        RECT 791.300 3267.410 791.560 3267.730 ;
        RECT 289.500 385.890 289.640 3267.410 ;
        RECT 791.360 3260.000 791.500 3267.410 ;
        RECT 791.250 3256.000 791.530 3260.000 ;
        RECT 289.440 385.570 289.700 385.890 ;
        RECT 303.700 385.570 303.960 385.890 ;
        RECT 303.760 283.890 303.900 385.570 ;
        RECT 278.860 283.570 279.120 283.890 ;
        RECT 303.700 283.570 303.960 283.890 ;
        RECT 278.920 58.130 279.060 283.570 ;
        RECT 278.860 57.810 279.120 58.130 ;
        RECT 1013.480 57.810 1013.740 58.130 ;
        RECT 1013.540 34.670 1013.680 57.810 ;
        RECT 1013.480 34.350 1013.740 34.670 ;
        RECT 1013.480 23.810 1013.740 24.130 ;
        RECT 1013.540 2.400 1013.680 23.810 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.390 259.660 295.710 259.720 ;
        RECT 1028.170 259.660 1028.490 259.720 ;
        RECT 295.390 259.520 1028.490 259.660 ;
        RECT 295.390 259.460 295.710 259.520 ;
        RECT 1028.170 259.460 1028.490 259.520 ;
        RECT 1028.170 2.960 1028.490 3.020 ;
        RECT 1031.390 2.960 1031.710 3.020 ;
        RECT 1028.170 2.820 1031.710 2.960 ;
        RECT 1028.170 2.760 1028.490 2.820 ;
        RECT 1031.390 2.760 1031.710 2.820 ;
      LAYER via ;
        RECT 295.420 259.460 295.680 259.720 ;
        RECT 1028.200 259.460 1028.460 259.720 ;
        RECT 1028.200 2.760 1028.460 3.020 ;
        RECT 1031.420 2.760 1031.680 3.020 ;
      LAYER met2 ;
        RECT 295.410 1996.635 295.690 1997.005 ;
        RECT 295.480 259.750 295.620 1996.635 ;
        RECT 295.420 259.430 295.680 259.750 ;
        RECT 1028.200 259.430 1028.460 259.750 ;
        RECT 1028.260 3.050 1028.400 259.430 ;
        RECT 1028.200 2.730 1028.460 3.050 ;
        RECT 1031.420 2.730 1031.680 3.050 ;
        RECT 1031.480 2.400 1031.620 2.730 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
      LAYER via2 ;
        RECT 295.410 1996.680 295.690 1996.960 ;
      LAYER met3 ;
        RECT 295.385 1996.970 295.715 1996.985 ;
        RECT 310.000 1996.970 314.000 1997.360 ;
        RECT 295.385 1996.760 314.000 1996.970 ;
        RECT 295.385 1996.670 310.500 1996.760 ;
        RECT 295.385 1996.655 295.715 1996.670 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2622.145 18.445 2622.315 19.635 ;
        RECT 2635.025 18.785 2635.195 19.635 ;
      LAYER mcon ;
        RECT 2622.145 19.465 2622.315 19.635 ;
        RECT 2635.025 19.465 2635.195 19.635 ;
      LAYER met1 ;
        RECT 2615.170 1393.900 2615.490 1393.960 ;
        RECT 2687.850 1393.900 2688.170 1393.960 ;
        RECT 2615.170 1393.760 2688.170 1393.900 ;
        RECT 2615.170 1393.700 2615.490 1393.760 ;
        RECT 2687.850 1393.700 2688.170 1393.760 ;
        RECT 2622.085 19.620 2622.375 19.665 ;
        RECT 2634.965 19.620 2635.255 19.665 ;
        RECT 2622.085 19.480 2635.255 19.620 ;
        RECT 2622.085 19.435 2622.375 19.480 ;
        RECT 2634.965 19.435 2635.255 19.480 ;
        RECT 2634.965 18.940 2635.255 18.985 ;
        RECT 2687.850 18.940 2688.170 19.000 ;
        RECT 2634.965 18.800 2688.170 18.940 ;
        RECT 2634.965 18.755 2635.255 18.800 ;
        RECT 2687.850 18.740 2688.170 18.800 ;
        RECT 1049.330 18.600 1049.650 18.660 ;
        RECT 2622.085 18.600 2622.375 18.645 ;
        RECT 1049.330 18.460 2622.375 18.600 ;
        RECT 1049.330 18.400 1049.650 18.460 ;
        RECT 2622.085 18.415 2622.375 18.460 ;
      LAYER via ;
        RECT 2615.200 1393.700 2615.460 1393.960 ;
        RECT 2687.880 1393.700 2688.140 1393.960 ;
        RECT 2687.880 18.740 2688.140 19.000 ;
        RECT 1049.360 18.400 1049.620 18.660 ;
      LAYER met2 ;
        RECT 2615.190 1395.515 2615.470 1395.885 ;
        RECT 2615.260 1393.990 2615.400 1395.515 ;
        RECT 2615.200 1393.670 2615.460 1393.990 ;
        RECT 2687.880 1393.670 2688.140 1393.990 ;
        RECT 2687.940 19.030 2688.080 1393.670 ;
        RECT 2687.880 18.710 2688.140 19.030 ;
        RECT 1049.360 18.370 1049.620 18.690 ;
        RECT 1049.420 2.400 1049.560 18.370 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1395.560 2615.470 1395.840 ;
      LAYER met3 ;
        RECT 2606.000 1395.850 2610.000 1396.240 ;
        RECT 2615.165 1395.850 2615.495 1395.865 ;
        RECT 2606.000 1395.640 2615.495 1395.850 ;
        RECT 2609.580 1395.550 2615.495 1395.640 ;
        RECT 2615.165 1395.535 2615.495 1395.550 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1062.745 48.365 1062.915 96.475 ;
      LAYER mcon ;
        RECT 1062.745 96.305 1062.915 96.475 ;
      LAYER met1 ;
        RECT 294.470 225.660 294.790 225.720 ;
        RECT 1062.670 225.660 1062.990 225.720 ;
        RECT 294.470 225.520 1062.990 225.660 ;
        RECT 294.470 225.460 294.790 225.520 ;
        RECT 1062.670 225.460 1062.990 225.520 ;
        RECT 1062.670 96.460 1062.990 96.520 ;
        RECT 1062.670 96.320 1063.185 96.460 ;
        RECT 1062.670 96.260 1062.990 96.320 ;
        RECT 1062.685 48.520 1062.975 48.565 ;
        RECT 1067.270 48.520 1067.590 48.580 ;
        RECT 1062.685 48.380 1067.590 48.520 ;
        RECT 1062.685 48.335 1062.975 48.380 ;
        RECT 1067.270 48.320 1067.590 48.380 ;
      LAYER via ;
        RECT 294.500 225.460 294.760 225.720 ;
        RECT 1062.700 225.460 1062.960 225.720 ;
        RECT 1062.700 96.260 1062.960 96.520 ;
        RECT 1067.300 48.320 1067.560 48.580 ;
      LAYER met2 ;
        RECT 294.490 1489.355 294.770 1489.725 ;
        RECT 294.560 225.750 294.700 1489.355 ;
        RECT 294.500 225.430 294.760 225.750 ;
        RECT 1062.700 225.430 1062.960 225.750 ;
        RECT 1062.760 96.550 1062.900 225.430 ;
        RECT 1062.700 96.230 1062.960 96.550 ;
        RECT 1067.300 48.290 1067.560 48.610 ;
        RECT 1067.360 2.400 1067.500 48.290 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
      LAYER via2 ;
        RECT 294.490 1489.400 294.770 1489.680 ;
      LAYER met3 ;
        RECT 294.465 1489.690 294.795 1489.705 ;
        RECT 310.000 1489.690 314.000 1490.080 ;
        RECT 294.465 1489.480 314.000 1489.690 ;
        RECT 294.465 1489.390 310.500 1489.480 ;
        RECT 294.465 1489.375 294.795 1489.390 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1085.210 14.860 1085.530 14.920 ;
        RECT 1089.810 14.860 1090.130 14.920 ;
        RECT 1085.210 14.720 1090.130 14.860 ;
        RECT 1085.210 14.660 1085.530 14.720 ;
        RECT 1089.810 14.660 1090.130 14.720 ;
      LAYER via ;
        RECT 1085.240 14.660 1085.500 14.920 ;
        RECT 1089.840 14.660 1090.100 14.920 ;
      LAYER met2 ;
        RECT 1089.830 204.155 1090.110 204.525 ;
        RECT 1089.900 14.950 1090.040 204.155 ;
        RECT 1085.240 14.630 1085.500 14.950 ;
        RECT 1089.840 14.630 1090.100 14.950 ;
        RECT 1085.300 2.400 1085.440 14.630 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
      LAYER via2 ;
        RECT 1089.830 204.200 1090.110 204.480 ;
      LAYER met3 ;
        RECT 2606.000 2980.250 2610.000 2980.640 ;
        RECT 2623.190 2980.250 2623.570 2980.260 ;
        RECT 2606.000 2980.040 2623.570 2980.250 ;
        RECT 2609.580 2979.950 2623.570 2980.040 ;
        RECT 2623.190 2979.940 2623.570 2979.950 ;
        RECT 1089.805 204.490 1090.135 204.505 ;
        RECT 2623.190 204.490 2623.570 204.500 ;
        RECT 1089.805 204.190 2623.570 204.490 ;
        RECT 1089.805 204.175 1090.135 204.190 ;
        RECT 2623.190 204.180 2623.570 204.190 ;
      LAYER via3 ;
        RECT 2623.220 2979.940 2623.540 2980.260 ;
        RECT 2623.220 204.180 2623.540 204.500 ;
      LAYER met4 ;
        RECT 2623.215 2979.935 2623.545 2980.265 ;
        RECT 2623.230 204.505 2623.530 2979.935 ;
        RECT 2623.215 204.175 2623.545 204.505 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.150 226.000 1103.470 226.060 ;
        RECT 2622.990 226.000 2623.310 226.060 ;
        RECT 1103.150 225.860 2623.310 226.000 ;
        RECT 1103.150 225.800 1103.470 225.860 ;
        RECT 2622.990 225.800 2623.310 225.860 ;
      LAYER via ;
        RECT 1103.180 225.800 1103.440 226.060 ;
        RECT 2623.020 225.800 2623.280 226.060 ;
      LAYER met2 ;
        RECT 2623.010 2135.355 2623.290 2135.725 ;
        RECT 2623.080 226.090 2623.220 2135.355 ;
        RECT 1103.180 225.770 1103.440 226.090 ;
        RECT 2623.020 225.770 2623.280 226.090 ;
        RECT 1103.240 3.130 1103.380 225.770 ;
        RECT 1102.780 2.990 1103.380 3.130 ;
        RECT 1102.780 2.400 1102.920 2.990 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 2623.010 2135.400 2623.290 2135.680 ;
      LAYER met3 ;
        RECT 2606.000 2135.690 2610.000 2136.080 ;
        RECT 2622.985 2135.690 2623.315 2135.705 ;
        RECT 2606.000 2135.480 2623.315 2135.690 ;
        RECT 2609.580 2135.390 2623.315 2135.480 ;
        RECT 2622.985 2135.375 2623.315 2135.390 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 312.870 2015.080 313.190 2015.140 ;
        RECT 314.710 2015.080 315.030 2015.140 ;
        RECT 312.870 2014.940 315.030 2015.080 ;
        RECT 312.870 2014.880 313.190 2014.940 ;
        RECT 314.710 2014.880 315.030 2014.940 ;
        RECT 314.710 337.320 315.030 337.580 ;
        RECT 314.800 337.180 314.940 337.320 ;
        RECT 314.340 337.040 314.940 337.180 ;
        RECT 314.340 336.900 314.480 337.040 ;
        RECT 314.250 336.640 314.570 336.900 ;
        RECT 314.710 259.320 315.030 259.380 ;
        RECT 1117.870 259.320 1118.190 259.380 ;
        RECT 314.710 259.180 1118.190 259.320 ;
        RECT 314.710 259.120 315.030 259.180 ;
        RECT 1117.870 259.120 1118.190 259.180 ;
        RECT 1117.870 2.960 1118.190 3.020 ;
        RECT 1120.630 2.960 1120.950 3.020 ;
        RECT 1117.870 2.820 1120.950 2.960 ;
        RECT 1117.870 2.760 1118.190 2.820 ;
        RECT 1120.630 2.760 1120.950 2.820 ;
      LAYER via ;
        RECT 312.900 2014.880 313.160 2015.140 ;
        RECT 314.740 2014.880 315.000 2015.140 ;
        RECT 314.740 337.320 315.000 337.580 ;
        RECT 314.280 336.640 314.540 336.900 ;
        RECT 314.740 259.120 315.000 259.380 ;
        RECT 1117.900 259.120 1118.160 259.380 ;
        RECT 1117.900 2.760 1118.160 3.020 ;
        RECT 1120.660 2.760 1120.920 3.020 ;
      LAYER met2 ;
        RECT 312.890 2015.675 313.170 2016.045 ;
        RECT 312.960 2015.170 313.100 2015.675 ;
        RECT 312.900 2014.850 313.160 2015.170 ;
        RECT 314.740 2014.850 315.000 2015.170 ;
        RECT 314.800 337.610 314.940 2014.850 ;
        RECT 314.740 337.290 315.000 337.610 ;
        RECT 314.280 336.610 314.540 336.930 ;
        RECT 314.340 313.890 314.480 336.610 ;
        RECT 314.340 313.750 314.940 313.890 ;
        RECT 314.800 259.410 314.940 313.750 ;
        RECT 314.740 259.090 315.000 259.410 ;
        RECT 1117.900 259.090 1118.160 259.410 ;
        RECT 1117.960 3.050 1118.100 259.090 ;
        RECT 1117.900 2.730 1118.160 3.050 ;
        RECT 1120.660 2.730 1120.920 3.050 ;
        RECT 1120.720 2.400 1120.860 2.730 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
      LAYER via2 ;
        RECT 312.890 2015.720 313.170 2016.000 ;
      LAYER met3 ;
        RECT 310.000 2018.520 314.000 2019.120 ;
        RECT 313.110 2016.025 313.410 2018.520 ;
        RECT 312.865 2015.710 313.410 2016.025 ;
        RECT 312.865 2015.695 313.195 2015.710 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1600.960 2615.490 1601.020 ;
        RECT 2695.210 1600.960 2695.530 1601.020 ;
        RECT 2615.170 1600.820 2695.530 1600.960 ;
        RECT 2615.170 1600.760 2615.490 1600.820 ;
        RECT 2695.210 1600.760 2695.530 1600.820 ;
        RECT 1145.010 232.120 1145.330 232.180 ;
        RECT 2695.210 232.120 2695.530 232.180 ;
        RECT 1145.010 231.980 2695.530 232.120 ;
        RECT 1145.010 231.920 1145.330 231.980 ;
        RECT 2695.210 231.920 2695.530 231.980 ;
        RECT 1138.570 16.900 1138.890 16.960 ;
        RECT 1145.010 16.900 1145.330 16.960 ;
        RECT 1138.570 16.760 1145.330 16.900 ;
        RECT 1138.570 16.700 1138.890 16.760 ;
        RECT 1145.010 16.700 1145.330 16.760 ;
      LAYER via ;
        RECT 2615.200 1600.760 2615.460 1601.020 ;
        RECT 2695.240 1600.760 2695.500 1601.020 ;
        RECT 1145.040 231.920 1145.300 232.180 ;
        RECT 2695.240 231.920 2695.500 232.180 ;
        RECT 1138.600 16.700 1138.860 16.960 ;
        RECT 1145.040 16.700 1145.300 16.960 ;
      LAYER met2 ;
        RECT 2615.190 1606.315 2615.470 1606.685 ;
        RECT 2615.260 1601.050 2615.400 1606.315 ;
        RECT 2615.200 1600.730 2615.460 1601.050 ;
        RECT 2695.240 1600.730 2695.500 1601.050 ;
        RECT 2695.300 232.210 2695.440 1600.730 ;
        RECT 1145.040 231.890 1145.300 232.210 ;
        RECT 2695.240 231.890 2695.500 232.210 ;
        RECT 1145.100 16.990 1145.240 231.890 ;
        RECT 1138.600 16.670 1138.860 16.990 ;
        RECT 1145.040 16.670 1145.300 16.990 ;
        RECT 1138.660 2.400 1138.800 16.670 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1606.360 2615.470 1606.640 ;
      LAYER met3 ;
        RECT 2606.000 1606.650 2610.000 1607.040 ;
        RECT 2615.165 1606.650 2615.495 1606.665 ;
        RECT 2606.000 1606.440 2615.495 1606.650 ;
        RECT 2609.580 1606.350 2615.495 1606.440 ;
        RECT 2615.165 1606.335 2615.495 1606.350 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 744.350 176.020 744.670 176.080 ;
        RECT 1152.370 176.020 1152.690 176.080 ;
        RECT 744.350 175.880 1152.690 176.020 ;
        RECT 744.350 175.820 744.670 175.880 ;
        RECT 1152.370 175.820 1152.690 175.880 ;
        RECT 1152.370 62.120 1152.690 62.180 ;
        RECT 1156.510 62.120 1156.830 62.180 ;
        RECT 1152.370 61.980 1156.830 62.120 ;
        RECT 1152.370 61.920 1152.690 61.980 ;
        RECT 1156.510 61.920 1156.830 61.980 ;
      LAYER via ;
        RECT 744.380 175.820 744.640 176.080 ;
        RECT 1152.400 175.820 1152.660 176.080 ;
        RECT 1152.400 61.920 1152.660 62.180 ;
        RECT 1156.540 61.920 1156.800 62.180 ;
      LAYER met2 ;
        RECT 741.570 260.170 741.850 264.000 ;
        RECT 741.570 260.030 744.580 260.170 ;
        RECT 741.570 260.000 741.850 260.030 ;
        RECT 744.440 176.110 744.580 260.030 ;
        RECT 744.380 175.790 744.640 176.110 ;
        RECT 1152.400 175.790 1152.660 176.110 ;
        RECT 1152.460 62.210 1152.600 175.790 ;
        RECT 1152.400 61.890 1152.660 62.210 ;
        RECT 1156.540 61.890 1156.800 62.210 ;
        RECT 1156.600 2.400 1156.740 61.890 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.830 258.555 676.110 258.925 ;
        RECT 675.900 3.130 676.040 258.555 ;
        RECT 674.520 2.990 676.040 3.130 ;
        RECT 674.520 2.400 674.660 2.990 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 675.830 258.600 676.110 258.880 ;
      LAYER met3 ;
        RECT 2606.000 1586.250 2610.000 1586.640 ;
        RECT 2618.590 1586.250 2618.970 1586.260 ;
        RECT 2606.000 1586.040 2618.970 1586.250 ;
        RECT 2609.580 1585.950 2618.970 1586.040 ;
        RECT 2618.590 1585.940 2618.970 1585.950 ;
        RECT 675.805 258.890 676.135 258.905 ;
        RECT 2618.590 258.890 2618.970 258.900 ;
        RECT 675.805 258.590 2618.970 258.890 ;
        RECT 675.805 258.575 676.135 258.590 ;
        RECT 2618.590 258.580 2618.970 258.590 ;
      LAYER via3 ;
        RECT 2618.620 1585.940 2618.940 1586.260 ;
        RECT 2618.620 258.580 2618.940 258.900 ;
      LAYER met4 ;
        RECT 2618.615 1585.935 2618.945 1586.265 ;
        RECT 2618.630 258.905 2618.930 1585.935 ;
        RECT 2618.615 258.575 2618.945 258.905 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1173.145 144.925 1173.315 193.035 ;
        RECT 1173.145 48.365 1173.315 137.955 ;
      LAYER mcon ;
        RECT 1173.145 192.865 1173.315 193.035 ;
        RECT 1173.145 137.785 1173.315 137.955 ;
      LAYER met1 ;
        RECT 295.850 217.840 296.170 217.900 ;
        RECT 1173.530 217.840 1173.850 217.900 ;
        RECT 295.850 217.700 1173.850 217.840 ;
        RECT 295.850 217.640 296.170 217.700 ;
        RECT 1173.530 217.640 1173.850 217.700 ;
        RECT 1173.070 193.020 1173.390 193.080 ;
        RECT 1172.875 192.880 1173.390 193.020 ;
        RECT 1173.070 192.820 1173.390 192.880 ;
        RECT 1173.070 145.080 1173.390 145.140 ;
        RECT 1172.875 144.940 1173.390 145.080 ;
        RECT 1173.070 144.880 1173.390 144.940 ;
        RECT 1173.070 137.940 1173.390 138.000 ;
        RECT 1172.875 137.800 1173.390 137.940 ;
        RECT 1173.070 137.740 1173.390 137.800 ;
        RECT 1173.085 48.520 1173.375 48.565 ;
        RECT 1173.990 48.520 1174.310 48.580 ;
        RECT 1173.085 48.380 1174.310 48.520 ;
        RECT 1173.085 48.335 1173.375 48.380 ;
        RECT 1173.990 48.320 1174.310 48.380 ;
      LAYER via ;
        RECT 295.880 217.640 296.140 217.900 ;
        RECT 1173.560 217.640 1173.820 217.900 ;
        RECT 1173.100 192.820 1173.360 193.080 ;
        RECT 1173.100 144.880 1173.360 145.140 ;
        RECT 1173.100 137.740 1173.360 138.000 ;
        RECT 1174.020 48.320 1174.280 48.580 ;
      LAYER met2 ;
        RECT 295.870 2038.795 296.150 2039.165 ;
        RECT 295.940 217.930 296.080 2038.795 ;
        RECT 295.880 217.610 296.140 217.930 ;
        RECT 1173.560 217.610 1173.820 217.930 ;
        RECT 1173.620 193.530 1173.760 217.610 ;
        RECT 1173.160 193.390 1173.760 193.530 ;
        RECT 1173.160 193.110 1173.300 193.390 ;
        RECT 1173.100 192.790 1173.360 193.110 ;
        RECT 1173.100 144.850 1173.360 145.170 ;
        RECT 1173.160 138.030 1173.300 144.850 ;
        RECT 1173.100 137.710 1173.360 138.030 ;
        RECT 1174.020 48.290 1174.280 48.610 ;
        RECT 1174.080 2.400 1174.220 48.290 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
      LAYER via2 ;
        RECT 295.870 2038.840 296.150 2039.120 ;
      LAYER met3 ;
        RECT 295.845 2039.130 296.175 2039.145 ;
        RECT 310.000 2039.130 314.000 2039.520 ;
        RECT 295.845 2038.920 314.000 2039.130 ;
        RECT 295.845 2038.830 310.500 2038.920 ;
        RECT 295.845 2038.815 296.175 2038.830 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 310.110 258.640 310.430 258.700 ;
        RECT 1186.870 258.640 1187.190 258.700 ;
        RECT 310.110 258.500 1187.190 258.640 ;
        RECT 310.110 258.440 310.430 258.500 ;
        RECT 1186.870 258.440 1187.190 258.500 ;
        RECT 1186.870 62.120 1187.190 62.180 ;
        RECT 1191.930 62.120 1192.250 62.180 ;
        RECT 1186.870 61.980 1192.250 62.120 ;
        RECT 1186.870 61.920 1187.190 61.980 ;
        RECT 1191.930 61.920 1192.250 61.980 ;
      LAYER via ;
        RECT 310.140 258.440 310.400 258.700 ;
        RECT 1186.900 258.440 1187.160 258.700 ;
        RECT 1186.900 61.920 1187.160 62.180 ;
        RECT 1191.960 61.920 1192.220 62.180 ;
      LAYER met2 ;
        RECT 310.130 283.035 310.410 283.405 ;
        RECT 310.200 258.730 310.340 283.035 ;
        RECT 310.140 258.410 310.400 258.730 ;
        RECT 1186.900 258.410 1187.160 258.730 ;
        RECT 1186.960 62.210 1187.100 258.410 ;
        RECT 1186.900 61.890 1187.160 62.210 ;
        RECT 1191.960 61.890 1192.220 62.210 ;
        RECT 1192.020 2.400 1192.160 61.890 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 310.130 283.080 310.410 283.360 ;
      LAYER met3 ;
        RECT 310.000 284.520 314.000 285.120 ;
        RECT 310.350 283.385 310.650 284.520 ;
        RECT 310.105 283.070 310.650 283.385 ;
        RECT 310.105 283.055 310.435 283.070 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1214.010 232.460 1214.330 232.520 ;
        RECT 2672.210 232.460 2672.530 232.520 ;
        RECT 1214.010 232.320 2672.530 232.460 ;
        RECT 1214.010 232.260 1214.330 232.320 ;
        RECT 2672.210 232.260 2672.530 232.320 ;
        RECT 1209.870 20.640 1210.190 20.700 ;
        RECT 1214.010 20.640 1214.330 20.700 ;
        RECT 1209.870 20.500 1214.330 20.640 ;
        RECT 1209.870 20.440 1210.190 20.500 ;
        RECT 1214.010 20.440 1214.330 20.500 ;
      LAYER via ;
        RECT 1214.040 232.260 1214.300 232.520 ;
        RECT 2672.240 232.260 2672.500 232.520 ;
        RECT 1209.900 20.440 1210.160 20.700 ;
        RECT 1214.040 20.440 1214.300 20.700 ;
      LAYER met2 ;
        RECT 1950.950 3260.755 1951.230 3261.125 ;
        RECT 1949.530 3259.650 1949.810 3260.000 ;
        RECT 1951.020 3259.650 1951.160 3260.755 ;
        RECT 1949.530 3259.510 1951.160 3259.650 ;
        RECT 1949.530 3256.000 1949.810 3259.510 ;
        RECT 2672.230 3251.235 2672.510 3251.605 ;
        RECT 2672.300 232.550 2672.440 3251.235 ;
        RECT 1214.040 232.230 1214.300 232.550 ;
        RECT 2672.240 232.230 2672.500 232.550 ;
        RECT 1214.100 20.730 1214.240 232.230 ;
        RECT 1209.900 20.410 1210.160 20.730 ;
        RECT 1214.040 20.410 1214.300 20.730 ;
        RECT 1209.960 2.400 1210.100 20.410 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
      LAYER via2 ;
        RECT 1950.950 3260.800 1951.230 3261.080 ;
        RECT 2672.230 3251.280 2672.510 3251.560 ;
      LAYER met3 ;
        RECT 1950.925 3261.090 1951.255 3261.105 ;
        RECT 1951.590 3261.090 1951.970 3261.100 ;
        RECT 1950.925 3260.790 1951.970 3261.090 ;
        RECT 1950.925 3260.775 1951.255 3260.790 ;
        RECT 1951.590 3260.780 1951.970 3260.790 ;
        RECT 1951.590 3251.570 1951.970 3251.580 ;
        RECT 2672.205 3251.570 2672.535 3251.585 ;
        RECT 1951.590 3251.270 2672.535 3251.570 ;
        RECT 1951.590 3251.260 1951.970 3251.270 ;
        RECT 2672.205 3251.255 2672.535 3251.270 ;
      LAYER via3 ;
        RECT 1951.620 3260.780 1951.940 3261.100 ;
        RECT 1951.620 3251.260 1951.940 3251.580 ;
      LAYER met4 ;
        RECT 1951.615 3260.775 1951.945 3261.105 ;
        RECT 1951.630 3251.585 1951.930 3260.775 ;
        RECT 1951.615 3251.255 1951.945 3251.585 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 155.280 1228.130 155.340 ;
        RECT 2620.230 155.280 2620.550 155.340 ;
        RECT 1227.810 155.140 2620.550 155.280 ;
        RECT 1227.810 155.080 1228.130 155.140 ;
        RECT 2620.230 155.080 2620.550 155.140 ;
      LAYER via ;
        RECT 1227.840 155.080 1228.100 155.340 ;
        RECT 2620.260 155.080 2620.520 155.340 ;
      LAYER met2 ;
        RECT 2620.250 571.355 2620.530 571.725 ;
        RECT 2620.320 155.370 2620.460 571.355 ;
        RECT 1227.840 155.050 1228.100 155.370 ;
        RECT 2620.260 155.050 2620.520 155.370 ;
        RECT 1227.900 2.400 1228.040 155.050 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
      LAYER via2 ;
        RECT 2620.250 571.400 2620.530 571.680 ;
      LAYER met3 ;
        RECT 2606.000 571.690 2610.000 572.080 ;
        RECT 2620.225 571.690 2620.555 571.705 ;
        RECT 2606.000 571.480 2620.555 571.690 ;
        RECT 2609.580 571.390 2620.555 571.480 ;
        RECT 2620.225 571.375 2620.555 571.390 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2620.690 1221.520 2621.010 1221.580 ;
        RECT 2652.430 1221.520 2652.750 1221.580 ;
        RECT 2620.690 1221.380 2652.750 1221.520 ;
        RECT 2620.690 1221.320 2621.010 1221.380 ;
        RECT 2652.430 1221.320 2652.750 1221.380 ;
        RECT 1248.510 226.340 1248.830 226.400 ;
        RECT 2652.430 226.340 2652.750 226.400 ;
        RECT 1248.510 226.200 2652.750 226.340 ;
        RECT 1248.510 226.140 1248.830 226.200 ;
        RECT 2652.430 226.140 2652.750 226.200 ;
        RECT 1245.750 20.640 1246.070 20.700 ;
        RECT 1248.510 20.640 1248.830 20.700 ;
        RECT 1245.750 20.500 1248.830 20.640 ;
        RECT 1245.750 20.440 1246.070 20.500 ;
        RECT 1248.510 20.440 1248.830 20.500 ;
      LAYER via ;
        RECT 2620.720 1221.320 2620.980 1221.580 ;
        RECT 2652.460 1221.320 2652.720 1221.580 ;
        RECT 1248.540 226.140 1248.800 226.400 ;
        RECT 2652.460 226.140 2652.720 226.400 ;
        RECT 1245.780 20.440 1246.040 20.700 ;
        RECT 1248.540 20.440 1248.800 20.700 ;
      LAYER met2 ;
        RECT 2620.710 1225.515 2620.990 1225.885 ;
        RECT 2620.780 1221.610 2620.920 1225.515 ;
        RECT 2620.720 1221.290 2620.980 1221.610 ;
        RECT 2652.460 1221.290 2652.720 1221.610 ;
        RECT 2652.520 226.430 2652.660 1221.290 ;
        RECT 1248.540 226.110 1248.800 226.430 ;
        RECT 2652.460 226.110 2652.720 226.430 ;
        RECT 1248.600 20.730 1248.740 226.110 ;
        RECT 1245.780 20.410 1246.040 20.730 ;
        RECT 1248.540 20.410 1248.800 20.730 ;
        RECT 1245.840 2.400 1245.980 20.410 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
      LAYER via2 ;
        RECT 2620.710 1225.560 2620.990 1225.840 ;
      LAYER met3 ;
        RECT 2606.000 1225.850 2610.000 1226.240 ;
        RECT 2620.685 1225.850 2621.015 1225.865 ;
        RECT 2606.000 1225.640 2621.015 1225.850 ;
        RECT 2609.580 1225.550 2621.015 1225.640 ;
        RECT 2620.685 1225.535 2621.015 1225.550 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 924.700 2615.490 924.760 ;
        RECT 2625.750 924.700 2626.070 924.760 ;
        RECT 2615.170 924.560 2626.070 924.700 ;
        RECT 2615.170 924.500 2615.490 924.560 ;
        RECT 2625.750 924.500 2626.070 924.560 ;
        RECT 1269.210 258.640 1269.530 258.700 ;
        RECT 2625.750 258.640 2626.070 258.700 ;
        RECT 1269.210 258.500 2626.070 258.640 ;
        RECT 1269.210 258.440 1269.530 258.500 ;
        RECT 2625.750 258.440 2626.070 258.500 ;
        RECT 1263.230 14.860 1263.550 14.920 ;
        RECT 1269.210 14.860 1269.530 14.920 ;
        RECT 1263.230 14.720 1269.530 14.860 ;
        RECT 1263.230 14.660 1263.550 14.720 ;
        RECT 1269.210 14.660 1269.530 14.720 ;
      LAYER via ;
        RECT 2615.200 924.500 2615.460 924.760 ;
        RECT 2625.780 924.500 2626.040 924.760 ;
        RECT 1269.240 258.440 1269.500 258.700 ;
        RECT 2625.780 258.440 2626.040 258.700 ;
        RECT 1263.260 14.660 1263.520 14.920 ;
        RECT 1269.240 14.660 1269.500 14.920 ;
      LAYER met2 ;
        RECT 2615.190 930.395 2615.470 930.765 ;
        RECT 2615.260 924.790 2615.400 930.395 ;
        RECT 2615.200 924.470 2615.460 924.790 ;
        RECT 2625.780 924.470 2626.040 924.790 ;
        RECT 2625.840 258.730 2625.980 924.470 ;
        RECT 1269.240 258.410 1269.500 258.730 ;
        RECT 2625.780 258.410 2626.040 258.730 ;
        RECT 1269.300 14.950 1269.440 258.410 ;
        RECT 1263.260 14.630 1263.520 14.950 ;
        RECT 1269.240 14.630 1269.500 14.950 ;
        RECT 1263.320 2.400 1263.460 14.630 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
      LAYER via2 ;
        RECT 2615.190 930.440 2615.470 930.720 ;
      LAYER met3 ;
        RECT 2606.000 930.730 2610.000 931.120 ;
        RECT 2615.165 930.730 2615.495 930.745 ;
        RECT 2606.000 930.520 2615.495 930.730 ;
        RECT 2609.580 930.430 2615.495 930.520 ;
        RECT 2615.165 930.415 2615.495 930.430 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1281.170 26.420 1281.490 26.480 ;
        RECT 1593.970 26.420 1594.290 26.480 ;
        RECT 1281.170 26.280 1594.290 26.420 ;
        RECT 1281.170 26.220 1281.490 26.280 ;
        RECT 1593.970 26.220 1594.290 26.280 ;
      LAYER via ;
        RECT 1281.200 26.220 1281.460 26.480 ;
        RECT 1594.000 26.220 1594.260 26.480 ;
      LAYER met2 ;
        RECT 1599.010 260.170 1599.290 264.000 ;
        RECT 1594.060 260.030 1599.290 260.170 ;
        RECT 1594.060 26.510 1594.200 260.030 ;
        RECT 1599.010 260.000 1599.290 260.030 ;
        RECT 1281.200 26.190 1281.460 26.510 ;
        RECT 1594.000 26.190 1594.260 26.510 ;
        RECT 1281.260 2.400 1281.400 26.190 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.110 15.880 1299.430 15.940 ;
        RECT 1303.710 15.880 1304.030 15.940 ;
        RECT 1299.110 15.740 1304.030 15.880 ;
        RECT 1299.110 15.680 1299.430 15.740 ;
        RECT 1303.710 15.680 1304.030 15.740 ;
      LAYER via ;
        RECT 1299.140 15.680 1299.400 15.940 ;
        RECT 1303.740 15.680 1304.000 15.940 ;
      LAYER met2 ;
        RECT 1303.730 79.035 1304.010 79.405 ;
        RECT 1303.800 15.970 1303.940 79.035 ;
        RECT 1299.140 15.650 1299.400 15.970 ;
        RECT 1303.740 15.650 1304.000 15.970 ;
        RECT 1299.200 2.400 1299.340 15.650 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
      LAYER via2 ;
        RECT 1303.730 79.080 1304.010 79.360 ;
      LAYER met3 ;
        RECT 2606.000 2472.970 2610.000 2473.360 ;
        RECT 2610.310 2472.970 2610.690 2472.980 ;
        RECT 2606.000 2472.760 2610.690 2472.970 ;
        RECT 2609.580 2472.670 2610.690 2472.760 ;
        RECT 2610.310 2472.660 2610.690 2472.670 ;
        RECT 1303.705 79.370 1304.035 79.385 ;
        RECT 2610.310 79.370 2610.690 79.380 ;
        RECT 1303.705 79.070 2610.690 79.370 ;
        RECT 1303.705 79.055 1304.035 79.070 ;
        RECT 2610.310 79.060 2610.690 79.070 ;
      LAYER via3 ;
        RECT 2610.340 2472.660 2610.660 2472.980 ;
        RECT 2610.340 79.060 2610.660 79.380 ;
      LAYER met4 ;
        RECT 2610.335 2472.655 2610.665 2472.985 ;
        RECT 2610.350 79.385 2610.650 2472.655 ;
        RECT 2610.335 79.055 2610.665 79.385 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 3257.100 240.970 3257.160 ;
        RECT 374.510 3257.100 374.830 3257.160 ;
        RECT 240.650 3256.960 374.830 3257.100 ;
        RECT 240.650 3256.900 240.970 3256.960 ;
        RECT 374.510 3256.900 374.830 3256.960 ;
        RECT 240.650 48.180 240.970 48.240 ;
        RECT 1317.050 48.180 1317.370 48.240 ;
        RECT 240.650 48.040 1317.370 48.180 ;
        RECT 240.650 47.980 240.970 48.040 ;
        RECT 1317.050 47.980 1317.370 48.040 ;
      LAYER via ;
        RECT 240.680 3256.900 240.940 3257.160 ;
        RECT 374.540 3256.900 374.800 3257.160 ;
        RECT 240.680 47.980 240.940 48.240 ;
        RECT 1317.080 47.980 1317.340 48.240 ;
      LAYER met2 ;
        RECT 240.680 3256.870 240.940 3257.190 ;
        RECT 374.540 3256.930 374.800 3257.190 ;
        RECT 376.330 3256.930 376.610 3260.000 ;
        RECT 374.540 3256.870 376.610 3256.930 ;
        RECT 240.740 48.270 240.880 3256.870 ;
        RECT 374.600 3256.790 376.610 3256.870 ;
        RECT 376.330 3256.000 376.610 3256.790 ;
        RECT 240.680 47.950 240.940 48.270 ;
        RECT 1317.080 47.950 1317.340 48.270 ;
        RECT 1317.140 2.400 1317.280 47.950 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1331.770 62.120 1332.090 62.180 ;
        RECT 1334.990 62.120 1335.310 62.180 ;
        RECT 1331.770 61.980 1335.310 62.120 ;
        RECT 1331.770 61.920 1332.090 61.980 ;
        RECT 1334.990 61.920 1335.310 61.980 ;
      LAYER via ;
        RECT 1331.800 61.920 1332.060 62.180 ;
        RECT 1335.020 61.920 1335.280 62.180 ;
      LAYER met2 ;
        RECT 317.490 259.915 317.770 260.285 ;
        RECT 1331.790 259.915 1332.070 260.285 ;
        RECT 317.560 258.245 317.700 259.915 ;
        RECT 317.490 257.875 317.770 258.245 ;
        RECT 1331.860 62.210 1332.000 259.915 ;
        RECT 1331.800 61.890 1332.060 62.210 ;
        RECT 1335.020 61.890 1335.280 62.210 ;
        RECT 1335.080 2.400 1335.220 61.890 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
      LAYER via2 ;
        RECT 317.490 259.960 317.770 260.240 ;
        RECT 1331.790 259.960 1332.070 260.240 ;
        RECT 317.490 257.920 317.770 258.200 ;
      LAYER met3 ;
        RECT 304.790 2905.450 305.170 2905.460 ;
        RECT 310.000 2905.450 314.000 2905.840 ;
        RECT 304.790 2905.240 314.000 2905.450 ;
        RECT 304.790 2905.150 310.500 2905.240 ;
        RECT 304.790 2905.140 305.170 2905.150 ;
        RECT 317.465 260.250 317.795 260.265 ;
        RECT 1331.765 260.250 1332.095 260.265 ;
        RECT 317.465 259.950 1332.095 260.250 ;
        RECT 317.465 259.935 317.795 259.950 ;
        RECT 1331.765 259.935 1332.095 259.950 ;
        RECT 304.790 258.210 305.170 258.220 ;
        RECT 317.465 258.210 317.795 258.225 ;
        RECT 304.790 257.910 317.795 258.210 ;
        RECT 304.790 257.900 305.170 257.910 ;
        RECT 317.465 257.895 317.795 257.910 ;
      LAYER via3 ;
        RECT 304.820 2905.140 305.140 2905.460 ;
        RECT 304.820 257.900 305.140 258.220 ;
      LAYER met4 ;
        RECT 304.815 2905.135 305.145 2905.465 ;
        RECT 304.830 258.225 305.130 2905.135 ;
        RECT 304.815 257.895 305.145 258.225 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 25.400 692.690 25.460 ;
        RECT 1324.870 25.400 1325.190 25.460 ;
        RECT 692.370 25.260 1325.190 25.400 ;
        RECT 692.370 25.200 692.690 25.260 ;
        RECT 1324.870 25.200 1325.190 25.260 ;
      LAYER via ;
        RECT 692.400 25.200 692.660 25.460 ;
        RECT 1324.900 25.200 1325.160 25.460 ;
      LAYER met2 ;
        RECT 1327.610 260.170 1327.890 264.000 ;
        RECT 1324.960 260.030 1327.890 260.170 ;
        RECT 1324.960 25.490 1325.100 260.030 ;
        RECT 1327.610 260.000 1327.890 260.030 ;
        RECT 692.400 25.170 692.660 25.490 ;
        RECT 1324.900 25.170 1325.160 25.490 ;
        RECT 692.460 2.400 692.600 25.170 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2035.110 3267.640 2035.430 3267.700 ;
        RECT 2685.550 3267.640 2685.870 3267.700 ;
        RECT 2035.110 3267.500 2685.870 3267.640 ;
        RECT 2035.110 3267.440 2035.430 3267.500 ;
        RECT 2685.550 3267.440 2685.870 3267.500 ;
        RECT 1358.910 233.480 1359.230 233.540 ;
        RECT 2685.550 233.480 2685.870 233.540 ;
        RECT 1358.910 233.340 2685.870 233.480 ;
        RECT 1358.910 233.280 1359.230 233.340 ;
        RECT 2685.550 233.280 2685.870 233.340 ;
        RECT 1352.470 20.640 1352.790 20.700 ;
        RECT 1358.910 20.640 1359.230 20.700 ;
        RECT 1352.470 20.500 1359.230 20.640 ;
        RECT 1352.470 20.440 1352.790 20.500 ;
        RECT 1358.910 20.440 1359.230 20.500 ;
      LAYER via ;
        RECT 2035.140 3267.440 2035.400 3267.700 ;
        RECT 2685.580 3267.440 2685.840 3267.700 ;
        RECT 1358.940 233.280 1359.200 233.540 ;
        RECT 2685.580 233.280 2685.840 233.540 ;
        RECT 1352.500 20.440 1352.760 20.700 ;
        RECT 1358.940 20.440 1359.200 20.700 ;
      LAYER met2 ;
        RECT 2035.140 3267.410 2035.400 3267.730 ;
        RECT 2685.580 3267.410 2685.840 3267.730 ;
        RECT 2035.200 3260.000 2035.340 3267.410 ;
        RECT 2035.090 3256.000 2035.370 3260.000 ;
        RECT 2685.640 233.570 2685.780 3267.410 ;
        RECT 1358.940 233.250 1359.200 233.570 ;
        RECT 2685.580 233.250 2685.840 233.570 ;
        RECT 1359.000 20.730 1359.140 233.250 ;
        RECT 1352.500 20.410 1352.760 20.730 ;
        RECT 1358.940 20.410 1359.200 20.730 ;
        RECT 1352.560 2.400 1352.700 20.410 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1876.870 3285.320 1877.190 3285.380 ;
        RECT 2704.870 3285.320 2705.190 3285.380 ;
        RECT 1876.870 3285.180 2705.190 3285.320 ;
        RECT 1876.870 3285.120 1877.190 3285.180 ;
        RECT 2704.870 3285.120 2705.190 3285.180 ;
        RECT 1372.710 233.140 1373.030 233.200 ;
        RECT 2704.870 233.140 2705.190 233.200 ;
        RECT 1372.710 233.000 2705.190 233.140 ;
        RECT 1372.710 232.940 1373.030 233.000 ;
        RECT 2704.870 232.940 2705.190 233.000 ;
        RECT 1370.410 20.640 1370.730 20.700 ;
        RECT 1372.710 20.640 1373.030 20.700 ;
        RECT 1370.410 20.500 1373.030 20.640 ;
        RECT 1370.410 20.440 1370.730 20.500 ;
        RECT 1372.710 20.440 1373.030 20.500 ;
      LAYER via ;
        RECT 1876.900 3285.120 1877.160 3285.380 ;
        RECT 2704.900 3285.120 2705.160 3285.380 ;
        RECT 1372.740 232.940 1373.000 233.200 ;
        RECT 2704.900 232.940 2705.160 233.200 ;
        RECT 1370.440 20.440 1370.700 20.700 ;
        RECT 1372.740 20.440 1373.000 20.700 ;
      LAYER met2 ;
        RECT 1876.900 3285.090 1877.160 3285.410 ;
        RECT 2704.900 3285.090 2705.160 3285.410 ;
        RECT 1876.960 3259.650 1877.100 3285.090 ;
        RECT 1877.770 3259.650 1878.050 3260.000 ;
        RECT 1876.960 3259.510 1878.050 3259.650 ;
        RECT 1877.770 3256.000 1878.050 3259.510 ;
        RECT 2704.960 233.230 2705.100 3285.090 ;
        RECT 1372.740 232.910 1373.000 233.230 ;
        RECT 2704.900 232.910 2705.160 233.230 ;
        RECT 1372.800 20.730 1372.940 232.910 ;
        RECT 1370.440 20.410 1370.700 20.730 ;
        RECT 1372.740 20.410 1373.000 20.730 ;
        RECT 1370.500 2.400 1370.640 20.410 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1388.350 15.200 1388.670 15.260 ;
        RECT 1393.410 15.200 1393.730 15.260 ;
        RECT 1388.350 15.060 1393.730 15.200 ;
        RECT 1388.350 15.000 1388.670 15.060 ;
        RECT 1393.410 15.000 1393.730 15.060 ;
      LAYER via ;
        RECT 1388.380 15.000 1388.640 15.260 ;
        RECT 1393.440 15.000 1393.700 15.260 ;
      LAYER met2 ;
        RECT 1393.430 232.035 1393.710 232.405 ;
        RECT 1393.500 15.290 1393.640 232.035 ;
        RECT 1388.380 14.970 1388.640 15.290 ;
        RECT 1393.440 14.970 1393.700 15.290 ;
        RECT 1388.440 2.400 1388.580 14.970 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
      LAYER via2 ;
        RECT 1393.430 232.080 1393.710 232.360 ;
      LAYER met3 ;
        RECT 2606.000 2156.090 2610.000 2156.480 ;
        RECT 2617.670 2156.090 2618.050 2156.100 ;
        RECT 2606.000 2155.880 2618.050 2156.090 ;
        RECT 2609.580 2155.790 2618.050 2155.880 ;
        RECT 2617.670 2155.780 2618.050 2155.790 ;
        RECT 1393.405 232.370 1393.735 232.385 ;
        RECT 2617.670 232.370 2618.050 232.380 ;
        RECT 1393.405 232.070 2618.050 232.370 ;
        RECT 1393.405 232.055 1393.735 232.070 ;
        RECT 2617.670 232.060 2618.050 232.070 ;
      LAYER via3 ;
        RECT 2617.700 2155.780 2618.020 2156.100 ;
        RECT 2617.700 232.060 2618.020 232.380 ;
      LAYER met4 ;
        RECT 2617.695 2155.775 2618.025 2156.105 ;
        RECT 2617.710 232.385 2618.010 2155.775 ;
        RECT 2617.695 232.055 2618.025 232.385 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 259.125 990.165 259.295 1014.135 ;
      LAYER mcon ;
        RECT 259.125 1013.965 259.295 1014.135 ;
      LAYER met1 ;
        RECT 259.050 3298.580 259.370 3298.640 ;
        RECT 959.170 3298.580 959.490 3298.640 ;
        RECT 259.050 3298.440 959.490 3298.580 ;
        RECT 259.050 3298.380 259.370 3298.440 ;
        RECT 959.170 3298.380 959.490 3298.440 ;
        RECT 259.050 1014.120 259.370 1014.180 ;
        RECT 259.050 1013.980 259.565 1014.120 ;
        RECT 259.050 1013.920 259.370 1013.980 ;
        RECT 259.050 990.320 259.370 990.380 ;
        RECT 258.855 990.180 259.370 990.320 ;
        RECT 259.050 990.120 259.370 990.180 ;
        RECT 237.890 503.780 238.210 503.840 ;
        RECT 259.050 503.780 259.370 503.840 ;
        RECT 237.890 503.640 259.370 503.780 ;
        RECT 237.890 503.580 238.210 503.640 ;
        RECT 259.050 503.580 259.370 503.640 ;
      LAYER via ;
        RECT 259.080 3298.380 259.340 3298.640 ;
        RECT 959.200 3298.380 959.460 3298.640 ;
        RECT 259.080 1013.920 259.340 1014.180 ;
        RECT 259.080 990.120 259.340 990.380 ;
        RECT 237.920 503.580 238.180 503.840 ;
        RECT 259.080 503.580 259.340 503.840 ;
      LAYER met2 ;
        RECT 259.080 3298.350 259.340 3298.670 ;
        RECT 959.200 3298.350 959.460 3298.670 ;
        RECT 259.140 1014.210 259.280 3298.350 ;
        RECT 959.260 3258.970 959.400 3298.350 ;
        RECT 962.370 3258.970 962.650 3260.000 ;
        RECT 959.260 3258.830 962.650 3258.970 ;
        RECT 962.370 3256.000 962.650 3258.830 ;
        RECT 259.080 1013.890 259.340 1014.210 ;
        RECT 259.080 990.090 259.340 990.410 ;
        RECT 259.140 503.870 259.280 990.090 ;
        RECT 237.920 503.550 238.180 503.870 ;
        RECT 259.080 503.550 259.340 503.870 ;
        RECT 237.980 60.365 238.120 503.550 ;
        RECT 237.910 59.995 238.190 60.365 ;
        RECT 1406.310 59.995 1406.590 60.365 ;
        RECT 1406.380 2.400 1406.520 59.995 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
      LAYER via2 ;
        RECT 237.910 60.040 238.190 60.320 ;
        RECT 1406.310 60.040 1406.590 60.320 ;
      LAYER met3 ;
        RECT 237.885 60.330 238.215 60.345 ;
        RECT 1406.285 60.330 1406.615 60.345 ;
        RECT 237.885 60.030 1406.615 60.330 ;
        RECT 237.885 60.015 238.215 60.030 ;
        RECT 1406.285 60.015 1406.615 60.030 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1144.550 176.360 1144.870 176.420 ;
        RECT 1421.930 176.360 1422.250 176.420 ;
        RECT 1144.550 176.220 1422.250 176.360 ;
        RECT 1144.550 176.160 1144.870 176.220 ;
        RECT 1421.930 176.160 1422.250 176.220 ;
      LAYER via ;
        RECT 1144.580 176.160 1144.840 176.420 ;
        RECT 1421.960 176.160 1422.220 176.420 ;
      LAYER met2 ;
        RECT 1141.770 260.170 1142.050 264.000 ;
        RECT 1141.770 260.030 1144.780 260.170 ;
        RECT 1141.770 260.000 1142.050 260.030 ;
        RECT 1144.640 176.450 1144.780 260.030 ;
        RECT 1144.580 176.130 1144.840 176.450 ;
        RECT 1421.960 176.130 1422.220 176.450 ;
        RECT 1422.020 3.130 1422.160 176.130 ;
        RECT 1422.020 2.990 1424.000 3.130 ;
        RECT 1423.860 2.400 1424.000 2.990 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 299.530 258.980 299.850 259.040 ;
        RECT 1435.270 258.980 1435.590 259.040 ;
        RECT 299.530 258.840 1435.590 258.980 ;
        RECT 299.530 258.780 299.850 258.840 ;
        RECT 1435.270 258.780 1435.590 258.840 ;
        RECT 1435.270 15.880 1435.590 15.940 ;
        RECT 1441.710 15.880 1442.030 15.940 ;
        RECT 1435.270 15.740 1442.030 15.880 ;
        RECT 1435.270 15.680 1435.590 15.740 ;
        RECT 1441.710 15.680 1442.030 15.740 ;
      LAYER via ;
        RECT 299.560 258.780 299.820 259.040 ;
        RECT 1435.300 258.780 1435.560 259.040 ;
        RECT 1435.300 15.680 1435.560 15.940 ;
        RECT 1441.740 15.680 1442.000 15.940 ;
      LAYER met2 ;
        RECT 299.550 1278.555 299.830 1278.925 ;
        RECT 299.620 259.070 299.760 1278.555 ;
        RECT 299.560 258.750 299.820 259.070 ;
        RECT 1435.300 258.750 1435.560 259.070 ;
        RECT 1435.360 15.970 1435.500 258.750 ;
        RECT 1435.300 15.650 1435.560 15.970 ;
        RECT 1441.740 15.650 1442.000 15.970 ;
        RECT 1441.800 2.400 1441.940 15.650 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
      LAYER via2 ;
        RECT 299.550 1278.600 299.830 1278.880 ;
      LAYER met3 ;
        RECT 299.525 1278.890 299.855 1278.905 ;
        RECT 310.000 1278.890 314.000 1279.280 ;
        RECT 299.525 1278.680 314.000 1278.890 ;
        RECT 299.525 1278.590 310.500 1278.680 ;
        RECT 299.525 1278.575 299.855 1278.590 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 424.190 3272.060 424.510 3272.120 ;
        RECT 1348.790 3272.060 1349.110 3272.120 ;
        RECT 424.190 3271.920 1349.110 3272.060 ;
        RECT 424.190 3271.860 424.510 3271.920 ;
        RECT 1348.790 3271.860 1349.110 3271.920 ;
        RECT 315.630 3268.320 315.950 3268.380 ;
        RECT 424.190 3268.320 424.510 3268.380 ;
        RECT 315.630 3268.180 424.510 3268.320 ;
        RECT 315.630 3268.120 315.950 3268.180 ;
        RECT 424.190 3268.120 424.510 3268.180 ;
        RECT 315.630 60.420 315.950 60.480 ;
        RECT 1455.970 60.420 1456.290 60.480 ;
        RECT 315.630 60.280 1456.290 60.420 ;
        RECT 315.630 60.220 315.950 60.280 ;
        RECT 1455.970 60.220 1456.290 60.280 ;
        RECT 1455.970 2.960 1456.290 3.020 ;
        RECT 1459.650 2.960 1459.970 3.020 ;
        RECT 1455.970 2.820 1459.970 2.960 ;
        RECT 1455.970 2.760 1456.290 2.820 ;
        RECT 1459.650 2.760 1459.970 2.820 ;
      LAYER via ;
        RECT 424.220 3271.860 424.480 3272.120 ;
        RECT 1348.820 3271.860 1349.080 3272.120 ;
        RECT 315.660 3268.120 315.920 3268.380 ;
        RECT 424.220 3268.120 424.480 3268.380 ;
        RECT 315.660 60.220 315.920 60.480 ;
        RECT 1456.000 60.220 1456.260 60.480 ;
        RECT 1456.000 2.760 1456.260 3.020 ;
        RECT 1459.680 2.760 1459.940 3.020 ;
      LAYER met2 ;
        RECT 424.220 3271.830 424.480 3272.150 ;
        RECT 1348.820 3271.830 1349.080 3272.150 ;
        RECT 424.280 3268.410 424.420 3271.830 ;
        RECT 315.660 3268.090 315.920 3268.410 ;
        RECT 424.220 3268.090 424.480 3268.410 ;
        RECT 315.720 60.510 315.860 3268.090 ;
        RECT 1348.880 3260.000 1349.020 3271.830 ;
        RECT 1348.770 3256.000 1349.050 3260.000 ;
        RECT 315.660 60.190 315.920 60.510 ;
        RECT 1456.000 60.190 1456.260 60.510 ;
        RECT 1456.060 3.050 1456.200 60.190 ;
        RECT 1456.000 2.730 1456.260 3.050 ;
        RECT 1459.680 2.730 1459.940 3.050 ;
        RECT 1459.740 2.400 1459.880 2.730 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.870 3272.400 2521.190 3272.460 ;
        RECT 2685.090 3272.400 2685.410 3272.460 ;
        RECT 2520.870 3272.260 2685.410 3272.400 ;
        RECT 2520.870 3272.200 2521.190 3272.260 ;
        RECT 2685.090 3272.200 2685.410 3272.260 ;
        RECT 1483.110 227.360 1483.430 227.420 ;
        RECT 2685.090 227.360 2685.410 227.420 ;
        RECT 1483.110 227.220 2685.410 227.360 ;
        RECT 1483.110 227.160 1483.430 227.220 ;
        RECT 2685.090 227.160 2685.410 227.220 ;
        RECT 1477.590 20.640 1477.910 20.700 ;
        RECT 1483.110 20.640 1483.430 20.700 ;
        RECT 1477.590 20.500 1483.430 20.640 ;
        RECT 1477.590 20.440 1477.910 20.500 ;
        RECT 1483.110 20.440 1483.430 20.500 ;
      LAYER via ;
        RECT 2520.900 3272.200 2521.160 3272.460 ;
        RECT 2685.120 3272.200 2685.380 3272.460 ;
        RECT 1483.140 227.160 1483.400 227.420 ;
        RECT 2685.120 227.160 2685.380 227.420 ;
        RECT 1477.620 20.440 1477.880 20.700 ;
        RECT 1483.140 20.440 1483.400 20.700 ;
      LAYER met2 ;
        RECT 2520.900 3272.170 2521.160 3272.490 ;
        RECT 2685.120 3272.170 2685.380 3272.490 ;
        RECT 2520.960 3260.000 2521.100 3272.170 ;
        RECT 2520.850 3256.000 2521.130 3260.000 ;
        RECT 2685.180 227.450 2685.320 3272.170 ;
        RECT 1483.140 227.130 1483.400 227.450 ;
        RECT 2685.120 227.130 2685.380 227.450 ;
        RECT 1483.200 20.730 1483.340 227.130 ;
        RECT 1477.620 20.410 1477.880 20.730 ;
        RECT 1483.140 20.410 1483.400 20.730 ;
        RECT 1477.680 2.400 1477.820 20.410 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 275.150 3274.780 275.470 3274.840 ;
        RECT 476.630 3274.780 476.950 3274.840 ;
        RECT 275.150 3274.640 476.950 3274.780 ;
        RECT 275.150 3274.580 275.470 3274.640 ;
        RECT 476.630 3274.580 476.950 3274.640 ;
      LAYER via ;
        RECT 275.180 3274.580 275.440 3274.840 ;
        RECT 476.660 3274.580 476.920 3274.840 ;
      LAYER met2 ;
        RECT 275.180 3274.550 275.440 3274.870 ;
        RECT 476.660 3274.550 476.920 3274.870 ;
        RECT 275.240 18.885 275.380 3274.550 ;
        RECT 476.720 3260.000 476.860 3274.550 ;
        RECT 476.610 3256.000 476.890 3260.000 ;
        RECT 275.170 18.515 275.450 18.885 ;
        RECT 1495.550 18.515 1495.830 18.885 ;
        RECT 1495.620 2.400 1495.760 18.515 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
      LAYER via2 ;
        RECT 275.170 18.560 275.450 18.840 ;
        RECT 1495.550 18.560 1495.830 18.840 ;
      LAYER met3 ;
        RECT 275.145 18.850 275.475 18.865 ;
        RECT 1495.525 18.850 1495.855 18.865 ;
        RECT 275.145 18.550 1495.855 18.850 ;
        RECT 275.145 18.535 275.475 18.550 ;
        RECT 1495.525 18.535 1495.855 18.550 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1513.010 25.060 1513.330 25.120 ;
        RECT 1580.170 25.060 1580.490 25.120 ;
        RECT 1513.010 24.920 1580.490 25.060 ;
        RECT 1513.010 24.860 1513.330 24.920 ;
        RECT 1580.170 24.860 1580.490 24.920 ;
      LAYER via ;
        RECT 1513.040 24.860 1513.300 25.120 ;
        RECT 1580.200 24.860 1580.460 25.120 ;
      LAYER met2 ;
        RECT 1585.210 260.170 1585.490 264.000 ;
        RECT 1580.260 260.030 1585.490 260.170 ;
        RECT 1580.260 25.150 1580.400 260.030 ;
        RECT 1585.210 260.000 1585.490 260.030 ;
        RECT 1513.040 24.830 1513.300 25.150 ;
        RECT 1580.200 24.830 1580.460 25.150 ;
        RECT 1513.100 2.400 1513.240 24.830 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 292.170 538.460 292.490 538.520 ;
        RECT 297.230 538.460 297.550 538.520 ;
        RECT 292.170 538.320 297.550 538.460 ;
        RECT 292.170 538.260 292.490 538.320 ;
        RECT 297.230 538.260 297.550 538.320 ;
        RECT 292.170 238.240 292.490 238.300 ;
        RECT 703.870 238.240 704.190 238.300 ;
        RECT 292.170 238.100 704.190 238.240 ;
        RECT 292.170 238.040 292.490 238.100 ;
        RECT 703.870 238.040 704.190 238.100 ;
        RECT 703.870 37.640 704.190 37.700 ;
        RECT 710.310 37.640 710.630 37.700 ;
        RECT 703.870 37.500 710.630 37.640 ;
        RECT 703.870 37.440 704.190 37.500 ;
        RECT 710.310 37.440 710.630 37.500 ;
      LAYER via ;
        RECT 292.200 538.260 292.460 538.520 ;
        RECT 297.260 538.260 297.520 538.520 ;
        RECT 292.200 238.040 292.460 238.300 ;
        RECT 703.900 238.040 704.160 238.300 ;
        RECT 703.900 37.440 704.160 37.700 ;
        RECT 710.340 37.440 710.600 37.700 ;
      LAYER met2 ;
        RECT 297.250 538.715 297.530 539.085 ;
        RECT 297.320 538.550 297.460 538.715 ;
        RECT 292.200 538.230 292.460 538.550 ;
        RECT 297.260 538.230 297.520 538.550 ;
        RECT 292.260 238.330 292.400 538.230 ;
        RECT 292.200 238.010 292.460 238.330 ;
        RECT 703.900 238.010 704.160 238.330 ;
        RECT 703.960 37.730 704.100 238.010 ;
        RECT 703.900 37.410 704.160 37.730 ;
        RECT 710.340 37.410 710.600 37.730 ;
        RECT 710.400 2.400 710.540 37.410 ;
        RECT 710.190 -4.800 710.750 2.400 ;
      LAYER via2 ;
        RECT 297.250 538.760 297.530 539.040 ;
      LAYER met3 ;
        RECT 297.225 539.050 297.555 539.065 ;
        RECT 310.000 539.050 314.000 539.440 ;
        RECT 297.225 538.840 314.000 539.050 ;
        RECT 297.225 538.750 310.500 538.840 ;
        RECT 297.225 538.735 297.555 538.750 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.550 227.020 293.870 227.080 ;
        RECT 1524.970 227.020 1525.290 227.080 ;
        RECT 293.550 226.880 1525.290 227.020 ;
        RECT 293.550 226.820 293.870 226.880 ;
        RECT 1524.970 226.820 1525.290 226.880 ;
        RECT 1524.970 37.640 1525.290 37.700 ;
        RECT 1530.950 37.640 1531.270 37.700 ;
        RECT 1524.970 37.500 1531.270 37.640 ;
        RECT 1524.970 37.440 1525.290 37.500 ;
        RECT 1530.950 37.440 1531.270 37.500 ;
      LAYER via ;
        RECT 293.580 226.820 293.840 227.080 ;
        RECT 1525.000 226.820 1525.260 227.080 ;
        RECT 1525.000 37.440 1525.260 37.700 ;
        RECT 1530.980 37.440 1531.240 37.700 ;
      LAYER met2 ;
        RECT 293.570 1256.795 293.850 1257.165 ;
        RECT 293.640 227.110 293.780 1256.795 ;
        RECT 293.580 226.790 293.840 227.110 ;
        RECT 1525.000 226.790 1525.260 227.110 ;
        RECT 1525.060 37.730 1525.200 226.790 ;
        RECT 1525.000 37.410 1525.260 37.730 ;
        RECT 1530.980 37.410 1531.240 37.730 ;
        RECT 1531.040 2.400 1531.180 37.410 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
      LAYER via2 ;
        RECT 293.570 1256.840 293.850 1257.120 ;
      LAYER met3 ;
        RECT 293.545 1257.130 293.875 1257.145 ;
        RECT 310.000 1257.130 314.000 1257.520 ;
        RECT 293.545 1256.920 314.000 1257.130 ;
        RECT 293.545 1256.830 310.500 1256.920 ;
        RECT 293.545 1256.815 293.875 1256.830 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 232.830 2670.600 233.150 2670.660 ;
        RECT 296.770 2670.600 297.090 2670.660 ;
        RECT 232.830 2670.460 297.090 2670.600 ;
        RECT 232.830 2670.400 233.150 2670.460 ;
        RECT 296.770 2670.400 297.090 2670.460 ;
      LAYER via ;
        RECT 232.860 2670.400 233.120 2670.660 ;
        RECT 296.800 2670.400 297.060 2670.660 ;
      LAYER met2 ;
        RECT 296.790 2672.555 297.070 2672.925 ;
        RECT 296.860 2670.690 297.000 2672.555 ;
        RECT 232.860 2670.370 233.120 2670.690 ;
        RECT 296.800 2670.370 297.060 2670.690 ;
        RECT 232.920 59.685 233.060 2670.370 ;
        RECT 232.850 59.315 233.130 59.685 ;
        RECT 1548.910 59.315 1549.190 59.685 ;
        RECT 1548.980 2.400 1549.120 59.315 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
      LAYER via2 ;
        RECT 296.790 2672.600 297.070 2672.880 ;
        RECT 232.850 59.360 233.130 59.640 ;
        RECT 1548.910 59.360 1549.190 59.640 ;
      LAYER met3 ;
        RECT 296.765 2672.890 297.095 2672.905 ;
        RECT 310.000 2672.890 314.000 2673.280 ;
        RECT 296.765 2672.680 314.000 2672.890 ;
        RECT 296.765 2672.590 310.500 2672.680 ;
        RECT 296.765 2672.575 297.095 2672.590 ;
        RECT 232.825 59.650 233.155 59.665 ;
        RECT 1548.885 59.650 1549.215 59.665 ;
        RECT 232.825 59.350 1549.215 59.650 ;
        RECT 232.825 59.335 233.155 59.350 ;
        RECT 1548.885 59.335 1549.215 59.350 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1566.445 48.365 1566.615 96.475 ;
      LAYER mcon ;
        RECT 1566.445 96.305 1566.615 96.475 ;
      LAYER met1 ;
        RECT 1357.990 129.100 1358.310 129.160 ;
        RECT 1566.370 129.100 1566.690 129.160 ;
        RECT 1357.990 128.960 1566.690 129.100 ;
        RECT 1357.990 128.900 1358.310 128.960 ;
        RECT 1566.370 128.900 1566.690 128.960 ;
        RECT 1566.370 96.460 1566.690 96.520 ;
        RECT 1566.175 96.320 1566.690 96.460 ;
        RECT 1566.370 96.260 1566.690 96.320 ;
        RECT 1566.385 48.520 1566.675 48.565 ;
        RECT 1566.830 48.520 1567.150 48.580 ;
        RECT 1566.385 48.380 1567.150 48.520 ;
        RECT 1566.385 48.335 1566.675 48.380 ;
        RECT 1566.830 48.320 1567.150 48.380 ;
      LAYER via ;
        RECT 1358.020 128.900 1358.280 129.160 ;
        RECT 1566.400 128.900 1566.660 129.160 ;
        RECT 1566.400 96.260 1566.660 96.520 ;
        RECT 1566.860 48.320 1567.120 48.580 ;
      LAYER met2 ;
        RECT 1356.130 260.170 1356.410 264.000 ;
        RECT 1356.130 260.030 1358.220 260.170 ;
        RECT 1356.130 260.000 1356.410 260.030 ;
        RECT 1358.080 129.190 1358.220 260.030 ;
        RECT 1358.020 128.870 1358.280 129.190 ;
        RECT 1566.400 128.870 1566.660 129.190 ;
        RECT 1566.460 96.550 1566.600 128.870 ;
        RECT 1566.400 96.230 1566.660 96.550 ;
        RECT 1566.860 48.290 1567.120 48.610 ;
        RECT 1566.920 2.400 1567.060 48.290 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.610 234.500 1586.930 234.560 ;
        RECT 2622.530 234.500 2622.850 234.560 ;
        RECT 1586.610 234.360 2622.850 234.500 ;
        RECT 1586.610 234.300 1586.930 234.360 ;
        RECT 2622.530 234.300 2622.850 234.360 ;
        RECT 1586.610 62.460 1586.930 62.520 ;
        RECT 1584.860 62.320 1586.930 62.460 ;
        RECT 1584.860 62.180 1585.000 62.320 ;
        RECT 1586.610 62.260 1586.930 62.320 ;
        RECT 1584.770 61.920 1585.090 62.180 ;
      LAYER via ;
        RECT 1586.640 234.300 1586.900 234.560 ;
        RECT 2622.560 234.300 2622.820 234.560 ;
        RECT 1586.640 62.260 1586.900 62.520 ;
        RECT 1584.800 61.920 1585.060 62.180 ;
      LAYER met2 ;
        RECT 2622.550 2811.275 2622.830 2811.645 ;
        RECT 2622.620 234.590 2622.760 2811.275 ;
        RECT 1586.640 234.270 1586.900 234.590 ;
        RECT 2622.560 234.270 2622.820 234.590 ;
        RECT 1586.700 62.550 1586.840 234.270 ;
        RECT 1586.640 62.230 1586.900 62.550 ;
        RECT 1584.800 61.890 1585.060 62.210 ;
        RECT 1584.860 2.400 1585.000 61.890 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
      LAYER via2 ;
        RECT 2622.550 2811.320 2622.830 2811.600 ;
      LAYER met3 ;
        RECT 2606.000 2811.610 2610.000 2812.000 ;
        RECT 2622.525 2811.610 2622.855 2811.625 ;
        RECT 2606.000 2811.400 2622.855 2811.610 ;
        RECT 2609.580 2811.310 2622.855 2811.400 ;
        RECT 2622.525 2811.295 2622.855 2811.310 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1602.325 2.805 1602.495 41.395 ;
      LAYER mcon ;
        RECT 1602.325 41.225 1602.495 41.395 ;
      LAYER met1 ;
        RECT 292.630 745.520 292.950 745.580 ;
        RECT 298.610 745.520 298.930 745.580 ;
        RECT 292.630 745.380 298.930 745.520 ;
        RECT 292.630 745.320 292.950 745.380 ;
        RECT 298.610 745.320 298.930 745.380 ;
        RECT 292.630 197.780 292.950 197.840 ;
        RECT 1600.870 197.780 1601.190 197.840 ;
        RECT 292.630 197.640 1601.190 197.780 ;
        RECT 292.630 197.580 292.950 197.640 ;
        RECT 1600.870 197.580 1601.190 197.640 ;
        RECT 1600.870 41.380 1601.190 41.440 ;
        RECT 1602.265 41.380 1602.555 41.425 ;
        RECT 1600.870 41.240 1602.555 41.380 ;
        RECT 1600.870 41.180 1601.190 41.240 ;
        RECT 1602.265 41.195 1602.555 41.240 ;
        RECT 1602.250 2.960 1602.570 3.020 ;
        RECT 1602.055 2.820 1602.570 2.960 ;
        RECT 1602.250 2.760 1602.570 2.820 ;
      LAYER via ;
        RECT 292.660 745.320 292.920 745.580 ;
        RECT 298.640 745.320 298.900 745.580 ;
        RECT 292.660 197.580 292.920 197.840 ;
        RECT 1600.900 197.580 1601.160 197.840 ;
        RECT 1600.900 41.180 1601.160 41.440 ;
        RECT 1602.280 2.760 1602.540 3.020 ;
      LAYER met2 ;
        RECT 298.630 749.515 298.910 749.885 ;
        RECT 298.700 745.610 298.840 749.515 ;
        RECT 292.660 745.290 292.920 745.610 ;
        RECT 298.640 745.290 298.900 745.610 ;
        RECT 292.720 197.870 292.860 745.290 ;
        RECT 292.660 197.550 292.920 197.870 ;
        RECT 1600.900 197.550 1601.160 197.870 ;
        RECT 1600.960 41.470 1601.100 197.550 ;
        RECT 1600.900 41.150 1601.160 41.470 ;
        RECT 1602.280 2.730 1602.540 3.050 ;
        RECT 1602.340 2.400 1602.480 2.730 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
      LAYER via2 ;
        RECT 298.630 749.560 298.910 749.840 ;
      LAYER met3 ;
        RECT 298.605 749.850 298.935 749.865 ;
        RECT 310.000 749.850 314.000 750.240 ;
        RECT 298.605 749.640 314.000 749.850 ;
        RECT 298.605 749.550 310.500 749.640 ;
        RECT 298.605 749.535 298.935 749.550 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1620.265 2.805 1620.435 14.195 ;
      LAYER mcon ;
        RECT 1620.265 14.025 1620.435 14.195 ;
      LAYER met1 ;
        RECT 2165.290 3260.160 2165.610 3260.220 ;
        RECT 2691.530 3260.160 2691.850 3260.220 ;
        RECT 2165.290 3260.020 2691.850 3260.160 ;
        RECT 2165.290 3259.960 2165.610 3260.020 ;
        RECT 2691.530 3259.960 2691.850 3260.020 ;
        RECT 1621.110 233.820 1621.430 233.880 ;
        RECT 2691.530 233.820 2691.850 233.880 ;
        RECT 1621.110 233.680 2691.850 233.820 ;
        RECT 1621.110 233.620 1621.430 233.680 ;
        RECT 2691.530 233.620 2691.850 233.680 ;
        RECT 1620.205 14.180 1620.495 14.225 ;
        RECT 1621.110 14.180 1621.430 14.240 ;
        RECT 1620.205 14.040 1621.430 14.180 ;
        RECT 1620.205 13.995 1620.495 14.040 ;
        RECT 1621.110 13.980 1621.430 14.040 ;
        RECT 1620.190 2.960 1620.510 3.020 ;
        RECT 1619.995 2.820 1620.510 2.960 ;
        RECT 1620.190 2.760 1620.510 2.820 ;
      LAYER via ;
        RECT 2165.320 3259.960 2165.580 3260.220 ;
        RECT 2691.560 3259.960 2691.820 3260.220 ;
        RECT 1621.140 233.620 1621.400 233.880 ;
        RECT 2691.560 233.620 2691.820 233.880 ;
        RECT 1621.140 13.980 1621.400 14.240 ;
        RECT 1620.220 2.760 1620.480 3.020 ;
      LAYER met2 ;
        RECT 2163.890 3259.650 2164.170 3260.000 ;
        RECT 2165.320 3259.930 2165.580 3260.250 ;
        RECT 2691.560 3259.930 2691.820 3260.250 ;
        RECT 2165.380 3259.650 2165.520 3259.930 ;
        RECT 2163.890 3259.510 2165.520 3259.650 ;
        RECT 2163.890 3256.000 2164.170 3259.510 ;
        RECT 2691.620 233.910 2691.760 3259.930 ;
        RECT 1621.140 233.590 1621.400 233.910 ;
        RECT 2691.560 233.590 2691.820 233.910 ;
        RECT 1621.200 14.270 1621.340 233.590 ;
        RECT 1621.140 13.950 1621.400 14.270 ;
        RECT 1620.220 2.730 1620.480 3.050 ;
        RECT 1620.280 2.400 1620.420 2.730 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2607.885 262.565 2608.055 272.935 ;
        RECT 2428.485 20.145 2429.115 20.315 ;
        RECT 2428.945 17.765 2429.115 20.145 ;
      LAYER mcon ;
        RECT 2607.885 272.765 2608.055 272.935 ;
      LAYER met1 ;
        RECT 1691.950 3265.260 1692.270 3265.320 ;
        RECT 2615.630 3265.260 2615.950 3265.320 ;
        RECT 1691.950 3265.120 2615.950 3265.260 ;
        RECT 1691.950 3265.060 1692.270 3265.120 ;
        RECT 2615.630 3265.060 2615.950 3265.120 ;
        RECT 2611.490 490.180 2611.810 490.240 ;
        RECT 2615.630 490.180 2615.950 490.240 ;
        RECT 2611.490 490.040 2615.950 490.180 ;
        RECT 2611.490 489.980 2611.810 490.040 ;
        RECT 2615.630 489.980 2615.950 490.040 ;
        RECT 2607.810 272.920 2608.130 272.980 ;
        RECT 2607.615 272.780 2608.130 272.920 ;
        RECT 2607.810 272.720 2608.130 272.780 ;
        RECT 2605.970 262.720 2606.290 262.780 ;
        RECT 2607.825 262.720 2608.115 262.765 ;
        RECT 2605.970 262.580 2608.115 262.720 ;
        RECT 2605.970 262.520 2606.290 262.580 ;
        RECT 2607.825 262.535 2608.115 262.580 ;
        RECT 1638.130 20.300 1638.450 20.360 ;
        RECT 2428.425 20.300 2428.715 20.345 ;
        RECT 1638.130 20.160 2428.715 20.300 ;
        RECT 1638.130 20.100 1638.450 20.160 ;
        RECT 2428.425 20.115 2428.715 20.160 ;
        RECT 2428.885 17.920 2429.175 17.965 ;
        RECT 2445.890 17.920 2446.210 17.980 ;
        RECT 2428.885 17.780 2446.210 17.920 ;
        RECT 2428.885 17.735 2429.175 17.780 ;
        RECT 2445.890 17.720 2446.210 17.780 ;
      LAYER via ;
        RECT 1691.980 3265.060 1692.240 3265.320 ;
        RECT 2615.660 3265.060 2615.920 3265.320 ;
        RECT 2611.520 489.980 2611.780 490.240 ;
        RECT 2615.660 489.980 2615.920 490.240 ;
        RECT 2607.840 272.720 2608.100 272.980 ;
        RECT 2606.000 262.520 2606.260 262.780 ;
        RECT 1638.160 20.100 1638.420 20.360 ;
        RECT 2445.920 17.720 2446.180 17.980 ;
      LAYER met2 ;
        RECT 1691.980 3265.030 1692.240 3265.350 ;
        RECT 2615.660 3265.030 2615.920 3265.350 ;
        RECT 1692.040 3260.000 1692.180 3265.030 ;
        RECT 1691.930 3256.000 1692.210 3260.000 ;
        RECT 2615.720 490.270 2615.860 3265.030 ;
        RECT 2611.520 489.950 2611.780 490.270 ;
        RECT 2615.660 489.950 2615.920 490.270 ;
        RECT 2611.580 352.085 2611.720 489.950 ;
        RECT 2611.510 351.715 2611.790 352.085 ;
        RECT 2607.830 280.315 2608.110 280.685 ;
        RECT 2607.900 273.010 2608.040 280.315 ;
        RECT 2607.840 272.690 2608.100 273.010 ;
        RECT 2605.990 262.635 2606.270 263.005 ;
        RECT 2606.000 262.490 2606.260 262.635 ;
        RECT 2445.910 234.075 2446.190 234.445 ;
        RECT 1638.160 20.070 1638.420 20.390 ;
        RECT 1638.220 2.400 1638.360 20.070 ;
        RECT 2445.980 18.010 2446.120 234.075 ;
        RECT 2445.920 17.690 2446.180 18.010 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
      LAYER via2 ;
        RECT 2611.510 351.760 2611.790 352.040 ;
        RECT 2607.830 280.360 2608.110 280.640 ;
        RECT 2605.990 262.680 2606.270 262.960 ;
        RECT 2445.910 234.120 2446.190 234.400 ;
      LAYER met3 ;
        RECT 2606.630 352.050 2607.010 352.060 ;
        RECT 2611.485 352.050 2611.815 352.065 ;
        RECT 2606.630 351.750 2611.815 352.050 ;
        RECT 2606.630 351.740 2607.010 351.750 ;
        RECT 2611.485 351.735 2611.815 351.750 ;
        RECT 2606.630 280.650 2607.010 280.660 ;
        RECT 2607.805 280.650 2608.135 280.665 ;
        RECT 2606.630 280.350 2608.135 280.650 ;
        RECT 2606.630 280.340 2607.010 280.350 ;
        RECT 2607.805 280.335 2608.135 280.350 ;
        RECT 2605.965 262.980 2606.295 262.985 ;
        RECT 2605.710 262.970 2606.295 262.980 ;
        RECT 2605.510 262.670 2606.295 262.970 ;
        RECT 2605.710 262.660 2606.295 262.670 ;
        RECT 2605.965 262.655 2606.295 262.660 ;
        RECT 2445.885 234.410 2446.215 234.425 ;
        RECT 2605.710 234.410 2606.090 234.420 ;
        RECT 2445.885 234.110 2606.090 234.410 ;
        RECT 2445.885 234.095 2446.215 234.110 ;
        RECT 2605.710 234.100 2606.090 234.110 ;
      LAYER via3 ;
        RECT 2606.660 351.740 2606.980 352.060 ;
        RECT 2606.660 280.340 2606.980 280.660 ;
        RECT 2605.740 262.660 2606.060 262.980 ;
        RECT 2605.740 234.100 2606.060 234.420 ;
      LAYER met4 ;
        RECT 2606.655 351.735 2606.985 352.065 ;
        RECT 2606.670 280.665 2606.970 351.735 ;
        RECT 2606.655 280.335 2606.985 280.665 ;
        RECT 2605.735 262.655 2606.065 262.985 ;
        RECT 2605.750 234.425 2606.050 262.655 ;
        RECT 2605.735 234.095 2606.065 234.425 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 258.980 1662.830 259.040 ;
        RECT 2623.910 258.980 2624.230 259.040 ;
        RECT 1662.510 258.840 2624.230 258.980 ;
        RECT 1662.510 258.780 1662.830 258.840 ;
        RECT 2623.910 258.780 2624.230 258.840 ;
        RECT 1656.070 15.880 1656.390 15.940 ;
        RECT 1662.510 15.880 1662.830 15.940 ;
        RECT 1656.070 15.740 1662.830 15.880 ;
        RECT 1656.070 15.680 1656.390 15.740 ;
        RECT 1662.510 15.680 1662.830 15.740 ;
      LAYER via ;
        RECT 1662.540 258.780 1662.800 259.040 ;
        RECT 2623.940 258.780 2624.200 259.040 ;
        RECT 1656.100 15.680 1656.360 15.940 ;
        RECT 1662.540 15.680 1662.800 15.940 ;
      LAYER met2 ;
        RECT 2623.930 1437.675 2624.210 1438.045 ;
        RECT 2624.000 259.070 2624.140 1437.675 ;
        RECT 1662.540 258.750 1662.800 259.070 ;
        RECT 2623.940 258.750 2624.200 259.070 ;
        RECT 1662.600 15.970 1662.740 258.750 ;
        RECT 1656.100 15.650 1656.360 15.970 ;
        RECT 1662.540 15.650 1662.800 15.970 ;
        RECT 1656.160 2.400 1656.300 15.650 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
      LAYER via2 ;
        RECT 2623.930 1437.720 2624.210 1438.000 ;
      LAYER met3 ;
        RECT 2606.000 1438.010 2610.000 1438.400 ;
        RECT 2623.905 1438.010 2624.235 1438.025 ;
        RECT 2606.000 1437.800 2624.235 1438.010 ;
        RECT 2609.580 1437.710 2624.235 1437.800 ;
        RECT 2623.905 1437.695 2624.235 1437.710 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1456.430 244.020 1456.750 244.080 ;
        RECT 1462.410 244.020 1462.730 244.080 ;
        RECT 1456.430 243.880 1462.730 244.020 ;
        RECT 1456.430 243.820 1456.750 243.880 ;
        RECT 1462.410 243.820 1462.730 243.880 ;
        RECT 1462.410 33.900 1462.730 33.960 ;
        RECT 1673.550 33.900 1673.870 33.960 ;
        RECT 1462.410 33.760 1673.870 33.900 ;
        RECT 1462.410 33.700 1462.730 33.760 ;
        RECT 1673.550 33.700 1673.870 33.760 ;
      LAYER via ;
        RECT 1456.460 243.820 1456.720 244.080 ;
        RECT 1462.440 243.820 1462.700 244.080 ;
        RECT 1462.440 33.700 1462.700 33.960 ;
        RECT 1673.580 33.700 1673.840 33.960 ;
      LAYER met2 ;
        RECT 1456.410 260.000 1456.690 264.000 ;
        RECT 1456.520 244.110 1456.660 260.000 ;
        RECT 1456.460 243.790 1456.720 244.110 ;
        RECT 1462.440 243.790 1462.700 244.110 ;
        RECT 1462.500 33.990 1462.640 243.790 ;
        RECT 1462.440 33.670 1462.700 33.990 ;
        RECT 1673.580 33.670 1673.840 33.990 ;
        RECT 1673.640 2.400 1673.780 33.670 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 260.890 766.260 261.210 766.320 ;
        RECT 296.770 766.260 297.090 766.320 ;
        RECT 260.890 766.120 297.090 766.260 ;
        RECT 260.890 766.060 261.210 766.120 ;
        RECT 296.770 766.060 297.090 766.120 ;
        RECT 260.890 60.080 261.210 60.140 ;
        RECT 1691.490 60.080 1691.810 60.140 ;
        RECT 260.890 59.940 1691.810 60.080 ;
        RECT 260.890 59.880 261.210 59.940 ;
        RECT 1691.490 59.880 1691.810 59.940 ;
      LAYER via ;
        RECT 260.920 766.060 261.180 766.320 ;
        RECT 296.800 766.060 297.060 766.320 ;
        RECT 260.920 59.880 261.180 60.140 ;
        RECT 1691.520 59.880 1691.780 60.140 ;
      LAYER met2 ;
        RECT 296.790 771.275 297.070 771.645 ;
        RECT 296.860 766.350 297.000 771.275 ;
        RECT 260.920 766.030 261.180 766.350 ;
        RECT 296.800 766.030 297.060 766.350 ;
        RECT 260.980 60.170 261.120 766.030 ;
        RECT 260.920 59.850 261.180 60.170 ;
        RECT 1691.520 59.850 1691.780 60.170 ;
        RECT 1691.580 2.400 1691.720 59.850 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
      LAYER via2 ;
        RECT 296.790 771.320 297.070 771.600 ;
      LAYER met3 ;
        RECT 296.765 771.610 297.095 771.625 ;
        RECT 310.000 771.610 314.000 772.000 ;
        RECT 296.765 771.400 314.000 771.610 ;
        RECT 296.765 771.310 310.500 771.400 ;
        RECT 296.765 771.295 297.095 771.310 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2656.660 2615.490 2656.720 ;
        RECT 2672.670 2656.660 2672.990 2656.720 ;
        RECT 2615.170 2656.520 2672.990 2656.660 ;
        RECT 2615.170 2656.460 2615.490 2656.520 ;
        RECT 2672.670 2656.460 2672.990 2656.520 ;
        RECT 731.010 224.300 731.330 224.360 ;
        RECT 2672.670 224.300 2672.990 224.360 ;
        RECT 731.010 224.160 2672.990 224.300 ;
        RECT 731.010 224.100 731.330 224.160 ;
        RECT 2672.670 224.100 2672.990 224.160 ;
        RECT 728.250 20.640 728.570 20.700 ;
        RECT 731.010 20.640 731.330 20.700 ;
        RECT 728.250 20.500 731.330 20.640 ;
        RECT 728.250 20.440 728.570 20.500 ;
        RECT 731.010 20.440 731.330 20.500 ;
      LAYER via ;
        RECT 2615.200 2656.460 2615.460 2656.720 ;
        RECT 2672.700 2656.460 2672.960 2656.720 ;
        RECT 731.040 224.100 731.300 224.360 ;
        RECT 2672.700 224.100 2672.960 224.360 ;
        RECT 728.280 20.440 728.540 20.700 ;
        RECT 731.040 20.440 731.300 20.700 ;
      LAYER met2 ;
        RECT 2615.190 2663.035 2615.470 2663.405 ;
        RECT 2615.260 2656.750 2615.400 2663.035 ;
        RECT 2615.200 2656.430 2615.460 2656.750 ;
        RECT 2672.700 2656.430 2672.960 2656.750 ;
        RECT 2672.760 224.390 2672.900 2656.430 ;
        RECT 731.040 224.070 731.300 224.390 ;
        RECT 2672.700 224.070 2672.960 224.390 ;
        RECT 731.100 20.730 731.240 224.070 ;
        RECT 728.280 20.410 728.540 20.730 ;
        RECT 731.040 20.410 731.300 20.730 ;
        RECT 728.340 2.400 728.480 20.410 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2663.080 2615.470 2663.360 ;
      LAYER met3 ;
        RECT 2606.000 2663.370 2610.000 2663.760 ;
        RECT 2615.165 2663.370 2615.495 2663.385 ;
        RECT 2606.000 2663.160 2615.495 2663.370 ;
        RECT 2609.580 2663.070 2615.495 2663.160 ;
        RECT 2615.165 2663.055 2615.495 2663.070 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1709.505 48.365 1709.675 62.475 ;
      LAYER mcon ;
        RECT 1709.505 62.305 1709.675 62.475 ;
      LAYER met1 ;
        RECT 1710.810 259.320 1711.130 259.380 ;
        RECT 2621.150 259.320 2621.470 259.380 ;
        RECT 1710.810 259.180 2621.470 259.320 ;
        RECT 1710.810 259.120 1711.130 259.180 ;
        RECT 2621.150 259.120 2621.470 259.180 ;
        RECT 1709.445 62.460 1709.735 62.505 ;
        RECT 1710.810 62.460 1711.130 62.520 ;
        RECT 1709.445 62.320 1711.130 62.460 ;
        RECT 1709.445 62.275 1709.735 62.320 ;
        RECT 1710.810 62.260 1711.130 62.320 ;
        RECT 1709.430 48.520 1709.750 48.580 ;
        RECT 1709.235 48.380 1709.750 48.520 ;
        RECT 1709.430 48.320 1709.750 48.380 ;
      LAYER via ;
        RECT 1710.840 259.120 1711.100 259.380 ;
        RECT 2621.180 259.120 2621.440 259.380 ;
        RECT 1710.840 62.260 1711.100 62.520 ;
        RECT 1709.460 48.320 1709.720 48.580 ;
      LAYER met2 ;
        RECT 2621.170 359.195 2621.450 359.565 ;
        RECT 2621.240 259.410 2621.380 359.195 ;
        RECT 1710.840 259.090 1711.100 259.410 ;
        RECT 2621.180 259.090 2621.440 259.410 ;
        RECT 1710.900 62.550 1711.040 259.090 ;
        RECT 1710.840 62.230 1711.100 62.550 ;
        RECT 1709.460 48.290 1709.720 48.610 ;
        RECT 1709.520 2.400 1709.660 48.290 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
      LAYER via2 ;
        RECT 2621.170 359.240 2621.450 359.520 ;
      LAYER met3 ;
        RECT 2606.000 359.530 2610.000 359.920 ;
        RECT 2621.145 359.530 2621.475 359.545 ;
        RECT 2606.000 359.320 2621.475 359.530 ;
        RECT 2609.580 359.230 2621.475 359.320 ;
        RECT 2621.145 359.215 2621.475 359.230 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1576.950 3272.400 1577.270 3272.460 ;
        RECT 2518.110 3272.400 2518.430 3272.460 ;
        RECT 1576.950 3272.260 2518.430 3272.400 ;
        RECT 1576.950 3272.200 1577.270 3272.260 ;
        RECT 2518.110 3272.200 2518.430 3272.260 ;
        RECT 1727.370 34.580 1727.690 34.640 ;
        RECT 1731.510 34.580 1731.830 34.640 ;
        RECT 1727.370 34.440 1731.830 34.580 ;
        RECT 1727.370 34.380 1727.690 34.440 ;
        RECT 1731.510 34.380 1731.830 34.440 ;
      LAYER via ;
        RECT 1576.980 3272.200 1577.240 3272.460 ;
        RECT 2518.140 3272.200 2518.400 3272.460 ;
        RECT 1727.400 34.380 1727.660 34.640 ;
        RECT 1731.540 34.380 1731.800 34.640 ;
      LAYER met2 ;
        RECT 1576.980 3272.170 1577.240 3272.490 ;
        RECT 2518.140 3272.170 2518.400 3272.490 ;
        RECT 1577.040 3260.000 1577.180 3272.170 ;
        RECT 2518.200 3261.125 2518.340 3272.170 ;
        RECT 2518.130 3260.755 2518.410 3261.125 ;
        RECT 1576.930 3256.000 1577.210 3260.000 ;
        RECT 1727.400 34.350 1727.660 34.670 ;
        RECT 1731.540 34.525 1731.800 34.670 ;
        RECT 1727.460 2.400 1727.600 34.350 ;
        RECT 1731.530 34.155 1731.810 34.525 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
      LAYER via2 ;
        RECT 2518.130 3260.800 2518.410 3261.080 ;
        RECT 1731.530 34.200 1731.810 34.480 ;
      LAYER met3 ;
        RECT 2518.105 3261.090 2518.435 3261.105 ;
        RECT 2590.990 3261.090 2591.370 3261.100 ;
        RECT 2518.105 3260.790 2591.370 3261.090 ;
        RECT 2518.105 3260.775 2518.435 3260.790 ;
        RECT 2590.990 3260.780 2591.370 3260.790 ;
        RECT 1731.505 34.490 1731.835 34.505 ;
        RECT 2590.990 34.490 2591.370 34.500 ;
        RECT 1731.505 34.190 2591.370 34.490 ;
        RECT 1731.505 34.175 1731.835 34.190 ;
        RECT 2590.990 34.180 2591.370 34.190 ;
      LAYER via3 ;
        RECT 2591.020 3260.780 2591.340 3261.100 ;
        RECT 2591.020 34.180 2591.340 34.500 ;
      LAYER met4 ;
        RECT 2591.015 3260.775 2591.345 3261.105 ;
        RECT 2591.030 34.505 2591.330 3260.775 ;
        RECT 2591.015 34.175 2591.345 34.505 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1897.780 2615.490 1897.840 ;
        RECT 2693.370 1897.780 2693.690 1897.840 ;
        RECT 2615.170 1897.640 2693.690 1897.780 ;
        RECT 2615.170 1897.580 2615.490 1897.640 ;
        RECT 2693.370 1897.580 2693.690 1897.640 ;
        RECT 1744.850 230.420 1745.170 230.480 ;
        RECT 2693.370 230.420 2693.690 230.480 ;
        RECT 1744.850 230.280 2693.690 230.420 ;
        RECT 1744.850 230.220 1745.170 230.280 ;
        RECT 2693.370 230.220 2693.690 230.280 ;
      LAYER via ;
        RECT 2615.200 1897.580 2615.460 1897.840 ;
        RECT 2693.400 1897.580 2693.660 1897.840 ;
        RECT 1744.880 230.220 1745.140 230.480 ;
        RECT 2693.400 230.220 2693.660 230.480 ;
      LAYER met2 ;
        RECT 2615.190 1902.795 2615.470 1903.165 ;
        RECT 2615.260 1897.870 2615.400 1902.795 ;
        RECT 2615.200 1897.550 2615.460 1897.870 ;
        RECT 2693.400 1897.550 2693.660 1897.870 ;
        RECT 2693.460 230.510 2693.600 1897.550 ;
        RECT 1744.880 230.190 1745.140 230.510 ;
        RECT 2693.400 230.190 2693.660 230.510 ;
        RECT 1744.940 7.890 1745.080 230.190 ;
        RECT 1744.940 7.750 1745.540 7.890 ;
        RECT 1745.400 2.400 1745.540 7.750 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1902.840 2615.470 1903.120 ;
      LAYER met3 ;
        RECT 2606.000 1903.130 2610.000 1903.520 ;
        RECT 2615.165 1903.130 2615.495 1903.145 ;
        RECT 2606.000 1902.920 2615.495 1903.130 ;
        RECT 2609.580 1902.830 2615.495 1902.920 ;
        RECT 2615.165 1902.815 2615.495 1902.830 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1013.985 30.345 1014.155 39.355 ;
      LAYER mcon ;
        RECT 1013.985 39.185 1014.155 39.355 ;
      LAYER met1 ;
        RECT 1013.910 39.340 1014.230 39.400 ;
        RECT 1013.715 39.200 1014.230 39.340 ;
        RECT 1013.910 39.140 1014.230 39.200 ;
        RECT 1013.925 30.500 1014.215 30.545 ;
        RECT 1762.790 30.500 1763.110 30.560 ;
        RECT 1013.925 30.360 1763.110 30.500 ;
        RECT 1013.925 30.315 1014.215 30.360 ;
        RECT 1762.790 30.300 1763.110 30.360 ;
      LAYER via ;
        RECT 1013.940 39.140 1014.200 39.400 ;
        RECT 1762.820 30.300 1763.080 30.560 ;
      LAYER met2 ;
        RECT 1012.970 260.170 1013.250 264.000 ;
        RECT 1012.970 260.030 1014.140 260.170 ;
        RECT 1012.970 260.000 1013.250 260.030 ;
        RECT 1014.000 39.430 1014.140 260.030 ;
        RECT 1013.940 39.110 1014.200 39.430 ;
        RECT 1762.820 30.270 1763.080 30.590 ;
        RECT 1762.880 2.400 1763.020 30.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1993.250 3256.220 1993.570 3256.480 ;
        RECT 1993.340 3254.380 1993.480 3256.220 ;
        RECT 2644.150 3254.380 2644.470 3254.440 ;
        RECT 1993.340 3254.240 2644.470 3254.380 ;
        RECT 2644.150 3254.180 2644.470 3254.240 ;
        RECT 2614.710 283.120 2615.030 283.180 ;
        RECT 2644.150 283.120 2644.470 283.180 ;
        RECT 2614.710 282.980 2644.470 283.120 ;
        RECT 2614.710 282.920 2615.030 282.980 ;
        RECT 2644.150 282.920 2644.470 282.980 ;
        RECT 2466.590 244.020 2466.910 244.080 ;
        RECT 2614.710 244.020 2615.030 244.080 ;
        RECT 2466.590 243.880 2615.030 244.020 ;
        RECT 2466.590 243.820 2466.910 243.880 ;
        RECT 2614.710 243.820 2615.030 243.880 ;
        RECT 2428.960 20.840 2435.540 20.980 ;
        RECT 1780.730 20.640 1781.050 20.700 ;
        RECT 2428.960 20.640 2429.100 20.840 ;
        RECT 1780.730 20.500 2429.100 20.640 ;
        RECT 1780.730 20.440 1781.050 20.500 ;
        RECT 2435.400 20.300 2435.540 20.840 ;
        RECT 2466.590 20.300 2466.910 20.360 ;
        RECT 2435.400 20.160 2466.910 20.300 ;
        RECT 2466.590 20.100 2466.910 20.160 ;
      LAYER via ;
        RECT 1993.280 3256.220 1993.540 3256.480 ;
        RECT 2644.180 3254.180 2644.440 3254.440 ;
        RECT 2614.740 282.920 2615.000 283.180 ;
        RECT 2644.180 282.920 2644.440 283.180 ;
        RECT 2466.620 243.820 2466.880 244.080 ;
        RECT 2614.740 243.820 2615.000 244.080 ;
        RECT 1780.760 20.440 1781.020 20.700 ;
        RECT 2466.620 20.100 2466.880 20.360 ;
      LAYER met2 ;
        RECT 1991.850 3256.930 1992.130 3260.000 ;
        RECT 1991.850 3256.790 1993.480 3256.930 ;
        RECT 1991.850 3256.000 1992.130 3256.790 ;
        RECT 1993.340 3256.510 1993.480 3256.790 ;
        RECT 1993.280 3256.190 1993.540 3256.510 ;
        RECT 2644.180 3254.150 2644.440 3254.470 ;
        RECT 2644.240 283.210 2644.380 3254.150 ;
        RECT 2614.740 282.890 2615.000 283.210 ;
        RECT 2644.180 282.890 2644.440 283.210 ;
        RECT 2614.800 244.110 2614.940 282.890 ;
        RECT 2466.620 243.790 2466.880 244.110 ;
        RECT 2614.740 243.790 2615.000 244.110 ;
        RECT 1780.760 20.410 1781.020 20.730 ;
        RECT 1780.820 2.400 1780.960 20.410 ;
        RECT 2466.680 20.390 2466.820 243.790 ;
        RECT 2466.620 20.070 2466.880 20.390 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 234.210 324.600 234.530 324.660 ;
        RECT 296.770 324.600 297.090 324.660 ;
        RECT 234.210 324.460 297.090 324.600 ;
        RECT 234.210 324.400 234.530 324.460 ;
        RECT 296.770 324.400 297.090 324.460 ;
        RECT 234.210 59.740 234.530 59.800 ;
        RECT 1798.670 59.740 1798.990 59.800 ;
        RECT 234.210 59.600 1798.990 59.740 ;
        RECT 234.210 59.540 234.530 59.600 ;
        RECT 1798.670 59.540 1798.990 59.600 ;
      LAYER via ;
        RECT 234.240 324.400 234.500 324.660 ;
        RECT 296.800 324.400 297.060 324.660 ;
        RECT 234.240 59.540 234.500 59.800 ;
        RECT 1798.700 59.540 1798.960 59.800 ;
      LAYER met2 ;
        RECT 296.790 326.555 297.070 326.925 ;
        RECT 296.860 324.690 297.000 326.555 ;
        RECT 234.240 324.370 234.500 324.690 ;
        RECT 296.800 324.370 297.060 324.690 ;
        RECT 234.300 59.830 234.440 324.370 ;
        RECT 234.240 59.510 234.500 59.830 ;
        RECT 1798.700 59.510 1798.960 59.830 ;
        RECT 1798.760 2.400 1798.900 59.510 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
      LAYER via2 ;
        RECT 296.790 326.600 297.070 326.880 ;
      LAYER met3 ;
        RECT 296.765 326.890 297.095 326.905 ;
        RECT 310.000 326.890 314.000 327.280 ;
        RECT 296.765 326.680 314.000 326.890 ;
        RECT 296.765 326.590 310.500 326.680 ;
        RECT 296.765 326.575 297.095 326.590 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1821.210 128.420 1821.530 128.480 ;
        RECT 1980.370 128.420 1980.690 128.480 ;
        RECT 1821.210 128.280 1980.690 128.420 ;
        RECT 1821.210 128.220 1821.530 128.280 ;
        RECT 1980.370 128.220 1980.690 128.280 ;
        RECT 1816.610 18.260 1816.930 18.320 ;
        RECT 1821.210 18.260 1821.530 18.320 ;
        RECT 1816.610 18.120 1821.530 18.260 ;
        RECT 1816.610 18.060 1816.930 18.120 ;
        RECT 1821.210 18.060 1821.530 18.120 ;
      LAYER via ;
        RECT 1821.240 128.220 1821.500 128.480 ;
        RECT 1980.400 128.220 1980.660 128.480 ;
        RECT 1816.640 18.060 1816.900 18.320 ;
        RECT 1821.240 18.060 1821.500 18.320 ;
      LAYER met2 ;
        RECT 1985.410 260.170 1985.690 264.000 ;
        RECT 1980.460 260.030 1985.690 260.170 ;
        RECT 1980.460 128.510 1980.600 260.030 ;
        RECT 1985.410 260.000 1985.690 260.030 ;
        RECT 1821.240 128.190 1821.500 128.510 ;
        RECT 1980.400 128.190 1980.660 128.510 ;
        RECT 1821.300 18.350 1821.440 128.190 ;
        RECT 1816.640 18.030 1816.900 18.350 ;
        RECT 1821.240 18.030 1821.500 18.350 ;
        RECT 1816.700 2.400 1816.840 18.030 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1172.610 190.300 1172.930 190.360 ;
        RECT 1828.570 190.300 1828.890 190.360 ;
        RECT 1172.610 190.160 1828.890 190.300 ;
        RECT 1172.610 190.100 1172.930 190.160 ;
        RECT 1828.570 190.100 1828.890 190.160 ;
        RECT 1828.570 37.640 1828.890 37.700 ;
        RECT 1834.550 37.640 1834.870 37.700 ;
        RECT 1828.570 37.500 1834.870 37.640 ;
        RECT 1828.570 37.440 1828.890 37.500 ;
        RECT 1834.550 37.440 1834.870 37.500 ;
      LAYER via ;
        RECT 1172.640 190.100 1172.900 190.360 ;
        RECT 1828.600 190.100 1828.860 190.360 ;
        RECT 1828.600 37.440 1828.860 37.700 ;
        RECT 1834.580 37.440 1834.840 37.700 ;
      LAYER met2 ;
        RECT 1170.290 260.170 1170.570 264.000 ;
        RECT 1170.290 260.030 1172.840 260.170 ;
        RECT 1170.290 260.000 1170.570 260.030 ;
        RECT 1172.700 190.390 1172.840 260.030 ;
        RECT 1172.640 190.070 1172.900 190.390 ;
        RECT 1828.600 190.070 1828.860 190.390 ;
        RECT 1828.660 37.730 1828.800 190.070 ;
        RECT 1828.600 37.410 1828.860 37.730 ;
        RECT 1834.580 37.410 1834.840 37.730 ;
        RECT 1834.640 2.400 1834.780 37.410 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 66.200 1856.030 66.260 ;
        RECT 2028.670 66.200 2028.990 66.260 ;
        RECT 1855.710 66.060 2028.990 66.200 ;
        RECT 1855.710 66.000 1856.030 66.060 ;
        RECT 2028.670 66.000 2028.990 66.060 ;
        RECT 1852.030 18.260 1852.350 18.320 ;
        RECT 1855.710 18.260 1856.030 18.320 ;
        RECT 1852.030 18.120 1856.030 18.260 ;
        RECT 1852.030 18.060 1852.350 18.120 ;
        RECT 1855.710 18.060 1856.030 18.120 ;
      LAYER via ;
        RECT 1855.740 66.000 1856.000 66.260 ;
        RECT 2028.700 66.000 2028.960 66.260 ;
        RECT 1852.060 18.060 1852.320 18.320 ;
        RECT 1855.740 18.060 1856.000 18.320 ;
      LAYER met2 ;
        RECT 2028.650 260.000 2028.930 264.000 ;
        RECT 2028.760 66.290 2028.900 260.000 ;
        RECT 1855.740 65.970 1856.000 66.290 ;
        RECT 2028.700 65.970 2028.960 66.290 ;
        RECT 1855.800 18.350 1855.940 65.970 ;
        RECT 1852.060 18.030 1852.320 18.350 ;
        RECT 1855.740 18.030 1856.000 18.350 ;
        RECT 1852.120 2.400 1852.260 18.030 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1875.950 93.740 1876.270 93.800 ;
        RECT 2256.370 93.740 2256.690 93.800 ;
        RECT 1875.950 93.600 2256.690 93.740 ;
        RECT 1875.950 93.540 1876.270 93.600 ;
        RECT 2256.370 93.540 2256.690 93.600 ;
        RECT 1869.970 18.260 1870.290 18.320 ;
        RECT 1875.950 18.260 1876.270 18.320 ;
        RECT 1869.970 18.120 1876.270 18.260 ;
        RECT 1869.970 18.060 1870.290 18.120 ;
        RECT 1875.950 18.060 1876.270 18.120 ;
      LAYER via ;
        RECT 1875.980 93.540 1876.240 93.800 ;
        RECT 2256.400 93.540 2256.660 93.800 ;
        RECT 1870.000 18.060 1870.260 18.320 ;
        RECT 1875.980 18.060 1876.240 18.320 ;
      LAYER met2 ;
        RECT 2256.810 260.170 2257.090 264.000 ;
        RECT 2256.460 260.030 2257.090 260.170 ;
        RECT 2256.460 93.830 2256.600 260.030 ;
        RECT 2256.810 260.000 2257.090 260.030 ;
        RECT 1875.980 93.510 1876.240 93.830 ;
        RECT 2256.400 93.510 2256.660 93.830 ;
        RECT 1876.040 18.350 1876.180 93.510 ;
        RECT 1870.000 18.030 1870.260 18.350 ;
        RECT 1875.980 18.030 1876.240 18.350 ;
        RECT 1870.060 2.400 1870.200 18.030 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1148.765 3253.885 1148.935 3255.415 ;
        RECT 745.345 57.205 745.515 88.655 ;
      LAYER mcon ;
        RECT 1148.765 3255.245 1148.935 3255.415 ;
        RECT 745.345 88.485 745.515 88.655 ;
      LAYER met1 ;
        RECT 1290.370 3256.420 1290.690 3256.480 ;
        RECT 1242.160 3256.280 1290.690 3256.420 ;
        RECT 1148.705 3255.400 1148.995 3255.445 ;
        RECT 1242.160 3255.400 1242.300 3256.280 ;
        RECT 1290.370 3256.220 1290.690 3256.280 ;
        RECT 1148.705 3255.260 1242.300 3255.400 ;
        RECT 1148.705 3255.215 1148.995 3255.260 ;
        RECT 1052.180 3254.240 1100.620 3254.380 ;
        RECT 239.270 3254.040 239.590 3254.100 ;
        RECT 1052.180 3254.040 1052.320 3254.240 ;
        RECT 239.270 3253.900 1052.320 3254.040 ;
        RECT 1100.480 3254.040 1100.620 3254.240 ;
        RECT 1148.705 3254.040 1148.995 3254.085 ;
        RECT 1100.480 3253.900 1148.995 3254.040 ;
        RECT 239.270 3253.840 239.590 3253.900 ;
        RECT 1148.705 3253.855 1148.995 3253.900 ;
        RECT 239.270 245.720 239.590 245.780 ;
        RECT 745.270 245.720 745.590 245.780 ;
        RECT 239.270 245.580 745.590 245.720 ;
        RECT 239.270 245.520 239.590 245.580 ;
        RECT 745.270 245.520 745.590 245.580 ;
        RECT 745.270 88.640 745.590 88.700 ;
        RECT 745.075 88.500 745.590 88.640 ;
        RECT 745.270 88.440 745.590 88.500 ;
        RECT 745.285 57.360 745.575 57.405 ;
        RECT 746.190 57.360 746.510 57.420 ;
        RECT 745.285 57.220 746.510 57.360 ;
        RECT 745.285 57.175 745.575 57.220 ;
        RECT 746.190 57.160 746.510 57.220 ;
      LAYER via ;
        RECT 1290.400 3256.220 1290.660 3256.480 ;
        RECT 239.300 3253.840 239.560 3254.100 ;
        RECT 239.300 245.520 239.560 245.780 ;
        RECT 745.300 245.520 745.560 245.780 ;
        RECT 745.300 88.440 745.560 88.700 ;
        RECT 746.220 57.160 746.480 57.420 ;
      LAYER met2 ;
        RECT 1291.730 3256.930 1292.010 3260.000 ;
        RECT 1290.460 3256.790 1292.010 3256.930 ;
        RECT 1290.460 3256.510 1290.600 3256.790 ;
        RECT 1290.400 3256.190 1290.660 3256.510 ;
        RECT 1291.730 3256.000 1292.010 3256.790 ;
        RECT 239.300 3253.810 239.560 3254.130 ;
        RECT 239.360 245.810 239.500 3253.810 ;
        RECT 239.300 245.490 239.560 245.810 ;
        RECT 745.300 245.490 745.560 245.810 ;
        RECT 745.360 88.730 745.500 245.490 ;
        RECT 745.300 88.410 745.560 88.730 ;
        RECT 746.220 57.130 746.480 57.450 ;
        RECT 746.280 2.400 746.420 57.130 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1883.845 48.365 1884.015 96.475 ;
      LAYER mcon ;
        RECT 1883.845 96.305 1884.015 96.475 ;
      LAYER met1 ;
        RECT 299.990 114.480 300.310 114.540 ;
        RECT 1883.770 114.480 1884.090 114.540 ;
        RECT 299.990 114.340 1884.090 114.480 ;
        RECT 299.990 114.280 300.310 114.340 ;
        RECT 1883.770 114.280 1884.090 114.340 ;
        RECT 1883.770 96.460 1884.090 96.520 ;
        RECT 1883.770 96.320 1884.285 96.460 ;
        RECT 1883.770 96.260 1884.090 96.320 ;
        RECT 1883.785 48.520 1884.075 48.565 ;
        RECT 1887.910 48.520 1888.230 48.580 ;
        RECT 1883.785 48.380 1888.230 48.520 ;
        RECT 1883.785 48.335 1884.075 48.380 ;
        RECT 1887.910 48.320 1888.230 48.380 ;
      LAYER via ;
        RECT 300.020 114.280 300.280 114.540 ;
        RECT 1883.800 114.280 1884.060 114.540 ;
        RECT 1883.800 96.260 1884.060 96.520 ;
        RECT 1887.940 48.320 1888.200 48.580 ;
      LAYER met2 ;
        RECT 300.010 368.715 300.290 369.085 ;
        RECT 300.080 114.570 300.220 368.715 ;
        RECT 300.020 114.250 300.280 114.570 ;
        RECT 1883.800 114.250 1884.060 114.570 ;
        RECT 1883.860 96.550 1884.000 114.250 ;
        RECT 1883.800 96.230 1884.060 96.550 ;
        RECT 1887.940 48.290 1888.200 48.610 ;
        RECT 1888.000 2.400 1888.140 48.290 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
      LAYER via2 ;
        RECT 300.010 368.760 300.290 369.040 ;
      LAYER met3 ;
        RECT 299.985 369.050 300.315 369.065 ;
        RECT 310.000 369.050 314.000 369.440 ;
        RECT 299.985 368.840 314.000 369.050 ;
        RECT 299.985 368.750 310.500 368.840 ;
        RECT 299.985 368.735 300.315 368.750 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1939.260 2615.490 1939.320 ;
        RECT 2680.030 1939.260 2680.350 1939.320 ;
        RECT 2615.170 1939.120 2680.350 1939.260 ;
        RECT 2615.170 1939.060 2615.490 1939.120 ;
        RECT 2680.030 1939.060 2680.350 1939.120 ;
        RECT 1910.910 245.720 1911.230 245.780 ;
        RECT 2680.030 245.720 2680.350 245.780 ;
        RECT 1910.910 245.580 2680.350 245.720 ;
        RECT 1910.910 245.520 1911.230 245.580 ;
        RECT 2680.030 245.520 2680.350 245.580 ;
        RECT 1905.850 15.200 1906.170 15.260 ;
        RECT 1910.910 15.200 1911.230 15.260 ;
        RECT 1905.850 15.060 1911.230 15.200 ;
        RECT 1905.850 15.000 1906.170 15.060 ;
        RECT 1910.910 15.000 1911.230 15.060 ;
      LAYER via ;
        RECT 2615.200 1939.060 2615.460 1939.320 ;
        RECT 2680.060 1939.060 2680.320 1939.320 ;
        RECT 1910.940 245.520 1911.200 245.780 ;
        RECT 2680.060 245.520 2680.320 245.780 ;
        RECT 1905.880 15.000 1906.140 15.260 ;
        RECT 1910.940 15.000 1911.200 15.260 ;
      LAYER met2 ;
        RECT 2615.190 1944.955 2615.470 1945.325 ;
        RECT 2615.260 1939.350 2615.400 1944.955 ;
        RECT 2615.200 1939.030 2615.460 1939.350 ;
        RECT 2680.060 1939.030 2680.320 1939.350 ;
        RECT 2680.120 245.810 2680.260 1939.030 ;
        RECT 1910.940 245.490 1911.200 245.810 ;
        RECT 2680.060 245.490 2680.320 245.810 ;
        RECT 1911.000 15.290 1911.140 245.490 ;
        RECT 1905.880 14.970 1906.140 15.290 ;
        RECT 1910.940 14.970 1911.200 15.290 ;
        RECT 1905.940 2.400 1906.080 14.970 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1945.000 2615.470 1945.280 ;
      LAYER met3 ;
        RECT 2606.000 1945.290 2610.000 1945.680 ;
        RECT 2615.165 1945.290 2615.495 1945.305 ;
        RECT 2606.000 1945.080 2615.495 1945.290 ;
        RECT 2609.580 1944.990 2615.495 1945.080 ;
        RECT 2615.165 1944.975 2615.495 1944.990 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 87.620 1925.030 87.680 ;
        RECT 2497.870 87.620 2498.190 87.680 ;
        RECT 1924.710 87.480 2498.190 87.620 ;
        RECT 1924.710 87.420 1925.030 87.480 ;
        RECT 2497.870 87.420 2498.190 87.480 ;
        RECT 1923.330 14.180 1923.650 14.240 ;
        RECT 1924.710 14.180 1925.030 14.240 ;
        RECT 1923.330 14.040 1925.030 14.180 ;
        RECT 1923.330 13.980 1923.650 14.040 ;
        RECT 1924.710 13.980 1925.030 14.040 ;
      LAYER via ;
        RECT 1924.740 87.420 1925.000 87.680 ;
        RECT 2497.900 87.420 2498.160 87.680 ;
        RECT 1923.360 13.980 1923.620 14.240 ;
        RECT 1924.740 13.980 1925.000 14.240 ;
      LAYER met2 ;
        RECT 2500.610 260.170 2500.890 264.000 ;
        RECT 2497.960 260.030 2500.890 260.170 ;
        RECT 2497.960 87.710 2498.100 260.030 ;
        RECT 2500.610 260.000 2500.890 260.030 ;
        RECT 1924.740 87.390 1925.000 87.710 ;
        RECT 2497.900 87.390 2498.160 87.710 ;
        RECT 1924.800 14.270 1924.940 87.390 ;
        RECT 1923.360 13.950 1923.620 14.270 ;
        RECT 1924.740 13.950 1925.000 14.270 ;
        RECT 1923.420 2.400 1923.560 13.950 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 697.240 2615.490 697.300 ;
        RECT 2660.710 697.240 2661.030 697.300 ;
        RECT 2615.170 697.100 2661.030 697.240 ;
        RECT 2615.170 697.040 2615.490 697.100 ;
        RECT 2660.710 697.040 2661.030 697.100 ;
        RECT 1945.410 227.020 1945.730 227.080 ;
        RECT 2660.710 227.020 2661.030 227.080 ;
        RECT 1945.410 226.880 2661.030 227.020 ;
        RECT 1945.410 226.820 1945.730 226.880 ;
        RECT 2660.710 226.820 2661.030 226.880 ;
        RECT 1941.270 16.900 1941.590 16.960 ;
        RECT 1945.410 16.900 1945.730 16.960 ;
        RECT 1941.270 16.760 1945.730 16.900 ;
        RECT 1941.270 16.700 1941.590 16.760 ;
        RECT 1945.410 16.700 1945.730 16.760 ;
      LAYER via ;
        RECT 2615.200 697.040 2615.460 697.300 ;
        RECT 2660.740 697.040 2661.000 697.300 ;
        RECT 1945.440 226.820 1945.700 227.080 ;
        RECT 2660.740 226.820 2661.000 227.080 ;
        RECT 1941.300 16.700 1941.560 16.960 ;
        RECT 1945.440 16.700 1945.700 16.960 ;
      LAYER met2 ;
        RECT 2615.190 697.835 2615.470 698.205 ;
        RECT 2615.260 697.330 2615.400 697.835 ;
        RECT 2615.200 697.010 2615.460 697.330 ;
        RECT 2660.740 697.010 2661.000 697.330 ;
        RECT 2660.800 227.110 2660.940 697.010 ;
        RECT 1945.440 226.790 1945.700 227.110 ;
        RECT 2660.740 226.790 2661.000 227.110 ;
        RECT 1945.500 16.990 1945.640 226.790 ;
        RECT 1941.300 16.670 1941.560 16.990 ;
        RECT 1945.440 16.670 1945.700 16.990 ;
        RECT 1941.360 2.400 1941.500 16.670 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
      LAYER via2 ;
        RECT 2615.190 697.880 2615.470 698.160 ;
      LAYER met3 ;
        RECT 2606.000 698.170 2610.000 698.560 ;
        RECT 2615.165 698.170 2615.495 698.185 ;
        RECT 2606.000 697.960 2615.495 698.170 ;
        RECT 2609.580 697.870 2615.495 697.960 ;
        RECT 2615.165 697.855 2615.495 697.870 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1959.210 259.660 1959.530 259.720 ;
        RECT 2616.090 259.660 2616.410 259.720 ;
        RECT 1959.210 259.520 2616.410 259.660 ;
        RECT 1959.210 259.460 1959.530 259.520 ;
        RECT 2616.090 259.460 2616.410 259.520 ;
      LAYER via ;
        RECT 1959.240 259.460 1959.500 259.720 ;
        RECT 2616.120 259.460 2616.380 259.720 ;
      LAYER met2 ;
        RECT 2616.110 338.795 2616.390 339.165 ;
        RECT 2616.180 259.750 2616.320 338.795 ;
        RECT 1959.240 259.430 1959.500 259.750 ;
        RECT 2616.120 259.430 2616.380 259.750 ;
        RECT 1959.300 2.400 1959.440 259.430 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
      LAYER via2 ;
        RECT 2616.110 338.840 2616.390 339.120 ;
      LAYER met3 ;
        RECT 2606.000 339.130 2610.000 339.520 ;
        RECT 2616.085 339.130 2616.415 339.145 ;
        RECT 2606.000 338.920 2616.415 339.130 ;
        RECT 2609.580 338.830 2616.415 338.920 ;
        RECT 2616.085 338.815 2616.415 338.830 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1973.545 48.365 1973.715 96.475 ;
      LAYER mcon ;
        RECT 1973.545 96.305 1973.715 96.475 ;
      LAYER met1 ;
        RECT 1973.470 96.460 1973.790 96.520 ;
        RECT 1973.275 96.320 1973.790 96.460 ;
        RECT 1973.470 96.260 1973.790 96.320 ;
        RECT 1973.485 48.520 1973.775 48.565 ;
        RECT 1977.150 48.520 1977.470 48.580 ;
        RECT 1973.485 48.380 1977.470 48.520 ;
        RECT 1973.485 48.335 1973.775 48.380 ;
        RECT 1977.150 48.320 1977.470 48.380 ;
      LAYER via ;
        RECT 1973.500 96.260 1973.760 96.520 ;
        RECT 1977.180 48.320 1977.440 48.580 ;
      LAYER met2 ;
        RECT 919.170 3271.635 919.450 3272.005 ;
        RECT 2529.170 3271.635 2529.450 3272.005 ;
        RECT 919.240 3260.000 919.380 3271.635 ;
        RECT 2529.240 3267.245 2529.380 3271.635 ;
        RECT 2529.170 3266.875 2529.450 3267.245 ;
        RECT 2613.350 3266.875 2613.630 3267.245 ;
        RECT 919.130 3256.000 919.410 3260.000 ;
        RECT 2613.420 376.565 2613.560 3266.875 ;
        RECT 2613.350 376.195 2613.630 376.565 ;
        RECT 1973.490 263.315 1973.770 263.685 ;
        RECT 1973.560 96.550 1973.700 263.315 ;
        RECT 1973.500 96.230 1973.760 96.550 ;
        RECT 1977.180 48.290 1977.440 48.610 ;
        RECT 1977.240 2.400 1977.380 48.290 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
      LAYER via2 ;
        RECT 919.170 3271.680 919.450 3271.960 ;
        RECT 2529.170 3271.680 2529.450 3271.960 ;
        RECT 2529.170 3266.920 2529.450 3267.200 ;
        RECT 2613.350 3266.920 2613.630 3267.200 ;
        RECT 2613.350 376.240 2613.630 376.520 ;
        RECT 1973.490 263.360 1973.770 263.640 ;
      LAYER met3 ;
        RECT 919.145 3271.970 919.475 3271.985 ;
        RECT 2529.145 3271.970 2529.475 3271.985 ;
        RECT 919.145 3271.670 2529.475 3271.970 ;
        RECT 919.145 3271.655 919.475 3271.670 ;
        RECT 2529.145 3271.655 2529.475 3271.670 ;
        RECT 2529.145 3267.210 2529.475 3267.225 ;
        RECT 2613.325 3267.210 2613.655 3267.225 ;
        RECT 2529.145 3266.910 2613.655 3267.210 ;
        RECT 2529.145 3266.895 2529.475 3266.910 ;
        RECT 2613.325 3266.895 2613.655 3266.910 ;
        RECT 2611.230 376.530 2611.610 376.540 ;
        RECT 2613.325 376.530 2613.655 376.545 ;
        RECT 2611.230 376.230 2613.655 376.530 ;
        RECT 2611.230 376.220 2611.610 376.230 ;
        RECT 2613.325 376.215 2613.655 376.230 ;
        RECT 1973.465 263.650 1973.795 263.665 ;
        RECT 2611.230 263.650 2611.610 263.660 ;
        RECT 1973.465 263.350 2611.610 263.650 ;
        RECT 1973.465 263.335 1973.795 263.350 ;
        RECT 2611.230 263.340 2611.610 263.350 ;
      LAYER via3 ;
        RECT 2611.260 376.220 2611.580 376.540 ;
        RECT 2611.260 263.340 2611.580 263.660 ;
      LAYER met4 ;
        RECT 2611.255 376.215 2611.585 376.545 ;
        RECT 2611.270 263.665 2611.570 376.215 ;
        RECT 2611.255 263.335 2611.585 263.665 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2463.830 3275.460 2464.150 3275.520 ;
        RECT 2636.790 3275.460 2637.110 3275.520 ;
        RECT 2463.830 3275.320 2637.110 3275.460 ;
        RECT 2463.830 3275.260 2464.150 3275.320 ;
        RECT 2636.790 3275.260 2637.110 3275.320 ;
        RECT 2000.610 239.940 2000.930 240.000 ;
        RECT 2636.790 239.940 2637.110 240.000 ;
        RECT 2000.610 239.800 2637.110 239.940 ;
        RECT 2000.610 239.740 2000.930 239.800 ;
        RECT 2636.790 239.740 2637.110 239.800 ;
        RECT 1995.090 16.900 1995.410 16.960 ;
        RECT 2000.610 16.900 2000.930 16.960 ;
        RECT 1995.090 16.760 2000.930 16.900 ;
        RECT 1995.090 16.700 1995.410 16.760 ;
        RECT 2000.610 16.700 2000.930 16.760 ;
      LAYER via ;
        RECT 2463.860 3275.260 2464.120 3275.520 ;
        RECT 2636.820 3275.260 2637.080 3275.520 ;
        RECT 2000.640 239.740 2000.900 240.000 ;
        RECT 2636.820 239.740 2637.080 240.000 ;
        RECT 1995.120 16.700 1995.380 16.960 ;
        RECT 2000.640 16.700 2000.900 16.960 ;
      LAYER met2 ;
        RECT 2463.860 3275.230 2464.120 3275.550 ;
        RECT 2636.820 3275.230 2637.080 3275.550 ;
        RECT 2463.920 3260.000 2464.060 3275.230 ;
        RECT 2463.810 3256.000 2464.090 3260.000 ;
        RECT 2636.880 240.030 2637.020 3275.230 ;
        RECT 2000.640 239.710 2000.900 240.030 ;
        RECT 2636.820 239.710 2637.080 240.030 ;
        RECT 2000.700 16.990 2000.840 239.710 ;
        RECT 1995.120 16.670 1995.380 16.990 ;
        RECT 2000.640 16.670 2000.900 16.990 ;
        RECT 1995.180 2.400 1995.320 16.670 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1372.250 121.960 1372.570 122.020 ;
        RECT 2007.970 121.960 2008.290 122.020 ;
        RECT 1372.250 121.820 2008.290 121.960 ;
        RECT 1372.250 121.760 1372.570 121.820 ;
        RECT 2007.970 121.760 2008.290 121.820 ;
        RECT 2007.970 14.180 2008.290 14.240 ;
        RECT 2007.970 14.040 2012.800 14.180 ;
        RECT 2007.970 13.980 2008.290 14.040 ;
        RECT 2012.660 13.900 2012.800 14.040 ;
        RECT 2012.570 13.640 2012.890 13.900 ;
      LAYER via ;
        RECT 1372.280 121.760 1372.540 122.020 ;
        RECT 2008.000 121.760 2008.260 122.020 ;
        RECT 2008.000 13.980 2008.260 14.240 ;
        RECT 2012.600 13.640 2012.860 13.900 ;
      LAYER met2 ;
        RECT 1370.850 260.170 1371.130 264.000 ;
        RECT 1370.850 260.030 1372.480 260.170 ;
        RECT 1370.850 260.000 1371.130 260.030 ;
        RECT 1372.340 122.050 1372.480 260.030 ;
        RECT 1372.280 121.730 1372.540 122.050 ;
        RECT 2008.000 121.730 2008.260 122.050 ;
        RECT 2008.060 14.270 2008.200 121.730 ;
        RECT 2008.000 13.950 2008.260 14.270 ;
        RECT 2012.600 13.610 2012.860 13.930 ;
        RECT 2012.660 2.400 2012.800 13.610 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2035.110 66.200 2035.430 66.260 ;
        RECT 2352.970 66.200 2353.290 66.260 ;
        RECT 2035.110 66.060 2353.290 66.200 ;
        RECT 2035.110 66.000 2035.430 66.060 ;
        RECT 2352.970 66.000 2353.290 66.060 ;
        RECT 2030.510 16.900 2030.830 16.960 ;
        RECT 2035.110 16.900 2035.430 16.960 ;
        RECT 2030.510 16.760 2035.430 16.900 ;
        RECT 2030.510 16.700 2030.830 16.760 ;
        RECT 2035.110 16.700 2035.430 16.760 ;
      LAYER via ;
        RECT 2035.140 66.000 2035.400 66.260 ;
        RECT 2353.000 66.000 2353.260 66.260 ;
        RECT 2030.540 16.700 2030.800 16.960 ;
        RECT 2035.140 16.700 2035.400 16.960 ;
      LAYER met2 ;
        RECT 2357.090 260.170 2357.370 264.000 ;
        RECT 2353.060 260.030 2357.370 260.170 ;
        RECT 2353.060 66.290 2353.200 260.030 ;
        RECT 2357.090 260.000 2357.370 260.030 ;
        RECT 2035.140 65.970 2035.400 66.290 ;
        RECT 2353.000 65.970 2353.260 66.290 ;
        RECT 2035.200 16.990 2035.340 65.970 ;
        RECT 2030.540 16.670 2030.800 16.990 ;
        RECT 2035.140 16.670 2035.400 16.990 ;
        RECT 2030.600 2.400 2030.740 16.670 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.610 100.540 413.930 100.600 ;
        RECT 2042.470 100.540 2042.790 100.600 ;
        RECT 413.610 100.400 2042.790 100.540 ;
        RECT 413.610 100.340 413.930 100.400 ;
        RECT 2042.470 100.340 2042.790 100.400 ;
        RECT 2042.470 37.640 2042.790 37.700 ;
        RECT 2048.450 37.640 2048.770 37.700 ;
        RECT 2042.470 37.500 2048.770 37.640 ;
        RECT 2042.470 37.440 2042.790 37.500 ;
        RECT 2048.450 37.440 2048.770 37.500 ;
      LAYER via ;
        RECT 413.640 100.340 413.900 100.600 ;
        RECT 2042.500 100.340 2042.760 100.600 ;
        RECT 2042.500 37.440 2042.760 37.700 ;
        RECT 2048.480 37.440 2048.740 37.700 ;
      LAYER met2 ;
        RECT 412.210 260.170 412.490 264.000 ;
        RECT 412.210 260.030 413.840 260.170 ;
        RECT 412.210 260.000 412.490 260.030 ;
        RECT 413.700 100.630 413.840 260.030 ;
        RECT 413.640 100.310 413.900 100.630 ;
        RECT 2042.500 100.310 2042.760 100.630 ;
        RECT 2042.560 37.730 2042.700 100.310 ;
        RECT 2042.500 37.410 2042.760 37.730 ;
        RECT 2048.480 37.410 2048.740 37.730 ;
        RECT 2048.540 2.400 2048.680 37.410 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.710 1263.000 2615.030 1263.060 ;
        RECT 2688.310 1263.000 2688.630 1263.060 ;
        RECT 2614.710 1262.860 2688.630 1263.000 ;
        RECT 2614.710 1262.800 2615.030 1262.860 ;
        RECT 2688.310 1262.800 2688.630 1262.860 ;
        RECT 765.510 231.440 765.830 231.500 ;
        RECT 2688.310 231.440 2688.630 231.500 ;
        RECT 765.510 231.300 2688.630 231.440 ;
        RECT 765.510 231.240 765.830 231.300 ;
        RECT 2688.310 231.240 2688.630 231.300 ;
      LAYER via ;
        RECT 2614.740 1262.800 2615.000 1263.060 ;
        RECT 2688.340 1262.800 2688.600 1263.060 ;
        RECT 765.540 231.240 765.800 231.500 ;
        RECT 2688.340 231.240 2688.600 231.500 ;
      LAYER met2 ;
        RECT 2614.730 1267.675 2615.010 1268.045 ;
        RECT 2614.800 1263.090 2614.940 1267.675 ;
        RECT 2614.740 1262.770 2615.000 1263.090 ;
        RECT 2688.340 1262.770 2688.600 1263.090 ;
        RECT 2688.400 231.530 2688.540 1262.770 ;
        RECT 765.540 231.210 765.800 231.530 ;
        RECT 2688.340 231.210 2688.600 231.530 ;
        RECT 765.600 12.650 765.740 231.210 ;
        RECT 763.760 12.510 765.740 12.650 ;
        RECT 763.760 2.400 763.900 12.510 ;
        RECT 763.550 -4.800 764.110 2.400 ;
      LAYER via2 ;
        RECT 2614.730 1267.720 2615.010 1268.000 ;
      LAYER met3 ;
        RECT 2606.000 1268.010 2610.000 1268.400 ;
        RECT 2614.705 1268.010 2615.035 1268.025 ;
        RECT 2606.000 1267.800 2615.035 1268.010 ;
        RECT 2609.580 1267.710 2615.035 1267.800 ;
        RECT 2614.705 1267.695 2615.035 1267.710 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 300.910 231.780 301.230 231.840 ;
        RECT 2063.170 231.780 2063.490 231.840 ;
        RECT 300.910 231.640 2063.490 231.780 ;
        RECT 300.910 231.580 301.230 231.640 ;
        RECT 2063.170 231.580 2063.490 231.640 ;
        RECT 2063.170 62.120 2063.490 62.180 ;
        RECT 2066.390 62.120 2066.710 62.180 ;
        RECT 2063.170 61.980 2066.710 62.120 ;
        RECT 2063.170 61.920 2063.490 61.980 ;
        RECT 2066.390 61.920 2066.710 61.980 ;
      LAYER via ;
        RECT 300.940 231.580 301.200 231.840 ;
        RECT 2063.200 231.580 2063.460 231.840 ;
        RECT 2063.200 61.920 2063.460 62.180 ;
        RECT 2066.420 61.920 2066.680 62.180 ;
      LAYER met2 ;
        RECT 300.930 623.035 301.210 623.405 ;
        RECT 301.000 231.870 301.140 623.035 ;
        RECT 300.940 231.550 301.200 231.870 ;
        RECT 2063.200 231.550 2063.460 231.870 ;
        RECT 2063.260 62.210 2063.400 231.550 ;
        RECT 2063.200 61.890 2063.460 62.210 ;
        RECT 2066.420 61.890 2066.680 62.210 ;
        RECT 2066.480 2.400 2066.620 61.890 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
      LAYER via2 ;
        RECT 300.930 623.080 301.210 623.360 ;
      LAYER met3 ;
        RECT 300.905 623.370 301.235 623.385 ;
        RECT 310.000 623.370 314.000 623.760 ;
        RECT 300.905 623.160 314.000 623.370 ;
        RECT 300.905 623.070 310.500 623.160 ;
        RECT 300.905 623.055 301.235 623.070 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 87.280 1159.130 87.340 ;
        RECT 2083.870 87.280 2084.190 87.340 ;
        RECT 1158.810 87.140 2084.190 87.280 ;
        RECT 1158.810 87.080 1159.130 87.140 ;
        RECT 2083.870 87.080 2084.190 87.140 ;
      LAYER via ;
        RECT 1158.840 87.080 1159.100 87.340 ;
        RECT 2083.900 87.080 2084.160 87.340 ;
      LAYER met2 ;
        RECT 1156.490 260.170 1156.770 264.000 ;
        RECT 1156.490 260.030 1159.040 260.170 ;
        RECT 1156.490 260.000 1156.770 260.030 ;
        RECT 1158.900 87.370 1159.040 260.030 ;
        RECT 1158.840 87.050 1159.100 87.370 ;
        RECT 2083.900 87.050 2084.160 87.370 ;
        RECT 2083.960 37.810 2084.100 87.050 ;
        RECT 2083.960 37.670 2084.560 37.810 ;
        RECT 2084.420 2.400 2084.560 37.670 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1885.150 244.360 1885.470 244.420 ;
        RECT 1890.210 244.360 1890.530 244.420 ;
        RECT 1885.150 244.220 1890.530 244.360 ;
        RECT 1885.150 244.160 1885.470 244.220 ;
        RECT 1890.210 244.160 1890.530 244.220 ;
        RECT 1890.210 114.480 1890.530 114.540 ;
        RECT 2097.670 114.480 2097.990 114.540 ;
        RECT 1890.210 114.340 2097.990 114.480 ;
        RECT 1890.210 114.280 1890.530 114.340 ;
        RECT 2097.670 114.280 2097.990 114.340 ;
        RECT 2097.670 62.120 2097.990 62.180 ;
        RECT 2101.810 62.120 2102.130 62.180 ;
        RECT 2097.670 61.980 2102.130 62.120 ;
        RECT 2097.670 61.920 2097.990 61.980 ;
        RECT 2101.810 61.920 2102.130 61.980 ;
      LAYER via ;
        RECT 1885.180 244.160 1885.440 244.420 ;
        RECT 1890.240 244.160 1890.500 244.420 ;
        RECT 1890.240 114.280 1890.500 114.540 ;
        RECT 2097.700 114.280 2097.960 114.540 ;
        RECT 2097.700 61.920 2097.960 62.180 ;
        RECT 2101.840 61.920 2102.100 62.180 ;
      LAYER met2 ;
        RECT 1885.130 260.000 1885.410 264.000 ;
        RECT 1885.240 244.450 1885.380 260.000 ;
        RECT 1885.180 244.130 1885.440 244.450 ;
        RECT 1890.240 244.130 1890.500 244.450 ;
        RECT 1890.300 114.570 1890.440 244.130 ;
        RECT 1890.240 114.250 1890.500 114.570 ;
        RECT 2097.700 114.250 2097.960 114.570 ;
        RECT 2097.760 62.210 2097.900 114.250 ;
        RECT 2097.700 61.890 2097.960 62.210 ;
        RECT 2101.840 61.890 2102.100 62.210 ;
        RECT 2101.900 2.400 2102.040 61.890 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2118.445 186.405 2118.615 193.715 ;
      LAYER mcon ;
        RECT 2118.445 193.545 2118.615 193.715 ;
      LAYER met1 ;
        RECT 2078.810 3256.220 2079.130 3256.480 ;
        RECT 2078.900 3254.720 2079.040 3256.220 ;
        RECT 2612.410 3254.720 2612.730 3254.780 ;
        RECT 2078.900 3254.580 2612.730 3254.720 ;
        RECT 2612.410 3254.520 2612.730 3254.580 ;
        RECT 2612.410 635.360 2612.730 635.420 ;
        RECT 2619.310 635.360 2619.630 635.420 ;
        RECT 2612.410 635.220 2619.630 635.360 ;
        RECT 2612.410 635.160 2612.730 635.220 ;
        RECT 2619.310 635.160 2619.630 635.220 ;
        RECT 2619.310 346.020 2619.630 346.080 ;
        RECT 2619.310 345.880 2637.940 346.020 ;
        RECT 2619.310 345.820 2619.630 345.880 ;
        RECT 2637.250 344.660 2637.570 344.720 ;
        RECT 2637.800 344.660 2637.940 345.880 ;
        RECT 2637.250 344.520 2637.940 344.660 ;
        RECT 2637.250 344.460 2637.570 344.520 ;
        RECT 2118.370 263.740 2118.690 263.800 ;
        RECT 2637.250 263.740 2637.570 263.800 ;
        RECT 2118.370 263.600 2637.570 263.740 ;
        RECT 2118.370 263.540 2118.690 263.600 ;
        RECT 2637.250 263.540 2637.570 263.600 ;
        RECT 2118.370 193.700 2118.690 193.760 ;
        RECT 2118.370 193.560 2118.885 193.700 ;
        RECT 2118.370 193.500 2118.690 193.560 ;
        RECT 2118.370 186.560 2118.690 186.620 ;
        RECT 2118.370 186.420 2118.885 186.560 ;
        RECT 2118.370 186.360 2118.690 186.420 ;
        RECT 2118.370 137.940 2118.690 138.000 ;
        RECT 2118.830 137.940 2119.150 138.000 ;
        RECT 2118.370 137.800 2119.150 137.940 ;
        RECT 2118.370 137.740 2118.690 137.800 ;
        RECT 2118.830 137.740 2119.150 137.800 ;
        RECT 2119.750 47.980 2120.070 48.240 ;
        RECT 2119.840 47.560 2119.980 47.980 ;
        RECT 2119.750 47.300 2120.070 47.560 ;
      LAYER via ;
        RECT 2078.840 3256.220 2079.100 3256.480 ;
        RECT 2612.440 3254.520 2612.700 3254.780 ;
        RECT 2612.440 635.160 2612.700 635.420 ;
        RECT 2619.340 635.160 2619.600 635.420 ;
        RECT 2619.340 345.820 2619.600 346.080 ;
        RECT 2637.280 344.460 2637.540 344.720 ;
        RECT 2118.400 263.540 2118.660 263.800 ;
        RECT 2637.280 263.540 2637.540 263.800 ;
        RECT 2118.400 193.500 2118.660 193.760 ;
        RECT 2118.400 186.360 2118.660 186.620 ;
        RECT 2118.400 137.740 2118.660 138.000 ;
        RECT 2118.860 137.740 2119.120 138.000 ;
        RECT 2119.780 47.980 2120.040 48.240 ;
        RECT 2119.780 47.300 2120.040 47.560 ;
      LAYER met2 ;
        RECT 2077.410 3256.930 2077.690 3260.000 ;
        RECT 2077.410 3256.790 2079.040 3256.930 ;
        RECT 2077.410 3256.000 2077.690 3256.790 ;
        RECT 2078.900 3256.510 2079.040 3256.790 ;
        RECT 2078.840 3256.190 2079.100 3256.510 ;
        RECT 2612.440 3254.490 2612.700 3254.810 ;
        RECT 2612.500 635.450 2612.640 3254.490 ;
        RECT 2612.440 635.130 2612.700 635.450 ;
        RECT 2619.340 635.130 2619.600 635.450 ;
        RECT 2619.400 346.110 2619.540 635.130 ;
        RECT 2619.340 345.790 2619.600 346.110 ;
        RECT 2637.280 344.430 2637.540 344.750 ;
        RECT 2637.340 263.830 2637.480 344.430 ;
        RECT 2118.400 263.510 2118.660 263.830 ;
        RECT 2637.280 263.510 2637.540 263.830 ;
        RECT 2118.460 193.790 2118.600 263.510 ;
        RECT 2118.400 193.470 2118.660 193.790 ;
        RECT 2118.400 186.330 2118.660 186.650 ;
        RECT 2118.460 138.030 2118.600 186.330 ;
        RECT 2118.400 137.710 2118.660 138.030 ;
        RECT 2118.860 137.710 2119.120 138.030 ;
        RECT 2118.920 48.805 2119.060 137.710 ;
        RECT 2118.850 48.435 2119.130 48.805 ;
        RECT 2119.770 48.435 2120.050 48.805 ;
        RECT 2119.840 48.270 2119.980 48.435 ;
        RECT 2119.780 47.950 2120.040 48.270 ;
        RECT 2119.780 47.270 2120.040 47.590 ;
        RECT 2119.840 2.400 2119.980 47.270 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
      LAYER via2 ;
        RECT 2118.850 48.480 2119.130 48.760 ;
        RECT 2119.770 48.480 2120.050 48.760 ;
      LAYER met3 ;
        RECT 2118.825 48.770 2119.155 48.785 ;
        RECT 2119.745 48.770 2120.075 48.785 ;
        RECT 2118.825 48.470 2120.075 48.770 ;
        RECT 2118.825 48.455 2119.155 48.470 ;
        RECT 2119.745 48.455 2120.075 48.470 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 237.430 1614.900 237.750 1614.960 ;
        RECT 296.770 1614.900 297.090 1614.960 ;
        RECT 237.430 1614.760 297.090 1614.900 ;
        RECT 237.430 1614.700 237.750 1614.760 ;
        RECT 296.770 1614.700 297.090 1614.760 ;
        RECT 237.430 59.400 237.750 59.460 ;
        RECT 2137.690 59.400 2138.010 59.460 ;
        RECT 237.430 59.260 2138.010 59.400 ;
        RECT 237.430 59.200 237.750 59.260 ;
        RECT 2137.690 59.200 2138.010 59.260 ;
      LAYER via ;
        RECT 237.460 1614.700 237.720 1614.960 ;
        RECT 296.800 1614.700 297.060 1614.960 ;
        RECT 237.460 59.200 237.720 59.460 ;
        RECT 2137.720 59.200 2137.980 59.460 ;
      LAYER met2 ;
        RECT 296.790 1615.835 297.070 1616.205 ;
        RECT 296.860 1614.990 297.000 1615.835 ;
        RECT 237.460 1614.670 237.720 1614.990 ;
        RECT 296.800 1614.670 297.060 1614.990 ;
        RECT 237.520 59.490 237.660 1614.670 ;
        RECT 237.460 59.170 237.720 59.490 ;
        RECT 2137.720 59.170 2137.980 59.490 ;
        RECT 2137.780 2.400 2137.920 59.170 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
      LAYER via2 ;
        RECT 296.790 1615.880 297.070 1616.160 ;
      LAYER met3 ;
        RECT 296.765 1616.170 297.095 1616.185 ;
        RECT 310.000 1616.170 314.000 1616.560 ;
        RECT 296.765 1615.960 314.000 1616.170 ;
        RECT 296.765 1615.870 310.500 1615.960 ;
        RECT 296.765 1615.855 297.095 1615.870 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2001.140 2615.490 2001.200 ;
        RECT 2692.910 2001.140 2693.230 2001.200 ;
        RECT 2615.170 2001.000 2693.230 2001.140 ;
        RECT 2615.170 2000.940 2615.490 2001.000 ;
        RECT 2692.910 2000.940 2693.230 2001.000 ;
        RECT 2159.310 251.160 2159.630 251.220 ;
        RECT 2692.910 251.160 2693.230 251.220 ;
        RECT 2159.310 251.020 2693.230 251.160 ;
        RECT 2159.310 250.960 2159.630 251.020 ;
        RECT 2692.910 250.960 2693.230 251.020 ;
        RECT 2155.630 18.940 2155.950 19.000 ;
        RECT 2159.310 18.940 2159.630 19.000 ;
        RECT 2155.630 18.800 2159.630 18.940 ;
        RECT 2155.630 18.740 2155.950 18.800 ;
        RECT 2159.310 18.740 2159.630 18.800 ;
      LAYER via ;
        RECT 2615.200 2000.940 2615.460 2001.200 ;
        RECT 2692.940 2000.940 2693.200 2001.200 ;
        RECT 2159.340 250.960 2159.600 251.220 ;
        RECT 2692.940 250.960 2693.200 251.220 ;
        RECT 2155.660 18.740 2155.920 19.000 ;
        RECT 2159.340 18.740 2159.600 19.000 ;
      LAYER met2 ;
        RECT 2615.190 2007.515 2615.470 2007.885 ;
        RECT 2615.260 2001.230 2615.400 2007.515 ;
        RECT 2615.200 2000.910 2615.460 2001.230 ;
        RECT 2692.940 2000.910 2693.200 2001.230 ;
        RECT 2693.000 251.250 2693.140 2000.910 ;
        RECT 2159.340 250.930 2159.600 251.250 ;
        RECT 2692.940 250.930 2693.200 251.250 ;
        RECT 2159.400 19.030 2159.540 250.930 ;
        RECT 2155.660 18.710 2155.920 19.030 ;
        RECT 2159.340 18.710 2159.600 19.030 ;
        RECT 2155.720 2.400 2155.860 18.710 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2007.560 2615.470 2007.840 ;
      LAYER met3 ;
        RECT 2606.000 2007.850 2610.000 2008.240 ;
        RECT 2615.165 2007.850 2615.495 2007.865 ;
        RECT 2606.000 2007.640 2615.495 2007.850 ;
        RECT 2609.580 2007.550 2615.495 2007.640 ;
        RECT 2615.165 2007.535 2615.495 2007.550 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1913.670 211.720 1913.990 211.780 ;
        RECT 2166.670 211.720 2166.990 211.780 ;
        RECT 1913.670 211.580 2166.990 211.720 ;
        RECT 1913.670 211.520 1913.990 211.580 ;
        RECT 2166.670 211.520 2166.990 211.580 ;
        RECT 2166.670 37.640 2166.990 37.700 ;
        RECT 2173.110 37.640 2173.430 37.700 ;
        RECT 2166.670 37.500 2173.430 37.640 ;
        RECT 2166.670 37.440 2166.990 37.500 ;
        RECT 2173.110 37.440 2173.430 37.500 ;
      LAYER via ;
        RECT 1913.700 211.520 1913.960 211.780 ;
        RECT 2166.700 211.520 2166.960 211.780 ;
        RECT 2166.700 37.440 2166.960 37.700 ;
        RECT 2173.140 37.440 2173.400 37.700 ;
      LAYER met2 ;
        RECT 1913.650 260.000 1913.930 264.000 ;
        RECT 1913.760 211.810 1913.900 260.000 ;
        RECT 1913.700 211.490 1913.960 211.810 ;
        RECT 2166.700 211.490 2166.960 211.810 ;
        RECT 2166.760 37.730 2166.900 211.490 ;
        RECT 2166.700 37.410 2166.960 37.730 ;
        RECT 2173.140 37.410 2173.400 37.730 ;
        RECT 2173.200 2.400 2173.340 37.410 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 231.450 2332.300 231.770 2332.360 ;
        RECT 296.770 2332.300 297.090 2332.360 ;
        RECT 231.450 2332.160 297.090 2332.300 ;
        RECT 231.450 2332.100 231.770 2332.160 ;
        RECT 296.770 2332.100 297.090 2332.160 ;
        RECT 231.450 32.540 231.770 32.600 ;
        RECT 2191.050 32.540 2191.370 32.600 ;
        RECT 231.450 32.400 2191.370 32.540 ;
        RECT 231.450 32.340 231.770 32.400 ;
        RECT 2191.050 32.340 2191.370 32.400 ;
      LAYER via ;
        RECT 231.480 2332.100 231.740 2332.360 ;
        RECT 296.800 2332.100 297.060 2332.360 ;
        RECT 231.480 32.340 231.740 32.600 ;
        RECT 2191.080 32.340 2191.340 32.600 ;
      LAYER met2 ;
        RECT 296.790 2335.275 297.070 2335.645 ;
        RECT 296.860 2332.390 297.000 2335.275 ;
        RECT 231.480 2332.070 231.740 2332.390 ;
        RECT 296.800 2332.070 297.060 2332.390 ;
        RECT 231.540 32.630 231.680 2332.070 ;
        RECT 231.480 32.310 231.740 32.630 ;
        RECT 2191.080 32.310 2191.340 32.630 ;
        RECT 2191.140 2.400 2191.280 32.310 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
      LAYER via2 ;
        RECT 296.790 2335.320 297.070 2335.600 ;
      LAYER met3 ;
        RECT 296.765 2335.610 297.095 2335.625 ;
        RECT 310.000 2335.610 314.000 2336.000 ;
        RECT 296.765 2335.400 314.000 2335.610 ;
        RECT 296.765 2335.310 310.500 2335.400 ;
        RECT 296.765 2335.295 297.095 2335.310 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2209.065 2.805 2209.235 48.195 ;
      LAYER mcon ;
        RECT 2209.065 48.025 2209.235 48.195 ;
      LAYER met1 ;
        RECT 2099.510 244.020 2099.830 244.080 ;
        RECT 2104.110 244.020 2104.430 244.080 ;
        RECT 2099.510 243.880 2104.430 244.020 ;
        RECT 2099.510 243.820 2099.830 243.880 ;
        RECT 2104.110 243.820 2104.430 243.880 ;
        RECT 2104.110 114.480 2104.430 114.540 ;
        RECT 2208.070 114.480 2208.390 114.540 ;
        RECT 2104.110 114.340 2208.390 114.480 ;
        RECT 2104.110 114.280 2104.430 114.340 ;
        RECT 2208.070 114.280 2208.390 114.340 ;
        RECT 2207.610 96.460 2207.930 96.520 ;
        RECT 2208.070 96.460 2208.390 96.520 ;
        RECT 2207.610 96.320 2208.390 96.460 ;
        RECT 2207.610 96.260 2207.930 96.320 ;
        RECT 2208.070 96.260 2208.390 96.320 ;
        RECT 2208.990 48.180 2209.310 48.240 ;
        RECT 2208.795 48.040 2209.310 48.180 ;
        RECT 2208.990 47.980 2209.310 48.040 ;
        RECT 2208.990 2.960 2209.310 3.020 ;
        RECT 2208.795 2.820 2209.310 2.960 ;
        RECT 2208.990 2.760 2209.310 2.820 ;
      LAYER via ;
        RECT 2099.540 243.820 2099.800 244.080 ;
        RECT 2104.140 243.820 2104.400 244.080 ;
        RECT 2104.140 114.280 2104.400 114.540 ;
        RECT 2208.100 114.280 2208.360 114.540 ;
        RECT 2207.640 96.260 2207.900 96.520 ;
        RECT 2208.100 96.260 2208.360 96.520 ;
        RECT 2209.020 47.980 2209.280 48.240 ;
        RECT 2209.020 2.760 2209.280 3.020 ;
      LAYER met2 ;
        RECT 2099.490 260.000 2099.770 264.000 ;
        RECT 2099.600 244.110 2099.740 260.000 ;
        RECT 2099.540 243.790 2099.800 244.110 ;
        RECT 2104.140 243.790 2104.400 244.110 ;
        RECT 2104.200 114.570 2104.340 243.790 ;
        RECT 2104.140 114.250 2104.400 114.570 ;
        RECT 2208.100 114.250 2208.360 114.570 ;
        RECT 2208.160 96.550 2208.300 114.250 ;
        RECT 2207.640 96.230 2207.900 96.550 ;
        RECT 2208.100 96.230 2208.360 96.550 ;
        RECT 2207.700 48.805 2207.840 96.230 ;
        RECT 2207.630 48.435 2207.910 48.805 ;
        RECT 2209.010 48.435 2209.290 48.805 ;
        RECT 2209.080 48.270 2209.220 48.435 ;
        RECT 2209.020 47.950 2209.280 48.270 ;
        RECT 2209.020 2.730 2209.280 3.050 ;
        RECT 2209.080 2.400 2209.220 2.730 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
      LAYER via2 ;
        RECT 2207.630 48.480 2207.910 48.760 ;
        RECT 2209.010 48.480 2209.290 48.760 ;
      LAYER met3 ;
        RECT 2207.605 48.770 2207.935 48.785 ;
        RECT 2208.985 48.770 2209.315 48.785 ;
        RECT 2207.605 48.470 2209.315 48.770 ;
        RECT 2207.605 48.455 2207.935 48.470 ;
        RECT 2208.985 48.455 2209.315 48.470 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 243.870 610.540 244.190 610.600 ;
        RECT 301.370 610.540 301.690 610.600 ;
        RECT 243.870 610.400 301.690 610.540 ;
        RECT 243.870 610.340 244.190 610.400 ;
        RECT 301.370 610.340 301.690 610.400 ;
        RECT 243.870 46.820 244.190 46.880 ;
        RECT 2226.930 46.820 2227.250 46.880 ;
        RECT 243.870 46.680 2227.250 46.820 ;
        RECT 243.870 46.620 244.190 46.680 ;
        RECT 2226.930 46.620 2227.250 46.680 ;
      LAYER via ;
        RECT 243.900 610.340 244.160 610.600 ;
        RECT 301.400 610.340 301.660 610.600 ;
        RECT 243.900 46.620 244.160 46.880 ;
        RECT 2226.960 46.620 2227.220 46.880 ;
      LAYER met2 ;
        RECT 301.390 1974.875 301.670 1975.245 ;
        RECT 301.460 610.630 301.600 1974.875 ;
        RECT 243.900 610.310 244.160 610.630 ;
        RECT 301.400 610.310 301.660 610.630 ;
        RECT 243.960 46.910 244.100 610.310 ;
        RECT 243.900 46.590 244.160 46.910 ;
        RECT 2226.960 46.590 2227.220 46.910 ;
        RECT 2227.020 2.400 2227.160 46.590 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
      LAYER via2 ;
        RECT 301.390 1974.920 301.670 1975.200 ;
      LAYER met3 ;
        RECT 301.365 1975.210 301.695 1975.225 ;
        RECT 310.000 1975.210 314.000 1975.600 ;
        RECT 301.365 1975.000 314.000 1975.210 ;
        RECT 301.365 1974.910 310.500 1975.000 ;
        RECT 301.365 1974.895 301.695 1974.910 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 779.845 96.645 780.015 144.755 ;
        RECT 779.845 48.365 780.015 96.135 ;
      LAYER mcon ;
        RECT 779.845 144.585 780.015 144.755 ;
        RECT 779.845 95.965 780.015 96.135 ;
      LAYER met1 ;
        RECT 288.490 2732.480 288.810 2732.540 ;
        RECT 296.770 2732.480 297.090 2732.540 ;
        RECT 288.490 2732.340 297.090 2732.480 ;
        RECT 288.490 2732.280 288.810 2732.340 ;
        RECT 296.770 2732.280 297.090 2732.340 ;
        RECT 288.490 169.560 288.810 169.620 ;
        RECT 779.770 169.560 780.090 169.620 ;
        RECT 288.490 169.420 780.090 169.560 ;
        RECT 288.490 169.360 288.810 169.420 ;
        RECT 779.770 169.360 780.090 169.420 ;
        RECT 779.770 144.740 780.090 144.800 ;
        RECT 779.575 144.600 780.090 144.740 ;
        RECT 779.770 144.540 780.090 144.600 ;
        RECT 779.770 96.800 780.090 96.860 ;
        RECT 779.575 96.660 780.090 96.800 ;
        RECT 779.770 96.600 780.090 96.660 ;
        RECT 779.770 96.120 780.090 96.180 ;
        RECT 779.575 95.980 780.090 96.120 ;
        RECT 779.770 95.920 780.090 95.980 ;
        RECT 779.785 48.520 780.075 48.565 ;
        RECT 781.610 48.520 781.930 48.580 ;
        RECT 779.785 48.380 781.930 48.520 ;
        RECT 779.785 48.335 780.075 48.380 ;
        RECT 781.610 48.320 781.930 48.380 ;
      LAYER via ;
        RECT 288.520 2732.280 288.780 2732.540 ;
        RECT 296.800 2732.280 297.060 2732.540 ;
        RECT 288.520 169.360 288.780 169.620 ;
        RECT 779.800 169.360 780.060 169.620 ;
        RECT 779.800 144.540 780.060 144.800 ;
        RECT 779.800 96.600 780.060 96.860 ;
        RECT 779.800 95.920 780.060 96.180 ;
        RECT 781.640 48.320 781.900 48.580 ;
      LAYER met2 ;
        RECT 296.790 2736.475 297.070 2736.845 ;
        RECT 296.860 2732.570 297.000 2736.475 ;
        RECT 288.520 2732.250 288.780 2732.570 ;
        RECT 296.800 2732.250 297.060 2732.570 ;
        RECT 288.580 169.650 288.720 2732.250 ;
        RECT 288.520 169.330 288.780 169.650 ;
        RECT 779.800 169.330 780.060 169.650 ;
        RECT 779.860 144.830 780.000 169.330 ;
        RECT 779.800 144.510 780.060 144.830 ;
        RECT 779.800 96.570 780.060 96.890 ;
        RECT 779.860 96.210 780.000 96.570 ;
        RECT 779.800 95.890 780.060 96.210 ;
        RECT 781.640 48.290 781.900 48.610 ;
        RECT 781.700 2.400 781.840 48.290 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 296.790 2736.520 297.070 2736.800 ;
      LAYER met3 ;
        RECT 296.765 2736.810 297.095 2736.825 ;
        RECT 310.000 2736.810 314.000 2737.200 ;
        RECT 296.765 2736.600 314.000 2736.810 ;
        RECT 296.765 2736.510 310.500 2736.600 ;
        RECT 296.765 2736.495 297.095 2736.510 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.890 51.835 2245.170 52.205 ;
        RECT 2244.960 2.400 2245.100 51.835 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
      LAYER via2 ;
        RECT 2244.890 51.880 2245.170 52.160 ;
      LAYER met3 ;
        RECT 288.230 2863.290 288.610 2863.300 ;
        RECT 310.000 2863.290 314.000 2863.680 ;
        RECT 288.230 2863.080 314.000 2863.290 ;
        RECT 288.230 2862.990 310.500 2863.080 ;
        RECT 288.230 2862.980 288.610 2862.990 ;
        RECT 288.230 52.170 288.610 52.180 ;
        RECT 2244.865 52.170 2245.195 52.185 ;
        RECT 288.230 51.870 2245.195 52.170 ;
        RECT 288.230 51.860 288.610 51.870 ;
        RECT 2244.865 51.855 2245.195 51.870 ;
      LAYER via3 ;
        RECT 288.260 2862.980 288.580 2863.300 ;
        RECT 288.260 51.860 288.580 52.180 ;
      LAYER met4 ;
        RECT 288.255 2862.975 288.585 2863.305 ;
        RECT 288.270 52.185 288.570 2862.975 ;
        RECT 288.255 51.855 288.585 52.185 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 298.610 72.320 298.930 72.380 ;
        RECT 2256.370 72.320 2256.690 72.380 ;
        RECT 298.610 72.180 2256.690 72.320 ;
        RECT 298.610 72.120 298.930 72.180 ;
        RECT 2256.370 72.120 2256.690 72.180 ;
        RECT 2256.370 37.640 2256.690 37.700 ;
        RECT 2262.350 37.640 2262.670 37.700 ;
        RECT 2256.370 37.500 2262.670 37.640 ;
        RECT 2256.370 37.440 2256.690 37.500 ;
        RECT 2262.350 37.440 2262.670 37.500 ;
      LAYER via ;
        RECT 298.640 72.120 298.900 72.380 ;
        RECT 2256.400 72.120 2256.660 72.380 ;
        RECT 2256.400 37.440 2256.660 37.700 ;
        RECT 2262.380 37.440 2262.640 37.700 ;
      LAYER met2 ;
        RECT 298.630 580.875 298.910 581.245 ;
        RECT 298.700 72.410 298.840 580.875 ;
        RECT 298.640 72.090 298.900 72.410 ;
        RECT 2256.400 72.090 2256.660 72.410 ;
        RECT 2256.460 37.730 2256.600 72.090 ;
        RECT 2256.400 37.410 2256.660 37.730 ;
        RECT 2262.380 37.410 2262.640 37.730 ;
        RECT 2262.440 2.400 2262.580 37.410 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
      LAYER via2 ;
        RECT 298.630 580.920 298.910 581.200 ;
      LAYER met3 ;
        RECT 298.605 581.210 298.935 581.225 ;
        RECT 310.000 581.210 314.000 581.600 ;
        RECT 298.605 581.000 314.000 581.210 ;
        RECT 298.605 580.910 310.500 581.000 ;
        RECT 298.605 580.895 298.935 580.910 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2283.510 260.340 2283.830 260.400 ;
        RECT 2610.570 260.340 2610.890 260.400 ;
        RECT 2283.510 260.200 2610.890 260.340 ;
        RECT 2283.510 260.140 2283.830 260.200 ;
        RECT 2610.570 260.140 2610.890 260.200 ;
        RECT 2280.290 17.920 2280.610 17.980 ;
        RECT 2283.510 17.920 2283.830 17.980 ;
        RECT 2280.290 17.780 2283.830 17.920 ;
        RECT 2280.290 17.720 2280.610 17.780 ;
        RECT 2283.510 17.720 2283.830 17.780 ;
      LAYER via ;
        RECT 2283.540 260.140 2283.800 260.400 ;
        RECT 2610.600 260.140 2610.860 260.400 ;
        RECT 2280.320 17.720 2280.580 17.980 ;
        RECT 2283.540 17.720 2283.800 17.980 ;
      LAYER met2 ;
        RECT 2610.590 1818.475 2610.870 1818.845 ;
        RECT 2610.660 260.430 2610.800 1818.475 ;
        RECT 2283.540 260.110 2283.800 260.430 ;
        RECT 2610.600 260.110 2610.860 260.430 ;
        RECT 2283.600 18.010 2283.740 260.110 ;
        RECT 2280.320 17.690 2280.580 18.010 ;
        RECT 2283.540 17.690 2283.800 18.010 ;
        RECT 2280.380 2.400 2280.520 17.690 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
      LAYER via2 ;
        RECT 2610.590 1818.520 2610.870 1818.800 ;
      LAYER met3 ;
        RECT 2606.000 1818.810 2610.000 1819.200 ;
        RECT 2610.565 1818.810 2610.895 1818.825 ;
        RECT 2606.000 1818.600 2610.895 1818.810 ;
        RECT 2609.580 1818.510 2610.895 1818.600 ;
        RECT 2610.565 1818.495 2610.895 1818.510 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.490 3257.440 978.810 3257.500 ;
        RECT 2664.390 3257.440 2664.710 3257.500 ;
        RECT 978.490 3257.300 2664.710 3257.440 ;
        RECT 978.490 3257.240 978.810 3257.300 ;
        RECT 2664.390 3257.240 2664.710 3257.300 ;
      LAYER via ;
        RECT 978.520 3257.240 978.780 3257.500 ;
        RECT 2664.420 3257.240 2664.680 3257.500 ;
      LAYER met2 ;
        RECT 977.090 3257.610 977.370 3260.000 ;
        RECT 977.090 3257.530 978.720 3257.610 ;
        RECT 977.090 3257.470 978.780 3257.530 ;
        RECT 977.090 3256.000 977.370 3257.470 ;
        RECT 978.520 3257.210 978.780 3257.470 ;
        RECT 2664.420 3257.210 2664.680 3257.530 ;
        RECT 2356.210 19.875 2356.490 20.245 ;
        RECT 2404.510 19.875 2404.790 20.245 ;
        RECT 2451.890 19.875 2452.170 20.245 ;
        RECT 2501.110 19.875 2501.390 20.245 ;
        RECT 2356.280 15.485 2356.420 19.875 ;
        RECT 2404.580 15.485 2404.720 19.875 ;
        RECT 2451.960 15.485 2452.100 19.875 ;
        RECT 2501.180 15.485 2501.320 19.875 ;
        RECT 2664.480 19.565 2664.620 3257.210 ;
        RECT 2586.210 19.195 2586.490 19.565 ;
        RECT 2664.410 19.195 2664.690 19.565 ;
        RECT 2586.280 16.845 2586.420 19.195 ;
        RECT 2549.410 16.475 2549.690 16.845 ;
        RECT 2586.210 16.475 2586.490 16.845 ;
        RECT 2549.480 15.485 2549.620 16.475 ;
        RECT 2298.250 15.115 2298.530 15.485 ;
        RECT 2356.210 15.115 2356.490 15.485 ;
        RECT 2404.510 15.115 2404.790 15.485 ;
        RECT 2451.890 15.115 2452.170 15.485 ;
        RECT 2501.110 15.115 2501.390 15.485 ;
        RECT 2549.410 15.115 2549.690 15.485 ;
        RECT 2298.320 2.400 2298.460 15.115 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
      LAYER via2 ;
        RECT 2356.210 19.920 2356.490 20.200 ;
        RECT 2404.510 19.920 2404.790 20.200 ;
        RECT 2451.890 19.920 2452.170 20.200 ;
        RECT 2501.110 19.920 2501.390 20.200 ;
        RECT 2586.210 19.240 2586.490 19.520 ;
        RECT 2664.410 19.240 2664.690 19.520 ;
        RECT 2549.410 16.520 2549.690 16.800 ;
        RECT 2586.210 16.520 2586.490 16.800 ;
        RECT 2298.250 15.160 2298.530 15.440 ;
        RECT 2356.210 15.160 2356.490 15.440 ;
        RECT 2404.510 15.160 2404.790 15.440 ;
        RECT 2451.890 15.160 2452.170 15.440 ;
        RECT 2501.110 15.160 2501.390 15.440 ;
        RECT 2549.410 15.160 2549.690 15.440 ;
      LAYER met3 ;
        RECT 2356.185 20.210 2356.515 20.225 ;
        RECT 2404.485 20.210 2404.815 20.225 ;
        RECT 2356.185 19.910 2404.815 20.210 ;
        RECT 2356.185 19.895 2356.515 19.910 ;
        RECT 2404.485 19.895 2404.815 19.910 ;
        RECT 2451.865 20.210 2452.195 20.225 ;
        RECT 2501.085 20.210 2501.415 20.225 ;
        RECT 2451.865 19.910 2501.415 20.210 ;
        RECT 2451.865 19.895 2452.195 19.910 ;
        RECT 2501.085 19.895 2501.415 19.910 ;
        RECT 2586.185 19.530 2586.515 19.545 ;
        RECT 2664.385 19.530 2664.715 19.545 ;
        RECT 2586.185 19.230 2664.715 19.530 ;
        RECT 2586.185 19.215 2586.515 19.230 ;
        RECT 2664.385 19.215 2664.715 19.230 ;
        RECT 2549.385 16.810 2549.715 16.825 ;
        RECT 2586.185 16.810 2586.515 16.825 ;
        RECT 2549.385 16.510 2586.515 16.810 ;
        RECT 2549.385 16.495 2549.715 16.510 ;
        RECT 2586.185 16.495 2586.515 16.510 ;
        RECT 2298.225 15.450 2298.555 15.465 ;
        RECT 2356.185 15.450 2356.515 15.465 ;
        RECT 2298.225 15.150 2356.515 15.450 ;
        RECT 2298.225 15.135 2298.555 15.150 ;
        RECT 2356.185 15.135 2356.515 15.150 ;
        RECT 2404.485 15.450 2404.815 15.465 ;
        RECT 2451.865 15.450 2452.195 15.465 ;
        RECT 2404.485 15.150 2452.195 15.450 ;
        RECT 2404.485 15.135 2404.815 15.150 ;
        RECT 2451.865 15.135 2452.195 15.150 ;
        RECT 2501.085 15.450 2501.415 15.465 ;
        RECT 2549.385 15.450 2549.715 15.465 ;
        RECT 2501.085 15.150 2549.715 15.450 ;
        RECT 2501.085 15.135 2501.415 15.150 ;
        RECT 2549.385 15.135 2549.715 15.150 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 223.960 2318.330 224.020 ;
        RECT 2606.890 223.960 2607.210 224.020 ;
        RECT 2318.010 223.820 2607.210 223.960 ;
        RECT 2318.010 223.760 2318.330 223.820 ;
        RECT 2606.890 223.760 2607.210 223.820 ;
        RECT 2316.170 2.960 2316.490 3.020 ;
        RECT 2318.010 2.960 2318.330 3.020 ;
        RECT 2316.170 2.820 2318.330 2.960 ;
        RECT 2316.170 2.760 2316.490 2.820 ;
        RECT 2318.010 2.760 2318.330 2.820 ;
      LAYER via ;
        RECT 2318.040 223.760 2318.300 224.020 ;
        RECT 2606.920 223.760 2607.180 224.020 ;
        RECT 2316.200 2.760 2316.460 3.020 ;
        RECT 2318.040 2.760 2318.300 3.020 ;
      LAYER met2 ;
        RECT 2606.910 1773.595 2607.190 1773.965 ;
        RECT 2606.980 224.050 2607.120 1773.595 ;
        RECT 2318.040 223.730 2318.300 224.050 ;
        RECT 2606.920 223.730 2607.180 224.050 ;
        RECT 2318.100 3.050 2318.240 223.730 ;
        RECT 2316.200 2.730 2316.460 3.050 ;
        RECT 2318.040 2.730 2318.300 3.050 ;
        RECT 2316.260 2.400 2316.400 2.730 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
      LAYER via2 ;
        RECT 2606.910 1773.640 2607.190 1773.920 ;
      LAYER met3 ;
        RECT 2606.000 1775.080 2610.000 1775.680 ;
        RECT 2606.670 1773.945 2606.970 1775.080 ;
        RECT 2606.670 1773.630 2607.215 1773.945 ;
        RECT 2606.885 1773.615 2607.215 1773.630 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2615.170 400.420 2615.490 400.480 ;
        RECT 2645.070 400.420 2645.390 400.480 ;
        RECT 2615.170 400.280 2645.390 400.420 ;
        RECT 2615.170 400.220 2615.490 400.280 ;
        RECT 2645.070 400.220 2645.390 400.280 ;
        RECT 2338.710 260.680 2339.030 260.740 ;
        RECT 2645.070 260.680 2645.390 260.740 ;
        RECT 2338.710 260.540 2645.390 260.680 ;
        RECT 2338.710 260.480 2339.030 260.540 ;
        RECT 2645.070 260.480 2645.390 260.540 ;
        RECT 2334.110 17.920 2334.430 17.980 ;
        RECT 2338.710 17.920 2339.030 17.980 ;
        RECT 2334.110 17.780 2339.030 17.920 ;
        RECT 2334.110 17.720 2334.430 17.780 ;
        RECT 2338.710 17.720 2339.030 17.780 ;
      LAYER via ;
        RECT 2615.200 400.220 2615.460 400.480 ;
        RECT 2645.100 400.220 2645.360 400.480 ;
        RECT 2338.740 260.480 2339.000 260.740 ;
        RECT 2645.100 260.480 2645.360 260.740 ;
        RECT 2334.140 17.720 2334.400 17.980 ;
        RECT 2338.740 17.720 2339.000 17.980 ;
      LAYER met2 ;
        RECT 2615.190 401.355 2615.470 401.725 ;
        RECT 2615.260 400.510 2615.400 401.355 ;
        RECT 2615.200 400.190 2615.460 400.510 ;
        RECT 2645.100 400.190 2645.360 400.510 ;
        RECT 2645.160 260.770 2645.300 400.190 ;
        RECT 2338.740 260.450 2339.000 260.770 ;
        RECT 2645.100 260.450 2645.360 260.770 ;
        RECT 2338.800 18.010 2338.940 260.450 ;
        RECT 2334.140 17.690 2334.400 18.010 ;
        RECT 2338.740 17.690 2339.000 18.010 ;
        RECT 2334.200 2.400 2334.340 17.690 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
      LAYER via2 ;
        RECT 2615.190 401.400 2615.470 401.680 ;
      LAYER met3 ;
        RECT 2606.000 401.690 2610.000 402.080 ;
        RECT 2615.165 401.690 2615.495 401.705 ;
        RECT 2606.000 401.480 2615.495 401.690 ;
        RECT 2609.580 401.390 2615.495 401.480 ;
        RECT 2615.165 401.375 2615.495 401.390 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 3259.395 457.610 3259.765 ;
        RECT 457.400 3258.970 457.540 3259.395 ;
        RECT 461.890 3258.970 462.170 3260.000 ;
        RECT 457.400 3258.830 462.170 3258.970 ;
        RECT 461.890 3256.000 462.170 3258.830 ;
        RECT 2351.610 15.795 2351.890 16.165 ;
        RECT 2351.680 2.400 2351.820 15.795 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
      LAYER via2 ;
        RECT 457.330 3259.440 457.610 3259.720 ;
        RECT 2351.610 15.840 2351.890 16.120 ;
      LAYER met3 ;
        RECT 247.750 3259.730 248.130 3259.740 ;
        RECT 457.305 3259.730 457.635 3259.745 ;
        RECT 247.750 3259.430 457.635 3259.730 ;
        RECT 247.750 3259.420 248.130 3259.430 ;
        RECT 457.305 3259.415 457.635 3259.430 ;
        RECT 1041.710 22.250 1042.090 22.260 ;
        RECT 1089.550 22.250 1089.930 22.260 ;
        RECT 1041.710 21.950 1089.930 22.250 ;
        RECT 1041.710 21.940 1042.090 21.950 ;
        RECT 1089.550 21.940 1089.930 21.950 ;
        RECT 1345.310 19.530 1345.690 19.540 ;
        RECT 1366.470 19.530 1366.850 19.540 ;
        RECT 1345.310 19.230 1366.850 19.530 ;
        RECT 1345.310 19.220 1345.690 19.230 ;
        RECT 1366.470 19.220 1366.850 19.230 ;
        RECT 1924.910 18.850 1925.290 18.860 ;
        RECT 1972.750 18.850 1973.130 18.860 ;
        RECT 1924.910 18.550 1973.130 18.850 ;
        RECT 1924.910 18.540 1925.290 18.550 ;
        RECT 1972.750 18.540 1973.130 18.550 ;
        RECT 1980.110 18.850 1980.490 18.860 ;
        RECT 2027.950 18.850 2028.330 18.860 ;
        RECT 1980.110 18.550 2028.330 18.850 ;
        RECT 1980.110 18.540 1980.490 18.550 ;
        RECT 2027.950 18.540 2028.330 18.550 ;
        RECT 2070.270 18.850 2070.650 18.860 ;
        RECT 2142.030 18.850 2142.410 18.860 ;
        RECT 2070.270 18.550 2142.410 18.850 ;
        RECT 2070.270 18.540 2070.650 18.550 ;
        RECT 2142.030 18.540 2142.410 18.550 ;
        RECT 2318.670 16.130 2319.050 16.140 ;
        RECT 2351.585 16.130 2351.915 16.145 ;
        RECT 2318.670 15.830 2351.915 16.130 ;
        RECT 2318.670 15.820 2319.050 15.830 ;
        RECT 2351.585 15.815 2351.915 15.830 ;
        RECT 444.630 15.450 445.010 15.460 ;
        RECT 468.550 15.450 468.930 15.460 ;
        RECT 444.630 15.150 468.930 15.450 ;
        RECT 444.630 15.140 445.010 15.150 ;
        RECT 468.550 15.140 468.930 15.150 ;
        RECT 589.990 15.450 590.370 15.460 ;
        RECT 596.430 15.450 596.810 15.460 ;
        RECT 589.990 15.150 596.810 15.450 ;
        RECT 589.990 15.140 590.370 15.150 ;
        RECT 596.430 15.140 596.810 15.150 ;
        RECT 613.910 15.450 614.290 15.460 ;
        RECT 661.750 15.450 662.130 15.460 ;
        RECT 613.910 15.150 662.130 15.450 ;
        RECT 613.910 15.140 614.290 15.150 ;
        RECT 661.750 15.140 662.130 15.150 ;
        RECT 807.110 15.450 807.490 15.460 ;
        RECT 896.350 15.450 896.730 15.460 ;
        RECT 807.110 15.150 896.730 15.450 ;
        RECT 807.110 15.140 807.490 15.150 ;
        RECT 896.350 15.140 896.730 15.150 ;
        RECT 1441.910 15.450 1442.290 15.460 ;
        RECT 1489.750 15.450 1490.130 15.460 ;
        RECT 1441.910 15.150 1490.130 15.450 ;
        RECT 1441.910 15.140 1442.290 15.150 ;
        RECT 1489.750 15.140 1490.130 15.150 ;
        RECT 1685.710 15.450 1686.090 15.460 ;
        RECT 1730.790 15.450 1731.170 15.460 ;
        RECT 1685.710 15.150 1731.170 15.450 ;
        RECT 1685.710 15.140 1686.090 15.150 ;
        RECT 1730.790 15.140 1731.170 15.150 ;
        RECT 1755.630 15.450 1756.010 15.460 ;
        RECT 1785.990 15.450 1786.370 15.460 ;
        RECT 1755.630 15.150 1786.370 15.450 ;
        RECT 1755.630 15.140 1756.010 15.150 ;
        RECT 1785.990 15.140 1786.370 15.150 ;
        RECT 1797.950 15.450 1798.330 15.460 ;
        RECT 1834.750 15.450 1835.130 15.460 ;
        RECT 1797.950 15.150 1835.130 15.450 ;
        RECT 1797.950 15.140 1798.330 15.150 ;
        RECT 1834.750 15.140 1835.130 15.150 ;
      LAYER via3 ;
        RECT 247.780 3259.420 248.100 3259.740 ;
        RECT 1041.740 21.940 1042.060 22.260 ;
        RECT 1089.580 21.940 1089.900 22.260 ;
        RECT 1345.340 19.220 1345.660 19.540 ;
        RECT 1366.500 19.220 1366.820 19.540 ;
        RECT 1924.940 18.540 1925.260 18.860 ;
        RECT 1972.780 18.540 1973.100 18.860 ;
        RECT 1980.140 18.540 1980.460 18.860 ;
        RECT 2027.980 18.540 2028.300 18.860 ;
        RECT 2070.300 18.540 2070.620 18.860 ;
        RECT 2142.060 18.540 2142.380 18.860 ;
        RECT 2318.700 15.820 2319.020 16.140 ;
        RECT 444.660 15.140 444.980 15.460 ;
        RECT 468.580 15.140 468.900 15.460 ;
        RECT 590.020 15.140 590.340 15.460 ;
        RECT 596.460 15.140 596.780 15.460 ;
        RECT 613.940 15.140 614.260 15.460 ;
        RECT 661.780 15.140 662.100 15.460 ;
        RECT 807.140 15.140 807.460 15.460 ;
        RECT 896.380 15.140 896.700 15.460 ;
        RECT 1441.940 15.140 1442.260 15.460 ;
        RECT 1489.780 15.140 1490.100 15.460 ;
        RECT 1685.740 15.140 1686.060 15.460 ;
        RECT 1730.820 15.140 1731.140 15.460 ;
        RECT 1755.660 15.140 1755.980 15.460 ;
        RECT 1786.020 15.140 1786.340 15.460 ;
        RECT 1797.980 15.140 1798.300 15.460 ;
        RECT 1834.780 15.140 1835.100 15.460 ;
      LAYER met4 ;
        RECT 247.775 3259.415 248.105 3259.745 ;
        RECT 247.790 15.890 248.090 3259.415 ;
        RECT 1041.310 21.510 1042.490 22.690 ;
        RECT 1089.575 21.935 1089.905 22.265 ;
        RECT 1096.510 22.250 1097.690 22.690 ;
        RECT 1096.510 21.950 1100.010 22.250 ;
        RECT 589.590 18.110 590.770 19.290 ;
        RECT 710.110 18.850 711.290 19.290 ;
        RECT 710.110 18.550 713.610 18.850 ;
        RECT 710.110 18.110 711.290 18.550 ;
        RECT 247.350 14.710 248.530 15.890 ;
        RECT 444.230 14.710 445.410 15.890 ;
        RECT 468.150 14.710 469.330 15.890 ;
        RECT 590.030 15.465 590.330 18.110 ;
        RECT 713.310 15.890 713.610 18.550 ;
        RECT 806.710 18.110 807.890 19.290 ;
        RECT 590.015 15.135 590.345 15.465 ;
        RECT 596.030 14.710 597.210 15.890 ;
        RECT 613.510 14.710 614.690 15.890 ;
        RECT 661.350 14.710 662.530 15.890 ;
        RECT 712.870 14.710 714.050 15.890 ;
        RECT 807.150 15.465 807.450 18.110 ;
        RECT 1089.590 15.890 1089.890 21.935 ;
        RECT 1096.510 21.510 1097.690 21.950 ;
        RECT 1099.710 19.290 1100.010 21.950 ;
        RECT 1730.390 21.510 1731.570 22.690 ;
        RECT 1755.230 21.510 1756.410 22.690 ;
        RECT 2141.630 21.510 2142.810 22.690 ;
        RECT 1345.335 19.290 1345.665 19.545 ;
        RECT 1366.495 19.290 1366.825 19.545 ;
        RECT 1099.270 18.110 1100.450 19.290 ;
        RECT 1344.910 18.110 1346.090 19.290 ;
        RECT 1366.070 18.110 1367.250 19.290 ;
        RECT 1441.510 18.110 1442.690 19.290 ;
        RECT 807.135 15.135 807.465 15.465 ;
        RECT 895.950 14.710 897.130 15.890 ;
        RECT 1089.150 14.710 1090.330 15.890 ;
        RECT 1441.950 15.465 1442.250 18.110 ;
        RECT 1441.935 15.135 1442.265 15.465 ;
        RECT 1489.350 14.710 1490.530 15.890 ;
        RECT 1685.310 14.710 1686.490 15.890 ;
        RECT 1730.830 15.465 1731.130 21.510 ;
        RECT 1755.670 15.465 1755.970 21.510 ;
        RECT 1834.350 18.110 1835.530 19.290 ;
        RECT 1924.510 18.110 1925.690 19.290 ;
        RECT 1972.350 18.110 1973.530 19.290 ;
        RECT 1979.710 18.110 1980.890 19.290 ;
        RECT 2142.070 18.865 2142.370 21.510 ;
        RECT 2027.975 18.535 2028.305 18.865 ;
        RECT 2070.295 18.535 2070.625 18.865 ;
        RECT 2142.055 18.535 2142.385 18.865 ;
        RECT 1730.815 15.135 1731.145 15.465 ;
        RECT 1755.655 15.135 1755.985 15.465 ;
        RECT 1785.590 14.710 1786.770 15.890 ;
        RECT 1797.550 14.710 1798.730 15.890 ;
        RECT 1834.790 15.465 1835.090 18.110 ;
        RECT 2027.990 15.890 2028.290 18.535 ;
        RECT 2070.310 15.890 2070.610 18.535 ;
        RECT 2175.670 18.110 2176.850 19.290 ;
        RECT 2318.270 18.110 2319.450 19.290 ;
        RECT 1834.775 15.135 1835.105 15.465 ;
        RECT 2027.550 14.710 2028.730 15.890 ;
        RECT 2069.870 14.710 2071.050 15.890 ;
        RECT 2172.910 15.450 2174.090 15.890 ;
        RECT 2176.110 15.450 2176.410 18.110 ;
        RECT 2318.710 16.145 2319.010 18.110 ;
        RECT 2318.695 15.815 2319.025 16.145 ;
        RECT 2172.910 15.150 2176.410 15.450 ;
        RECT 2172.910 14.710 2174.090 15.150 ;
      LAYER met5 ;
        RECT 944.500 21.300 993.940 22.900 ;
        RECT 330.860 17.900 375.700 19.500 ;
        RECT 330.860 16.100 332.460 17.900 ;
        RECT 247.140 14.500 332.460 16.100 ;
        RECT 374.100 16.100 375.700 17.900 ;
        RECT 419.180 16.100 421.700 18.140 ;
        RECT 496.460 17.900 590.980 19.500 ;
        RECT 685.980 17.900 711.500 19.500 ;
        RECT 758.660 17.900 808.100 19.500 ;
        RECT 496.460 16.100 498.060 17.900 ;
        RECT 685.980 16.100 687.580 17.900 ;
        RECT 758.660 16.100 760.260 17.900 ;
        RECT 944.500 16.100 946.100 21.300 ;
        RECT 374.100 14.500 445.620 16.100 ;
        RECT 467.940 14.500 498.060 16.100 ;
        RECT 595.820 14.500 614.900 16.100 ;
        RECT 661.140 14.500 687.580 16.100 ;
        RECT 712.660 14.500 760.260 16.100 ;
        RECT 895.740 14.500 946.100 16.100 ;
        RECT 992.340 16.100 993.940 21.300 ;
        RECT 1001.540 21.300 1042.700 22.900 ;
        RECT 1095.380 21.300 1098.680 22.900 ;
        RECT 1497.420 21.300 1545.940 22.900 ;
        RECT 1730.180 21.300 1756.620 22.900 ;
        RECT 2141.420 21.300 2166.940 22.900 ;
        RECT 1001.540 16.100 1003.140 21.300 ;
        RECT 1095.380 16.100 1096.980 21.300 ;
        RECT 1099.060 17.900 1174.260 19.500 ;
        RECT 992.340 14.500 1003.140 16.100 ;
        RECT 1088.940 14.500 1096.980 16.100 ;
        RECT 1172.660 16.100 1174.260 17.900 ;
        RECT 1220.500 17.900 1346.300 19.500 ;
        RECT 1365.860 17.900 1394.140 19.500 ;
        RECT 1220.500 16.100 1222.100 17.900 ;
        RECT 1172.660 14.500 1222.100 16.100 ;
        RECT 1392.540 16.100 1394.140 17.900 ;
        RECT 1414.620 17.900 1442.900 19.500 ;
        RECT 1414.620 16.100 1416.220 17.900 ;
        RECT 1497.420 16.100 1499.020 21.300 ;
        RECT 1392.540 14.500 1416.220 16.100 ;
        RECT 1489.140 14.500 1499.020 16.100 ;
        RECT 1544.340 16.100 1545.940 21.300 ;
        RECT 1606.900 17.900 1660.020 19.500 ;
        RECT 1834.140 17.900 1925.900 19.500 ;
        RECT 1972.140 17.900 1981.100 19.500 ;
        RECT 1606.900 16.100 1608.500 17.900 ;
        RECT 1544.340 14.500 1608.500 16.100 ;
        RECT 1658.420 16.100 1660.020 17.900 ;
        RECT 2165.340 16.100 2166.940 21.300 ;
        RECT 2175.460 17.900 2319.660 19.500 ;
        RECT 1658.420 14.500 1686.700 16.100 ;
        RECT 1785.380 14.500 1798.940 16.100 ;
        RECT 2027.340 14.500 2071.260 16.100 ;
        RECT 2165.340 14.500 2174.300 16.100 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2369.605 2.805 2369.775 48.195 ;
      LAYER mcon ;
        RECT 2369.605 48.025 2369.775 48.195 ;
      LAYER met1 ;
        RECT 386.010 65.520 386.330 65.580 ;
        RECT 2367.230 65.520 2367.550 65.580 ;
        RECT 386.010 65.380 2367.550 65.520 ;
        RECT 386.010 65.320 386.330 65.380 ;
        RECT 2367.230 65.320 2367.550 65.380 ;
        RECT 2367.230 48.180 2367.550 48.240 ;
        RECT 2369.545 48.180 2369.835 48.225 ;
        RECT 2367.230 48.040 2369.835 48.180 ;
        RECT 2367.230 47.980 2367.550 48.040 ;
        RECT 2369.545 47.995 2369.835 48.040 ;
        RECT 2369.530 2.960 2369.850 3.020 ;
        RECT 2369.335 2.820 2369.850 2.960 ;
        RECT 2369.530 2.760 2369.850 2.820 ;
      LAYER via ;
        RECT 386.040 65.320 386.300 65.580 ;
        RECT 2367.260 65.320 2367.520 65.580 ;
        RECT 2367.260 47.980 2367.520 48.240 ;
        RECT 2369.560 2.760 2369.820 3.020 ;
      LAYER met2 ;
        RECT 383.690 260.170 383.970 264.000 ;
        RECT 383.690 260.030 386.240 260.170 ;
        RECT 383.690 260.000 383.970 260.030 ;
        RECT 386.100 65.610 386.240 260.030 ;
        RECT 386.040 65.290 386.300 65.610 ;
        RECT 2367.260 65.290 2367.520 65.610 ;
        RECT 2367.320 48.270 2367.460 65.290 ;
        RECT 2367.260 47.950 2367.520 48.270 ;
        RECT 2369.560 2.730 2369.820 3.050 ;
        RECT 2369.620 2.400 2369.760 2.730 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2392.070 3273.760 2392.390 3273.820 ;
        RECT 2661.170 3273.760 2661.490 3273.820 ;
        RECT 2392.070 3273.620 2661.490 3273.760 ;
        RECT 2392.070 3273.560 2392.390 3273.620 ;
        RECT 2661.170 3273.560 2661.490 3273.620 ;
        RECT 2387.470 17.920 2387.790 17.980 ;
        RECT 2393.910 17.920 2394.230 17.980 ;
        RECT 2387.470 17.780 2394.230 17.920 ;
        RECT 2387.470 17.720 2387.790 17.780 ;
        RECT 2393.910 17.720 2394.230 17.780 ;
      LAYER via ;
        RECT 2392.100 3273.560 2392.360 3273.820 ;
        RECT 2661.200 3273.560 2661.460 3273.820 ;
        RECT 2387.500 17.720 2387.760 17.980 ;
        RECT 2393.940 17.720 2394.200 17.980 ;
      LAYER met2 ;
        RECT 2392.100 3273.530 2392.360 3273.850 ;
        RECT 2661.200 3273.530 2661.460 3273.850 ;
        RECT 2392.160 3260.000 2392.300 3273.530 ;
        RECT 2392.050 3256.000 2392.330 3260.000 ;
        RECT 2661.260 260.965 2661.400 3273.530 ;
        RECT 2393.930 260.595 2394.210 260.965 ;
        RECT 2661.190 260.595 2661.470 260.965 ;
        RECT 2394.000 18.010 2394.140 260.595 ;
        RECT 2387.500 17.690 2387.760 18.010 ;
        RECT 2393.940 17.690 2394.200 18.010 ;
        RECT 2387.560 2.400 2387.700 17.690 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
      LAYER via2 ;
        RECT 2393.930 260.640 2394.210 260.920 ;
        RECT 2661.190 260.640 2661.470 260.920 ;
      LAYER met3 ;
        RECT 2393.905 260.930 2394.235 260.945 ;
        RECT 2661.165 260.930 2661.495 260.945 ;
        RECT 2393.905 260.630 2661.495 260.930 ;
        RECT 2393.905 260.615 2394.235 260.630 ;
        RECT 2661.165 260.615 2661.495 260.630 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2456.085 7.565 2456.255 16.235 ;
        RECT 2463.905 15.895 2464.075 16.235 ;
        RECT 2463.445 15.725 2464.075 15.895 ;
        RECT 2504.845 15.045 2505.015 16.235 ;
        RECT 2552.685 15.045 2552.855 16.235 ;
      LAYER mcon ;
        RECT 2456.085 16.065 2456.255 16.235 ;
        RECT 2463.905 16.065 2464.075 16.235 ;
        RECT 2504.845 16.065 2505.015 16.235 ;
        RECT 2552.685 16.065 2552.855 16.235 ;
      LAYER met1 ;
        RECT 2306.510 3275.120 2306.830 3275.180 ;
        RECT 2635.870 3275.120 2636.190 3275.180 ;
        RECT 2306.510 3274.980 2636.190 3275.120 ;
        RECT 2306.510 3274.920 2306.830 3274.980 ;
        RECT 2635.870 3274.920 2636.190 3274.980 ;
        RECT 2456.025 16.220 2456.315 16.265 ;
        RECT 2463.845 16.220 2464.135 16.265 ;
        RECT 2504.785 16.220 2505.075 16.265 ;
        RECT 2456.025 16.080 2463.600 16.220 ;
        RECT 2456.025 16.035 2456.315 16.080 ;
        RECT 2463.460 15.925 2463.600 16.080 ;
        RECT 2463.845 16.080 2505.075 16.220 ;
        RECT 2463.845 16.035 2464.135 16.080 ;
        RECT 2504.785 16.035 2505.075 16.080 ;
        RECT 2552.625 16.220 2552.915 16.265 ;
        RECT 2559.970 16.220 2560.290 16.280 ;
        RECT 2552.625 16.080 2560.290 16.220 ;
        RECT 2552.625 16.035 2552.915 16.080 ;
        RECT 2559.970 16.020 2560.290 16.080 ;
        RECT 2560.890 16.220 2561.210 16.280 ;
        RECT 2635.870 16.220 2636.190 16.280 ;
        RECT 2560.890 16.080 2636.190 16.220 ;
        RECT 2560.890 16.020 2561.210 16.080 ;
        RECT 2635.870 16.020 2636.190 16.080 ;
        RECT 2463.385 15.695 2463.675 15.925 ;
        RECT 2504.785 15.200 2505.075 15.245 ;
        RECT 2552.625 15.200 2552.915 15.245 ;
        RECT 2504.785 15.060 2552.915 15.200 ;
        RECT 2504.785 15.015 2505.075 15.060 ;
        RECT 2552.625 15.015 2552.915 15.060 ;
        RECT 2405.410 7.720 2405.730 7.780 ;
        RECT 2456.025 7.720 2456.315 7.765 ;
        RECT 2405.410 7.580 2456.315 7.720 ;
        RECT 2405.410 7.520 2405.730 7.580 ;
        RECT 2456.025 7.535 2456.315 7.580 ;
      LAYER via ;
        RECT 2306.540 3274.920 2306.800 3275.180 ;
        RECT 2635.900 3274.920 2636.160 3275.180 ;
        RECT 2560.000 16.020 2560.260 16.280 ;
        RECT 2560.920 16.020 2561.180 16.280 ;
        RECT 2635.900 16.020 2636.160 16.280 ;
        RECT 2405.440 7.520 2405.700 7.780 ;
      LAYER met2 ;
        RECT 2306.540 3274.890 2306.800 3275.210 ;
        RECT 2635.900 3274.890 2636.160 3275.210 ;
        RECT 2306.600 3260.000 2306.740 3274.890 ;
        RECT 2306.490 3256.000 2306.770 3260.000 ;
        RECT 2635.960 16.310 2636.100 3274.890 ;
        RECT 2560.000 16.050 2560.260 16.310 ;
        RECT 2560.920 16.050 2561.180 16.310 ;
        RECT 2560.000 15.990 2561.180 16.050 ;
        RECT 2635.900 15.990 2636.160 16.310 ;
        RECT 2560.060 15.910 2561.120 15.990 ;
        RECT 2405.440 7.490 2405.700 7.810 ;
        RECT 2405.500 2.400 2405.640 7.490 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 3029.300 289.270 3029.360 ;
        RECT 296.770 3029.300 297.090 3029.360 ;
        RECT 288.950 3029.160 297.090 3029.300 ;
        RECT 288.950 3029.100 289.270 3029.160 ;
        RECT 296.770 3029.100 297.090 3029.160 ;
        RECT 288.950 204.240 289.270 204.300 ;
        RECT 793.570 204.240 793.890 204.300 ;
        RECT 288.950 204.100 793.890 204.240 ;
        RECT 288.950 204.040 289.270 204.100 ;
        RECT 793.570 204.040 793.890 204.100 ;
        RECT 793.570 49.200 793.890 49.260 ;
        RECT 799.550 49.200 799.870 49.260 ;
        RECT 793.570 49.060 799.870 49.200 ;
        RECT 793.570 49.000 793.890 49.060 ;
        RECT 799.550 49.000 799.870 49.060 ;
      LAYER via ;
        RECT 288.980 3029.100 289.240 3029.360 ;
        RECT 296.800 3029.100 297.060 3029.360 ;
        RECT 288.980 204.040 289.240 204.300 ;
        RECT 793.600 204.040 793.860 204.300 ;
        RECT 793.600 49.000 793.860 49.260 ;
        RECT 799.580 49.000 799.840 49.260 ;
      LAYER met2 ;
        RECT 296.790 3032.955 297.070 3033.325 ;
        RECT 296.860 3029.390 297.000 3032.955 ;
        RECT 288.980 3029.070 289.240 3029.390 ;
        RECT 296.800 3029.070 297.060 3029.390 ;
        RECT 289.040 204.330 289.180 3029.070 ;
        RECT 288.980 204.010 289.240 204.330 ;
        RECT 793.600 204.010 793.860 204.330 ;
        RECT 793.660 49.290 793.800 204.010 ;
        RECT 793.600 48.970 793.860 49.290 ;
        RECT 799.580 48.970 799.840 49.290 ;
        RECT 799.640 2.400 799.780 48.970 ;
        RECT 799.430 -4.800 799.990 2.400 ;
      LAYER via2 ;
        RECT 296.790 3033.000 297.070 3033.280 ;
      LAYER met3 ;
        RECT 296.765 3033.290 297.095 3033.305 ;
        RECT 310.000 3033.290 314.000 3033.680 ;
        RECT 296.765 3033.080 314.000 3033.290 ;
        RECT 296.765 3032.990 310.500 3033.080 ;
        RECT 296.765 3032.975 297.095 3032.990 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 641.845 145.265 642.015 234.515 ;
        RECT 641.845 89.845 642.015 137.955 ;
      LAYER mcon ;
        RECT 641.845 234.345 642.015 234.515 ;
        RECT 641.845 137.785 642.015 137.955 ;
      LAYER met1 ;
        RECT 288.030 2291.160 288.350 2291.220 ;
        RECT 296.770 2291.160 297.090 2291.220 ;
        RECT 288.030 2291.020 297.090 2291.160 ;
        RECT 288.030 2290.960 288.350 2291.020 ;
        RECT 296.770 2290.960 297.090 2291.020 ;
        RECT 288.030 247.080 288.350 247.140 ;
        RECT 642.230 247.080 642.550 247.140 ;
        RECT 288.030 246.940 642.550 247.080 ;
        RECT 288.030 246.880 288.350 246.940 ;
        RECT 642.230 246.880 642.550 246.940 ;
        RECT 641.770 234.500 642.090 234.560 ;
        RECT 641.575 234.360 642.090 234.500 ;
        RECT 641.770 234.300 642.090 234.360 ;
        RECT 641.770 145.420 642.090 145.480 ;
        RECT 641.575 145.280 642.090 145.420 ;
        RECT 641.770 145.220 642.090 145.280 ;
        RECT 641.770 137.940 642.090 138.000 ;
        RECT 641.575 137.800 642.090 137.940 ;
        RECT 641.770 137.740 642.090 137.800 ;
        RECT 641.770 90.000 642.090 90.060 ;
        RECT 641.575 89.860 642.090 90.000 ;
        RECT 641.770 89.800 642.090 89.860 ;
        RECT 642.690 57.360 643.010 57.420 ;
        RECT 644.990 57.360 645.310 57.420 ;
        RECT 642.690 57.220 645.310 57.360 ;
        RECT 642.690 57.160 643.010 57.220 ;
        RECT 644.990 57.160 645.310 57.220 ;
      LAYER via ;
        RECT 288.060 2290.960 288.320 2291.220 ;
        RECT 296.800 2290.960 297.060 2291.220 ;
        RECT 288.060 246.880 288.320 247.140 ;
        RECT 642.260 246.880 642.520 247.140 ;
        RECT 641.800 234.300 642.060 234.560 ;
        RECT 641.800 145.220 642.060 145.480 ;
        RECT 641.800 137.740 642.060 138.000 ;
        RECT 641.800 89.800 642.060 90.060 ;
        RECT 642.720 57.160 642.980 57.420 ;
        RECT 645.020 57.160 645.280 57.420 ;
      LAYER met2 ;
        RECT 296.790 2293.115 297.070 2293.485 ;
        RECT 296.860 2291.250 297.000 2293.115 ;
        RECT 288.060 2290.930 288.320 2291.250 ;
        RECT 296.800 2290.930 297.060 2291.250 ;
        RECT 288.120 247.170 288.260 2290.930 ;
        RECT 288.060 246.850 288.320 247.170 ;
        RECT 642.260 246.850 642.520 247.170 ;
        RECT 642.320 241.810 642.460 246.850 ;
        RECT 641.860 241.670 642.460 241.810 ;
        RECT 641.860 234.590 642.000 241.670 ;
        RECT 641.800 234.270 642.060 234.590 ;
        RECT 641.800 145.190 642.060 145.510 ;
        RECT 641.860 138.030 642.000 145.190 ;
        RECT 641.800 137.710 642.060 138.030 ;
        RECT 641.800 89.770 642.060 90.090 ;
        RECT 641.860 72.490 642.000 89.770 ;
        RECT 641.860 72.350 642.920 72.490 ;
        RECT 642.780 57.450 642.920 72.350 ;
        RECT 642.720 57.130 642.980 57.450 ;
        RECT 645.020 57.130 645.280 57.450 ;
        RECT 645.080 2.400 645.220 57.130 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 296.790 2293.160 297.070 2293.440 ;
      LAYER met3 ;
        RECT 296.765 2293.450 297.095 2293.465 ;
        RECT 310.000 2293.450 314.000 2293.840 ;
        RECT 296.765 2293.240 314.000 2293.450 ;
        RECT 296.765 2293.150 310.500 2293.240 ;
        RECT 296.765 2293.135 297.095 2293.150 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2597.160 2615.490 2597.220 ;
        RECT 2633.570 2597.160 2633.890 2597.220 ;
        RECT 2615.170 2597.020 2633.890 2597.160 ;
        RECT 2615.170 2596.960 2615.490 2597.020 ;
        RECT 2633.570 2596.960 2633.890 2597.020 ;
        RECT 2434.850 244.700 2435.170 244.760 ;
        RECT 2633.570 244.700 2633.890 244.760 ;
        RECT 2434.850 244.560 2633.890 244.700 ;
        RECT 2434.850 244.500 2435.170 244.560 ;
        RECT 2633.570 244.500 2633.890 244.560 ;
        RECT 2428.870 20.300 2429.190 20.360 ;
        RECT 2434.850 20.300 2435.170 20.360 ;
        RECT 2428.870 20.160 2435.170 20.300 ;
        RECT 2428.870 20.100 2429.190 20.160 ;
        RECT 2434.850 20.100 2435.170 20.160 ;
      LAYER via ;
        RECT 2615.200 2596.960 2615.460 2597.220 ;
        RECT 2633.600 2596.960 2633.860 2597.220 ;
        RECT 2434.880 244.500 2435.140 244.760 ;
        RECT 2633.600 244.500 2633.860 244.760 ;
        RECT 2428.900 20.100 2429.160 20.360 ;
        RECT 2434.880 20.100 2435.140 20.360 ;
      LAYER met2 ;
        RECT 2615.190 2600.475 2615.470 2600.845 ;
        RECT 2615.260 2597.250 2615.400 2600.475 ;
        RECT 2615.200 2596.930 2615.460 2597.250 ;
        RECT 2633.600 2596.930 2633.860 2597.250 ;
        RECT 2633.660 244.790 2633.800 2596.930 ;
        RECT 2434.880 244.470 2435.140 244.790 ;
        RECT 2633.600 244.470 2633.860 244.790 ;
        RECT 2434.940 20.390 2435.080 244.470 ;
        RECT 2428.900 20.070 2429.160 20.390 ;
        RECT 2434.880 20.070 2435.140 20.390 ;
        RECT 2428.960 2.400 2429.100 20.070 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2600.520 2615.470 2600.800 ;
      LAYER met3 ;
        RECT 2606.000 2600.810 2610.000 2601.200 ;
        RECT 2615.165 2600.810 2615.495 2600.825 ;
        RECT 2606.000 2600.600 2615.495 2600.810 ;
        RECT 2609.580 2600.510 2615.495 2600.600 ;
        RECT 2615.165 2600.495 2615.495 2600.510 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1320.290 3274.355 1320.570 3274.725 ;
        RECT 2650.610 3274.355 2650.890 3274.725 ;
        RECT 1320.360 3260.000 1320.500 3274.355 ;
        RECT 1320.250 3256.000 1320.530 3260.000 ;
        RECT 2650.680 16.165 2650.820 3274.355 ;
        RECT 2446.830 15.795 2447.110 16.165 ;
        RECT 2650.610 15.795 2650.890 16.165 ;
        RECT 2446.900 2.400 2447.040 15.795 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
      LAYER via2 ;
        RECT 1320.290 3274.400 1320.570 3274.680 ;
        RECT 2650.610 3274.400 2650.890 3274.680 ;
        RECT 2446.830 15.840 2447.110 16.120 ;
        RECT 2650.610 15.840 2650.890 16.120 ;
      LAYER met3 ;
        RECT 1320.265 3274.690 1320.595 3274.705 ;
        RECT 2650.585 3274.690 2650.915 3274.705 ;
        RECT 1320.265 3274.390 2650.915 3274.690 ;
        RECT 1320.265 3274.375 1320.595 3274.390 ;
        RECT 2650.585 3274.375 2650.915 3274.390 ;
        RECT 2446.805 16.130 2447.135 16.145 ;
        RECT 2650.585 16.130 2650.915 16.145 ;
        RECT 2446.805 15.830 2650.915 16.130 ;
        RECT 2446.805 15.815 2447.135 15.830 ;
        RECT 2650.585 15.815 2650.915 15.830 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1199.750 79.460 1200.070 79.520 ;
        RECT 2463.370 79.460 2463.690 79.520 ;
        RECT 1199.750 79.320 2463.690 79.460 ;
        RECT 1199.750 79.260 1200.070 79.320 ;
        RECT 2463.370 79.260 2463.690 79.320 ;
      LAYER via ;
        RECT 1199.780 79.260 1200.040 79.520 ;
        RECT 2463.400 79.260 2463.660 79.520 ;
      LAYER met2 ;
        RECT 1198.810 260.170 1199.090 264.000 ;
        RECT 1198.810 260.030 1199.980 260.170 ;
        RECT 1198.810 260.000 1199.090 260.030 ;
        RECT 1199.840 79.550 1199.980 260.030 ;
        RECT 1199.780 79.230 1200.040 79.550 ;
        RECT 2463.400 79.230 2463.660 79.550 ;
        RECT 2463.460 19.620 2463.600 79.230 ;
        RECT 2463.460 19.480 2464.520 19.620 ;
        RECT 2464.380 13.840 2464.520 19.480 ;
        RECT 2464.380 13.700 2464.980 13.840 ;
        RECT 2464.840 2.400 2464.980 13.700 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1270.590 244.020 1270.910 244.080 ;
        RECT 1276.110 244.020 1276.430 244.080 ;
        RECT 1270.590 243.880 1276.430 244.020 ;
        RECT 1270.590 243.820 1270.910 243.880 ;
        RECT 1276.110 243.820 1276.430 243.880 ;
        RECT 1276.110 162.760 1276.430 162.820 ;
        RECT 2477.170 162.760 2477.490 162.820 ;
        RECT 1276.110 162.620 2477.490 162.760 ;
        RECT 1276.110 162.560 1276.430 162.620 ;
        RECT 2477.170 162.560 2477.490 162.620 ;
        RECT 2477.170 37.640 2477.490 37.700 ;
        RECT 2482.690 37.640 2483.010 37.700 ;
        RECT 2477.170 37.500 2483.010 37.640 ;
        RECT 2477.170 37.440 2477.490 37.500 ;
        RECT 2482.690 37.440 2483.010 37.500 ;
      LAYER via ;
        RECT 1270.620 243.820 1270.880 244.080 ;
        RECT 1276.140 243.820 1276.400 244.080 ;
        RECT 1276.140 162.560 1276.400 162.820 ;
        RECT 2477.200 162.560 2477.460 162.820 ;
        RECT 2477.200 37.440 2477.460 37.700 ;
        RECT 2482.720 37.440 2482.980 37.700 ;
      LAYER met2 ;
        RECT 1270.570 260.000 1270.850 264.000 ;
        RECT 1270.680 244.110 1270.820 260.000 ;
        RECT 1270.620 243.790 1270.880 244.110 ;
        RECT 1276.140 243.790 1276.400 244.110 ;
        RECT 1276.200 162.850 1276.340 243.790 ;
        RECT 1276.140 162.530 1276.400 162.850 ;
        RECT 2477.200 162.530 2477.460 162.850 ;
        RECT 2477.260 37.730 2477.400 162.530 ;
        RECT 2477.200 37.410 2477.460 37.730 ;
        RECT 2482.720 37.410 2482.980 37.730 ;
        RECT 2482.780 2.400 2482.920 37.410 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2504.310 257.620 2504.630 257.680 ;
        RECT 2609.190 257.620 2609.510 257.680 ;
        RECT 2504.310 257.480 2609.510 257.620 ;
        RECT 2504.310 257.420 2504.630 257.480 ;
        RECT 2609.190 257.420 2609.510 257.480 ;
        RECT 2500.630 22.000 2500.950 22.060 ;
        RECT 2504.310 22.000 2504.630 22.060 ;
        RECT 2500.630 21.860 2504.630 22.000 ;
        RECT 2500.630 21.800 2500.950 21.860 ;
        RECT 2504.310 21.800 2504.630 21.860 ;
      LAYER via ;
        RECT 2504.340 257.420 2504.600 257.680 ;
        RECT 2609.220 257.420 2609.480 257.680 ;
        RECT 2500.660 21.800 2500.920 22.060 ;
        RECT 2504.340 21.800 2504.600 22.060 ;
      LAYER met2 ;
        RECT 2609.210 2070.075 2609.490 2070.445 ;
        RECT 2609.280 257.710 2609.420 2070.075 ;
        RECT 2504.340 257.390 2504.600 257.710 ;
        RECT 2609.220 257.390 2609.480 257.710 ;
        RECT 2504.400 22.090 2504.540 257.390 ;
        RECT 2500.660 21.770 2500.920 22.090 ;
        RECT 2504.340 21.770 2504.600 22.090 ;
        RECT 2500.720 2.400 2500.860 21.770 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
      LAYER via2 ;
        RECT 2609.210 2070.120 2609.490 2070.400 ;
      LAYER met3 ;
        RECT 2606.000 2071.560 2610.000 2072.160 ;
        RECT 2609.430 2070.425 2609.730 2071.560 ;
        RECT 2609.185 2070.110 2609.730 2070.425 ;
        RECT 2609.185 2070.095 2609.515 2070.110 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2518.130 217.075 2518.410 217.445 ;
        RECT 2518.200 2.400 2518.340 217.075 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
      LAYER via2 ;
        RECT 2518.130 217.120 2518.410 217.400 ;
      LAYER met3 ;
        RECT 2606.000 1670.360 2610.000 1670.960 ;
        RECT 2607.590 1667.860 2607.890 1670.360 ;
        RECT 2607.550 1667.540 2607.930 1667.860 ;
        RECT 2518.105 217.410 2518.435 217.425 ;
        RECT 2596.510 217.410 2596.890 217.420 ;
        RECT 2518.105 217.110 2596.890 217.410 ;
        RECT 2518.105 217.095 2518.435 217.110 ;
        RECT 2596.510 217.100 2596.890 217.110 ;
      LAYER via3 ;
        RECT 2607.580 1667.540 2607.900 1667.860 ;
        RECT 2596.540 217.100 2596.860 217.420 ;
      LAYER met4 ;
        RECT 2607.575 1667.535 2607.905 1667.865 ;
        RECT 2607.590 1647.450 2607.890 1667.535 ;
        RECT 2606.670 1647.150 2607.890 1647.450 ;
        RECT 2606.670 1637.690 2606.970 1647.150 ;
        RECT 2596.110 1636.510 2597.290 1637.690 ;
        RECT 2606.230 1636.510 2607.410 1637.690 ;
        RECT 2596.550 957.250 2596.850 1636.510 ;
        RECT 2595.630 956.950 2596.850 957.250 ;
        RECT 2595.630 913.050 2595.930 956.950 ;
        RECT 2595.630 912.750 2596.850 913.050 ;
        RECT 2596.550 732.850 2596.850 912.750 ;
        RECT 2592.870 732.550 2596.850 732.850 ;
        RECT 2592.870 705.650 2593.170 732.550 ;
        RECT 2592.870 705.350 2596.850 705.650 ;
        RECT 2596.550 566.250 2596.850 705.350 ;
        RECT 2595.630 565.950 2596.850 566.250 ;
        RECT 2595.630 556.050 2595.930 565.950 ;
        RECT 2595.630 555.750 2596.850 556.050 ;
        RECT 2596.550 515.250 2596.850 555.750 ;
        RECT 2595.630 514.950 2596.850 515.250 ;
        RECT 2595.630 501.650 2595.930 514.950 ;
        RECT 2595.630 501.350 2596.850 501.650 ;
        RECT 2596.550 484.650 2596.850 501.350 ;
        RECT 2596.550 484.350 2597.770 484.650 ;
        RECT 2597.470 477.850 2597.770 484.350 ;
        RECT 2596.550 477.550 2597.770 477.850 ;
        RECT 2596.550 217.425 2596.850 477.550 ;
        RECT 2596.535 217.095 2596.865 217.425 ;
      LAYER met5 ;
        RECT 2595.900 1636.300 2607.620 1637.900 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 399.810 93.060 400.130 93.120 ;
        RECT 2532.370 93.060 2532.690 93.120 ;
        RECT 399.810 92.920 2532.690 93.060 ;
        RECT 399.810 92.860 400.130 92.920 ;
        RECT 2532.370 92.860 2532.690 92.920 ;
        RECT 2532.370 14.180 2532.690 14.240 ;
        RECT 2532.370 14.040 2536.280 14.180 ;
        RECT 2532.370 13.980 2532.690 14.040 ;
        RECT 2536.140 13.900 2536.280 14.040 ;
        RECT 2536.050 13.640 2536.370 13.900 ;
      LAYER via ;
        RECT 399.840 92.860 400.100 93.120 ;
        RECT 2532.400 92.860 2532.660 93.120 ;
        RECT 2532.400 13.980 2532.660 14.240 ;
        RECT 2536.080 13.640 2536.340 13.900 ;
      LAYER met2 ;
        RECT 398.410 260.170 398.690 264.000 ;
        RECT 398.410 260.030 400.040 260.170 ;
        RECT 398.410 260.000 398.690 260.030 ;
        RECT 399.900 93.150 400.040 260.030 ;
        RECT 399.840 92.830 400.100 93.150 ;
        RECT 2532.400 92.830 2532.660 93.150 ;
        RECT 2532.460 14.270 2532.600 92.830 ;
        RECT 2532.400 13.950 2532.660 14.270 ;
        RECT 2536.080 13.610 2536.340 13.930 ;
        RECT 2536.140 2.400 2536.280 13.610 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.110 33.560 1414.430 33.620 ;
        RECT 2553.990 33.560 2554.310 33.620 ;
        RECT 1414.110 33.420 2554.310 33.560 ;
        RECT 1414.110 33.360 1414.430 33.420 ;
        RECT 2553.990 33.360 2554.310 33.420 ;
      LAYER via ;
        RECT 1414.140 33.360 1414.400 33.620 ;
        RECT 2554.020 33.360 2554.280 33.620 ;
      LAYER met2 ;
        RECT 1413.170 260.170 1413.450 264.000 ;
        RECT 1413.170 260.030 1414.340 260.170 ;
        RECT 1413.170 260.000 1413.450 260.030 ;
        RECT 1414.200 33.650 1414.340 260.030 ;
        RECT 1414.140 33.330 1414.400 33.650 ;
        RECT 2554.020 33.330 2554.280 33.650 ;
        RECT 2554.080 2.400 2554.220 33.330 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2607.350 1858.000 2607.670 1858.060 ;
        RECT 2617.010 1858.000 2617.330 1858.060 ;
        RECT 2607.350 1857.860 2617.330 1858.000 ;
        RECT 2607.350 1857.800 2607.670 1857.860 ;
        RECT 2617.010 1857.800 2617.330 1857.860 ;
        RECT 2571.930 20.640 2572.250 20.700 ;
        RECT 2607.350 20.640 2607.670 20.700 ;
        RECT 2571.930 20.500 2607.670 20.640 ;
        RECT 2571.930 20.440 2572.250 20.500 ;
        RECT 2607.350 20.440 2607.670 20.500 ;
      LAYER via ;
        RECT 2607.380 1857.800 2607.640 1858.060 ;
        RECT 2617.040 1857.800 2617.300 1858.060 ;
        RECT 2571.960 20.440 2572.220 20.700 ;
        RECT 2607.380 20.440 2607.640 20.700 ;
      LAYER met2 ;
        RECT 2617.030 2726.955 2617.310 2727.325 ;
        RECT 2617.100 1858.090 2617.240 2726.955 ;
        RECT 2607.380 1857.770 2607.640 1858.090 ;
        RECT 2617.040 1857.770 2617.300 1858.090 ;
        RECT 2607.440 20.730 2607.580 1857.770 ;
        RECT 2571.960 20.410 2572.220 20.730 ;
        RECT 2607.380 20.410 2607.640 20.730 ;
        RECT 2572.020 2.400 2572.160 20.410 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
      LAYER via2 ;
        RECT 2617.030 2727.000 2617.310 2727.280 ;
      LAYER met3 ;
        RECT 2606.000 2727.290 2610.000 2727.680 ;
        RECT 2617.005 2727.290 2617.335 2727.305 ;
        RECT 2606.000 2727.080 2617.335 2727.290 ;
        RECT 2609.580 2726.990 2617.335 2727.080 ;
        RECT 2617.005 2726.975 2617.335 2726.990 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1192.850 3258.460 1193.170 3258.520 ;
        RECT 2691.070 3258.460 2691.390 3258.520 ;
        RECT 1192.850 3258.320 2691.390 3258.460 ;
        RECT 1192.850 3258.260 1193.170 3258.320 ;
        RECT 2691.070 3258.260 2691.390 3258.320 ;
        RECT 2589.410 19.960 2589.730 20.020 ;
        RECT 2691.070 19.960 2691.390 20.020 ;
        RECT 2589.410 19.820 2691.390 19.960 ;
        RECT 2589.410 19.760 2589.730 19.820 ;
        RECT 2691.070 19.760 2691.390 19.820 ;
      LAYER via ;
        RECT 1192.880 3258.260 1193.140 3258.520 ;
        RECT 2691.100 3258.260 2691.360 3258.520 ;
        RECT 2589.440 19.760 2589.700 20.020 ;
        RECT 2691.100 19.760 2691.360 20.020 ;
      LAYER met2 ;
        RECT 1191.450 3258.290 1191.730 3260.000 ;
        RECT 1192.880 3258.290 1193.140 3258.550 ;
        RECT 1191.450 3258.230 1193.140 3258.290 ;
        RECT 2691.100 3258.230 2691.360 3258.550 ;
        RECT 1191.450 3258.150 1193.080 3258.230 ;
        RECT 1191.450 3256.000 1191.730 3258.150 ;
        RECT 2691.160 20.050 2691.300 3258.230 ;
        RECT 2589.440 19.730 2589.700 20.050 ;
        RECT 2691.100 19.730 2691.360 20.050 ;
        RECT 2589.500 2.400 2589.640 19.730 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 211.380 827.930 211.440 ;
        RECT 2630.810 211.380 2631.130 211.440 ;
        RECT 827.610 211.240 2631.130 211.380 ;
        RECT 827.610 211.180 827.930 211.240 ;
        RECT 2630.810 211.180 2631.130 211.240 ;
        RECT 823.470 14.520 823.790 14.580 ;
        RECT 827.610 14.520 827.930 14.580 ;
        RECT 823.470 14.380 827.930 14.520 ;
        RECT 823.470 14.320 823.790 14.380 ;
        RECT 827.610 14.320 827.930 14.380 ;
      LAYER via ;
        RECT 827.640 211.180 827.900 211.440 ;
        RECT 2630.840 211.180 2631.100 211.440 ;
        RECT 823.500 14.320 823.760 14.580 ;
        RECT 827.640 14.320 827.900 14.580 ;
      LAYER met2 ;
        RECT 2630.830 2303.995 2631.110 2304.365 ;
        RECT 2630.900 211.470 2631.040 2303.995 ;
        RECT 827.640 211.150 827.900 211.470 ;
        RECT 2630.840 211.150 2631.100 211.470 ;
        RECT 827.700 14.610 827.840 211.150 ;
        RECT 823.500 14.290 823.760 14.610 ;
        RECT 827.640 14.290 827.900 14.610 ;
        RECT 823.560 2.400 823.700 14.290 ;
        RECT 823.350 -4.800 823.910 2.400 ;
      LAYER via2 ;
        RECT 2630.830 2304.040 2631.110 2304.320 ;
      LAYER met3 ;
        RECT 2606.000 2304.330 2610.000 2304.720 ;
        RECT 2630.805 2304.330 2631.135 2304.345 ;
        RECT 2606.000 2304.120 2631.135 2304.330 ;
        RECT 2609.580 2304.030 2631.135 2304.120 ;
        RECT 2630.805 2304.015 2631.135 2304.030 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1205.290 3272.995 1205.570 3273.365 ;
        RECT 1205.360 3260.000 1205.500 3272.995 ;
        RECT 1205.250 3256.000 1205.530 3260.000 ;
        RECT 2607.370 16.475 2607.650 16.845 ;
        RECT 2607.440 2.400 2607.580 16.475 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
      LAYER via2 ;
        RECT 1205.290 3273.040 1205.570 3273.320 ;
        RECT 2607.370 16.520 2607.650 16.800 ;
      LAYER met3 ;
        RECT 1205.265 3273.330 1205.595 3273.345 ;
        RECT 2691.270 3273.330 2691.650 3273.340 ;
        RECT 1205.265 3273.030 2691.650 3273.330 ;
        RECT 1205.265 3273.015 1205.595 3273.030 ;
        RECT 2691.270 3273.020 2691.650 3273.030 ;
        RECT 2607.345 16.810 2607.675 16.825 ;
        RECT 2691.270 16.810 2691.650 16.820 ;
        RECT 2607.345 16.510 2691.650 16.810 ;
        RECT 2607.345 16.495 2607.675 16.510 ;
        RECT 2691.270 16.500 2691.650 16.510 ;
      LAYER via3 ;
        RECT 2691.300 3273.020 2691.620 3273.340 ;
        RECT 2691.300 16.500 2691.620 16.820 ;
      LAYER met4 ;
        RECT 2691.295 3273.015 2691.625 3273.345 ;
        RECT 2691.310 16.825 2691.610 3273.015 ;
        RECT 2691.295 16.495 2691.625 16.825 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1835.010 3259.820 1835.330 3259.880 ;
        RECT 2684.630 3259.820 2684.950 3259.880 ;
        RECT 1835.010 3259.680 2684.950 3259.820 ;
        RECT 1835.010 3259.620 1835.330 3259.680 ;
        RECT 2684.630 3259.620 2684.950 3259.680 ;
        RECT 2625.290 19.280 2625.610 19.340 ;
        RECT 2684.170 19.280 2684.490 19.340 ;
        RECT 2625.290 19.140 2684.490 19.280 ;
        RECT 2625.290 19.080 2625.610 19.140 ;
        RECT 2684.170 19.080 2684.490 19.140 ;
      LAYER via ;
        RECT 1835.040 3259.620 1835.300 3259.880 ;
        RECT 2684.660 3259.620 2684.920 3259.880 ;
        RECT 2625.320 19.080 2625.580 19.340 ;
        RECT 2684.200 19.080 2684.460 19.340 ;
      LAYER met2 ;
        RECT 1834.530 3259.650 1834.810 3260.000 ;
        RECT 1835.040 3259.650 1835.300 3259.910 ;
        RECT 1834.530 3259.590 1835.300 3259.650 ;
        RECT 2684.660 3259.590 2684.920 3259.910 ;
        RECT 1834.530 3259.510 1835.240 3259.590 ;
        RECT 1834.530 3256.000 1834.810 3259.510 ;
        RECT 2684.720 36.450 2684.860 3259.590 ;
        RECT 2684.260 36.310 2684.860 36.450 ;
        RECT 2684.260 19.370 2684.400 36.310 ;
        RECT 2625.320 19.050 2625.580 19.370 ;
        RECT 2684.200 19.050 2684.460 19.370 ;
        RECT 2625.380 2.400 2625.520 19.050 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2000.150 148.820 2000.470 148.880 ;
        RECT 2625.290 148.820 2625.610 148.880 ;
        RECT 2000.150 148.680 2625.610 148.820 ;
        RECT 2000.150 148.620 2000.470 148.680 ;
        RECT 2625.290 148.620 2625.610 148.680 ;
        RECT 2625.290 20.640 2625.610 20.700 ;
        RECT 2643.230 20.640 2643.550 20.700 ;
        RECT 2625.290 20.500 2643.550 20.640 ;
        RECT 2625.290 20.440 2625.610 20.500 ;
        RECT 2643.230 20.440 2643.550 20.500 ;
      LAYER via ;
        RECT 2000.180 148.620 2000.440 148.880 ;
        RECT 2625.320 148.620 2625.580 148.880 ;
        RECT 2625.320 20.440 2625.580 20.700 ;
        RECT 2643.260 20.440 2643.520 20.700 ;
      LAYER met2 ;
        RECT 2000.130 260.000 2000.410 264.000 ;
        RECT 2000.240 148.910 2000.380 260.000 ;
        RECT 2000.180 148.590 2000.440 148.910 ;
        RECT 2625.320 148.590 2625.580 148.910 ;
        RECT 2625.380 20.730 2625.520 148.590 ;
        RECT 2625.320 20.410 2625.580 20.730 ;
        RECT 2643.260 20.410 2643.520 20.730 ;
        RECT 2643.320 2.400 2643.460 20.410 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1470.230 244.020 1470.550 244.080 ;
        RECT 1476.210 244.020 1476.530 244.080 ;
        RECT 1470.230 243.880 1476.530 244.020 ;
        RECT 1470.230 243.820 1470.550 243.880 ;
        RECT 1476.210 243.820 1476.530 243.880 ;
        RECT 1476.210 169.560 1476.530 169.620 ;
        RECT 2657.030 169.560 2657.350 169.620 ;
        RECT 1476.210 169.420 2657.350 169.560 ;
        RECT 1476.210 169.360 1476.530 169.420 ;
        RECT 2657.030 169.360 2657.350 169.420 ;
        RECT 2657.030 62.120 2657.350 62.180 ;
        RECT 2661.170 62.120 2661.490 62.180 ;
        RECT 2657.030 61.980 2661.490 62.120 ;
        RECT 2657.030 61.920 2657.350 61.980 ;
        RECT 2661.170 61.920 2661.490 61.980 ;
      LAYER via ;
        RECT 1470.260 243.820 1470.520 244.080 ;
        RECT 1476.240 243.820 1476.500 244.080 ;
        RECT 1476.240 169.360 1476.500 169.620 ;
        RECT 2657.060 169.360 2657.320 169.620 ;
        RECT 2657.060 61.920 2657.320 62.180 ;
        RECT 2661.200 61.920 2661.460 62.180 ;
      LAYER met2 ;
        RECT 1470.210 260.000 1470.490 264.000 ;
        RECT 1470.320 244.110 1470.460 260.000 ;
        RECT 1470.260 243.790 1470.520 244.110 ;
        RECT 1476.240 243.790 1476.500 244.110 ;
        RECT 1476.300 169.650 1476.440 243.790 ;
        RECT 1476.240 169.330 1476.500 169.650 ;
        RECT 2657.060 169.330 2657.320 169.650 ;
        RECT 2657.120 62.210 2657.260 169.330 ;
        RECT 2657.060 61.890 2657.320 62.210 ;
        RECT 2661.200 61.890 2661.460 62.210 ;
        RECT 2661.260 2.400 2661.400 61.890 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2677.345 48.365 2677.515 96.475 ;
      LAYER mcon ;
        RECT 2677.345 96.305 2677.515 96.475 ;
      LAYER met1 ;
        RECT 2676.350 144.740 2676.670 144.800 ;
        RECT 2677.270 144.740 2677.590 144.800 ;
        RECT 2676.350 144.600 2677.590 144.740 ;
        RECT 2676.350 144.540 2676.670 144.600 ;
        RECT 2677.270 144.540 2677.590 144.600 ;
        RECT 2677.270 96.460 2677.590 96.520 ;
        RECT 2677.075 96.320 2677.590 96.460 ;
        RECT 2677.270 96.260 2677.590 96.320 ;
        RECT 2677.270 48.520 2677.590 48.580 ;
        RECT 2677.075 48.380 2677.590 48.520 ;
        RECT 2677.270 48.320 2677.590 48.380 ;
        RECT 2677.270 14.180 2677.590 14.240 ;
        RECT 2677.270 14.040 2678.880 14.180 ;
        RECT 2677.270 13.980 2677.590 14.040 ;
        RECT 2678.740 13.900 2678.880 14.040 ;
        RECT 2678.650 13.640 2678.970 13.900 ;
      LAYER via ;
        RECT 2676.380 144.540 2676.640 144.800 ;
        RECT 2677.300 144.540 2677.560 144.800 ;
        RECT 2677.300 96.260 2677.560 96.520 ;
        RECT 2677.300 48.320 2677.560 48.580 ;
        RECT 2677.300 13.980 2677.560 14.240 ;
        RECT 2678.680 13.640 2678.940 13.900 ;
      LAYER met2 ;
        RECT 2677.290 202.795 2677.570 203.165 ;
        RECT 2677.360 144.830 2677.500 202.795 ;
        RECT 2676.380 144.510 2676.640 144.830 ;
        RECT 2677.300 144.510 2677.560 144.830 ;
        RECT 2676.440 97.085 2676.580 144.510 ;
        RECT 2676.370 96.715 2676.650 97.085 ;
        RECT 2677.290 96.715 2677.570 97.085 ;
        RECT 2677.360 96.550 2677.500 96.715 ;
        RECT 2677.300 96.230 2677.560 96.550 ;
        RECT 2677.300 48.290 2677.560 48.610 ;
        RECT 2677.360 14.270 2677.500 48.290 ;
        RECT 2677.300 13.950 2677.560 14.270 ;
        RECT 2678.680 13.610 2678.940 13.930 ;
        RECT 2678.740 2.400 2678.880 13.610 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
      LAYER via2 ;
        RECT 2677.290 202.840 2677.570 203.120 ;
        RECT 2676.370 96.760 2676.650 97.040 ;
        RECT 2677.290 96.760 2677.570 97.040 ;
      LAYER met3 ;
        RECT 287.310 2694.650 287.690 2694.660 ;
        RECT 310.000 2694.650 314.000 2695.040 ;
        RECT 287.310 2694.440 314.000 2694.650 ;
        RECT 287.310 2694.350 310.500 2694.440 ;
        RECT 287.310 2694.340 287.690 2694.350 ;
        RECT 287.310 203.130 287.690 203.140 ;
        RECT 2677.265 203.130 2677.595 203.145 ;
        RECT 287.310 202.830 2677.595 203.130 ;
        RECT 287.310 202.820 287.690 202.830 ;
        RECT 2677.265 202.815 2677.595 202.830 ;
        RECT 2676.345 97.050 2676.675 97.065 ;
        RECT 2677.265 97.050 2677.595 97.065 ;
        RECT 2676.345 96.750 2677.595 97.050 ;
        RECT 2676.345 96.735 2676.675 96.750 ;
        RECT 2677.265 96.735 2677.595 96.750 ;
      LAYER via3 ;
        RECT 287.340 2694.340 287.660 2694.660 ;
        RECT 287.340 202.820 287.660 203.140 ;
      LAYER met4 ;
        RECT 287.335 2694.335 287.665 2694.665 ;
        RECT 287.350 203.145 287.650 2694.335 ;
        RECT 287.335 202.815 287.665 203.145 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 302.750 58.720 303.070 58.780 ;
        RECT 2696.590 58.720 2696.910 58.780 ;
        RECT 302.750 58.580 2696.910 58.720 ;
        RECT 302.750 58.520 303.070 58.580 ;
        RECT 2696.590 58.520 2696.910 58.580 ;
      LAYER via ;
        RECT 302.780 58.520 303.040 58.780 ;
        RECT 2696.620 58.520 2696.880 58.780 ;
      LAYER met2 ;
        RECT 302.770 432.635 303.050 433.005 ;
        RECT 302.840 58.810 302.980 432.635 ;
        RECT 302.780 58.490 303.040 58.810 ;
        RECT 2696.620 58.490 2696.880 58.810 ;
        RECT 2696.680 2.400 2696.820 58.490 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 302.770 432.680 303.050 432.960 ;
      LAYER met3 ;
        RECT 302.745 432.970 303.075 432.985 ;
        RECT 310.000 432.970 314.000 433.360 ;
        RECT 302.745 432.760 314.000 432.970 ;
        RECT 302.745 432.670 310.500 432.760 ;
        RECT 302.745 432.655 303.075 432.670 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2711.845 3181.125 2712.015 3229.235 ;
        RECT 2711.845 3084.225 2712.015 3132.675 ;
        RECT 2711.845 2408.305 2712.015 2456.415 ;
        RECT 2711.845 2311.745 2712.015 2359.855 ;
        RECT 2711.845 2214.845 2712.015 2262.955 ;
        RECT 2711.845 2118.285 2712.015 2166.395 ;
        RECT 2711.845 2021.725 2712.015 2069.835 ;
        RECT 2711.845 1925.165 2712.015 1973.275 ;
        RECT 2711.845 1828.605 2712.015 1876.715 ;
        RECT 2711.845 1732.045 2712.015 1780.155 ;
        RECT 2711.845 1635.825 2712.015 1683.595 ;
        RECT 2711.845 1490.985 2712.015 1538.755 ;
        RECT 2712.305 1007.505 2712.475 1055.615 ;
        RECT 2712.305 910.945 2712.475 959.055 ;
        RECT 2711.845 766.105 2712.015 814.215 ;
        RECT 2711.385 717.825 2711.555 765.595 ;
        RECT 2711.845 669.545 2712.015 717.655 ;
        RECT 2711.845 572.985 2712.015 620.755 ;
        RECT 2711.845 476.425 2712.015 524.195 ;
        RECT 2711.845 379.865 2712.015 427.635 ;
        RECT 2711.845 283.305 2712.015 331.075 ;
        RECT 2711.845 186.745 2712.015 234.515 ;
        RECT 2711.845 138.465 2712.015 186.235 ;
        RECT 2711.845 90.185 2712.015 137.955 ;
        RECT 2711.845 41.905 2712.015 89.675 ;
        RECT 2714.605 2.805 2714.775 41.395 ;
      LAYER mcon ;
        RECT 2711.845 3229.065 2712.015 3229.235 ;
        RECT 2711.845 3132.505 2712.015 3132.675 ;
        RECT 2711.845 2456.245 2712.015 2456.415 ;
        RECT 2711.845 2359.685 2712.015 2359.855 ;
        RECT 2711.845 2262.785 2712.015 2262.955 ;
        RECT 2711.845 2166.225 2712.015 2166.395 ;
        RECT 2711.845 2069.665 2712.015 2069.835 ;
        RECT 2711.845 1973.105 2712.015 1973.275 ;
        RECT 2711.845 1876.545 2712.015 1876.715 ;
        RECT 2711.845 1779.985 2712.015 1780.155 ;
        RECT 2711.845 1683.425 2712.015 1683.595 ;
        RECT 2711.845 1538.585 2712.015 1538.755 ;
        RECT 2712.305 1055.445 2712.475 1055.615 ;
        RECT 2712.305 958.885 2712.475 959.055 ;
        RECT 2711.845 814.045 2712.015 814.215 ;
        RECT 2711.385 765.425 2711.555 765.595 ;
        RECT 2711.845 717.485 2712.015 717.655 ;
        RECT 2711.845 620.585 2712.015 620.755 ;
        RECT 2711.845 524.025 2712.015 524.195 ;
        RECT 2711.845 427.465 2712.015 427.635 ;
        RECT 2711.845 330.905 2712.015 331.075 ;
        RECT 2711.845 234.345 2712.015 234.515 ;
        RECT 2711.845 186.065 2712.015 186.235 ;
        RECT 2711.845 137.785 2712.015 137.955 ;
        RECT 2711.845 89.505 2712.015 89.675 ;
        RECT 2714.605 41.225 2714.775 41.395 ;
      LAYER met1 ;
        RECT 2711.770 3229.220 2712.090 3229.280 ;
        RECT 2711.575 3229.080 2712.090 3229.220 ;
        RECT 2711.770 3229.020 2712.090 3229.080 ;
        RECT 2711.770 3181.280 2712.090 3181.340 ;
        RECT 2711.575 3181.140 2712.090 3181.280 ;
        RECT 2711.770 3181.080 2712.090 3181.140 ;
        RECT 2711.770 3132.660 2712.090 3132.720 ;
        RECT 2711.575 3132.520 2712.090 3132.660 ;
        RECT 2711.770 3132.460 2712.090 3132.520 ;
        RECT 2711.770 3084.380 2712.090 3084.440 ;
        RECT 2711.575 3084.240 2712.090 3084.380 ;
        RECT 2711.770 3084.180 2712.090 3084.240 ;
        RECT 2710.850 2987.820 2711.170 2987.880 ;
        RECT 2711.770 2987.820 2712.090 2987.880 ;
        RECT 2710.850 2987.680 2712.090 2987.820 ;
        RECT 2710.850 2987.620 2711.170 2987.680 ;
        RECT 2711.770 2987.620 2712.090 2987.680 ;
        RECT 2710.850 2891.260 2711.170 2891.320 ;
        RECT 2711.770 2891.260 2712.090 2891.320 ;
        RECT 2710.850 2891.120 2712.090 2891.260 ;
        RECT 2710.850 2891.060 2711.170 2891.120 ;
        RECT 2711.770 2891.060 2712.090 2891.120 ;
        RECT 2710.850 2794.700 2711.170 2794.760 ;
        RECT 2711.770 2794.700 2712.090 2794.760 ;
        RECT 2710.850 2794.560 2712.090 2794.700 ;
        RECT 2710.850 2794.500 2711.170 2794.560 ;
        RECT 2711.770 2794.500 2712.090 2794.560 ;
        RECT 2710.850 2649.520 2711.170 2649.580 ;
        RECT 2711.770 2649.520 2712.090 2649.580 ;
        RECT 2710.850 2649.380 2712.090 2649.520 ;
        RECT 2710.850 2649.320 2711.170 2649.380 ;
        RECT 2711.770 2649.320 2712.090 2649.380 ;
        RECT 2710.850 2552.960 2711.170 2553.020 ;
        RECT 2711.770 2552.960 2712.090 2553.020 ;
        RECT 2710.850 2552.820 2712.090 2552.960 ;
        RECT 2710.850 2552.760 2711.170 2552.820 ;
        RECT 2711.770 2552.760 2712.090 2552.820 ;
        RECT 2711.770 2456.400 2712.090 2456.460 ;
        RECT 2711.575 2456.260 2712.090 2456.400 ;
        RECT 2711.770 2456.200 2712.090 2456.260 ;
        RECT 2711.770 2408.460 2712.090 2408.520 ;
        RECT 2711.575 2408.320 2712.090 2408.460 ;
        RECT 2711.770 2408.260 2712.090 2408.320 ;
        RECT 2711.770 2359.840 2712.090 2359.900 ;
        RECT 2711.575 2359.700 2712.090 2359.840 ;
        RECT 2711.770 2359.640 2712.090 2359.700 ;
        RECT 2711.770 2311.900 2712.090 2311.960 ;
        RECT 2711.575 2311.760 2712.090 2311.900 ;
        RECT 2711.770 2311.700 2712.090 2311.760 ;
        RECT 2711.770 2262.940 2712.090 2263.000 ;
        RECT 2711.575 2262.800 2712.090 2262.940 ;
        RECT 2711.770 2262.740 2712.090 2262.800 ;
        RECT 2711.770 2215.000 2712.090 2215.060 ;
        RECT 2711.575 2214.860 2712.090 2215.000 ;
        RECT 2711.770 2214.800 2712.090 2214.860 ;
        RECT 2711.770 2166.380 2712.090 2166.440 ;
        RECT 2711.575 2166.240 2712.090 2166.380 ;
        RECT 2711.770 2166.180 2712.090 2166.240 ;
        RECT 2711.770 2118.440 2712.090 2118.500 ;
        RECT 2711.575 2118.300 2712.090 2118.440 ;
        RECT 2711.770 2118.240 2712.090 2118.300 ;
        RECT 2711.770 2069.820 2712.090 2069.880 ;
        RECT 2711.575 2069.680 2712.090 2069.820 ;
        RECT 2711.770 2069.620 2712.090 2069.680 ;
        RECT 2711.770 2021.880 2712.090 2021.940 ;
        RECT 2711.575 2021.740 2712.090 2021.880 ;
        RECT 2711.770 2021.680 2712.090 2021.740 ;
        RECT 2711.770 1973.260 2712.090 1973.320 ;
        RECT 2711.575 1973.120 2712.090 1973.260 ;
        RECT 2711.770 1973.060 2712.090 1973.120 ;
        RECT 2711.770 1925.320 2712.090 1925.380 ;
        RECT 2711.575 1925.180 2712.090 1925.320 ;
        RECT 2711.770 1925.120 2712.090 1925.180 ;
        RECT 2711.770 1876.700 2712.090 1876.760 ;
        RECT 2711.575 1876.560 2712.090 1876.700 ;
        RECT 2711.770 1876.500 2712.090 1876.560 ;
        RECT 2711.770 1828.760 2712.090 1828.820 ;
        RECT 2711.575 1828.620 2712.090 1828.760 ;
        RECT 2711.770 1828.560 2712.090 1828.620 ;
        RECT 2711.770 1780.140 2712.090 1780.200 ;
        RECT 2711.575 1780.000 2712.090 1780.140 ;
        RECT 2711.770 1779.940 2712.090 1780.000 ;
        RECT 2711.770 1732.200 2712.090 1732.260 ;
        RECT 2711.575 1732.060 2712.090 1732.200 ;
        RECT 2711.770 1732.000 2712.090 1732.060 ;
        RECT 2711.770 1691.540 2712.090 1691.800 ;
        RECT 2711.860 1690.780 2712.000 1691.540 ;
        RECT 2711.770 1690.520 2712.090 1690.780 ;
        RECT 2711.770 1683.580 2712.090 1683.640 ;
        RECT 2711.575 1683.440 2712.090 1683.580 ;
        RECT 2711.770 1683.380 2712.090 1683.440 ;
        RECT 2711.310 1635.980 2711.630 1636.040 ;
        RECT 2711.785 1635.980 2712.075 1636.025 ;
        RECT 2711.310 1635.840 2712.075 1635.980 ;
        RECT 2711.310 1635.780 2711.630 1635.840 ;
        RECT 2711.785 1635.795 2712.075 1635.840 ;
        RECT 2711.770 1538.740 2712.090 1538.800 ;
        RECT 2711.575 1538.600 2712.090 1538.740 ;
        RECT 2711.770 1538.540 2712.090 1538.600 ;
        RECT 2711.770 1491.140 2712.090 1491.200 ;
        RECT 2711.575 1491.000 2712.090 1491.140 ;
        RECT 2711.770 1490.940 2712.090 1491.000 ;
        RECT 2711.770 1490.460 2712.090 1490.520 ;
        RECT 2713.150 1490.460 2713.470 1490.520 ;
        RECT 2711.770 1490.320 2713.470 1490.460 ;
        RECT 2711.770 1490.260 2712.090 1490.320 ;
        RECT 2713.150 1490.260 2713.470 1490.320 ;
        RECT 2710.850 1393.900 2711.170 1393.960 ;
        RECT 2711.770 1393.900 2712.090 1393.960 ;
        RECT 2710.850 1393.760 2712.090 1393.900 ;
        RECT 2710.850 1393.700 2711.170 1393.760 ;
        RECT 2711.770 1393.700 2712.090 1393.760 ;
        RECT 2710.850 1346.300 2711.170 1346.360 ;
        RECT 2711.770 1346.300 2712.090 1346.360 ;
        RECT 2710.850 1346.160 2712.090 1346.300 ;
        RECT 2710.850 1346.100 2711.170 1346.160 ;
        RECT 2711.770 1346.100 2712.090 1346.160 ;
        RECT 2710.850 1297.340 2711.170 1297.400 ;
        RECT 2711.770 1297.340 2712.090 1297.400 ;
        RECT 2710.850 1297.200 2712.090 1297.340 ;
        RECT 2710.850 1297.140 2711.170 1297.200 ;
        RECT 2711.770 1297.140 2712.090 1297.200 ;
        RECT 2710.850 1249.740 2711.170 1249.800 ;
        RECT 2711.770 1249.740 2712.090 1249.800 ;
        RECT 2710.850 1249.600 2712.090 1249.740 ;
        RECT 2710.850 1249.540 2711.170 1249.600 ;
        RECT 2711.770 1249.540 2712.090 1249.600 ;
        RECT 2710.850 1200.780 2711.170 1200.840 ;
        RECT 2711.770 1200.780 2712.090 1200.840 ;
        RECT 2710.850 1200.640 2712.090 1200.780 ;
        RECT 2710.850 1200.580 2711.170 1200.640 ;
        RECT 2711.770 1200.580 2712.090 1200.640 ;
        RECT 2710.850 1104.220 2711.170 1104.280 ;
        RECT 2711.770 1104.220 2712.090 1104.280 ;
        RECT 2710.850 1104.080 2712.090 1104.220 ;
        RECT 2710.850 1104.020 2711.170 1104.080 ;
        RECT 2711.770 1104.020 2712.090 1104.080 ;
        RECT 2712.230 1055.600 2712.550 1055.660 ;
        RECT 2712.035 1055.460 2712.550 1055.600 ;
        RECT 2712.230 1055.400 2712.550 1055.460 ;
        RECT 2711.310 1007.660 2711.630 1007.720 ;
        RECT 2712.245 1007.660 2712.535 1007.705 ;
        RECT 2711.310 1007.520 2712.535 1007.660 ;
        RECT 2711.310 1007.460 2711.630 1007.520 ;
        RECT 2712.245 1007.475 2712.535 1007.520 ;
        RECT 2711.770 1007.320 2712.090 1007.380 ;
        RECT 2713.150 1007.320 2713.470 1007.380 ;
        RECT 2711.770 1007.180 2713.470 1007.320 ;
        RECT 2711.770 1007.120 2712.090 1007.180 ;
        RECT 2713.150 1007.120 2713.470 1007.180 ;
        RECT 2712.230 959.040 2712.550 959.100 ;
        RECT 2712.035 958.900 2712.550 959.040 ;
        RECT 2712.230 958.840 2712.550 958.900 ;
        RECT 2711.310 911.100 2711.630 911.160 ;
        RECT 2712.245 911.100 2712.535 911.145 ;
        RECT 2711.310 910.960 2712.535 911.100 ;
        RECT 2711.310 910.900 2711.630 910.960 ;
        RECT 2712.245 910.915 2712.535 910.960 ;
        RECT 2711.770 910.760 2712.090 910.820 ;
        RECT 2713.150 910.760 2713.470 910.820 ;
        RECT 2711.770 910.620 2713.470 910.760 ;
        RECT 2711.770 910.560 2712.090 910.620 ;
        RECT 2713.150 910.560 2713.470 910.620 ;
        RECT 2710.850 862.480 2711.170 862.540 ;
        RECT 2712.230 862.480 2712.550 862.540 ;
        RECT 2710.850 862.340 2712.550 862.480 ;
        RECT 2710.850 862.280 2711.170 862.340 ;
        RECT 2712.230 862.280 2712.550 862.340 ;
        RECT 2711.770 814.200 2712.090 814.260 ;
        RECT 2711.575 814.060 2712.090 814.200 ;
        RECT 2711.770 814.000 2712.090 814.060 ;
        RECT 2711.785 766.260 2712.075 766.305 ;
        RECT 2712.230 766.260 2712.550 766.320 ;
        RECT 2711.785 766.120 2712.550 766.260 ;
        RECT 2711.785 766.075 2712.075 766.120 ;
        RECT 2712.230 766.060 2712.550 766.120 ;
        RECT 2711.325 765.580 2711.615 765.625 ;
        RECT 2711.770 765.580 2712.090 765.640 ;
        RECT 2711.325 765.440 2712.090 765.580 ;
        RECT 2711.325 765.395 2711.615 765.440 ;
        RECT 2711.770 765.380 2712.090 765.440 ;
        RECT 2711.310 717.980 2711.630 718.040 ;
        RECT 2711.115 717.840 2711.630 717.980 ;
        RECT 2711.310 717.780 2711.630 717.840 ;
        RECT 2711.770 717.640 2712.090 717.700 ;
        RECT 2711.575 717.500 2712.090 717.640 ;
        RECT 2711.770 717.440 2712.090 717.500 ;
        RECT 2711.310 669.700 2711.630 669.760 ;
        RECT 2711.785 669.700 2712.075 669.745 ;
        RECT 2711.310 669.560 2712.075 669.700 ;
        RECT 2711.310 669.500 2711.630 669.560 ;
        RECT 2711.785 669.515 2712.075 669.560 ;
        RECT 2710.850 669.020 2711.170 669.080 ;
        RECT 2711.770 669.020 2712.090 669.080 ;
        RECT 2710.850 668.880 2712.090 669.020 ;
        RECT 2710.850 668.820 2711.170 668.880 ;
        RECT 2711.770 668.820 2712.090 668.880 ;
        RECT 2711.770 620.740 2712.090 620.800 ;
        RECT 2711.575 620.600 2712.090 620.740 ;
        RECT 2711.770 620.540 2712.090 620.600 ;
        RECT 2711.310 573.140 2711.630 573.200 ;
        RECT 2711.785 573.140 2712.075 573.185 ;
        RECT 2711.310 573.000 2712.075 573.140 ;
        RECT 2711.310 572.940 2711.630 573.000 ;
        RECT 2711.785 572.955 2712.075 573.000 ;
        RECT 2711.770 572.460 2712.090 572.520 ;
        RECT 2712.690 572.460 2713.010 572.520 ;
        RECT 2711.770 572.320 2713.010 572.460 ;
        RECT 2711.770 572.260 2712.090 572.320 ;
        RECT 2712.690 572.260 2713.010 572.320 ;
        RECT 2711.770 524.180 2712.090 524.240 ;
        RECT 2711.575 524.040 2712.090 524.180 ;
        RECT 2711.770 523.980 2712.090 524.040 ;
        RECT 2711.310 476.580 2711.630 476.640 ;
        RECT 2711.785 476.580 2712.075 476.625 ;
        RECT 2711.310 476.440 2712.075 476.580 ;
        RECT 2711.310 476.380 2711.630 476.440 ;
        RECT 2711.785 476.395 2712.075 476.440 ;
        RECT 2711.770 475.900 2712.090 475.960 ;
        RECT 2712.690 475.900 2713.010 475.960 ;
        RECT 2711.770 475.760 2713.010 475.900 ;
        RECT 2711.770 475.700 2712.090 475.760 ;
        RECT 2712.690 475.700 2713.010 475.760 ;
        RECT 2711.770 427.620 2712.090 427.680 ;
        RECT 2711.575 427.480 2712.090 427.620 ;
        RECT 2711.770 427.420 2712.090 427.480 ;
        RECT 2711.310 380.020 2711.630 380.080 ;
        RECT 2711.785 380.020 2712.075 380.065 ;
        RECT 2711.310 379.880 2712.075 380.020 ;
        RECT 2711.310 379.820 2711.630 379.880 ;
        RECT 2711.785 379.835 2712.075 379.880 ;
        RECT 2711.770 379.340 2712.090 379.400 ;
        RECT 2712.690 379.340 2713.010 379.400 ;
        RECT 2711.770 379.200 2713.010 379.340 ;
        RECT 2711.770 379.140 2712.090 379.200 ;
        RECT 2712.690 379.140 2713.010 379.200 ;
        RECT 2711.770 331.060 2712.090 331.120 ;
        RECT 2711.575 330.920 2712.090 331.060 ;
        RECT 2711.770 330.860 2712.090 330.920 ;
        RECT 2711.310 283.460 2711.630 283.520 ;
        RECT 2711.785 283.460 2712.075 283.505 ;
        RECT 2711.310 283.320 2712.075 283.460 ;
        RECT 2711.310 283.260 2711.630 283.320 ;
        RECT 2711.785 283.275 2712.075 283.320 ;
        RECT 2711.770 282.780 2712.090 282.840 ;
        RECT 2712.690 282.780 2713.010 282.840 ;
        RECT 2711.770 282.640 2713.010 282.780 ;
        RECT 2711.770 282.580 2712.090 282.640 ;
        RECT 2712.690 282.580 2713.010 282.640 ;
        RECT 2711.770 234.500 2712.090 234.560 ;
        RECT 2711.575 234.360 2712.090 234.500 ;
        RECT 2711.770 234.300 2712.090 234.360 ;
        RECT 2711.310 186.900 2711.630 186.960 ;
        RECT 2711.785 186.900 2712.075 186.945 ;
        RECT 2711.310 186.760 2712.075 186.900 ;
        RECT 2711.310 186.700 2711.630 186.760 ;
        RECT 2711.785 186.715 2712.075 186.760 ;
        RECT 2711.770 186.220 2712.090 186.280 ;
        RECT 2711.575 186.080 2712.090 186.220 ;
        RECT 2711.770 186.020 2712.090 186.080 ;
        RECT 2711.770 138.620 2712.090 138.680 ;
        RECT 2711.575 138.480 2712.090 138.620 ;
        RECT 2711.770 138.420 2712.090 138.480 ;
        RECT 2711.770 137.940 2712.090 138.000 ;
        RECT 2711.575 137.800 2712.090 137.940 ;
        RECT 2711.770 137.740 2712.090 137.800 ;
        RECT 2711.310 90.340 2711.630 90.400 ;
        RECT 2711.785 90.340 2712.075 90.385 ;
        RECT 2711.310 90.200 2712.075 90.340 ;
        RECT 2711.310 90.140 2711.630 90.200 ;
        RECT 2711.785 90.155 2712.075 90.200 ;
        RECT 2711.770 89.660 2712.090 89.720 ;
        RECT 2711.575 89.520 2712.090 89.660 ;
        RECT 2711.770 89.460 2712.090 89.520 ;
        RECT 2711.770 42.060 2712.090 42.120 ;
        RECT 2711.575 41.920 2712.090 42.060 ;
        RECT 2711.770 41.860 2712.090 41.920 ;
        RECT 2711.770 41.380 2712.090 41.440 ;
        RECT 2714.545 41.380 2714.835 41.425 ;
        RECT 2711.770 41.240 2714.835 41.380 ;
        RECT 2711.770 41.180 2712.090 41.240 ;
        RECT 2714.545 41.195 2714.835 41.240 ;
        RECT 2714.530 2.960 2714.850 3.020 ;
        RECT 2714.335 2.820 2714.850 2.960 ;
        RECT 2714.530 2.760 2714.850 2.820 ;
      LAYER via ;
        RECT 2711.800 3229.020 2712.060 3229.280 ;
        RECT 2711.800 3181.080 2712.060 3181.340 ;
        RECT 2711.800 3132.460 2712.060 3132.720 ;
        RECT 2711.800 3084.180 2712.060 3084.440 ;
        RECT 2710.880 2987.620 2711.140 2987.880 ;
        RECT 2711.800 2987.620 2712.060 2987.880 ;
        RECT 2710.880 2891.060 2711.140 2891.320 ;
        RECT 2711.800 2891.060 2712.060 2891.320 ;
        RECT 2710.880 2794.500 2711.140 2794.760 ;
        RECT 2711.800 2794.500 2712.060 2794.760 ;
        RECT 2710.880 2649.320 2711.140 2649.580 ;
        RECT 2711.800 2649.320 2712.060 2649.580 ;
        RECT 2710.880 2552.760 2711.140 2553.020 ;
        RECT 2711.800 2552.760 2712.060 2553.020 ;
        RECT 2711.800 2456.200 2712.060 2456.460 ;
        RECT 2711.800 2408.260 2712.060 2408.520 ;
        RECT 2711.800 2359.640 2712.060 2359.900 ;
        RECT 2711.800 2311.700 2712.060 2311.960 ;
        RECT 2711.800 2262.740 2712.060 2263.000 ;
        RECT 2711.800 2214.800 2712.060 2215.060 ;
        RECT 2711.800 2166.180 2712.060 2166.440 ;
        RECT 2711.800 2118.240 2712.060 2118.500 ;
        RECT 2711.800 2069.620 2712.060 2069.880 ;
        RECT 2711.800 2021.680 2712.060 2021.940 ;
        RECT 2711.800 1973.060 2712.060 1973.320 ;
        RECT 2711.800 1925.120 2712.060 1925.380 ;
        RECT 2711.800 1876.500 2712.060 1876.760 ;
        RECT 2711.800 1828.560 2712.060 1828.820 ;
        RECT 2711.800 1779.940 2712.060 1780.200 ;
        RECT 2711.800 1732.000 2712.060 1732.260 ;
        RECT 2711.800 1691.540 2712.060 1691.800 ;
        RECT 2711.800 1690.520 2712.060 1690.780 ;
        RECT 2711.800 1683.380 2712.060 1683.640 ;
        RECT 2711.340 1635.780 2711.600 1636.040 ;
        RECT 2711.800 1538.540 2712.060 1538.800 ;
        RECT 2711.800 1490.940 2712.060 1491.200 ;
        RECT 2711.800 1490.260 2712.060 1490.520 ;
        RECT 2713.180 1490.260 2713.440 1490.520 ;
        RECT 2710.880 1393.700 2711.140 1393.960 ;
        RECT 2711.800 1393.700 2712.060 1393.960 ;
        RECT 2710.880 1346.100 2711.140 1346.360 ;
        RECT 2711.800 1346.100 2712.060 1346.360 ;
        RECT 2710.880 1297.140 2711.140 1297.400 ;
        RECT 2711.800 1297.140 2712.060 1297.400 ;
        RECT 2710.880 1249.540 2711.140 1249.800 ;
        RECT 2711.800 1249.540 2712.060 1249.800 ;
        RECT 2710.880 1200.580 2711.140 1200.840 ;
        RECT 2711.800 1200.580 2712.060 1200.840 ;
        RECT 2710.880 1104.020 2711.140 1104.280 ;
        RECT 2711.800 1104.020 2712.060 1104.280 ;
        RECT 2712.260 1055.400 2712.520 1055.660 ;
        RECT 2711.340 1007.460 2711.600 1007.720 ;
        RECT 2711.800 1007.120 2712.060 1007.380 ;
        RECT 2713.180 1007.120 2713.440 1007.380 ;
        RECT 2712.260 958.840 2712.520 959.100 ;
        RECT 2711.340 910.900 2711.600 911.160 ;
        RECT 2711.800 910.560 2712.060 910.820 ;
        RECT 2713.180 910.560 2713.440 910.820 ;
        RECT 2710.880 862.280 2711.140 862.540 ;
        RECT 2712.260 862.280 2712.520 862.540 ;
        RECT 2711.800 814.000 2712.060 814.260 ;
        RECT 2712.260 766.060 2712.520 766.320 ;
        RECT 2711.800 765.380 2712.060 765.640 ;
        RECT 2711.340 717.780 2711.600 718.040 ;
        RECT 2711.800 717.440 2712.060 717.700 ;
        RECT 2711.340 669.500 2711.600 669.760 ;
        RECT 2710.880 668.820 2711.140 669.080 ;
        RECT 2711.800 668.820 2712.060 669.080 ;
        RECT 2711.800 620.540 2712.060 620.800 ;
        RECT 2711.340 572.940 2711.600 573.200 ;
        RECT 2711.800 572.260 2712.060 572.520 ;
        RECT 2712.720 572.260 2712.980 572.520 ;
        RECT 2711.800 523.980 2712.060 524.240 ;
        RECT 2711.340 476.380 2711.600 476.640 ;
        RECT 2711.800 475.700 2712.060 475.960 ;
        RECT 2712.720 475.700 2712.980 475.960 ;
        RECT 2711.800 427.420 2712.060 427.680 ;
        RECT 2711.340 379.820 2711.600 380.080 ;
        RECT 2711.800 379.140 2712.060 379.400 ;
        RECT 2712.720 379.140 2712.980 379.400 ;
        RECT 2711.800 330.860 2712.060 331.120 ;
        RECT 2711.340 283.260 2711.600 283.520 ;
        RECT 2711.800 282.580 2712.060 282.840 ;
        RECT 2712.720 282.580 2712.980 282.840 ;
        RECT 2711.800 234.300 2712.060 234.560 ;
        RECT 2711.340 186.700 2711.600 186.960 ;
        RECT 2711.800 186.020 2712.060 186.280 ;
        RECT 2711.800 138.420 2712.060 138.680 ;
        RECT 2711.800 137.740 2712.060 138.000 ;
        RECT 2711.340 90.140 2711.600 90.400 ;
        RECT 2711.800 89.460 2712.060 89.720 ;
        RECT 2711.800 41.860 2712.060 42.120 ;
        RECT 2711.800 41.180 2712.060 41.440 ;
        RECT 2714.560 2.760 2714.820 3.020 ;
      LAYER met2 ;
        RECT 890.610 3258.290 890.890 3260.000 ;
        RECT 892.030 3258.290 892.310 3258.405 ;
        RECT 890.610 3258.150 892.310 3258.290 ;
        RECT 890.610 3256.000 890.890 3258.150 ;
        RECT 892.030 3258.035 892.310 3258.150 ;
        RECT 2711.790 3258.035 2712.070 3258.405 ;
        RECT 2711.860 3229.310 2712.000 3258.035 ;
        RECT 2711.800 3228.990 2712.060 3229.310 ;
        RECT 2711.800 3181.050 2712.060 3181.370 ;
        RECT 2711.860 3132.750 2712.000 3181.050 ;
        RECT 2711.800 3132.430 2712.060 3132.750 ;
        RECT 2711.800 3084.150 2712.060 3084.470 ;
        RECT 2711.860 3036.045 2712.000 3084.150 ;
        RECT 2710.870 3035.675 2711.150 3036.045 ;
        RECT 2711.790 3035.675 2712.070 3036.045 ;
        RECT 2710.940 2987.910 2711.080 3035.675 ;
        RECT 2710.880 2987.590 2711.140 2987.910 ;
        RECT 2711.800 2987.590 2712.060 2987.910 ;
        RECT 2711.860 2939.485 2712.000 2987.590 ;
        RECT 2710.870 2939.115 2711.150 2939.485 ;
        RECT 2711.790 2939.115 2712.070 2939.485 ;
        RECT 2710.940 2891.350 2711.080 2939.115 ;
        RECT 2710.880 2891.030 2711.140 2891.350 ;
        RECT 2711.800 2891.030 2712.060 2891.350 ;
        RECT 2711.860 2851.085 2712.000 2891.030 ;
        RECT 2711.790 2850.715 2712.070 2851.085 ;
        RECT 2711.790 2850.035 2712.070 2850.405 ;
        RECT 2711.860 2842.925 2712.000 2850.035 ;
        RECT 2710.870 2842.555 2711.150 2842.925 ;
        RECT 2711.790 2842.555 2712.070 2842.925 ;
        RECT 2710.940 2794.790 2711.080 2842.555 ;
        RECT 2710.880 2794.470 2711.140 2794.790 ;
        RECT 2711.800 2794.470 2712.060 2794.790 ;
        RECT 2711.860 2746.365 2712.000 2794.470 ;
        RECT 2710.870 2745.995 2711.150 2746.365 ;
        RECT 2711.790 2745.995 2712.070 2746.365 ;
        RECT 2710.940 2698.085 2711.080 2745.995 ;
        RECT 2710.870 2697.715 2711.150 2698.085 ;
        RECT 2711.790 2697.715 2712.070 2698.085 ;
        RECT 2711.860 2649.610 2712.000 2697.715 ;
        RECT 2710.880 2649.290 2711.140 2649.610 ;
        RECT 2711.800 2649.290 2712.060 2649.610 ;
        RECT 2710.940 2601.525 2711.080 2649.290 ;
        RECT 2710.870 2601.155 2711.150 2601.525 ;
        RECT 2711.790 2601.155 2712.070 2601.525 ;
        RECT 2711.860 2553.050 2712.000 2601.155 ;
        RECT 2710.880 2552.730 2711.140 2553.050 ;
        RECT 2711.800 2552.730 2712.060 2553.050 ;
        RECT 2710.940 2504.965 2711.080 2552.730 ;
        RECT 2710.870 2504.595 2711.150 2504.965 ;
        RECT 2711.790 2504.595 2712.070 2504.965 ;
        RECT 2711.860 2456.490 2712.000 2504.595 ;
        RECT 2711.800 2456.170 2712.060 2456.490 ;
        RECT 2711.800 2408.230 2712.060 2408.550 ;
        RECT 2711.860 2359.930 2712.000 2408.230 ;
        RECT 2711.800 2359.610 2712.060 2359.930 ;
        RECT 2711.800 2311.670 2712.060 2311.990 ;
        RECT 2711.860 2263.030 2712.000 2311.670 ;
        RECT 2711.800 2262.710 2712.060 2263.030 ;
        RECT 2711.800 2214.770 2712.060 2215.090 ;
        RECT 2711.860 2166.470 2712.000 2214.770 ;
        RECT 2711.800 2166.150 2712.060 2166.470 ;
        RECT 2711.800 2118.210 2712.060 2118.530 ;
        RECT 2711.860 2069.910 2712.000 2118.210 ;
        RECT 2711.800 2069.590 2712.060 2069.910 ;
        RECT 2711.800 2021.650 2712.060 2021.970 ;
        RECT 2711.860 1973.350 2712.000 2021.650 ;
        RECT 2711.800 1973.030 2712.060 1973.350 ;
        RECT 2711.800 1925.090 2712.060 1925.410 ;
        RECT 2711.860 1876.790 2712.000 1925.090 ;
        RECT 2711.800 1876.470 2712.060 1876.790 ;
        RECT 2711.800 1828.530 2712.060 1828.850 ;
        RECT 2711.860 1780.230 2712.000 1828.530 ;
        RECT 2711.800 1779.910 2712.060 1780.230 ;
        RECT 2711.800 1731.970 2712.060 1732.290 ;
        RECT 2711.860 1691.830 2712.000 1731.970 ;
        RECT 2711.800 1691.510 2712.060 1691.830 ;
        RECT 2711.800 1690.490 2712.060 1690.810 ;
        RECT 2711.860 1683.670 2712.000 1690.490 ;
        RECT 2711.800 1683.350 2712.060 1683.670 ;
        RECT 2711.340 1635.810 2711.600 1636.070 ;
        RECT 2711.340 1635.750 2712.000 1635.810 ;
        RECT 2711.400 1635.670 2712.000 1635.750 ;
        RECT 2711.860 1538.830 2712.000 1635.670 ;
        RECT 2711.800 1538.510 2712.060 1538.830 ;
        RECT 2711.800 1490.910 2712.060 1491.230 ;
        RECT 2711.860 1490.550 2712.000 1490.910 ;
        RECT 2711.800 1490.230 2712.060 1490.550 ;
        RECT 2713.180 1490.230 2713.440 1490.550 ;
        RECT 2713.240 1442.805 2713.380 1490.230 ;
        RECT 2711.790 1442.435 2712.070 1442.805 ;
        RECT 2713.170 1442.435 2713.450 1442.805 ;
        RECT 2711.860 1442.125 2712.000 1442.435 ;
        RECT 2710.870 1441.755 2711.150 1442.125 ;
        RECT 2711.790 1441.755 2712.070 1442.125 ;
        RECT 2710.940 1393.990 2711.080 1441.755 ;
        RECT 2710.880 1393.845 2711.140 1393.990 ;
        RECT 2711.800 1393.845 2712.060 1393.990 ;
        RECT 2710.870 1393.475 2711.150 1393.845 ;
        RECT 2711.790 1393.475 2712.070 1393.845 ;
        RECT 2710.940 1346.390 2711.080 1393.475 ;
        RECT 2710.880 1346.070 2711.140 1346.390 ;
        RECT 2711.800 1346.070 2712.060 1346.390 ;
        RECT 2711.860 1345.565 2712.000 1346.070 ;
        RECT 2710.870 1345.195 2711.150 1345.565 ;
        RECT 2711.790 1345.195 2712.070 1345.565 ;
        RECT 2710.940 1297.430 2711.080 1345.195 ;
        RECT 2710.880 1297.285 2711.140 1297.430 ;
        RECT 2711.800 1297.285 2712.060 1297.430 ;
        RECT 2710.870 1296.915 2711.150 1297.285 ;
        RECT 2711.790 1296.915 2712.070 1297.285 ;
        RECT 2710.940 1249.830 2711.080 1296.915 ;
        RECT 2710.880 1249.510 2711.140 1249.830 ;
        RECT 2711.800 1249.510 2712.060 1249.830 ;
        RECT 2711.860 1249.005 2712.000 1249.510 ;
        RECT 2710.870 1248.635 2711.150 1249.005 ;
        RECT 2711.790 1248.635 2712.070 1249.005 ;
        RECT 2710.940 1200.870 2711.080 1248.635 ;
        RECT 2710.880 1200.550 2711.140 1200.870 ;
        RECT 2711.800 1200.550 2712.060 1200.870 ;
        RECT 2711.860 1152.445 2712.000 1200.550 ;
        RECT 2710.870 1152.075 2711.150 1152.445 ;
        RECT 2711.790 1152.075 2712.070 1152.445 ;
        RECT 2710.940 1104.310 2711.080 1152.075 ;
        RECT 2710.880 1103.990 2711.140 1104.310 ;
        RECT 2711.800 1104.165 2712.060 1104.310 ;
        RECT 2711.790 1103.795 2712.070 1104.165 ;
        RECT 2713.170 1103.795 2713.450 1104.165 ;
        RECT 2713.240 1055.885 2713.380 1103.795 ;
        RECT 2712.250 1055.515 2712.530 1055.885 ;
        RECT 2713.170 1055.515 2713.450 1055.885 ;
        RECT 2712.260 1055.370 2712.520 1055.515 ;
        RECT 2711.340 1007.490 2711.600 1007.750 ;
        RECT 2711.340 1007.430 2712.000 1007.490 ;
        RECT 2711.400 1007.410 2712.000 1007.430 ;
        RECT 2711.400 1007.350 2712.060 1007.410 ;
        RECT 2711.800 1007.090 2712.060 1007.350 ;
        RECT 2713.180 1007.090 2713.440 1007.410 ;
        RECT 2713.240 959.325 2713.380 1007.090 ;
        RECT 2712.250 958.955 2712.530 959.325 ;
        RECT 2713.170 958.955 2713.450 959.325 ;
        RECT 2712.260 958.810 2712.520 958.955 ;
        RECT 2711.340 910.930 2711.600 911.190 ;
        RECT 2711.340 910.870 2712.000 910.930 ;
        RECT 2711.400 910.850 2712.000 910.870 ;
        RECT 2711.400 910.790 2712.060 910.850 ;
        RECT 2711.800 910.530 2712.060 910.790 ;
        RECT 2713.180 910.530 2713.440 910.850 ;
        RECT 2713.240 862.765 2713.380 910.530 ;
        RECT 2710.880 862.250 2711.140 862.570 ;
        RECT 2712.250 862.395 2712.530 862.765 ;
        RECT 2713.170 862.395 2713.450 862.765 ;
        RECT 2712.260 862.250 2712.520 862.395 ;
        RECT 2710.940 814.485 2711.080 862.250 ;
        RECT 2710.870 814.115 2711.150 814.485 ;
        RECT 2711.790 814.115 2712.070 814.485 ;
        RECT 2711.800 813.970 2712.060 814.115 ;
        RECT 2712.260 766.090 2712.520 766.350 ;
        RECT 2711.860 766.030 2712.520 766.090 ;
        RECT 2711.860 765.950 2712.460 766.030 ;
        RECT 2711.860 765.670 2712.000 765.950 ;
        RECT 2711.800 765.350 2712.060 765.670 ;
        RECT 2711.340 717.810 2711.600 718.070 ;
        RECT 2711.340 717.750 2712.000 717.810 ;
        RECT 2711.400 717.730 2712.000 717.750 ;
        RECT 2711.400 717.670 2712.060 717.730 ;
        RECT 2711.800 717.410 2712.060 717.670 ;
        RECT 2711.340 669.530 2711.600 669.790 ;
        RECT 2711.340 669.470 2712.000 669.530 ;
        RECT 2711.400 669.390 2712.000 669.470 ;
        RECT 2711.860 669.110 2712.000 669.390 ;
        RECT 2710.880 668.790 2711.140 669.110 ;
        RECT 2711.800 668.790 2712.060 669.110 ;
        RECT 2710.940 621.365 2711.080 668.790 ;
        RECT 2710.870 620.995 2711.150 621.365 ;
        RECT 2711.790 620.995 2712.070 621.365 ;
        RECT 2711.860 620.830 2712.000 620.995 ;
        RECT 2711.800 620.510 2712.060 620.830 ;
        RECT 2711.340 572.970 2711.600 573.230 ;
        RECT 2711.340 572.910 2712.000 572.970 ;
        RECT 2711.400 572.830 2712.000 572.910 ;
        RECT 2711.860 572.550 2712.000 572.830 ;
        RECT 2711.800 572.230 2712.060 572.550 ;
        RECT 2712.720 572.230 2712.980 572.550 ;
        RECT 2712.780 524.805 2712.920 572.230 ;
        RECT 2711.790 524.435 2712.070 524.805 ;
        RECT 2712.710 524.435 2712.990 524.805 ;
        RECT 2711.860 524.270 2712.000 524.435 ;
        RECT 2711.800 523.950 2712.060 524.270 ;
        RECT 2711.340 476.410 2711.600 476.670 ;
        RECT 2711.340 476.350 2712.000 476.410 ;
        RECT 2711.400 476.270 2712.000 476.350 ;
        RECT 2711.860 475.990 2712.000 476.270 ;
        RECT 2711.800 475.670 2712.060 475.990 ;
        RECT 2712.720 475.670 2712.980 475.990 ;
        RECT 2712.780 428.245 2712.920 475.670 ;
        RECT 2711.790 427.875 2712.070 428.245 ;
        RECT 2712.710 427.875 2712.990 428.245 ;
        RECT 2711.860 427.710 2712.000 427.875 ;
        RECT 2711.800 427.390 2712.060 427.710 ;
        RECT 2711.340 379.850 2711.600 380.110 ;
        RECT 2711.340 379.790 2712.000 379.850 ;
        RECT 2711.400 379.710 2712.000 379.790 ;
        RECT 2711.860 379.430 2712.000 379.710 ;
        RECT 2711.800 379.110 2712.060 379.430 ;
        RECT 2712.720 379.110 2712.980 379.430 ;
        RECT 2712.780 331.685 2712.920 379.110 ;
        RECT 2711.790 331.315 2712.070 331.685 ;
        RECT 2712.710 331.315 2712.990 331.685 ;
        RECT 2711.860 331.150 2712.000 331.315 ;
        RECT 2711.800 330.830 2712.060 331.150 ;
        RECT 2711.340 283.290 2711.600 283.550 ;
        RECT 2711.340 283.230 2712.000 283.290 ;
        RECT 2711.400 283.150 2712.000 283.230 ;
        RECT 2711.860 282.870 2712.000 283.150 ;
        RECT 2711.800 282.550 2712.060 282.870 ;
        RECT 2712.720 282.550 2712.980 282.870 ;
        RECT 2712.780 235.125 2712.920 282.550 ;
        RECT 2711.790 234.755 2712.070 235.125 ;
        RECT 2712.710 234.755 2712.990 235.125 ;
        RECT 2711.860 234.590 2712.000 234.755 ;
        RECT 2711.800 234.270 2712.060 234.590 ;
        RECT 2711.340 186.730 2711.600 186.990 ;
        RECT 2711.340 186.670 2712.000 186.730 ;
        RECT 2711.400 186.590 2712.000 186.670 ;
        RECT 2711.860 186.310 2712.000 186.590 ;
        RECT 2711.800 185.990 2712.060 186.310 ;
        RECT 2711.800 138.390 2712.060 138.710 ;
        RECT 2711.860 138.030 2712.000 138.390 ;
        RECT 2711.800 137.710 2712.060 138.030 ;
        RECT 2711.340 90.170 2711.600 90.430 ;
        RECT 2711.340 90.110 2712.000 90.170 ;
        RECT 2711.400 90.030 2712.000 90.110 ;
        RECT 2711.860 89.750 2712.000 90.030 ;
        RECT 2711.800 89.430 2712.060 89.750 ;
        RECT 2711.800 41.830 2712.060 42.150 ;
        RECT 2711.860 41.470 2712.000 41.830 ;
        RECT 2711.800 41.150 2712.060 41.470 ;
        RECT 2714.560 2.730 2714.820 3.050 ;
        RECT 2714.620 2.400 2714.760 2.730 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
      LAYER via2 ;
        RECT 892.030 3258.080 892.310 3258.360 ;
        RECT 2711.790 3258.080 2712.070 3258.360 ;
        RECT 2710.870 3035.720 2711.150 3036.000 ;
        RECT 2711.790 3035.720 2712.070 3036.000 ;
        RECT 2710.870 2939.160 2711.150 2939.440 ;
        RECT 2711.790 2939.160 2712.070 2939.440 ;
        RECT 2711.790 2850.760 2712.070 2851.040 ;
        RECT 2711.790 2850.080 2712.070 2850.360 ;
        RECT 2710.870 2842.600 2711.150 2842.880 ;
        RECT 2711.790 2842.600 2712.070 2842.880 ;
        RECT 2710.870 2746.040 2711.150 2746.320 ;
        RECT 2711.790 2746.040 2712.070 2746.320 ;
        RECT 2710.870 2697.760 2711.150 2698.040 ;
        RECT 2711.790 2697.760 2712.070 2698.040 ;
        RECT 2710.870 2601.200 2711.150 2601.480 ;
        RECT 2711.790 2601.200 2712.070 2601.480 ;
        RECT 2710.870 2504.640 2711.150 2504.920 ;
        RECT 2711.790 2504.640 2712.070 2504.920 ;
        RECT 2711.790 1442.480 2712.070 1442.760 ;
        RECT 2713.170 1442.480 2713.450 1442.760 ;
        RECT 2710.870 1441.800 2711.150 1442.080 ;
        RECT 2711.790 1441.800 2712.070 1442.080 ;
        RECT 2710.870 1393.520 2711.150 1393.800 ;
        RECT 2711.790 1393.520 2712.070 1393.800 ;
        RECT 2710.870 1345.240 2711.150 1345.520 ;
        RECT 2711.790 1345.240 2712.070 1345.520 ;
        RECT 2710.870 1296.960 2711.150 1297.240 ;
        RECT 2711.790 1296.960 2712.070 1297.240 ;
        RECT 2710.870 1248.680 2711.150 1248.960 ;
        RECT 2711.790 1248.680 2712.070 1248.960 ;
        RECT 2710.870 1152.120 2711.150 1152.400 ;
        RECT 2711.790 1152.120 2712.070 1152.400 ;
        RECT 2711.790 1103.840 2712.070 1104.120 ;
        RECT 2713.170 1103.840 2713.450 1104.120 ;
        RECT 2712.250 1055.560 2712.530 1055.840 ;
        RECT 2713.170 1055.560 2713.450 1055.840 ;
        RECT 2712.250 959.000 2712.530 959.280 ;
        RECT 2713.170 959.000 2713.450 959.280 ;
        RECT 2712.250 862.440 2712.530 862.720 ;
        RECT 2713.170 862.440 2713.450 862.720 ;
        RECT 2710.870 814.160 2711.150 814.440 ;
        RECT 2711.790 814.160 2712.070 814.440 ;
        RECT 2710.870 621.040 2711.150 621.320 ;
        RECT 2711.790 621.040 2712.070 621.320 ;
        RECT 2711.790 524.480 2712.070 524.760 ;
        RECT 2712.710 524.480 2712.990 524.760 ;
        RECT 2711.790 427.920 2712.070 428.200 ;
        RECT 2712.710 427.920 2712.990 428.200 ;
        RECT 2711.790 331.360 2712.070 331.640 ;
        RECT 2712.710 331.360 2712.990 331.640 ;
        RECT 2711.790 234.800 2712.070 235.080 ;
        RECT 2712.710 234.800 2712.990 235.080 ;
      LAYER met3 ;
        RECT 892.005 3258.370 892.335 3258.385 ;
        RECT 2711.765 3258.370 2712.095 3258.385 ;
        RECT 892.005 3258.070 2712.095 3258.370 ;
        RECT 892.005 3258.055 892.335 3258.070 ;
        RECT 2711.765 3258.055 2712.095 3258.070 ;
        RECT 2710.845 3036.010 2711.175 3036.025 ;
        RECT 2711.765 3036.010 2712.095 3036.025 ;
        RECT 2710.845 3035.710 2712.095 3036.010 ;
        RECT 2710.845 3035.695 2711.175 3035.710 ;
        RECT 2711.765 3035.695 2712.095 3035.710 ;
        RECT 2710.845 2939.450 2711.175 2939.465 ;
        RECT 2711.765 2939.450 2712.095 2939.465 ;
        RECT 2710.845 2939.150 2712.095 2939.450 ;
        RECT 2710.845 2939.135 2711.175 2939.150 ;
        RECT 2711.765 2939.135 2712.095 2939.150 ;
        RECT 2711.765 2851.050 2712.095 2851.065 ;
        RECT 2711.765 2850.750 2712.770 2851.050 ;
        RECT 2711.765 2850.735 2712.095 2850.750 ;
        RECT 2711.765 2850.370 2712.095 2850.385 ;
        RECT 2712.470 2850.370 2712.770 2850.750 ;
        RECT 2711.765 2850.070 2712.770 2850.370 ;
        RECT 2711.765 2850.055 2712.095 2850.070 ;
        RECT 2710.845 2842.890 2711.175 2842.905 ;
        RECT 2711.765 2842.890 2712.095 2842.905 ;
        RECT 2710.845 2842.590 2712.095 2842.890 ;
        RECT 2710.845 2842.575 2711.175 2842.590 ;
        RECT 2711.765 2842.575 2712.095 2842.590 ;
        RECT 2710.845 2746.330 2711.175 2746.345 ;
        RECT 2711.765 2746.330 2712.095 2746.345 ;
        RECT 2710.845 2746.030 2712.095 2746.330 ;
        RECT 2710.845 2746.015 2711.175 2746.030 ;
        RECT 2711.765 2746.015 2712.095 2746.030 ;
        RECT 2710.845 2698.050 2711.175 2698.065 ;
        RECT 2711.765 2698.050 2712.095 2698.065 ;
        RECT 2710.845 2697.750 2712.095 2698.050 ;
        RECT 2710.845 2697.735 2711.175 2697.750 ;
        RECT 2711.765 2697.735 2712.095 2697.750 ;
        RECT 2710.845 2601.490 2711.175 2601.505 ;
        RECT 2711.765 2601.490 2712.095 2601.505 ;
        RECT 2710.845 2601.190 2712.095 2601.490 ;
        RECT 2710.845 2601.175 2711.175 2601.190 ;
        RECT 2711.765 2601.175 2712.095 2601.190 ;
        RECT 2710.845 2504.930 2711.175 2504.945 ;
        RECT 2711.765 2504.930 2712.095 2504.945 ;
        RECT 2710.845 2504.630 2712.095 2504.930 ;
        RECT 2710.845 2504.615 2711.175 2504.630 ;
        RECT 2711.765 2504.615 2712.095 2504.630 ;
        RECT 2711.765 1442.770 2712.095 1442.785 ;
        RECT 2713.145 1442.770 2713.475 1442.785 ;
        RECT 2711.765 1442.470 2713.475 1442.770 ;
        RECT 2711.765 1442.455 2712.095 1442.470 ;
        RECT 2713.145 1442.455 2713.475 1442.470 ;
        RECT 2710.845 1442.090 2711.175 1442.105 ;
        RECT 2711.765 1442.090 2712.095 1442.105 ;
        RECT 2710.845 1441.790 2712.095 1442.090 ;
        RECT 2710.845 1441.775 2711.175 1441.790 ;
        RECT 2711.765 1441.775 2712.095 1441.790 ;
        RECT 2710.845 1393.810 2711.175 1393.825 ;
        RECT 2711.765 1393.810 2712.095 1393.825 ;
        RECT 2710.845 1393.510 2712.095 1393.810 ;
        RECT 2710.845 1393.495 2711.175 1393.510 ;
        RECT 2711.765 1393.495 2712.095 1393.510 ;
        RECT 2710.845 1345.530 2711.175 1345.545 ;
        RECT 2711.765 1345.530 2712.095 1345.545 ;
        RECT 2710.845 1345.230 2712.095 1345.530 ;
        RECT 2710.845 1345.215 2711.175 1345.230 ;
        RECT 2711.765 1345.215 2712.095 1345.230 ;
        RECT 2710.845 1297.250 2711.175 1297.265 ;
        RECT 2711.765 1297.250 2712.095 1297.265 ;
        RECT 2710.845 1296.950 2712.095 1297.250 ;
        RECT 2710.845 1296.935 2711.175 1296.950 ;
        RECT 2711.765 1296.935 2712.095 1296.950 ;
        RECT 2710.845 1248.970 2711.175 1248.985 ;
        RECT 2711.765 1248.970 2712.095 1248.985 ;
        RECT 2710.845 1248.670 2712.095 1248.970 ;
        RECT 2710.845 1248.655 2711.175 1248.670 ;
        RECT 2711.765 1248.655 2712.095 1248.670 ;
        RECT 2710.845 1152.410 2711.175 1152.425 ;
        RECT 2711.765 1152.410 2712.095 1152.425 ;
        RECT 2710.845 1152.110 2712.095 1152.410 ;
        RECT 2710.845 1152.095 2711.175 1152.110 ;
        RECT 2711.765 1152.095 2712.095 1152.110 ;
        RECT 2711.765 1104.130 2712.095 1104.145 ;
        RECT 2713.145 1104.130 2713.475 1104.145 ;
        RECT 2711.765 1103.830 2713.475 1104.130 ;
        RECT 2711.765 1103.815 2712.095 1103.830 ;
        RECT 2713.145 1103.815 2713.475 1103.830 ;
        RECT 2712.225 1055.850 2712.555 1055.865 ;
        RECT 2713.145 1055.850 2713.475 1055.865 ;
        RECT 2712.225 1055.550 2713.475 1055.850 ;
        RECT 2712.225 1055.535 2712.555 1055.550 ;
        RECT 2713.145 1055.535 2713.475 1055.550 ;
        RECT 2712.225 959.290 2712.555 959.305 ;
        RECT 2713.145 959.290 2713.475 959.305 ;
        RECT 2712.225 958.990 2713.475 959.290 ;
        RECT 2712.225 958.975 2712.555 958.990 ;
        RECT 2713.145 958.975 2713.475 958.990 ;
        RECT 2712.225 862.730 2712.555 862.745 ;
        RECT 2713.145 862.730 2713.475 862.745 ;
        RECT 2712.225 862.430 2713.475 862.730 ;
        RECT 2712.225 862.415 2712.555 862.430 ;
        RECT 2713.145 862.415 2713.475 862.430 ;
        RECT 2710.845 814.450 2711.175 814.465 ;
        RECT 2711.765 814.450 2712.095 814.465 ;
        RECT 2710.845 814.150 2712.095 814.450 ;
        RECT 2710.845 814.135 2711.175 814.150 ;
        RECT 2711.765 814.135 2712.095 814.150 ;
        RECT 2710.845 621.330 2711.175 621.345 ;
        RECT 2711.765 621.330 2712.095 621.345 ;
        RECT 2710.845 621.030 2712.095 621.330 ;
        RECT 2710.845 621.015 2711.175 621.030 ;
        RECT 2711.765 621.015 2712.095 621.030 ;
        RECT 2711.765 524.770 2712.095 524.785 ;
        RECT 2712.685 524.770 2713.015 524.785 ;
        RECT 2711.765 524.470 2713.015 524.770 ;
        RECT 2711.765 524.455 2712.095 524.470 ;
        RECT 2712.685 524.455 2713.015 524.470 ;
        RECT 2711.765 428.210 2712.095 428.225 ;
        RECT 2712.685 428.210 2713.015 428.225 ;
        RECT 2711.765 427.910 2713.015 428.210 ;
        RECT 2711.765 427.895 2712.095 427.910 ;
        RECT 2712.685 427.895 2713.015 427.910 ;
        RECT 2711.765 331.650 2712.095 331.665 ;
        RECT 2712.685 331.650 2713.015 331.665 ;
        RECT 2711.765 331.350 2713.015 331.650 ;
        RECT 2711.765 331.335 2712.095 331.350 ;
        RECT 2712.685 331.335 2713.015 331.350 ;
        RECT 2711.765 235.090 2712.095 235.105 ;
        RECT 2712.685 235.090 2713.015 235.105 ;
        RECT 2711.765 234.790 2713.015 235.090 ;
        RECT 2711.765 234.775 2712.095 234.790 ;
        RECT 2712.685 234.775 2713.015 234.790 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1434.830 3260.075 1435.110 3260.445 ;
        RECT 1434.330 3259.650 1434.610 3260.000 ;
        RECT 1434.900 3259.650 1435.040 3260.075 ;
        RECT 1434.330 3259.510 1435.040 3259.650 ;
        RECT 1434.330 3256.000 1434.610 3259.510 ;
        RECT 2732.490 17.155 2732.770 17.525 ;
        RECT 2732.560 2.400 2732.700 17.155 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 1434.830 3260.120 1435.110 3260.400 ;
        RECT 2732.490 17.200 2732.770 17.480 ;
      LAYER met3 ;
        RECT 1434.805 3260.410 1435.135 3260.425 ;
        RECT 2680.230 3260.410 2680.610 3260.420 ;
        RECT 1434.805 3260.110 2680.610 3260.410 ;
        RECT 1434.805 3260.095 1435.135 3260.110 ;
        RECT 2680.230 3260.100 2680.610 3260.110 ;
        RECT 2680.230 17.490 2680.610 17.500 ;
        RECT 2732.465 17.490 2732.795 17.505 ;
        RECT 2680.230 17.190 2732.795 17.490 ;
        RECT 2680.230 17.180 2680.610 17.190 ;
        RECT 2732.465 17.175 2732.795 17.190 ;
      LAYER via3 ;
        RECT 2680.260 3260.100 2680.580 3260.420 ;
        RECT 2680.260 17.180 2680.580 17.500 ;
      LAYER met4 ;
        RECT 2680.255 3260.095 2680.585 3260.425 ;
        RECT 2680.270 17.505 2680.570 3260.095 ;
        RECT 2680.255 17.175 2680.585 17.505 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1283.740 2615.490 1283.800 ;
        RECT 2746.270 1283.740 2746.590 1283.800 ;
        RECT 2615.170 1283.600 2746.590 1283.740 ;
        RECT 2615.170 1283.540 2615.490 1283.600 ;
        RECT 2746.270 1283.540 2746.590 1283.600 ;
        RECT 2746.270 62.120 2746.590 62.180 ;
        RECT 2750.410 62.120 2750.730 62.180 ;
        RECT 2746.270 61.980 2750.730 62.120 ;
        RECT 2746.270 61.920 2746.590 61.980 ;
        RECT 2750.410 61.920 2750.730 61.980 ;
      LAYER via ;
        RECT 2615.200 1283.540 2615.460 1283.800 ;
        RECT 2746.300 1283.540 2746.560 1283.800 ;
        RECT 2746.300 61.920 2746.560 62.180 ;
        RECT 2750.440 61.920 2750.700 62.180 ;
      LAYER met2 ;
        RECT 2615.190 1289.435 2615.470 1289.805 ;
        RECT 2615.260 1283.830 2615.400 1289.435 ;
        RECT 2615.200 1283.510 2615.460 1283.830 ;
        RECT 2746.300 1283.510 2746.560 1283.830 ;
        RECT 2746.360 62.210 2746.500 1283.510 ;
        RECT 2746.300 61.890 2746.560 62.210 ;
        RECT 2750.440 61.890 2750.700 62.210 ;
        RECT 2750.500 2.400 2750.640 61.890 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1289.480 2615.470 1289.760 ;
      LAYER met3 ;
        RECT 2606.000 1289.770 2610.000 1290.160 ;
        RECT 2615.165 1289.770 2615.495 1289.785 ;
        RECT 2606.000 1289.560 2615.495 1289.770 ;
        RECT 2609.580 1289.470 2615.495 1289.560 ;
        RECT 2615.165 1289.455 2615.495 1289.470 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2767.045 48.365 2767.215 96.475 ;
      LAYER mcon ;
        RECT 2767.045 96.305 2767.215 96.475 ;
      LAYER met1 ;
        RECT 286.650 1145.700 286.970 1145.760 ;
        RECT 296.770 1145.700 297.090 1145.760 ;
        RECT 286.650 1145.560 297.090 1145.700 ;
        RECT 286.650 1145.500 286.970 1145.560 ;
        RECT 296.770 1145.500 297.090 1145.560 ;
        RECT 286.650 134.540 286.970 134.600 ;
        RECT 2766.970 134.540 2767.290 134.600 ;
        RECT 286.650 134.400 2767.290 134.540 ;
        RECT 286.650 134.340 286.970 134.400 ;
        RECT 2766.970 134.340 2767.290 134.400 ;
        RECT 2766.970 96.460 2767.290 96.520 ;
        RECT 2766.775 96.320 2767.290 96.460 ;
        RECT 2766.970 96.260 2767.290 96.320 ;
        RECT 2766.985 48.520 2767.275 48.565 ;
        RECT 2767.890 48.520 2768.210 48.580 ;
        RECT 2766.985 48.380 2768.210 48.520 ;
        RECT 2766.985 48.335 2767.275 48.380 ;
        RECT 2767.890 48.320 2768.210 48.380 ;
      LAYER via ;
        RECT 286.680 1145.500 286.940 1145.760 ;
        RECT 296.800 1145.500 297.060 1145.760 ;
        RECT 286.680 134.340 286.940 134.600 ;
        RECT 2767.000 134.340 2767.260 134.600 ;
        RECT 2767.000 96.260 2767.260 96.520 ;
        RECT 2767.920 48.320 2768.180 48.580 ;
      LAYER met2 ;
        RECT 296.790 1150.715 297.070 1151.085 ;
        RECT 296.860 1145.790 297.000 1150.715 ;
        RECT 286.680 1145.470 286.940 1145.790 ;
        RECT 296.800 1145.470 297.060 1145.790 ;
        RECT 286.740 134.630 286.880 1145.470 ;
        RECT 286.680 134.310 286.940 134.630 ;
        RECT 2767.000 134.310 2767.260 134.630 ;
        RECT 2767.060 96.550 2767.200 134.310 ;
        RECT 2767.000 96.230 2767.260 96.550 ;
        RECT 2767.920 48.290 2768.180 48.610 ;
        RECT 2767.980 2.400 2768.120 48.290 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
      LAYER via2 ;
        RECT 296.790 1150.760 297.070 1151.040 ;
      LAYER met3 ;
        RECT 296.765 1151.050 297.095 1151.065 ;
        RECT 310.000 1151.050 314.000 1151.440 ;
        RECT 296.765 1150.840 314.000 1151.050 ;
        RECT 296.765 1150.750 310.500 1150.840 ;
        RECT 296.765 1150.735 297.095 1150.750 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.190 3268.660 240.510 3268.720 ;
        RECT 748.030 3268.660 748.350 3268.720 ;
        RECT 240.190 3268.520 748.350 3268.660 ;
        RECT 240.190 3268.460 240.510 3268.520 ;
        RECT 748.030 3268.460 748.350 3268.520 ;
        RECT 240.190 57.700 240.510 57.760 ;
        RECT 840.950 57.700 841.270 57.760 ;
        RECT 240.190 57.560 841.270 57.700 ;
        RECT 240.190 57.500 240.510 57.560 ;
        RECT 840.950 57.500 841.270 57.560 ;
      LAYER via ;
        RECT 240.220 3268.460 240.480 3268.720 ;
        RECT 748.060 3268.460 748.320 3268.720 ;
        RECT 240.220 57.500 240.480 57.760 ;
        RECT 840.980 57.500 841.240 57.760 ;
      LAYER met2 ;
        RECT 240.220 3268.430 240.480 3268.750 ;
        RECT 748.060 3268.430 748.320 3268.750 ;
        RECT 240.280 57.790 240.420 3268.430 ;
        RECT 748.120 3260.000 748.260 3268.430 ;
        RECT 748.010 3256.000 748.290 3260.000 ;
        RECT 240.220 57.470 240.480 57.790 ;
        RECT 840.980 57.470 841.240 57.790 ;
        RECT 841.040 2.400 841.180 57.470 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1764.170 3259.480 1764.490 3259.540 ;
        RECT 2780.770 3259.480 2781.090 3259.540 ;
        RECT 1764.170 3259.340 2781.090 3259.480 ;
        RECT 1764.170 3259.280 1764.490 3259.340 ;
        RECT 2780.770 3259.280 2781.090 3259.340 ;
        RECT 2780.770 62.120 2781.090 62.180 ;
        RECT 2785.830 62.120 2786.150 62.180 ;
        RECT 2780.770 61.980 2786.150 62.120 ;
        RECT 2780.770 61.920 2781.090 61.980 ;
        RECT 2785.830 61.920 2786.150 61.980 ;
      LAYER via ;
        RECT 1764.200 3259.280 1764.460 3259.540 ;
        RECT 2780.800 3259.280 2781.060 3259.540 ;
        RECT 2780.800 61.920 2781.060 62.180 ;
        RECT 2785.860 61.920 2786.120 62.180 ;
      LAYER met2 ;
        RECT 1762.770 3259.650 1763.050 3260.000 ;
        RECT 1762.770 3259.570 1764.400 3259.650 ;
        RECT 1762.770 3259.510 1764.460 3259.570 ;
        RECT 1762.770 3256.000 1763.050 3259.510 ;
        RECT 1764.200 3259.250 1764.460 3259.510 ;
        RECT 2780.800 3259.250 2781.060 3259.570 ;
        RECT 2780.860 62.210 2781.000 3259.250 ;
        RECT 2780.800 61.890 2781.060 62.210 ;
        RECT 2785.860 61.890 2786.120 62.210 ;
        RECT 2785.920 2.400 2786.060 61.890 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 348.365 16.065 348.535 17.255 ;
        RECT 2560.505 17.085 2561.135 17.255 ;
      LAYER mcon ;
        RECT 348.365 17.085 348.535 17.255 ;
        RECT 2560.965 17.085 2561.135 17.255 ;
      LAYER met1 ;
        RECT 299.990 379.340 300.310 379.400 ;
        RECT 307.350 379.340 307.670 379.400 ;
        RECT 299.990 379.200 307.670 379.340 ;
        RECT 299.990 379.140 300.310 379.200 ;
        RECT 307.350 379.140 307.670 379.200 ;
        RECT 348.305 17.240 348.595 17.285 ;
        RECT 2560.445 17.240 2560.735 17.285 ;
        RECT 348.305 17.100 2560.735 17.240 ;
        RECT 348.305 17.055 348.595 17.100 ;
        RECT 2560.445 17.055 2560.735 17.100 ;
        RECT 2560.905 17.240 2561.195 17.285 ;
        RECT 2803.770 17.240 2804.090 17.300 ;
        RECT 2560.905 17.100 2804.090 17.240 ;
        RECT 2560.905 17.055 2561.195 17.100 ;
        RECT 2803.770 17.040 2804.090 17.100 ;
        RECT 307.350 16.220 307.670 16.280 ;
        RECT 348.305 16.220 348.595 16.265 ;
        RECT 307.350 16.080 348.595 16.220 ;
        RECT 307.350 16.020 307.670 16.080 ;
        RECT 348.305 16.035 348.595 16.080 ;
      LAYER via ;
        RECT 300.020 379.140 300.280 379.400 ;
        RECT 307.380 379.140 307.640 379.400 ;
        RECT 2803.800 17.040 2804.060 17.300 ;
        RECT 307.380 16.020 307.640 16.280 ;
      LAYER met2 ;
        RECT 300.010 601.275 300.290 601.645 ;
        RECT 300.080 379.430 300.220 601.275 ;
        RECT 300.020 379.110 300.280 379.430 ;
        RECT 307.380 379.110 307.640 379.430 ;
        RECT 307.440 16.310 307.580 379.110 ;
        RECT 2803.800 17.010 2804.060 17.330 ;
        RECT 307.380 15.990 307.640 16.310 ;
        RECT 2803.860 2.400 2804.000 17.010 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 300.010 601.320 300.290 601.600 ;
      LAYER met3 ;
        RECT 299.985 601.610 300.315 601.625 ;
        RECT 310.000 601.610 314.000 602.000 ;
        RECT 299.985 601.400 314.000 601.610 ;
        RECT 299.985 601.310 310.500 601.400 ;
        RECT 299.985 601.295 300.315 601.310 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 738.380 2615.490 738.440 ;
        RECT 2815.270 738.380 2815.590 738.440 ;
        RECT 2615.170 738.240 2815.590 738.380 ;
        RECT 2615.170 738.180 2615.490 738.240 ;
        RECT 2815.270 738.180 2815.590 738.240 ;
        RECT 2815.270 37.980 2815.590 38.040 ;
        RECT 2821.710 37.980 2822.030 38.040 ;
        RECT 2815.270 37.840 2822.030 37.980 ;
        RECT 2815.270 37.780 2815.590 37.840 ;
        RECT 2821.710 37.780 2822.030 37.840 ;
      LAYER via ;
        RECT 2615.200 738.180 2615.460 738.440 ;
        RECT 2815.300 738.180 2815.560 738.440 ;
        RECT 2815.300 37.780 2815.560 38.040 ;
        RECT 2821.740 37.780 2822.000 38.040 ;
      LAYER met2 ;
        RECT 2615.190 739.995 2615.470 740.365 ;
        RECT 2615.260 738.470 2615.400 739.995 ;
        RECT 2615.200 738.150 2615.460 738.470 ;
        RECT 2815.300 738.150 2815.560 738.470 ;
        RECT 2815.360 38.070 2815.500 738.150 ;
        RECT 2815.300 37.750 2815.560 38.070 ;
        RECT 2821.740 37.750 2822.000 38.070 ;
        RECT 2821.800 2.400 2821.940 37.750 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
      LAYER via2 ;
        RECT 2615.190 740.040 2615.470 740.320 ;
      LAYER met3 ;
        RECT 2606.000 740.330 2610.000 740.720 ;
        RECT 2615.165 740.330 2615.495 740.345 ;
        RECT 2606.000 740.120 2615.495 740.330 ;
        RECT 2609.580 740.030 2615.495 740.120 ;
        RECT 2615.165 740.015 2615.495 740.030 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1407.210 3258.800 1407.530 3258.860 ;
        RECT 2835.970 3258.800 2836.290 3258.860 ;
        RECT 1407.210 3258.660 2836.290 3258.800 ;
        RECT 1407.210 3258.600 1407.530 3258.660 ;
        RECT 2835.970 3258.600 2836.290 3258.660 ;
        RECT 2835.970 62.120 2836.290 62.180 ;
        RECT 2839.190 62.120 2839.510 62.180 ;
        RECT 2835.970 61.980 2839.510 62.120 ;
        RECT 2835.970 61.920 2836.290 61.980 ;
        RECT 2839.190 61.920 2839.510 61.980 ;
      LAYER via ;
        RECT 1407.240 3258.600 1407.500 3258.860 ;
        RECT 2836.000 3258.600 2836.260 3258.860 ;
        RECT 2836.000 61.920 2836.260 62.180 ;
        RECT 2839.220 61.920 2839.480 62.180 ;
      LAYER met2 ;
        RECT 1405.810 3258.970 1406.090 3260.000 ;
        RECT 1405.810 3258.890 1407.440 3258.970 ;
        RECT 1405.810 3258.830 1407.500 3258.890 ;
        RECT 1405.810 3256.000 1406.090 3258.830 ;
        RECT 1407.240 3258.570 1407.500 3258.830 ;
        RECT 2836.000 3258.570 2836.260 3258.890 ;
        RECT 2836.060 62.210 2836.200 3258.570 ;
        RECT 2836.000 61.890 2836.260 62.210 ;
        RECT 2839.220 61.890 2839.480 62.210 ;
        RECT 2839.280 2.400 2839.420 61.890 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 462.640 2615.490 462.700 ;
        RECT 2857.130 462.640 2857.450 462.700 ;
        RECT 2615.170 462.500 2857.450 462.640 ;
        RECT 2615.170 462.440 2615.490 462.500 ;
        RECT 2857.130 462.440 2857.450 462.500 ;
      LAYER via ;
        RECT 2615.200 462.440 2615.460 462.700 ;
        RECT 2857.160 462.440 2857.420 462.700 ;
      LAYER met2 ;
        RECT 2615.190 465.275 2615.470 465.645 ;
        RECT 2615.260 462.730 2615.400 465.275 ;
        RECT 2615.200 462.410 2615.460 462.730 ;
        RECT 2857.160 462.410 2857.420 462.730 ;
        RECT 2857.220 2.400 2857.360 462.410 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
      LAYER via2 ;
        RECT 2615.190 465.320 2615.470 465.600 ;
      LAYER met3 ;
        RECT 2606.000 465.610 2610.000 466.000 ;
        RECT 2615.165 465.610 2615.495 465.625 ;
        RECT 2606.000 465.400 2615.495 465.610 ;
        RECT 2609.580 465.310 2615.495 465.400 ;
        RECT 2615.165 465.295 2615.495 465.310 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 3229.560 2615.490 3229.620 ;
        RECT 2870.470 3229.560 2870.790 3229.620 ;
        RECT 2615.170 3229.420 2870.790 3229.560 ;
        RECT 2615.170 3229.360 2615.490 3229.420 ;
        RECT 2870.470 3229.360 2870.790 3229.420 ;
      LAYER via ;
        RECT 2615.200 3229.360 2615.460 3229.620 ;
        RECT 2870.500 3229.360 2870.760 3229.620 ;
      LAYER met2 ;
        RECT 2615.190 3234.235 2615.470 3234.605 ;
        RECT 2615.260 3229.650 2615.400 3234.235 ;
        RECT 2615.200 3229.330 2615.460 3229.650 ;
        RECT 2870.500 3229.330 2870.760 3229.650 ;
        RECT 2870.560 20.130 2870.700 3229.330 ;
        RECT 2870.560 19.990 2875.300 20.130 ;
        RECT 2875.160 2.400 2875.300 19.990 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 2615.190 3234.280 2615.470 3234.560 ;
      LAYER met3 ;
        RECT 2606.000 3234.570 2610.000 3234.960 ;
        RECT 2615.165 3234.570 2615.495 3234.585 ;
        RECT 2606.000 3234.360 2615.495 3234.570 ;
        RECT 2609.580 3234.270 2615.495 3234.360 ;
        RECT 2615.165 3234.255 2615.495 3234.270 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 945.440 2615.490 945.500 ;
        RECT 2860.350 945.440 2860.670 945.500 ;
        RECT 2615.170 945.300 2860.670 945.440 ;
        RECT 2615.170 945.240 2615.490 945.300 ;
        RECT 2860.350 945.240 2860.670 945.300 ;
        RECT 2860.350 16.220 2860.670 16.280 ;
        RECT 2893.010 16.220 2893.330 16.280 ;
        RECT 2860.350 16.080 2893.330 16.220 ;
        RECT 2860.350 16.020 2860.670 16.080 ;
        RECT 2893.010 16.020 2893.330 16.080 ;
      LAYER via ;
        RECT 2615.200 945.240 2615.460 945.500 ;
        RECT 2860.380 945.240 2860.640 945.500 ;
        RECT 2860.380 16.020 2860.640 16.280 ;
        RECT 2893.040 16.020 2893.300 16.280 ;
      LAYER met2 ;
        RECT 2615.190 950.795 2615.470 951.165 ;
        RECT 2615.260 945.530 2615.400 950.795 ;
        RECT 2615.200 945.210 2615.460 945.530 ;
        RECT 2860.380 945.210 2860.640 945.530 ;
        RECT 2860.440 16.310 2860.580 945.210 ;
        RECT 2860.380 15.990 2860.640 16.310 ;
        RECT 2893.040 15.990 2893.300 16.310 ;
        RECT 2893.100 2.400 2893.240 15.990 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 2615.190 950.840 2615.470 951.120 ;
      LAYER met3 ;
        RECT 2606.000 951.130 2610.000 951.520 ;
        RECT 2615.165 951.130 2615.495 951.145 ;
        RECT 2606.000 950.920 2615.495 951.130 ;
        RECT 2609.580 950.830 2615.495 950.920 ;
        RECT 2615.165 950.815 2615.495 950.830 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 669.830 244.020 670.150 244.080 ;
        RECT 675.350 244.020 675.670 244.080 ;
        RECT 669.830 243.880 675.670 244.020 ;
        RECT 669.830 243.820 670.150 243.880 ;
        RECT 675.350 243.820 675.670 243.880 ;
        RECT 675.350 120.940 675.670 121.000 ;
        RECT 2866.790 120.940 2867.110 121.000 ;
        RECT 675.350 120.800 2867.110 120.940 ;
        RECT 675.350 120.740 675.670 120.800 ;
        RECT 2866.790 120.740 2867.110 120.800 ;
        RECT 2866.790 20.300 2867.110 20.360 ;
        RECT 2910.950 20.300 2911.270 20.360 ;
        RECT 2866.790 20.160 2911.270 20.300 ;
        RECT 2866.790 20.100 2867.110 20.160 ;
        RECT 2910.950 20.100 2911.270 20.160 ;
      LAYER via ;
        RECT 669.860 243.820 670.120 244.080 ;
        RECT 675.380 243.820 675.640 244.080 ;
        RECT 675.380 120.740 675.640 121.000 ;
        RECT 2866.820 120.740 2867.080 121.000 ;
        RECT 2866.820 20.100 2867.080 20.360 ;
        RECT 2910.980 20.100 2911.240 20.360 ;
      LAYER met2 ;
        RECT 669.810 260.000 670.090 264.000 ;
        RECT 669.920 244.110 670.060 260.000 ;
        RECT 669.860 243.790 670.120 244.110 ;
        RECT 675.380 243.790 675.640 244.110 ;
        RECT 675.440 121.030 675.580 243.790 ;
        RECT 675.380 120.710 675.640 121.030 ;
        RECT 2866.820 120.710 2867.080 121.030 ;
        RECT 2866.880 20.390 2867.020 120.710 ;
        RECT 2866.820 20.070 2867.080 20.390 ;
        RECT 2910.980 20.070 2911.240 20.390 ;
        RECT 2911.040 2.400 2911.180 20.070 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 285.730 1235.460 286.050 1235.520 ;
        RECT 296.770 1235.460 297.090 1235.520 ;
        RECT 285.730 1235.320 297.090 1235.460 ;
        RECT 285.730 1235.260 286.050 1235.320 ;
        RECT 296.770 1235.260 297.090 1235.320 ;
        RECT 285.730 237.900 286.050 237.960 ;
        RECT 855.670 237.900 855.990 237.960 ;
        RECT 285.730 237.760 855.990 237.900 ;
        RECT 285.730 237.700 286.050 237.760 ;
        RECT 855.670 237.700 855.990 237.760 ;
        RECT 854.750 193.020 855.070 193.080 ;
        RECT 855.670 193.020 855.990 193.080 ;
        RECT 854.750 192.880 855.990 193.020 ;
        RECT 854.750 192.820 855.070 192.880 ;
        RECT 855.670 192.820 855.990 192.880 ;
        RECT 855.670 137.940 855.990 138.000 ;
        RECT 856.130 137.940 856.450 138.000 ;
        RECT 855.670 137.800 856.450 137.940 ;
        RECT 855.670 137.740 855.990 137.800 ;
        RECT 856.130 137.740 856.450 137.800 ;
        RECT 855.670 14.180 855.990 14.240 ;
        RECT 855.670 14.040 859.120 14.180 ;
        RECT 855.670 13.980 855.990 14.040 ;
        RECT 858.980 13.900 859.120 14.040 ;
        RECT 858.890 13.640 859.210 13.900 ;
      LAYER via ;
        RECT 285.760 1235.260 286.020 1235.520 ;
        RECT 296.800 1235.260 297.060 1235.520 ;
        RECT 285.760 237.700 286.020 237.960 ;
        RECT 855.700 237.700 855.960 237.960 ;
        RECT 854.780 192.820 855.040 193.080 ;
        RECT 855.700 192.820 855.960 193.080 ;
        RECT 855.700 137.740 855.960 138.000 ;
        RECT 856.160 137.740 856.420 138.000 ;
        RECT 855.700 13.980 855.960 14.240 ;
        RECT 858.920 13.640 859.180 13.900 ;
      LAYER met2 ;
        RECT 285.760 1235.230 286.020 1235.550 ;
        RECT 296.800 1235.405 297.060 1235.550 ;
        RECT 285.820 237.990 285.960 1235.230 ;
        RECT 296.790 1235.035 297.070 1235.405 ;
        RECT 285.760 237.670 286.020 237.990 ;
        RECT 855.700 237.670 855.960 237.990 ;
        RECT 855.760 193.110 855.900 237.670 ;
        RECT 854.780 192.790 855.040 193.110 ;
        RECT 855.700 192.790 855.960 193.110 ;
        RECT 854.840 145.365 854.980 192.790 ;
        RECT 854.770 144.995 855.050 145.365 ;
        RECT 855.690 144.995 855.970 145.365 ;
        RECT 855.760 138.030 855.900 144.995 ;
        RECT 855.700 137.710 855.960 138.030 ;
        RECT 856.160 137.710 856.420 138.030 ;
        RECT 856.220 48.690 856.360 137.710 ;
        RECT 855.760 48.550 856.360 48.690 ;
        RECT 855.760 14.270 855.900 48.550 ;
        RECT 855.700 13.950 855.960 14.270 ;
        RECT 858.920 13.610 859.180 13.930 ;
        RECT 858.980 2.400 859.120 13.610 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 296.790 1235.080 297.070 1235.360 ;
        RECT 854.770 145.040 855.050 145.320 ;
        RECT 855.690 145.040 855.970 145.320 ;
      LAYER met3 ;
        RECT 296.765 1235.370 297.095 1235.385 ;
        RECT 310.000 1235.370 314.000 1235.760 ;
        RECT 296.765 1235.160 314.000 1235.370 ;
        RECT 296.765 1235.070 310.500 1235.160 ;
        RECT 296.765 1235.055 297.095 1235.070 ;
        RECT 854.745 145.330 855.075 145.345 ;
        RECT 855.665 145.330 855.995 145.345 ;
        RECT 854.745 145.030 855.995 145.330 ;
        RECT 854.745 145.015 855.075 145.030 ;
        RECT 855.665 145.015 855.995 145.030 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.830 15.880 877.150 15.940 ;
        RECT 882.810 15.880 883.130 15.940 ;
        RECT 876.830 15.740 883.130 15.880 ;
        RECT 876.830 15.680 877.150 15.740 ;
        RECT 882.810 15.680 883.130 15.740 ;
      LAYER via ;
        RECT 876.860 15.680 877.120 15.940 ;
        RECT 882.840 15.680 883.100 15.940 ;
      LAYER met2 ;
        RECT 2105.970 3260.755 2106.250 3261.125 ;
        RECT 2106.040 3260.000 2106.180 3260.755 ;
        RECT 2105.930 3256.000 2106.210 3260.000 ;
        RECT 882.830 244.955 883.110 245.325 ;
        RECT 882.900 15.970 883.040 244.955 ;
        RECT 876.860 15.650 877.120 15.970 ;
        RECT 882.840 15.650 883.100 15.970 ;
        RECT 876.920 2.400 877.060 15.650 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 2105.970 3260.800 2106.250 3261.080 ;
        RECT 882.830 245.000 883.110 245.280 ;
      LAYER met3 ;
        RECT 2105.945 3261.100 2106.275 3261.105 ;
        RECT 2105.945 3261.090 2106.530 3261.100 ;
        RECT 2105.945 3260.790 2106.730 3261.090 ;
        RECT 2105.945 3260.780 2106.530 3260.790 ;
        RECT 2105.945 3260.775 2106.275 3260.780 ;
        RECT 2106.150 3252.250 2106.530 3252.260 ;
        RECT 2683.910 3252.250 2684.290 3252.260 ;
        RECT 2106.150 3251.950 2684.290 3252.250 ;
        RECT 2106.150 3251.940 2106.530 3251.950 ;
        RECT 2683.910 3251.940 2684.290 3251.950 ;
        RECT 882.805 245.290 883.135 245.305 ;
        RECT 2683.910 245.290 2684.290 245.300 ;
        RECT 882.805 244.990 2684.290 245.290 ;
        RECT 882.805 244.975 883.135 244.990 ;
        RECT 2683.910 244.980 2684.290 244.990 ;
      LAYER via3 ;
        RECT 2106.180 3260.780 2106.500 3261.100 ;
        RECT 2106.180 3251.940 2106.500 3252.260 ;
        RECT 2683.940 3251.940 2684.260 3252.260 ;
        RECT 2683.940 244.980 2684.260 245.300 ;
      LAYER met4 ;
        RECT 2106.175 3260.775 2106.505 3261.105 ;
        RECT 2106.190 3252.265 2106.490 3260.775 ;
        RECT 2106.175 3251.935 2106.505 3252.265 ;
        RECT 2683.935 3251.935 2684.265 3252.265 ;
        RECT 2683.950 245.305 2684.250 3251.935 ;
        RECT 2683.935 244.975 2684.265 245.305 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2011.190 247.760 2011.510 247.820 ;
        RECT 2400.350 247.760 2400.670 247.820 ;
        RECT 2011.190 247.620 2400.670 247.760 ;
        RECT 2011.190 247.560 2011.510 247.620 ;
        RECT 2400.350 247.560 2400.670 247.620 ;
        RECT 896.610 86.940 896.930 87.000 ;
        RECT 2011.190 86.940 2011.510 87.000 ;
        RECT 896.610 86.800 2011.510 86.940 ;
        RECT 896.610 86.740 896.930 86.800 ;
        RECT 2011.190 86.740 2011.510 86.800 ;
        RECT 894.770 14.180 895.090 14.240 ;
        RECT 896.610 14.180 896.930 14.240 ;
        RECT 894.770 14.040 896.930 14.180 ;
        RECT 894.770 13.980 895.090 14.040 ;
        RECT 896.610 13.980 896.930 14.040 ;
      LAYER via ;
        RECT 2011.220 247.560 2011.480 247.820 ;
        RECT 2400.380 247.560 2400.640 247.820 ;
        RECT 896.640 86.740 896.900 87.000 ;
        RECT 2011.220 86.740 2011.480 87.000 ;
        RECT 894.800 13.980 895.060 14.240 ;
        RECT 896.640 13.980 896.900 14.240 ;
      LAYER met2 ;
        RECT 2400.330 260.000 2400.610 264.000 ;
        RECT 2400.440 247.850 2400.580 260.000 ;
        RECT 2011.220 247.530 2011.480 247.850 ;
        RECT 2400.380 247.530 2400.640 247.850 ;
        RECT 2011.280 87.030 2011.420 247.530 ;
        RECT 896.640 86.710 896.900 87.030 ;
        RECT 2011.220 86.710 2011.480 87.030 ;
        RECT 896.700 14.270 896.840 86.710 ;
        RECT 894.800 13.950 895.060 14.270 ;
        RECT 896.640 13.950 896.900 14.270 ;
        RECT 894.860 2.400 895.000 13.950 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 15.880 913.030 15.940 ;
        RECT 917.310 15.880 917.630 15.940 ;
        RECT 912.710 15.740 917.630 15.880 ;
        RECT 912.710 15.680 913.030 15.740 ;
        RECT 917.310 15.680 917.630 15.740 ;
      LAYER via ;
        RECT 912.740 15.680 913.000 15.940 ;
        RECT 917.340 15.680 917.600 15.940 ;
      LAYER met2 ;
        RECT 2608.290 1211.915 2608.570 1212.285 ;
        RECT 2608.360 1159.130 2608.500 1211.915 ;
        RECT 2607.900 1158.990 2608.500 1159.130 ;
        RECT 2607.900 1083.085 2608.040 1158.990 ;
        RECT 2607.830 1082.715 2608.110 1083.085 ;
        RECT 2602.770 262.635 2603.050 263.005 ;
        RECT 2602.840 193.645 2602.980 262.635 ;
        RECT 2602.770 193.275 2603.050 193.645 ;
        RECT 2603.230 192.595 2603.510 192.965 ;
        RECT 2603.300 180.725 2603.440 192.595 ;
        RECT 2603.230 180.355 2603.510 180.725 ;
        RECT 917.330 99.435 917.610 99.805 ;
        RECT 917.400 15.970 917.540 99.435 ;
        RECT 912.740 15.650 913.000 15.970 ;
        RECT 917.340 15.650 917.600 15.970 ;
        RECT 912.800 2.400 912.940 15.650 ;
        RECT 912.590 -4.800 913.150 2.400 ;
      LAYER via2 ;
        RECT 2608.290 1211.960 2608.570 1212.240 ;
        RECT 2607.830 1082.760 2608.110 1083.040 ;
        RECT 2602.770 262.680 2603.050 262.960 ;
        RECT 2602.770 193.320 2603.050 193.600 ;
        RECT 2603.230 192.640 2603.510 192.920 ;
        RECT 2603.230 180.400 2603.510 180.680 ;
        RECT 917.330 99.480 917.610 99.760 ;
      LAYER met3 ;
        RECT 2606.000 1311.320 2610.000 1311.920 ;
        RECT 2606.670 1310.860 2606.970 1311.320 ;
        RECT 2606.630 1310.540 2607.010 1310.860 ;
        RECT 2606.630 1212.250 2607.010 1212.260 ;
        RECT 2608.265 1212.250 2608.595 1212.265 ;
        RECT 2606.630 1211.950 2608.595 1212.250 ;
        RECT 2606.630 1211.940 2607.010 1211.950 ;
        RECT 2608.265 1211.935 2608.595 1211.950 ;
        RECT 2607.805 1083.050 2608.135 1083.065 ;
        RECT 2612.150 1083.050 2612.530 1083.060 ;
        RECT 2607.805 1082.750 2612.530 1083.050 ;
        RECT 2607.805 1082.735 2608.135 1082.750 ;
        RECT 2612.150 1082.740 2612.530 1082.750 ;
        RECT 2602.745 262.970 2603.075 262.985 ;
        RECT 2603.870 262.970 2604.250 262.980 ;
        RECT 2602.745 262.670 2604.250 262.970 ;
        RECT 2602.745 262.655 2603.075 262.670 ;
        RECT 2603.870 262.660 2604.250 262.670 ;
        RECT 2602.745 193.610 2603.075 193.625 ;
        RECT 2602.745 193.295 2603.290 193.610 ;
        RECT 2602.990 192.945 2603.290 193.295 ;
        RECT 2602.990 192.630 2603.535 192.945 ;
        RECT 2603.205 192.615 2603.535 192.630 ;
        RECT 2603.205 180.690 2603.535 180.705 ;
        RECT 2603.870 180.690 2604.250 180.700 ;
        RECT 2603.205 180.390 2604.250 180.690 ;
        RECT 2603.205 180.375 2603.535 180.390 ;
        RECT 2603.870 180.380 2604.250 180.390 ;
        RECT 917.305 99.770 917.635 99.785 ;
        RECT 2603.870 99.770 2604.250 99.780 ;
        RECT 917.305 99.470 2604.250 99.770 ;
        RECT 917.305 99.455 917.635 99.470 ;
        RECT 2603.870 99.460 2604.250 99.470 ;
      LAYER via3 ;
        RECT 2606.660 1310.540 2606.980 1310.860 ;
        RECT 2606.660 1211.940 2606.980 1212.260 ;
        RECT 2612.180 1082.740 2612.500 1083.060 ;
        RECT 2603.900 262.660 2604.220 262.980 ;
        RECT 2603.900 180.380 2604.220 180.700 ;
        RECT 2603.900 99.460 2604.220 99.780 ;
      LAYER met4 ;
        RECT 2606.655 1310.850 2606.985 1310.865 ;
        RECT 2601.150 1310.550 2606.985 1310.850 ;
        RECT 2601.150 1246.250 2601.450 1310.550 ;
        RECT 2606.655 1310.535 2606.985 1310.550 ;
        RECT 2601.150 1245.950 2605.130 1246.250 ;
        RECT 2604.830 1212.250 2605.130 1245.950 ;
        RECT 2606.655 1212.250 2606.985 1212.265 ;
        RECT 2604.830 1211.950 2606.985 1212.250 ;
        RECT 2606.655 1211.935 2606.985 1211.950 ;
        RECT 2601.630 1082.310 2602.810 1083.490 ;
        RECT 2611.750 1082.310 2612.930 1083.490 ;
        RECT 2602.070 1038.850 2602.370 1082.310 ;
        RECT 2602.070 1038.550 2605.130 1038.850 ;
        RECT 2604.830 981.050 2605.130 1038.550 ;
        RECT 2602.070 980.750 2605.130 981.050 ;
        RECT 2602.070 977.650 2602.370 980.750 ;
        RECT 2602.070 977.350 2603.290 977.650 ;
        RECT 2602.990 943.650 2603.290 977.350 ;
        RECT 2601.150 943.350 2603.290 943.650 ;
        RECT 2601.150 821.250 2601.450 943.350 ;
        RECT 2601.150 820.950 2604.210 821.250 ;
        RECT 2603.910 811.050 2604.210 820.950 ;
        RECT 2602.070 810.750 2604.210 811.050 ;
        RECT 2602.070 780.450 2602.370 810.750 ;
        RECT 2602.070 780.150 2603.290 780.450 ;
        RECT 2592.430 684.510 2593.610 685.690 ;
        RECT 2592.870 556.490 2593.170 684.510 ;
        RECT 2602.990 682.290 2603.290 780.150 ;
        RECT 2602.550 681.110 2603.730 682.290 ;
        RECT 2592.430 555.310 2593.610 556.490 ;
        RECT 2605.310 555.310 2606.490 556.490 ;
        RECT 2605.750 508.450 2606.050 555.310 ;
        RECT 2605.750 508.150 2607.890 508.450 ;
        RECT 2607.590 498.250 2607.890 508.150 ;
        RECT 2606.670 497.950 2607.890 498.250 ;
        RECT 2606.670 474.450 2606.970 497.950 ;
        RECT 2605.750 474.150 2606.970 474.450 ;
        RECT 2605.750 447.690 2606.050 474.150 ;
        RECT 2605.310 446.510 2606.490 447.690 ;
        RECT 2601.630 439.710 2602.810 440.890 ;
        RECT 2602.070 426.850 2602.370 439.710 ;
        RECT 2601.150 426.550 2602.370 426.850 ;
        RECT 2601.150 383.090 2601.450 426.550 ;
        RECT 2600.710 381.910 2601.890 383.090 ;
        RECT 2606.230 381.910 2607.410 383.090 ;
        RECT 2606.670 362.250 2606.970 381.910 ;
        RECT 2605.750 361.950 2606.970 362.250 ;
        RECT 2605.750 328.250 2606.050 361.950 ;
        RECT 2604.830 327.950 2606.050 328.250 ;
        RECT 2604.830 324.850 2605.130 327.950 ;
        RECT 2603.910 324.550 2605.130 324.850 ;
        RECT 2603.910 304.450 2604.210 324.550 ;
        RECT 2603.910 304.150 2605.130 304.450 ;
        RECT 2604.830 273.850 2605.130 304.150 ;
        RECT 2603.910 273.550 2605.130 273.850 ;
        RECT 2603.910 262.985 2604.210 273.550 ;
        RECT 2603.895 262.655 2604.225 262.985 ;
        RECT 2603.895 180.375 2604.225 180.705 ;
        RECT 2603.910 99.785 2604.210 180.375 ;
        RECT 2603.895 99.455 2604.225 99.785 ;
      LAYER met5 ;
        RECT 2601.420 1082.100 2613.140 1083.700 ;
        RECT 2592.220 684.300 2603.940 685.900 ;
        RECT 2602.340 680.900 2603.940 684.300 ;
        RECT 2592.220 555.100 2606.700 556.700 ;
        RECT 2597.740 446.300 2606.700 447.900 ;
        RECT 2597.740 441.100 2599.340 446.300 ;
        RECT 2597.740 439.500 2603.020 441.100 ;
        RECT 2600.500 381.700 2607.620 383.300 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 931.185 41.565 931.355 89.675 ;
      LAYER mcon ;
        RECT 931.185 89.505 931.355 89.675 ;
      LAYER met1 ;
        RECT 931.110 197.100 931.430 197.160 ;
        RECT 2623.450 197.100 2623.770 197.160 ;
        RECT 931.110 196.960 2623.770 197.100 ;
        RECT 931.110 196.900 931.430 196.960 ;
        RECT 2623.450 196.900 2623.770 196.960 ;
        RECT 931.110 89.660 931.430 89.720 ;
        RECT 930.915 89.520 931.430 89.660 ;
        RECT 931.110 89.460 931.430 89.520 ;
        RECT 931.110 41.720 931.430 41.780 ;
        RECT 930.915 41.580 931.430 41.720 ;
        RECT 931.110 41.520 931.430 41.580 ;
        RECT 931.110 14.180 931.430 14.240 ;
        RECT 930.280 14.040 931.430 14.180 ;
        RECT 930.280 13.900 930.420 14.040 ;
        RECT 931.110 13.980 931.430 14.040 ;
        RECT 930.190 13.640 930.510 13.900 ;
      LAYER via ;
        RECT 931.140 196.900 931.400 197.160 ;
        RECT 2623.480 196.900 2623.740 197.160 ;
        RECT 931.140 89.460 931.400 89.720 ;
        RECT 931.140 41.520 931.400 41.780 ;
        RECT 931.140 13.980 931.400 14.240 ;
        RECT 930.220 13.640 930.480 13.900 ;
      LAYER met2 ;
        RECT 2623.470 1415.915 2623.750 1416.285 ;
        RECT 2623.540 197.190 2623.680 1415.915 ;
        RECT 931.140 196.870 931.400 197.190 ;
        RECT 2623.480 196.870 2623.740 197.190 ;
        RECT 931.200 90.850 931.340 196.870 ;
        RECT 931.200 90.710 931.800 90.850 ;
        RECT 931.660 90.170 931.800 90.710 ;
        RECT 931.200 90.030 931.800 90.170 ;
        RECT 931.200 89.750 931.340 90.030 ;
        RECT 931.140 89.430 931.400 89.750 ;
        RECT 931.140 41.490 931.400 41.810 ;
        RECT 931.200 14.270 931.340 41.490 ;
        RECT 931.140 13.950 931.400 14.270 ;
        RECT 930.220 13.610 930.480 13.930 ;
        RECT 930.280 2.400 930.420 13.610 ;
        RECT 930.070 -4.800 930.630 2.400 ;
      LAYER via2 ;
        RECT 2623.470 1415.960 2623.750 1416.240 ;
      LAYER met3 ;
        RECT 2606.000 1416.250 2610.000 1416.640 ;
        RECT 2623.445 1416.250 2623.775 1416.265 ;
        RECT 2606.000 1416.040 2623.775 1416.250 ;
        RECT 2609.580 1415.950 2623.775 1416.040 ;
        RECT 2623.445 1415.935 2623.775 1415.950 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 14.520 948.450 14.580 ;
        RECT 951.810 14.520 952.130 14.580 ;
        RECT 948.130 14.380 952.130 14.520 ;
        RECT 948.130 14.320 948.450 14.380 ;
        RECT 951.810 14.320 952.130 14.380 ;
      LAYER via ;
        RECT 948.160 14.320 948.420 14.580 ;
        RECT 951.840 14.320 952.100 14.580 ;
      LAYER met2 ;
        RECT 951.830 182.395 952.110 182.765 ;
        RECT 951.900 14.610 952.040 182.395 ;
        RECT 948.160 14.290 948.420 14.610 ;
        RECT 951.840 14.290 952.100 14.610 ;
        RECT 948.220 2.400 948.360 14.290 ;
        RECT 948.010 -4.800 948.570 2.400 ;
      LAYER via2 ;
        RECT 951.830 182.440 952.110 182.720 ;
      LAYER met3 ;
        RECT 2606.000 2558.650 2610.000 2559.040 ;
        RECT 2629.630 2558.650 2630.010 2558.660 ;
        RECT 2606.000 2558.440 2630.010 2558.650 ;
        RECT 2609.580 2558.350 2630.010 2558.440 ;
        RECT 2629.630 2558.340 2630.010 2558.350 ;
        RECT 951.805 182.730 952.135 182.745 ;
        RECT 2629.630 182.730 2630.010 182.740 ;
        RECT 951.805 182.430 2630.010 182.730 ;
        RECT 951.805 182.415 952.135 182.430 ;
        RECT 2629.630 182.420 2630.010 182.430 ;
      LAYER via3 ;
        RECT 2629.660 2558.340 2629.980 2558.660 ;
        RECT 2629.660 182.420 2629.980 182.740 ;
      LAYER met4 ;
        RECT 2629.655 2558.335 2629.985 2558.665 ;
        RECT 2629.670 182.745 2629.970 2558.335 ;
        RECT 2629.655 182.415 2629.985 182.745 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 347.905 17.085 348.075 18.615 ;
      LAYER mcon ;
        RECT 347.905 18.445 348.075 18.615 ;
      LAYER met1 ;
        RECT 233.750 3265.260 234.070 3265.320 ;
        RECT 1534.630 3265.260 1534.950 3265.320 ;
        RECT 233.750 3265.120 1534.950 3265.260 ;
        RECT 233.750 3265.060 234.070 3265.120 ;
        RECT 1534.630 3265.060 1534.950 3265.120 ;
        RECT 229.610 262.720 229.930 262.780 ;
        RECT 233.750 262.720 234.070 262.780 ;
        RECT 229.610 262.580 234.070 262.720 ;
        RECT 229.610 262.520 229.930 262.580 ;
        RECT 233.750 262.520 234.070 262.580 ;
        RECT 229.610 244.360 229.930 244.420 ;
        RECT 334.490 244.360 334.810 244.420 ;
        RECT 229.610 244.220 334.810 244.360 ;
        RECT 229.610 244.160 229.930 244.220 ;
        RECT 334.490 244.160 334.810 244.220 ;
        RECT 347.845 18.600 348.135 18.645 ;
        RECT 966.070 18.600 966.390 18.660 ;
        RECT 347.845 18.460 966.390 18.600 ;
        RECT 347.845 18.415 348.135 18.460 ;
        RECT 966.070 18.400 966.390 18.460 ;
        RECT 334.490 17.240 334.810 17.300 ;
        RECT 347.845 17.240 348.135 17.285 ;
        RECT 334.490 17.100 348.135 17.240 ;
        RECT 334.490 17.040 334.810 17.100 ;
        RECT 347.845 17.055 348.135 17.100 ;
      LAYER via ;
        RECT 233.780 3265.060 234.040 3265.320 ;
        RECT 1534.660 3265.060 1534.920 3265.320 ;
        RECT 229.640 262.520 229.900 262.780 ;
        RECT 233.780 262.520 234.040 262.780 ;
        RECT 229.640 244.160 229.900 244.420 ;
        RECT 334.520 244.160 334.780 244.420 ;
        RECT 966.100 18.400 966.360 18.660 ;
        RECT 334.520 17.040 334.780 17.300 ;
      LAYER met2 ;
        RECT 233.780 3265.030 234.040 3265.350 ;
        RECT 1534.660 3265.030 1534.920 3265.350 ;
        RECT 233.840 262.810 233.980 3265.030 ;
        RECT 1534.720 3260.000 1534.860 3265.030 ;
        RECT 1534.610 3256.000 1534.890 3260.000 ;
        RECT 229.640 262.490 229.900 262.810 ;
        RECT 233.780 262.490 234.040 262.810 ;
        RECT 229.700 244.450 229.840 262.490 ;
        RECT 229.640 244.130 229.900 244.450 ;
        RECT 334.520 244.130 334.780 244.450 ;
        RECT 334.580 17.330 334.720 244.130 ;
        RECT 966.100 18.370 966.360 18.690 ;
        RECT 334.520 17.010 334.780 17.330 ;
        RECT 966.160 2.400 966.300 18.370 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 230.530 641.820 230.850 641.880 ;
        RECT 296.770 641.820 297.090 641.880 ;
        RECT 230.530 641.680 297.090 641.820 ;
        RECT 230.530 641.620 230.850 641.680 ;
        RECT 296.770 641.620 297.090 641.680 ;
        RECT 230.530 58.380 230.850 58.440 ;
        RECT 984.010 58.380 984.330 58.440 ;
        RECT 230.530 58.240 984.330 58.380 ;
        RECT 230.530 58.180 230.850 58.240 ;
        RECT 984.010 58.180 984.330 58.240 ;
      LAYER via ;
        RECT 230.560 641.620 230.820 641.880 ;
        RECT 296.800 641.620 297.060 641.880 ;
        RECT 230.560 58.180 230.820 58.440 ;
        RECT 984.040 58.180 984.300 58.440 ;
      LAYER met2 ;
        RECT 296.790 643.435 297.070 643.805 ;
        RECT 296.860 641.910 297.000 643.435 ;
        RECT 230.560 641.590 230.820 641.910 ;
        RECT 296.800 641.590 297.060 641.910 ;
        RECT 230.620 58.470 230.760 641.590 ;
        RECT 230.560 58.150 230.820 58.470 ;
        RECT 984.040 58.150 984.300 58.470 ;
        RECT 984.100 2.400 984.240 58.150 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 296.790 643.480 297.070 643.760 ;
      LAYER met3 ;
        RECT 296.765 643.770 297.095 643.785 ;
        RECT 310.000 643.770 314.000 644.160 ;
        RECT 296.765 643.560 314.000 643.770 ;
        RECT 296.765 643.470 310.500 643.560 ;
        RECT 296.765 643.455 297.095 643.470 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 287.570 1780.480 287.890 1780.540 ;
        RECT 299.530 1780.480 299.850 1780.540 ;
        RECT 287.570 1780.340 299.850 1780.480 ;
        RECT 287.570 1780.280 287.890 1780.340 ;
        RECT 299.530 1780.280 299.850 1780.340 ;
        RECT 287.570 238.580 287.890 238.640 ;
        RECT 662.470 238.580 662.790 238.640 ;
        RECT 287.570 238.440 662.790 238.580 ;
        RECT 287.570 238.380 287.890 238.440 ;
        RECT 662.470 238.380 662.790 238.440 ;
      LAYER via ;
        RECT 287.600 1780.280 287.860 1780.540 ;
        RECT 299.560 1780.280 299.820 1780.540 ;
        RECT 287.600 238.380 287.860 238.640 ;
        RECT 662.500 238.380 662.760 238.640 ;
      LAYER met2 ;
        RECT 299.550 1785.835 299.830 1786.205 ;
        RECT 299.620 1780.570 299.760 1785.835 ;
        RECT 287.600 1780.250 287.860 1780.570 ;
        RECT 299.560 1780.250 299.820 1780.570 ;
        RECT 287.660 238.670 287.800 1780.250 ;
        RECT 287.600 238.350 287.860 238.670 ;
        RECT 662.500 238.350 662.760 238.670 ;
        RECT 662.560 3.130 662.700 238.350 ;
        RECT 662.560 2.990 663.160 3.130 ;
        RECT 663.020 2.400 663.160 2.990 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 299.550 1785.880 299.830 1786.160 ;
      LAYER met3 ;
        RECT 299.525 1786.170 299.855 1786.185 ;
        RECT 310.000 1786.170 314.000 1786.560 ;
        RECT 299.525 1785.960 314.000 1786.170 ;
        RECT 299.525 1785.870 310.500 1785.960 ;
        RECT 299.525 1785.855 299.855 1785.870 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 169.220 1007.330 169.280 ;
        RECT 1421.470 169.220 1421.790 169.280 ;
        RECT 1007.010 169.080 1421.790 169.220 ;
        RECT 1007.010 169.020 1007.330 169.080 ;
        RECT 1421.470 169.020 1421.790 169.080 ;
        RECT 1001.950 15.540 1002.270 15.600 ;
        RECT 1007.010 15.540 1007.330 15.600 ;
        RECT 1001.950 15.400 1007.330 15.540 ;
        RECT 1001.950 15.340 1002.270 15.400 ;
        RECT 1007.010 15.340 1007.330 15.400 ;
      LAYER via ;
        RECT 1007.040 169.020 1007.300 169.280 ;
        RECT 1421.500 169.020 1421.760 169.280 ;
        RECT 1001.980 15.340 1002.240 15.600 ;
        RECT 1007.040 15.340 1007.300 15.600 ;
      LAYER met2 ;
        RECT 1427.890 260.170 1428.170 264.000 ;
        RECT 1421.560 260.030 1428.170 260.170 ;
        RECT 1421.560 169.310 1421.700 260.030 ;
        RECT 1427.890 260.000 1428.170 260.030 ;
        RECT 1007.040 168.990 1007.300 169.310 ;
        RECT 1421.500 168.990 1421.760 169.310 ;
        RECT 1007.100 15.630 1007.240 168.990 ;
        RECT 1001.980 15.310 1002.240 15.630 ;
        RECT 1007.040 15.310 1007.300 15.630 ;
        RECT 1002.040 2.400 1002.180 15.310 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1987.540 2615.490 1987.600 ;
        RECT 2631.270 1987.540 2631.590 1987.600 ;
        RECT 2615.170 1987.400 2631.590 1987.540 ;
        RECT 2615.170 1987.340 2615.490 1987.400 ;
        RECT 2631.270 1987.340 2631.590 1987.400 ;
        RECT 1020.810 114.140 1021.130 114.200 ;
        RECT 2631.270 114.140 2631.590 114.200 ;
        RECT 1020.810 114.000 2631.590 114.140 ;
        RECT 1020.810 113.940 1021.130 114.000 ;
        RECT 2631.270 113.940 2631.590 114.000 ;
      LAYER via ;
        RECT 2615.200 1987.340 2615.460 1987.600 ;
        RECT 2631.300 1987.340 2631.560 1987.600 ;
        RECT 1020.840 113.940 1021.100 114.200 ;
        RECT 2631.300 113.940 2631.560 114.200 ;
      LAYER met2 ;
        RECT 2615.200 1987.485 2615.460 1987.630 ;
        RECT 2615.190 1987.115 2615.470 1987.485 ;
        RECT 2631.300 1987.310 2631.560 1987.630 ;
        RECT 2631.360 114.230 2631.500 1987.310 ;
        RECT 1020.840 113.910 1021.100 114.230 ;
        RECT 2631.300 113.910 2631.560 114.230 ;
        RECT 1020.900 2.960 1021.040 113.910 ;
        RECT 1019.520 2.820 1021.040 2.960 ;
        RECT 1019.520 2.400 1019.660 2.820 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1987.160 2615.470 1987.440 ;
      LAYER met3 ;
        RECT 2606.000 1987.450 2610.000 1987.840 ;
        RECT 2615.165 1987.450 2615.495 1987.465 ;
        RECT 2606.000 1987.240 2615.495 1987.450 ;
        RECT 2609.580 1987.150 2615.495 1987.240 ;
        RECT 2615.165 1987.135 2615.495 1987.150 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1035.605 186.405 1035.775 234.515 ;
      LAYER mcon ;
        RECT 1035.605 234.345 1035.775 234.515 ;
      LAYER met1 ;
        RECT 315.170 3265.600 315.490 3265.660 ;
        RECT 1491.390 3265.600 1491.710 3265.660 ;
        RECT 315.170 3265.460 1491.710 3265.600 ;
        RECT 315.170 3265.400 315.490 3265.460 ;
        RECT 1491.390 3265.400 1491.710 3265.460 ;
        RECT 314.710 336.300 315.030 336.560 ;
        RECT 314.800 335.880 314.940 336.300 ;
        RECT 314.710 335.620 315.030 335.880 ;
        RECT 315.170 252.520 315.490 252.580 ;
        RECT 1035.990 252.520 1036.310 252.580 ;
        RECT 315.170 252.380 1036.310 252.520 ;
        RECT 315.170 252.320 315.490 252.380 ;
        RECT 1035.990 252.320 1036.310 252.380 ;
        RECT 1035.530 234.500 1035.850 234.560 ;
        RECT 1035.335 234.360 1035.850 234.500 ;
        RECT 1035.530 234.300 1035.850 234.360 ;
        RECT 1035.530 186.560 1035.850 186.620 ;
        RECT 1035.335 186.420 1035.850 186.560 ;
        RECT 1035.530 186.360 1035.850 186.420 ;
        RECT 1035.530 137.940 1035.850 138.000 ;
        RECT 1037.370 137.940 1037.690 138.000 ;
        RECT 1035.530 137.800 1037.690 137.940 ;
        RECT 1035.530 137.740 1035.850 137.800 ;
        RECT 1037.370 137.740 1037.690 137.800 ;
      LAYER via ;
        RECT 315.200 3265.400 315.460 3265.660 ;
        RECT 1491.420 3265.400 1491.680 3265.660 ;
        RECT 314.740 336.300 315.000 336.560 ;
        RECT 314.740 335.620 315.000 335.880 ;
        RECT 315.200 252.320 315.460 252.580 ;
        RECT 1036.020 252.320 1036.280 252.580 ;
        RECT 1035.560 234.300 1035.820 234.560 ;
        RECT 1035.560 186.360 1035.820 186.620 ;
        RECT 1035.560 137.740 1035.820 138.000 ;
        RECT 1037.400 137.740 1037.660 138.000 ;
      LAYER met2 ;
        RECT 315.200 3265.370 315.460 3265.690 ;
        RECT 1491.420 3265.370 1491.680 3265.690 ;
        RECT 315.260 337.010 315.400 3265.370 ;
        RECT 1491.480 3260.000 1491.620 3265.370 ;
        RECT 1491.370 3256.000 1491.650 3260.000 ;
        RECT 314.800 336.870 315.400 337.010 ;
        RECT 314.800 336.590 314.940 336.870 ;
        RECT 314.740 336.270 315.000 336.590 ;
        RECT 314.740 335.590 315.000 335.910 ;
        RECT 314.800 314.570 314.940 335.590 ;
        RECT 314.800 314.430 315.400 314.570 ;
        RECT 315.260 252.610 315.400 314.430 ;
        RECT 315.200 252.290 315.460 252.610 ;
        RECT 1036.020 252.290 1036.280 252.610 ;
        RECT 1036.080 241.810 1036.220 252.290 ;
        RECT 1035.620 241.670 1036.220 241.810 ;
        RECT 1035.620 234.590 1035.760 241.670 ;
        RECT 1035.560 234.270 1035.820 234.590 ;
        RECT 1035.560 186.330 1035.820 186.650 ;
        RECT 1035.620 138.030 1035.760 186.330 ;
        RECT 1035.560 137.710 1035.820 138.030 ;
        RECT 1037.400 137.710 1037.660 138.030 ;
        RECT 1037.460 2.400 1037.600 137.710 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.310 128.080 1055.630 128.140 ;
        RECT 2624.830 128.080 2625.150 128.140 ;
        RECT 1055.310 127.940 2625.150 128.080 ;
        RECT 1055.310 127.880 1055.630 127.940 ;
        RECT 2624.830 127.880 2625.150 127.940 ;
      LAYER via ;
        RECT 1055.340 127.880 1055.600 128.140 ;
        RECT 2624.860 127.880 2625.120 128.140 ;
      LAYER met2 ;
        RECT 2624.850 1035.115 2625.130 1035.485 ;
        RECT 2624.920 128.170 2625.060 1035.115 ;
        RECT 1055.340 127.850 1055.600 128.170 ;
        RECT 2624.860 127.850 2625.120 128.170 ;
        RECT 1055.400 2.400 1055.540 127.850 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
      LAYER via2 ;
        RECT 2624.850 1035.160 2625.130 1035.440 ;
      LAYER met3 ;
        RECT 2606.000 1035.450 2610.000 1035.840 ;
        RECT 2624.825 1035.450 2625.155 1035.465 ;
        RECT 2606.000 1035.240 2625.155 1035.450 ;
        RECT 2609.580 1035.150 2625.155 1035.240 ;
        RECT 2624.825 1035.135 2625.155 1035.150 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 224.550 2249.680 224.870 2249.740 ;
        RECT 296.770 2249.680 297.090 2249.740 ;
        RECT 224.550 2249.540 297.090 2249.680 ;
        RECT 224.550 2249.480 224.870 2249.540 ;
        RECT 296.770 2249.480 297.090 2249.540 ;
        RECT 224.550 62.120 224.870 62.180 ;
        RECT 1073.250 62.120 1073.570 62.180 ;
        RECT 224.550 61.980 1073.570 62.120 ;
        RECT 224.550 61.920 224.870 61.980 ;
        RECT 1073.250 61.920 1073.570 61.980 ;
      LAYER via ;
        RECT 224.580 2249.480 224.840 2249.740 ;
        RECT 296.800 2249.480 297.060 2249.740 ;
        RECT 224.580 61.920 224.840 62.180 ;
        RECT 1073.280 61.920 1073.540 62.180 ;
      LAYER met2 ;
        RECT 296.790 2250.955 297.070 2251.325 ;
        RECT 296.860 2249.770 297.000 2250.955 ;
        RECT 224.580 2249.450 224.840 2249.770 ;
        RECT 296.800 2249.450 297.060 2249.770 ;
        RECT 224.640 62.210 224.780 2249.450 ;
        RECT 224.580 61.890 224.840 62.210 ;
        RECT 1073.280 61.890 1073.540 62.210 ;
        RECT 1073.340 2.400 1073.480 61.890 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 296.790 2251.000 297.070 2251.280 ;
      LAYER met3 ;
        RECT 296.765 2251.290 297.095 2251.305 ;
        RECT 310.000 2251.290 314.000 2251.680 ;
        RECT 296.765 2251.080 314.000 2251.290 ;
        RECT 296.765 2250.990 310.500 2251.080 ;
        RECT 296.765 2250.975 297.095 2250.990 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2450.960 2615.490 2451.020 ;
        RECT 2630.350 2450.960 2630.670 2451.020 ;
        RECT 2615.170 2450.820 2630.670 2450.960 ;
        RECT 2615.170 2450.760 2615.490 2450.820 ;
        RECT 2630.350 2450.760 2630.670 2450.820 ;
        RECT 1096.710 225.660 1097.030 225.720 ;
        RECT 2630.350 225.660 2630.670 225.720 ;
        RECT 1096.710 225.520 2630.670 225.660 ;
        RECT 1096.710 225.460 1097.030 225.520 ;
        RECT 2630.350 225.460 2630.670 225.520 ;
        RECT 1090.730 16.560 1091.050 16.620 ;
        RECT 1096.710 16.560 1097.030 16.620 ;
        RECT 1090.730 16.420 1097.030 16.560 ;
        RECT 1090.730 16.360 1091.050 16.420 ;
        RECT 1096.710 16.360 1097.030 16.420 ;
      LAYER via ;
        RECT 2615.200 2450.760 2615.460 2451.020 ;
        RECT 2630.380 2450.760 2630.640 2451.020 ;
        RECT 1096.740 225.460 1097.000 225.720 ;
        RECT 2630.380 225.460 2630.640 225.720 ;
        RECT 1090.760 16.360 1091.020 16.620 ;
        RECT 1096.740 16.360 1097.000 16.620 ;
      LAYER met2 ;
        RECT 2615.190 2452.235 2615.470 2452.605 ;
        RECT 2615.260 2451.050 2615.400 2452.235 ;
        RECT 2615.200 2450.730 2615.460 2451.050 ;
        RECT 2630.380 2450.730 2630.640 2451.050 ;
        RECT 2630.440 225.750 2630.580 2450.730 ;
        RECT 1096.740 225.430 1097.000 225.750 ;
        RECT 2630.380 225.430 2630.640 225.750 ;
        RECT 1096.800 16.650 1096.940 225.430 ;
        RECT 1090.760 16.330 1091.020 16.650 ;
        RECT 1096.740 16.330 1097.000 16.650 ;
        RECT 1090.820 2.400 1090.960 16.330 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2452.280 2615.470 2452.560 ;
      LAYER met3 ;
        RECT 2606.000 2452.570 2610.000 2452.960 ;
        RECT 2615.165 2452.570 2615.495 2452.585 ;
        RECT 2606.000 2452.360 2615.495 2452.570 ;
        RECT 2609.580 2452.270 2615.495 2452.360 ;
        RECT 2615.165 2452.255 2615.495 2452.270 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1108.670 34.240 1108.990 34.300 ;
        RECT 1393.870 34.240 1394.190 34.300 ;
        RECT 1108.670 34.100 1394.190 34.240 ;
        RECT 1108.670 34.040 1108.990 34.100 ;
        RECT 1393.870 34.040 1394.190 34.100 ;
      LAYER via ;
        RECT 1108.700 34.040 1108.960 34.300 ;
        RECT 1393.900 34.040 1394.160 34.300 ;
      LAYER met2 ;
        RECT 1399.370 260.170 1399.650 264.000 ;
        RECT 1393.960 260.030 1399.650 260.170 ;
        RECT 1393.960 34.330 1394.100 260.030 ;
        RECT 1399.370 260.000 1399.650 260.030 ;
        RECT 1108.700 34.010 1108.960 34.330 ;
        RECT 1393.900 34.010 1394.160 34.330 ;
        RECT 1108.760 2.400 1108.900 34.010 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.710 190.300 1028.030 190.360 ;
        RECT 1124.770 190.300 1125.090 190.360 ;
        RECT 1027.710 190.160 1125.090 190.300 ;
        RECT 1027.710 190.100 1028.030 190.160 ;
        RECT 1124.770 190.100 1125.090 190.160 ;
      LAYER via ;
        RECT 1027.740 190.100 1028.000 190.360 ;
        RECT 1124.800 190.100 1125.060 190.360 ;
      LAYER met2 ;
        RECT 1027.690 260.000 1027.970 264.000 ;
        RECT 1027.800 190.390 1027.940 260.000 ;
        RECT 1027.740 190.070 1028.000 190.390 ;
        RECT 1124.800 190.070 1125.060 190.390 ;
        RECT 1124.860 3.130 1125.000 190.070 ;
        RECT 1124.860 2.990 1126.840 3.130 ;
        RECT 1126.700 2.400 1126.840 2.990 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1144.550 148.480 1144.870 148.540 ;
        RECT 2617.930 148.480 2618.250 148.540 ;
        RECT 1144.550 148.340 2618.250 148.480 ;
        RECT 1144.550 148.280 1144.870 148.340 ;
        RECT 2617.930 148.280 2618.250 148.340 ;
      LAYER via ;
        RECT 1144.580 148.280 1144.840 148.540 ;
        RECT 2617.960 148.280 2618.220 148.540 ;
      LAYER met2 ;
        RECT 2617.950 655.675 2618.230 656.045 ;
        RECT 2618.020 148.570 2618.160 655.675 ;
        RECT 1144.580 148.250 1144.840 148.570 ;
        RECT 2617.960 148.250 2618.220 148.570 ;
        RECT 1144.640 2.400 1144.780 148.250 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
      LAYER via2 ;
        RECT 2617.950 655.720 2618.230 656.000 ;
      LAYER met3 ;
        RECT 2606.000 656.010 2610.000 656.400 ;
        RECT 2617.925 656.010 2618.255 656.025 ;
        RECT 2606.000 655.800 2618.255 656.010 ;
        RECT 2609.580 655.710 2618.255 655.800 ;
        RECT 2617.925 655.695 2618.255 655.710 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 61.440 1162.810 61.500 ;
        RECT 1621.570 61.440 1621.890 61.500 ;
        RECT 1162.490 61.300 1621.890 61.440 ;
        RECT 1162.490 61.240 1162.810 61.300 ;
        RECT 1621.570 61.240 1621.890 61.300 ;
      LAYER via ;
        RECT 1162.520 61.240 1162.780 61.500 ;
        RECT 1621.600 61.240 1621.860 61.500 ;
      LAYER met2 ;
        RECT 1627.530 260.170 1627.810 264.000 ;
        RECT 1621.660 260.030 1627.810 260.170 ;
        RECT 1621.660 61.530 1621.800 260.030 ;
        RECT 1627.530 260.000 1627.810 260.030 ;
        RECT 1162.520 61.210 1162.780 61.530 ;
        RECT 1621.600 61.210 1621.860 61.530 ;
        RECT 1162.580 2.400 1162.720 61.210 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 189.960 683.030 190.020 ;
        RECT 2617.470 189.960 2617.790 190.020 ;
        RECT 682.710 189.820 2617.790 189.960 ;
        RECT 682.710 189.760 683.030 189.820 ;
        RECT 2617.470 189.760 2617.790 189.820 ;
        RECT 680.410 20.640 680.730 20.700 ;
        RECT 682.710 20.640 683.030 20.700 ;
        RECT 680.410 20.500 683.030 20.640 ;
        RECT 680.410 20.440 680.730 20.500 ;
        RECT 682.710 20.440 683.030 20.500 ;
      LAYER via ;
        RECT 682.740 189.760 683.000 190.020 ;
        RECT 2617.500 189.760 2617.760 190.020 ;
        RECT 680.440 20.440 680.700 20.700 ;
        RECT 682.740 20.440 683.000 20.700 ;
      LAYER met2 ;
        RECT 2617.490 888.235 2617.770 888.605 ;
        RECT 2617.560 190.050 2617.700 888.235 ;
        RECT 682.740 189.730 683.000 190.050 ;
        RECT 2617.500 189.730 2617.760 190.050 ;
        RECT 682.800 20.730 682.940 189.730 ;
        RECT 680.440 20.410 680.700 20.730 ;
        RECT 682.740 20.410 683.000 20.730 ;
        RECT 680.500 2.400 680.640 20.410 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 2617.490 888.280 2617.770 888.560 ;
      LAYER met3 ;
        RECT 2606.000 888.570 2610.000 888.960 ;
        RECT 2617.465 888.570 2617.795 888.585 ;
        RECT 2606.000 888.360 2617.795 888.570 ;
        RECT 2609.580 888.270 2617.795 888.360 ;
        RECT 2617.465 888.255 2617.795 888.270 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 176.020 1186.730 176.080 ;
        RECT 1642.270 176.020 1642.590 176.080 ;
        RECT 1186.410 175.880 1642.590 176.020 ;
        RECT 1186.410 175.820 1186.730 175.880 ;
        RECT 1642.270 175.820 1642.590 175.880 ;
        RECT 1179.970 16.900 1180.290 16.960 ;
        RECT 1186.410 16.900 1186.730 16.960 ;
        RECT 1179.970 16.760 1186.730 16.900 ;
        RECT 1179.970 16.700 1180.290 16.760 ;
        RECT 1186.410 16.700 1186.730 16.760 ;
      LAYER via ;
        RECT 1186.440 175.820 1186.700 176.080 ;
        RECT 1642.300 175.820 1642.560 176.080 ;
        RECT 1180.000 16.700 1180.260 16.960 ;
        RECT 1186.440 16.700 1186.700 16.960 ;
      LAYER met2 ;
        RECT 1642.250 260.000 1642.530 264.000 ;
        RECT 1642.360 176.110 1642.500 260.000 ;
        RECT 1186.440 175.790 1186.700 176.110 ;
        RECT 1642.300 175.790 1642.560 176.110 ;
        RECT 1186.500 16.990 1186.640 175.790 ;
        RECT 1180.000 16.670 1180.260 16.990 ;
        RECT 1186.440 16.670 1186.700 16.990 ;
        RECT 1180.060 2.400 1180.200 16.670 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 246.060 1200.530 246.120 ;
        RECT 2070.990 246.060 2071.310 246.120 ;
        RECT 1200.210 245.920 2071.310 246.060 ;
        RECT 1200.210 245.860 1200.530 245.920 ;
        RECT 2070.990 245.860 2071.310 245.920 ;
        RECT 1197.910 20.640 1198.230 20.700 ;
        RECT 1200.210 20.640 1200.530 20.700 ;
        RECT 1197.910 20.500 1200.530 20.640 ;
        RECT 1197.910 20.440 1198.230 20.500 ;
        RECT 1200.210 20.440 1200.530 20.500 ;
      LAYER via ;
        RECT 1200.240 245.860 1200.500 246.120 ;
        RECT 2071.020 245.860 2071.280 246.120 ;
        RECT 1197.940 20.440 1198.200 20.700 ;
        RECT 1200.240 20.440 1200.500 20.700 ;
      LAYER met2 ;
        RECT 2070.970 260.000 2071.250 264.000 ;
        RECT 2071.080 246.150 2071.220 260.000 ;
        RECT 1200.240 245.830 1200.500 246.150 ;
        RECT 2071.020 245.830 2071.280 246.150 ;
        RECT 1200.300 20.730 1200.440 245.830 ;
        RECT 1197.940 20.410 1198.200 20.730 ;
        RECT 1200.240 20.410 1200.500 20.730 ;
        RECT 1198.000 2.400 1198.140 20.410 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1215.925 48.365 1216.095 80.155 ;
      LAYER mcon ;
        RECT 1215.925 79.985 1216.095 80.155 ;
      LAYER met1 ;
        RECT 326.670 241.640 326.990 241.700 ;
        RECT 334.950 241.640 335.270 241.700 ;
        RECT 326.670 241.500 335.270 241.640 ;
        RECT 326.670 241.440 326.990 241.500 ;
        RECT 334.950 241.440 335.270 241.500 ;
        RECT 334.950 80.140 335.270 80.200 ;
        RECT 1215.865 80.140 1216.155 80.185 ;
        RECT 334.950 80.000 1216.155 80.140 ;
        RECT 334.950 79.940 335.270 80.000 ;
        RECT 1215.865 79.955 1216.155 80.000 ;
        RECT 1215.850 48.520 1216.170 48.580 ;
        RECT 1215.655 48.380 1216.170 48.520 ;
        RECT 1215.850 48.320 1216.170 48.380 ;
      LAYER via ;
        RECT 326.700 241.440 326.960 241.700 ;
        RECT 334.980 241.440 335.240 241.700 ;
        RECT 334.980 79.940 335.240 80.200 ;
        RECT 1215.880 48.320 1216.140 48.580 ;
      LAYER met2 ;
        RECT 326.650 260.000 326.930 264.000 ;
        RECT 326.760 241.730 326.900 260.000 ;
        RECT 326.700 241.410 326.960 241.730 ;
        RECT 334.980 241.410 335.240 241.730 ;
        RECT 335.040 80.230 335.180 241.410 ;
        RECT 334.980 79.910 335.240 80.230 ;
        RECT 1215.880 48.290 1216.140 48.610 ;
        RECT 1215.940 2.400 1216.080 48.290 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1997.390 246.740 1997.710 246.800 ;
        RECT 2514.430 246.740 2514.750 246.800 ;
        RECT 1997.390 246.600 2514.750 246.740 ;
        RECT 1997.390 246.540 1997.710 246.600 ;
        RECT 2514.430 246.540 2514.750 246.600 ;
        RECT 1233.790 51.920 1234.110 51.980 ;
        RECT 1997.390 51.920 1997.710 51.980 ;
        RECT 1233.790 51.780 1997.710 51.920 ;
        RECT 1233.790 51.720 1234.110 51.780 ;
        RECT 1997.390 51.720 1997.710 51.780 ;
      LAYER via ;
        RECT 1997.420 246.540 1997.680 246.800 ;
        RECT 2514.460 246.540 2514.720 246.800 ;
        RECT 1233.820 51.720 1234.080 51.980 ;
        RECT 1997.420 51.720 1997.680 51.980 ;
      LAYER met2 ;
        RECT 2514.410 260.000 2514.690 264.000 ;
        RECT 2514.520 246.830 2514.660 260.000 ;
        RECT 1997.420 246.510 1997.680 246.830 ;
        RECT 2514.460 246.510 2514.720 246.830 ;
        RECT 1997.480 52.010 1997.620 246.510 ;
        RECT 1233.820 51.690 1234.080 52.010 ;
        RECT 1997.420 51.690 1997.680 52.010 ;
        RECT 1233.880 2.400 1234.020 51.690 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 217.840 1255.730 217.900 ;
        RECT 2618.390 217.840 2618.710 217.900 ;
        RECT 1255.410 217.700 2618.710 217.840 ;
        RECT 1255.410 217.640 1255.730 217.700 ;
        RECT 2618.390 217.640 2618.710 217.700 ;
        RECT 1251.730 20.640 1252.050 20.700 ;
        RECT 1255.410 20.640 1255.730 20.700 ;
        RECT 1251.730 20.500 1255.730 20.640 ;
        RECT 1251.730 20.440 1252.050 20.500 ;
        RECT 1255.410 20.440 1255.730 20.500 ;
      LAYER via ;
        RECT 1255.440 217.640 1255.700 217.900 ;
        RECT 2618.420 217.640 2618.680 217.900 ;
        RECT 1251.760 20.440 1252.020 20.700 ;
        RECT 1255.440 20.440 1255.700 20.700 ;
      LAYER met2 ;
        RECT 2618.410 549.595 2618.690 549.965 ;
        RECT 2618.480 217.930 2618.620 549.595 ;
        RECT 1255.440 217.610 1255.700 217.930 ;
        RECT 2618.420 217.610 2618.680 217.930 ;
        RECT 1255.500 20.730 1255.640 217.610 ;
        RECT 1251.760 20.410 1252.020 20.730 ;
        RECT 1255.440 20.410 1255.700 20.730 ;
        RECT 1251.820 2.400 1251.960 20.410 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
      LAYER via2 ;
        RECT 2618.410 549.640 2618.690 549.920 ;
      LAYER met3 ;
        RECT 2606.000 549.930 2610.000 550.320 ;
        RECT 2618.385 549.930 2618.715 549.945 ;
        RECT 2606.000 549.720 2618.715 549.930 ;
        RECT 2609.580 549.630 2618.715 549.720 ;
        RECT 2618.385 549.615 2618.715 549.630 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 254.450 3275.460 254.770 3275.520 ;
        RECT 633.950 3275.460 634.270 3275.520 ;
        RECT 254.450 3275.320 634.270 3275.460 ;
        RECT 254.450 3275.260 254.770 3275.320 ;
        RECT 633.950 3275.260 634.270 3275.320 ;
        RECT 254.450 44.440 254.770 44.500 ;
        RECT 1268.290 44.440 1268.610 44.500 ;
        RECT 254.450 44.300 1268.610 44.440 ;
        RECT 254.450 44.240 254.770 44.300 ;
        RECT 1268.290 44.240 1268.610 44.300 ;
      LAYER via ;
        RECT 254.480 3275.260 254.740 3275.520 ;
        RECT 633.980 3275.260 634.240 3275.520 ;
        RECT 254.480 44.240 254.740 44.500 ;
        RECT 1268.320 44.240 1268.580 44.500 ;
      LAYER met2 ;
        RECT 254.480 3275.230 254.740 3275.550 ;
        RECT 633.980 3275.230 634.240 3275.550 ;
        RECT 254.540 44.530 254.680 3275.230 ;
        RECT 634.040 3260.000 634.180 3275.230 ;
        RECT 633.930 3256.000 634.210 3260.000 ;
        RECT 254.480 44.210 254.740 44.530 ;
        RECT 1268.320 44.210 1268.580 44.530 ;
        RECT 1268.380 14.010 1268.520 44.210 ;
        RECT 1268.380 13.870 1269.440 14.010 ;
        RECT 1269.300 2.400 1269.440 13.870 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 3260.500 264.430 3260.560 ;
        RECT 433.390 3260.500 433.710 3260.560 ;
        RECT 264.110 3260.360 433.710 3260.500 ;
        RECT 264.110 3260.300 264.430 3260.360 ;
        RECT 433.390 3260.300 433.710 3260.360 ;
      LAYER via ;
        RECT 264.140 3260.300 264.400 3260.560 ;
        RECT 433.420 3260.300 433.680 3260.560 ;
      LAYER met2 ;
        RECT 264.140 3260.270 264.400 3260.590 ;
        RECT 433.420 3260.270 433.680 3260.590 ;
        RECT 264.200 61.045 264.340 3260.270 ;
        RECT 433.480 3260.000 433.620 3260.270 ;
        RECT 433.370 3256.000 433.650 3260.000 ;
        RECT 264.130 60.675 264.410 61.045 ;
        RECT 1287.170 60.675 1287.450 61.045 ;
        RECT 1287.240 2.400 1287.380 60.675 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
      LAYER via2 ;
        RECT 264.130 60.720 264.410 61.000 ;
        RECT 1287.170 60.720 1287.450 61.000 ;
      LAYER met3 ;
        RECT 264.105 61.010 264.435 61.025 ;
        RECT 1287.145 61.010 1287.475 61.025 ;
        RECT 264.105 60.710 1287.475 61.010 ;
        RECT 264.105 60.695 264.435 60.710 ;
        RECT 1287.145 60.695 1287.475 60.710 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.170 14.180 1304.490 14.240 ;
        RECT 1304.170 14.040 1305.320 14.180 ;
        RECT 1304.170 13.980 1304.490 14.040 ;
        RECT 1305.180 13.900 1305.320 14.040 ;
        RECT 1305.090 13.640 1305.410 13.900 ;
      LAYER via ;
        RECT 1304.200 13.980 1304.460 14.240 ;
        RECT 1305.120 13.640 1305.380 13.900 ;
      LAYER met2 ;
        RECT 1304.190 154.515 1304.470 154.885 ;
        RECT 1304.260 14.270 1304.400 154.515 ;
        RECT 1304.200 13.950 1304.460 14.270 ;
        RECT 1305.120 13.610 1305.380 13.930 ;
        RECT 1305.180 2.400 1305.320 13.610 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
      LAYER via2 ;
        RECT 1304.190 154.560 1304.470 154.840 ;
      LAYER met3 ;
        RECT 289.150 3053.690 289.530 3053.700 ;
        RECT 310.000 3053.690 314.000 3054.080 ;
        RECT 289.150 3053.480 314.000 3053.690 ;
        RECT 289.150 3053.390 310.500 3053.480 ;
        RECT 289.150 3053.380 289.530 3053.390 ;
        RECT 289.150 154.850 289.530 154.860 ;
        RECT 1304.165 154.850 1304.495 154.865 ;
        RECT 289.150 154.550 1304.495 154.850 ;
        RECT 289.150 154.540 289.530 154.550 ;
        RECT 1304.165 154.535 1304.495 154.550 ;
      LAYER via3 ;
        RECT 289.180 3053.380 289.500 3053.700 ;
        RECT 289.180 154.540 289.500 154.860 ;
      LAYER met4 ;
        RECT 289.175 3053.375 289.505 3053.705 ;
        RECT 289.190 154.865 289.490 3053.375 ;
        RECT 289.175 154.535 289.505 154.865 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 238.350 2139.180 238.670 2139.240 ;
        RECT 296.770 2139.180 297.090 2139.240 ;
        RECT 238.350 2139.040 297.090 2139.180 ;
        RECT 238.350 2138.980 238.670 2139.040 ;
        RECT 296.770 2138.980 297.090 2139.040 ;
        RECT 238.350 60.760 238.670 60.820 ;
        RECT 1323.030 60.760 1323.350 60.820 ;
        RECT 238.350 60.620 1323.350 60.760 ;
        RECT 238.350 60.560 238.670 60.620 ;
        RECT 1323.030 60.560 1323.350 60.620 ;
      LAYER via ;
        RECT 238.380 2138.980 238.640 2139.240 ;
        RECT 296.800 2138.980 297.060 2139.240 ;
        RECT 238.380 60.560 238.640 60.820 ;
        RECT 1323.060 60.560 1323.320 60.820 ;
      LAYER met2 ;
        RECT 296.790 2144.875 297.070 2145.245 ;
        RECT 296.860 2139.270 297.000 2144.875 ;
        RECT 238.380 2138.950 238.640 2139.270 ;
        RECT 296.800 2138.950 297.060 2139.270 ;
        RECT 238.440 60.850 238.580 2138.950 ;
        RECT 238.380 60.530 238.640 60.850 ;
        RECT 1323.060 60.530 1323.320 60.850 ;
        RECT 1323.120 2.400 1323.260 60.530 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
      LAYER via2 ;
        RECT 296.790 2144.920 297.070 2145.200 ;
      LAYER met3 ;
        RECT 296.765 2145.210 297.095 2145.225 ;
        RECT 310.000 2145.210 314.000 2145.600 ;
        RECT 296.765 2145.000 314.000 2145.210 ;
        RECT 296.765 2144.910 310.500 2145.000 ;
        RECT 296.765 2144.895 297.095 2144.910 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1338.745 144.925 1338.915 193.035 ;
        RECT 1338.745 48.365 1338.915 96.475 ;
      LAYER mcon ;
        RECT 1338.745 192.865 1338.915 193.035 ;
        RECT 1338.745 96.305 1338.915 96.475 ;
      LAYER met1 ;
        RECT 280.210 1573.420 280.530 1573.480 ;
        RECT 296.770 1573.420 297.090 1573.480 ;
        RECT 280.210 1573.280 297.090 1573.420 ;
        RECT 280.210 1573.220 280.530 1573.280 ;
        RECT 296.770 1573.220 297.090 1573.280 ;
        RECT 280.210 212.400 280.530 212.460 ;
        RECT 1338.670 212.400 1338.990 212.460 ;
        RECT 280.210 212.260 1338.990 212.400 ;
        RECT 280.210 212.200 280.530 212.260 ;
        RECT 1338.670 212.200 1338.990 212.260 ;
        RECT 1338.670 193.020 1338.990 193.080 ;
        RECT 1338.475 192.880 1338.990 193.020 ;
        RECT 1338.670 192.820 1338.990 192.880 ;
        RECT 1338.670 145.080 1338.990 145.140 ;
        RECT 1338.475 144.940 1338.990 145.080 ;
        RECT 1338.670 144.880 1338.990 144.940 ;
        RECT 1338.670 96.460 1338.990 96.520 ;
        RECT 1338.475 96.320 1338.990 96.460 ;
        RECT 1338.670 96.260 1338.990 96.320 ;
        RECT 1338.670 48.520 1338.990 48.580 ;
        RECT 1338.475 48.380 1338.990 48.520 ;
        RECT 1338.670 48.320 1338.990 48.380 ;
      LAYER via ;
        RECT 280.240 1573.220 280.500 1573.480 ;
        RECT 296.800 1573.220 297.060 1573.480 ;
        RECT 280.240 212.200 280.500 212.460 ;
        RECT 1338.700 212.200 1338.960 212.460 ;
        RECT 1338.700 192.820 1338.960 193.080 ;
        RECT 1338.700 144.880 1338.960 145.140 ;
        RECT 1338.700 96.260 1338.960 96.520 ;
        RECT 1338.700 48.320 1338.960 48.580 ;
      LAYER met2 ;
        RECT 296.790 1573.675 297.070 1574.045 ;
        RECT 296.860 1573.510 297.000 1573.675 ;
        RECT 280.240 1573.190 280.500 1573.510 ;
        RECT 296.800 1573.190 297.060 1573.510 ;
        RECT 280.300 212.490 280.440 1573.190 ;
        RECT 280.240 212.170 280.500 212.490 ;
        RECT 1338.700 212.170 1338.960 212.490 ;
        RECT 1338.760 193.110 1338.900 212.170 ;
        RECT 1338.700 192.790 1338.960 193.110 ;
        RECT 1338.700 144.850 1338.960 145.170 ;
        RECT 1338.760 96.550 1338.900 144.850 ;
        RECT 1338.700 96.230 1338.960 96.550 ;
        RECT 1338.700 48.290 1338.960 48.610 ;
        RECT 1338.760 12.650 1338.900 48.290 ;
        RECT 1338.760 12.510 1340.740 12.650 ;
        RECT 1340.600 2.400 1340.740 12.510 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
      LAYER via2 ;
        RECT 296.790 1573.720 297.070 1574.000 ;
      LAYER met3 ;
        RECT 296.765 1574.010 297.095 1574.025 ;
        RECT 310.000 1574.010 314.000 1574.400 ;
        RECT 296.765 1573.800 314.000 1574.010 ;
        RECT 296.765 1573.710 310.500 1573.800 ;
        RECT 296.765 1573.695 297.095 1573.710 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2606.910 2456.995 2607.190 2457.365 ;
        RECT 2606.980 2409.085 2607.120 2456.995 ;
        RECT 2606.910 2408.715 2607.190 2409.085 ;
        RECT 2607.830 1341.115 2608.110 1341.485 ;
        RECT 2607.900 1304.085 2608.040 1341.115 ;
        RECT 2607.830 1303.715 2608.110 1304.085 ;
        RECT 2607.830 1249.315 2608.110 1249.685 ;
        RECT 2607.900 1211.605 2608.040 1249.315 ;
        RECT 2607.830 1211.235 2608.110 1211.605 ;
        RECT 698.370 32.795 698.650 33.165 ;
        RECT 1011.170 33.050 1011.450 33.165 ;
        RECT 1013.930 33.050 1014.210 33.165 ;
        RECT 1011.170 32.910 1014.210 33.050 ;
        RECT 1011.170 32.795 1011.450 32.910 ;
        RECT 1013.930 32.795 1014.210 32.910 ;
        RECT 698.440 2.400 698.580 32.795 ;
        RECT 698.230 -4.800 698.790 2.400 ;
      LAYER via2 ;
        RECT 2606.910 2457.040 2607.190 2457.320 ;
        RECT 2606.910 2408.760 2607.190 2409.040 ;
        RECT 2607.830 1341.160 2608.110 1341.440 ;
        RECT 2607.830 1303.760 2608.110 1304.040 ;
        RECT 2607.830 1249.360 2608.110 1249.640 ;
        RECT 2607.830 1211.280 2608.110 1211.560 ;
        RECT 698.370 32.840 698.650 33.120 ;
        RECT 1011.170 32.840 1011.450 33.120 ;
        RECT 1013.930 32.840 1014.210 33.120 ;
      LAYER met3 ;
        RECT 2606.000 2494.520 2610.000 2495.120 ;
        RECT 2607.590 2492.020 2607.890 2494.520 ;
        RECT 2607.550 2491.700 2607.930 2492.020 ;
        RECT 2606.885 2457.330 2607.215 2457.345 ;
        RECT 2607.550 2457.330 2607.930 2457.340 ;
        RECT 2606.885 2457.030 2607.930 2457.330 ;
        RECT 2606.885 2457.015 2607.215 2457.030 ;
        RECT 2607.550 2457.020 2607.930 2457.030 ;
        RECT 2606.885 2409.060 2607.215 2409.065 ;
        RECT 2606.630 2409.050 2607.215 2409.060 ;
        RECT 2606.430 2408.750 2607.215 2409.050 ;
        RECT 2606.630 2408.740 2607.215 2408.750 ;
        RECT 2606.885 2408.735 2607.215 2408.740 ;
        RECT 2606.630 1341.450 2607.010 1341.460 ;
        RECT 2607.805 1341.450 2608.135 1341.465 ;
        RECT 2606.630 1341.150 2608.135 1341.450 ;
        RECT 2606.630 1341.140 2607.010 1341.150 ;
        RECT 2607.805 1341.135 2608.135 1341.150 ;
        RECT 2606.630 1304.050 2607.010 1304.060 ;
        RECT 2607.805 1304.050 2608.135 1304.065 ;
        RECT 2606.630 1303.750 2608.135 1304.050 ;
        RECT 2606.630 1303.740 2607.010 1303.750 ;
        RECT 2607.805 1303.735 2608.135 1303.750 ;
        RECT 2606.630 1249.650 2607.010 1249.660 ;
        RECT 2607.805 1249.650 2608.135 1249.665 ;
        RECT 2606.630 1249.350 2608.135 1249.650 ;
        RECT 2606.630 1249.340 2607.010 1249.350 ;
        RECT 2607.805 1249.335 2608.135 1249.350 ;
        RECT 2607.805 1211.570 2608.135 1211.585 ;
        RECT 2606.670 1211.270 2608.135 1211.570 ;
        RECT 2606.670 1210.900 2606.970 1211.270 ;
        RECT 2607.805 1211.255 2608.135 1211.270 ;
        RECT 2606.630 1210.580 2607.010 1210.900 ;
        RECT 2606.630 1120.450 2607.010 1120.460 ;
        RECT 2612.150 1120.450 2612.530 1120.460 ;
        RECT 2606.630 1120.150 2612.530 1120.450 ;
        RECT 2606.630 1120.140 2607.010 1120.150 ;
        RECT 2612.150 1120.140 2612.530 1120.150 ;
        RECT 2601.110 243.250 2601.490 243.260 ;
        RECT 2604.790 243.250 2605.170 243.260 ;
        RECT 2601.110 242.950 2605.170 243.250 ;
        RECT 2601.110 242.940 2601.490 242.950 ;
        RECT 2604.790 242.940 2605.170 242.950 ;
        RECT 2601.110 181.370 2601.490 181.380 ;
        RECT 2603.870 181.370 2604.250 181.380 ;
        RECT 2601.110 181.070 2604.250 181.370 ;
        RECT 2601.110 181.060 2601.490 181.070 ;
        RECT 2603.870 181.060 2604.250 181.070 ;
        RECT 1707.830 33.510 1730.210 33.810 ;
        RECT 698.345 33.130 698.675 33.145 ;
        RECT 1011.145 33.130 1011.475 33.145 ;
        RECT 698.345 32.830 1011.475 33.130 ;
        RECT 698.345 32.815 698.675 32.830 ;
        RECT 1011.145 32.815 1011.475 32.830 ;
        RECT 1013.905 33.130 1014.235 33.145 ;
        RECT 1707.830 33.130 1708.130 33.510 ;
        RECT 1013.905 32.830 1708.130 33.130 ;
        RECT 1729.910 33.130 1730.210 33.510 ;
        RECT 2602.030 33.130 2602.410 33.140 ;
        RECT 1729.910 32.830 2602.410 33.130 ;
        RECT 1013.905 32.815 1014.235 32.830 ;
        RECT 2602.030 32.820 2602.410 32.830 ;
      LAYER via3 ;
        RECT 2607.580 2491.700 2607.900 2492.020 ;
        RECT 2607.580 2457.020 2607.900 2457.340 ;
        RECT 2606.660 2408.740 2606.980 2409.060 ;
        RECT 2606.660 1341.140 2606.980 1341.460 ;
        RECT 2606.660 1303.740 2606.980 1304.060 ;
        RECT 2606.660 1249.340 2606.980 1249.660 ;
        RECT 2606.660 1210.580 2606.980 1210.900 ;
        RECT 2606.660 1120.140 2606.980 1120.460 ;
        RECT 2612.180 1120.140 2612.500 1120.460 ;
        RECT 2601.140 242.940 2601.460 243.260 ;
        RECT 2604.820 242.940 2605.140 243.260 ;
        RECT 2601.140 181.060 2601.460 181.380 ;
        RECT 2603.900 181.060 2604.220 181.380 ;
        RECT 2602.060 32.820 2602.380 33.140 ;
      LAYER met4 ;
        RECT 2607.575 2491.695 2607.905 2492.025 ;
        RECT 2607.590 2457.345 2607.890 2491.695 ;
        RECT 2607.575 2457.015 2607.905 2457.345 ;
        RECT 2600.710 2408.310 2601.890 2409.490 ;
        RECT 2606.230 2408.310 2607.410 2409.490 ;
        RECT 2601.150 2344.450 2601.450 2408.310 ;
        RECT 2601.150 2344.150 2602.370 2344.450 ;
        RECT 2602.070 2341.050 2602.370 2344.150 ;
        RECT 2602.070 2340.750 2603.290 2341.050 ;
        RECT 2602.990 2279.850 2603.290 2340.750 ;
        RECT 2602.070 2279.550 2603.290 2279.850 ;
        RECT 2602.070 2225.450 2602.370 2279.550 ;
        RECT 2602.070 2225.150 2604.210 2225.450 ;
        RECT 2603.910 2215.250 2604.210 2225.150 ;
        RECT 2602.070 2214.950 2604.210 2215.250 ;
        RECT 2602.070 2140.450 2602.370 2214.950 ;
        RECT 2602.070 2140.150 2603.290 2140.450 ;
        RECT 2602.990 2065.650 2603.290 2140.150 ;
        RECT 2601.150 2065.350 2603.290 2065.650 ;
        RECT 2601.150 2014.650 2601.450 2065.350 ;
        RECT 2601.150 2014.350 2602.370 2014.650 ;
        RECT 2602.070 1913.090 2602.370 2014.350 ;
        RECT 2601.630 1911.910 2602.810 1913.090 ;
        RECT 2606.230 1911.910 2607.410 1913.090 ;
        RECT 2606.670 1872.290 2606.970 1911.910 ;
        RECT 2600.710 1871.110 2601.890 1872.290 ;
        RECT 2606.230 1871.110 2607.410 1872.290 ;
        RECT 2601.150 1841.250 2601.450 1871.110 ;
        RECT 2601.150 1840.950 2602.370 1841.250 ;
        RECT 2602.070 1810.650 2602.370 1840.950 ;
        RECT 2601.150 1810.350 2602.370 1810.650 ;
        RECT 2601.150 1766.450 2601.450 1810.350 ;
        RECT 2601.150 1766.150 2602.370 1766.450 ;
        RECT 2602.070 1715.450 2602.370 1766.150 ;
        RECT 2599.310 1715.150 2602.370 1715.450 ;
        RECT 2599.310 1674.650 2599.610 1715.150 ;
        RECT 2599.310 1674.350 2602.370 1674.650 ;
        RECT 2602.070 1661.050 2602.370 1674.350 ;
        RECT 2601.150 1660.750 2602.370 1661.050 ;
        RECT 2601.150 1603.250 2601.450 1660.750 ;
        RECT 2601.150 1602.950 2602.370 1603.250 ;
        RECT 2602.070 1528.450 2602.370 1602.950 ;
        RECT 2602.070 1528.150 2603.290 1528.450 ;
        RECT 2602.990 1463.850 2603.290 1528.150 ;
        RECT 2602.990 1463.550 2604.210 1463.850 ;
        RECT 2603.910 1460.450 2604.210 1463.550 ;
        RECT 2602.070 1460.150 2604.210 1460.450 ;
        RECT 2602.070 1426.890 2602.370 1460.150 ;
        RECT 2597.950 1425.710 2599.130 1426.890 ;
        RECT 2601.630 1425.710 2602.810 1426.890 ;
        RECT 2598.390 1406.050 2598.690 1425.710 ;
        RECT 2598.390 1405.750 2599.610 1406.050 ;
        RECT 2599.310 1395.850 2599.610 1405.750 ;
        RECT 2597.470 1395.550 2599.610 1395.850 ;
        RECT 2597.470 1392.450 2597.770 1395.550 ;
        RECT 2597.470 1392.150 2598.690 1392.450 ;
        RECT 2598.390 1389.490 2598.690 1392.150 ;
        RECT 2597.950 1388.310 2599.130 1389.490 ;
        RECT 2604.390 1388.310 2605.570 1389.490 ;
        RECT 2604.830 1361.850 2605.130 1388.310 ;
        RECT 2604.830 1361.550 2606.050 1361.850 ;
        RECT 2605.750 1341.450 2606.050 1361.550 ;
        RECT 2606.655 1341.450 2606.985 1341.465 ;
        RECT 2605.750 1341.150 2606.985 1341.450 ;
        RECT 2606.655 1341.135 2606.985 1341.150 ;
        RECT 2606.655 1304.050 2606.985 1304.065 ;
        RECT 2604.830 1303.750 2606.985 1304.050 ;
        RECT 2604.830 1270.050 2605.130 1303.750 ;
        RECT 2606.655 1303.735 2606.985 1303.750 ;
        RECT 2602.990 1269.750 2605.130 1270.050 ;
        RECT 2602.990 1249.650 2603.290 1269.750 ;
        RECT 2606.655 1249.650 2606.985 1249.665 ;
        RECT 2602.990 1249.350 2606.985 1249.650 ;
        RECT 2606.655 1249.335 2606.985 1249.350 ;
        RECT 2606.655 1210.890 2606.985 1210.905 ;
        RECT 2605.750 1210.590 2606.985 1210.890 ;
        RECT 2605.750 1208.850 2606.050 1210.590 ;
        RECT 2606.655 1210.575 2606.985 1210.590 ;
        RECT 2603.910 1208.550 2606.050 1208.850 ;
        RECT 2603.910 1195.250 2604.210 1208.550 ;
        RECT 2603.910 1194.950 2606.050 1195.250 ;
        RECT 2605.750 1192.290 2606.050 1194.950 ;
        RECT 2605.310 1191.110 2606.490 1192.290 ;
        RECT 2601.630 1187.710 2602.810 1188.890 ;
        RECT 2602.070 1178.250 2602.370 1187.710 ;
        RECT 2599.310 1177.950 2602.370 1178.250 ;
        RECT 2599.310 1154.890 2599.610 1177.950 ;
        RECT 2598.870 1153.710 2600.050 1154.890 ;
        RECT 2605.310 1153.710 2606.490 1154.890 ;
        RECT 2605.750 1120.450 2606.050 1153.710 ;
        RECT 2606.655 1120.450 2606.985 1120.465 ;
        RECT 2605.750 1120.150 2606.985 1120.450 ;
        RECT 2606.655 1120.135 2606.985 1120.150 ;
        RECT 2612.175 1120.135 2612.505 1120.465 ;
        RECT 2612.190 1103.890 2612.490 1120.135 ;
        RECT 2597.950 1102.710 2599.130 1103.890 ;
        RECT 2611.750 1102.710 2612.930 1103.890 ;
        RECT 2598.390 1100.050 2598.690 1102.710 ;
        RECT 2598.390 1099.750 2599.610 1100.050 ;
        RECT 2599.310 1052.450 2599.610 1099.750 ;
        RECT 2598.390 1052.150 2599.610 1052.450 ;
        RECT 2598.390 981.050 2598.690 1052.150 ;
        RECT 2597.470 980.750 2598.690 981.050 ;
        RECT 2597.470 967.450 2597.770 980.750 ;
        RECT 2597.470 967.150 2599.610 967.450 ;
        RECT 2599.310 950.450 2599.610 967.150 ;
        RECT 2597.470 950.150 2599.610 950.450 ;
        RECT 2597.470 913.050 2597.770 950.150 ;
        RECT 2597.470 912.750 2599.610 913.050 ;
        RECT 2599.310 841.650 2599.610 912.750 ;
        RECT 2598.390 841.350 2599.610 841.650 ;
        RECT 2598.390 790.650 2598.690 841.350 ;
        RECT 2597.470 790.350 2598.690 790.650 ;
        RECT 2597.470 787.250 2597.770 790.350 ;
        RECT 2597.470 786.950 2599.610 787.250 ;
        RECT 2599.310 746.450 2599.610 786.950 ;
        RECT 2599.310 746.150 2600.530 746.450 ;
        RECT 2600.230 739.650 2600.530 746.150 ;
        RECT 2599.310 739.350 2600.530 739.650 ;
        RECT 2599.310 726.050 2599.610 739.350 ;
        RECT 2595.630 725.750 2599.610 726.050 ;
        RECT 2595.630 716.290 2595.930 725.750 ;
        RECT 2595.190 715.110 2596.370 716.290 ;
        RECT 2599.790 715.110 2600.970 716.290 ;
        RECT 2600.230 709.050 2600.530 715.110 ;
        RECT 2600.230 708.750 2601.450 709.050 ;
        RECT 2601.150 651.250 2601.450 708.750 ;
        RECT 2601.150 650.950 2603.290 651.250 ;
        RECT 2602.990 644.450 2603.290 650.950 ;
        RECT 2601.150 644.150 2603.290 644.450 ;
        RECT 2601.150 634.250 2601.450 644.150 ;
        RECT 2601.150 633.950 2602.370 634.250 ;
        RECT 2602.070 627.450 2602.370 633.950 ;
        RECT 2602.070 627.150 2604.210 627.450 ;
        RECT 2603.910 583.250 2604.210 627.150 ;
        RECT 2601.150 582.950 2604.210 583.250 ;
        RECT 2601.150 447.250 2601.450 582.950 ;
        RECT 2601.150 446.950 2602.370 447.250 ;
        RECT 2602.070 444.290 2602.370 446.950 ;
        RECT 2601.630 443.110 2602.810 444.290 ;
        RECT 2605.310 443.110 2606.490 444.290 ;
        RECT 2605.750 406.450 2606.050 443.110 ;
        RECT 2603.910 406.150 2606.050 406.450 ;
        RECT 2603.910 379.930 2604.210 406.150 ;
        RECT 2601.150 379.630 2604.210 379.930 ;
        RECT 2601.150 243.265 2601.450 379.630 ;
        RECT 2601.135 242.935 2601.465 243.265 ;
        RECT 2604.815 242.935 2605.145 243.265 ;
        RECT 2604.830 209.250 2605.130 242.935 ;
        RECT 2604.830 208.950 2606.050 209.250 ;
        RECT 2605.750 205.850 2606.050 208.950 ;
        RECT 2603.910 205.550 2606.050 205.850 ;
        RECT 2603.910 181.385 2604.210 205.550 ;
        RECT 2601.135 181.055 2601.465 181.385 ;
        RECT 2603.895 181.055 2604.225 181.385 ;
        RECT 2601.150 131.050 2601.450 181.055 ;
        RECT 2601.150 130.750 2603.290 131.050 ;
        RECT 2602.990 63.050 2603.290 130.750 ;
        RECT 2602.070 62.750 2603.290 63.050 ;
        RECT 2602.070 33.145 2602.370 62.750 ;
        RECT 2602.055 32.815 2602.385 33.145 ;
      LAYER met5 ;
        RECT 2600.500 2408.100 2607.620 2409.700 ;
        RECT 2601.420 1911.700 2607.620 1913.300 ;
        RECT 2600.500 1870.900 2607.620 1872.500 ;
        RECT 2597.740 1425.500 2603.020 1427.100 ;
        RECT 2597.740 1388.100 2605.780 1389.700 ;
        RECT 2605.100 1189.100 2606.700 1192.500 ;
        RECT 2601.420 1187.500 2606.700 1189.100 ;
        RECT 2598.660 1153.500 2606.700 1155.100 ;
        RECT 2597.740 1102.500 2613.140 1104.100 ;
        RECT 2594.980 714.900 2601.180 716.500 ;
        RECT 2601.420 442.900 2606.700 444.500 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.470 154.515 1358.750 154.885 ;
        RECT 1358.540 2.400 1358.680 154.515 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
      LAYER via2 ;
        RECT 1358.470 154.560 1358.750 154.840 ;
      LAYER met3 ;
        RECT 2606.000 2895.930 2610.000 2896.320 ;
        RECT 2628.710 2895.930 2629.090 2895.940 ;
        RECT 2606.000 2895.720 2629.090 2895.930 ;
        RECT 2609.580 2895.630 2629.090 2895.720 ;
        RECT 2628.710 2895.620 2629.090 2895.630 ;
        RECT 1358.445 154.850 1358.775 154.865 ;
        RECT 2628.710 154.850 2629.090 154.860 ;
        RECT 1358.445 154.550 2629.090 154.850 ;
        RECT 1358.445 154.535 1358.775 154.550 ;
        RECT 2628.710 154.540 2629.090 154.550 ;
      LAYER via3 ;
        RECT 2628.740 2895.620 2629.060 2895.940 ;
        RECT 2628.740 154.540 2629.060 154.860 ;
      LAYER met4 ;
        RECT 2628.735 2895.615 2629.065 2895.945 ;
        RECT 2628.750 154.865 2629.050 2895.615 ;
        RECT 2628.735 154.535 2629.065 154.865 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1376.390 20.640 1376.710 20.700 ;
        RECT 1379.610 20.640 1379.930 20.700 ;
        RECT 1376.390 20.500 1379.930 20.640 ;
        RECT 1376.390 20.440 1376.710 20.500 ;
        RECT 1379.610 20.440 1379.930 20.500 ;
      LAYER via ;
        RECT 1376.420 20.440 1376.680 20.700 ;
        RECT 1379.640 20.440 1379.900 20.700 ;
      LAYER met2 ;
        RECT 2249.450 3256.930 2249.730 3260.000 ;
        RECT 2250.870 3256.930 2251.150 3257.045 ;
        RECT 2249.450 3256.790 2251.150 3256.930 ;
        RECT 2249.450 3256.000 2249.730 3256.790 ;
        RECT 2250.870 3256.675 2251.150 3256.790 ;
        RECT 1379.630 245.635 1379.910 246.005 ;
        RECT 1379.700 20.730 1379.840 245.635 ;
        RECT 1376.420 20.410 1376.680 20.730 ;
        RECT 1379.640 20.410 1379.900 20.730 ;
        RECT 1376.480 2.400 1376.620 20.410 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
      LAYER via2 ;
        RECT 2250.870 3256.720 2251.150 3257.000 ;
        RECT 1379.630 245.680 1379.910 245.960 ;
      LAYER met3 ;
        RECT 2250.845 3257.010 2251.175 3257.025 ;
        RECT 2677.470 3257.010 2677.850 3257.020 ;
        RECT 2250.845 3256.710 2677.850 3257.010 ;
        RECT 2250.845 3256.695 2251.175 3256.710 ;
        RECT 2677.470 3256.700 2677.850 3256.710 ;
        RECT 1379.605 245.970 1379.935 245.985 ;
        RECT 2677.470 245.970 2677.850 245.980 ;
        RECT 1379.605 245.670 2677.850 245.970 ;
        RECT 1379.605 245.655 1379.935 245.670 ;
        RECT 2677.470 245.660 2677.850 245.670 ;
      LAYER via3 ;
        RECT 2677.500 3256.700 2677.820 3257.020 ;
        RECT 2677.500 245.660 2677.820 245.980 ;
      LAYER met4 ;
        RECT 2677.495 3256.695 2677.825 3257.025 ;
        RECT 2677.510 245.985 2677.810 3256.695 ;
        RECT 2677.495 245.655 2677.825 245.985 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2532.560 2615.490 2532.620 ;
        RECT 2628.970 2532.560 2629.290 2532.620 ;
        RECT 2615.170 2532.420 2629.290 2532.560 ;
        RECT 2615.170 2532.360 2615.490 2532.420 ;
        RECT 2628.970 2532.360 2629.290 2532.420 ;
        RECT 1400.310 162.420 1400.630 162.480 ;
        RECT 2628.970 162.420 2629.290 162.480 ;
        RECT 1400.310 162.280 2629.290 162.420 ;
        RECT 1400.310 162.220 1400.630 162.280 ;
        RECT 2628.970 162.220 2629.290 162.280 ;
        RECT 1394.330 16.560 1394.650 16.620 ;
        RECT 1400.310 16.560 1400.630 16.620 ;
        RECT 1394.330 16.420 1400.630 16.560 ;
        RECT 1394.330 16.360 1394.650 16.420 ;
        RECT 1400.310 16.360 1400.630 16.420 ;
      LAYER via ;
        RECT 2615.200 2532.360 2615.460 2532.620 ;
        RECT 2629.000 2532.360 2629.260 2532.620 ;
        RECT 1400.340 162.220 1400.600 162.480 ;
        RECT 2629.000 162.220 2629.260 162.480 ;
        RECT 1394.360 16.360 1394.620 16.620 ;
        RECT 1400.340 16.360 1400.600 16.620 ;
      LAYER met2 ;
        RECT 2615.190 2536.555 2615.470 2536.925 ;
        RECT 2615.260 2532.650 2615.400 2536.555 ;
        RECT 2615.200 2532.330 2615.460 2532.650 ;
        RECT 2629.000 2532.330 2629.260 2532.650 ;
        RECT 2629.060 162.510 2629.200 2532.330 ;
        RECT 1400.340 162.190 1400.600 162.510 ;
        RECT 2629.000 162.190 2629.260 162.510 ;
        RECT 1400.400 16.650 1400.540 162.190 ;
        RECT 1394.360 16.330 1394.620 16.650 ;
        RECT 1400.340 16.330 1400.600 16.650 ;
        RECT 1394.420 2.400 1394.560 16.330 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2536.600 2615.470 2536.880 ;
      LAYER met3 ;
        RECT 2606.000 2536.890 2610.000 2537.280 ;
        RECT 2615.165 2536.890 2615.495 2536.905 ;
        RECT 2606.000 2536.680 2615.495 2536.890 ;
        RECT 2609.580 2536.590 2615.495 2536.680 ;
        RECT 2615.165 2536.575 2615.495 2536.590 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 2836.180 282.370 2836.240 ;
        RECT 296.770 2836.180 297.090 2836.240 ;
        RECT 282.050 2836.040 297.090 2836.180 ;
        RECT 282.050 2835.980 282.370 2836.040 ;
        RECT 296.770 2835.980 297.090 2836.040 ;
        RECT 282.050 86.600 282.370 86.660 ;
        RECT 1407.670 86.600 1407.990 86.660 ;
        RECT 282.050 86.460 1407.990 86.600 ;
        RECT 282.050 86.400 282.370 86.460 ;
        RECT 1407.670 86.400 1407.990 86.460 ;
        RECT 1407.670 2.960 1407.990 3.020 ;
        RECT 1412.270 2.960 1412.590 3.020 ;
        RECT 1407.670 2.820 1412.590 2.960 ;
        RECT 1407.670 2.760 1407.990 2.820 ;
        RECT 1412.270 2.760 1412.590 2.820 ;
      LAYER via ;
        RECT 282.080 2835.980 282.340 2836.240 ;
        RECT 296.800 2835.980 297.060 2836.240 ;
        RECT 282.080 86.400 282.340 86.660 ;
        RECT 1407.700 86.400 1407.960 86.660 ;
        RECT 1407.700 2.760 1407.960 3.020 ;
        RECT 1412.300 2.760 1412.560 3.020 ;
      LAYER met2 ;
        RECT 296.790 2842.555 297.070 2842.925 ;
        RECT 296.860 2836.270 297.000 2842.555 ;
        RECT 282.080 2835.950 282.340 2836.270 ;
        RECT 296.800 2835.950 297.060 2836.270 ;
        RECT 282.140 86.690 282.280 2835.950 ;
        RECT 282.080 86.370 282.340 86.690 ;
        RECT 1407.700 86.370 1407.960 86.690 ;
        RECT 1407.760 3.050 1407.900 86.370 ;
        RECT 1407.700 2.730 1407.960 3.050 ;
        RECT 1412.300 2.730 1412.560 3.050 ;
        RECT 1412.360 2.400 1412.500 2.730 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
      LAYER via2 ;
        RECT 296.790 2842.600 297.070 2842.880 ;
      LAYER met3 ;
        RECT 296.765 2842.890 297.095 2842.905 ;
        RECT 310.000 2842.890 314.000 2843.280 ;
        RECT 296.765 2842.680 314.000 2842.890 ;
        RECT 296.765 2842.590 310.500 2842.680 ;
        RECT 296.765 2842.575 297.095 2842.590 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 779.860 2615.490 779.920 ;
        RECT 2667.150 779.860 2667.470 779.920 ;
        RECT 2615.170 779.720 2667.470 779.860 ;
        RECT 2615.170 779.660 2615.490 779.720 ;
        RECT 2667.150 779.660 2667.470 779.720 ;
        RECT 1434.810 226.680 1435.130 226.740 ;
        RECT 2667.150 226.680 2667.470 226.740 ;
        RECT 1434.810 226.540 2667.470 226.680 ;
        RECT 1434.810 226.480 1435.130 226.540 ;
        RECT 2667.150 226.480 2667.470 226.540 ;
        RECT 1429.750 20.640 1430.070 20.700 ;
        RECT 1434.810 20.640 1435.130 20.700 ;
        RECT 1429.750 20.500 1435.130 20.640 ;
        RECT 1429.750 20.440 1430.070 20.500 ;
        RECT 1434.810 20.440 1435.130 20.500 ;
      LAYER via ;
        RECT 2615.200 779.660 2615.460 779.920 ;
        RECT 2667.180 779.660 2667.440 779.920 ;
        RECT 1434.840 226.480 1435.100 226.740 ;
        RECT 2667.180 226.480 2667.440 226.740 ;
        RECT 1429.780 20.440 1430.040 20.700 ;
        RECT 1434.840 20.440 1435.100 20.700 ;
      LAYER met2 ;
        RECT 2615.190 782.155 2615.470 782.525 ;
        RECT 2615.260 779.950 2615.400 782.155 ;
        RECT 2615.200 779.630 2615.460 779.950 ;
        RECT 2667.180 779.630 2667.440 779.950 ;
        RECT 2667.240 226.770 2667.380 779.630 ;
        RECT 1434.840 226.450 1435.100 226.770 ;
        RECT 2667.180 226.450 2667.440 226.770 ;
        RECT 1434.900 20.730 1435.040 226.450 ;
        RECT 1429.780 20.410 1430.040 20.730 ;
        RECT 1434.840 20.410 1435.100 20.730 ;
        RECT 1429.840 2.400 1429.980 20.410 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
      LAYER via2 ;
        RECT 2615.190 782.200 2615.470 782.480 ;
      LAYER met3 ;
        RECT 2606.000 782.490 2610.000 782.880 ;
        RECT 2615.165 782.490 2615.495 782.505 ;
        RECT 2606.000 782.280 2615.495 782.490 ;
        RECT 2609.580 782.190 2615.495 782.280 ;
        RECT 2615.165 782.175 2615.495 782.190 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1447.690 2.960 1448.010 3.020 ;
        RECT 1448.610 2.960 1448.930 3.020 ;
        RECT 1447.690 2.820 1448.930 2.960 ;
        RECT 1447.690 2.760 1448.010 2.820 ;
        RECT 1448.610 2.760 1448.930 2.820 ;
      LAYER via ;
        RECT 1447.720 2.760 1447.980 3.020 ;
        RECT 1448.640 2.760 1448.900 3.020 ;
      LAYER met2 ;
        RECT 2177.690 3257.610 2177.970 3260.000 ;
        RECT 2178.650 3257.610 2178.930 3257.725 ;
        RECT 2177.690 3257.470 2178.930 3257.610 ;
        RECT 2177.690 3256.000 2177.970 3257.470 ;
        RECT 2178.650 3257.355 2178.930 3257.470 ;
        RECT 2677.750 3252.595 2678.030 3252.965 ;
        RECT 2677.820 246.685 2677.960 3252.595 ;
        RECT 1448.630 246.315 1448.910 246.685 ;
        RECT 2677.750 246.315 2678.030 246.685 ;
        RECT 1448.700 3.050 1448.840 246.315 ;
        RECT 1447.720 2.730 1447.980 3.050 ;
        RECT 1448.640 2.730 1448.900 3.050 ;
        RECT 1447.780 2.400 1447.920 2.730 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
      LAYER via2 ;
        RECT 2178.650 3257.400 2178.930 3257.680 ;
        RECT 2677.750 3252.640 2678.030 3252.920 ;
        RECT 1448.630 246.360 1448.910 246.640 ;
        RECT 2677.750 246.360 2678.030 246.640 ;
      LAYER met3 ;
        RECT 2178.625 3257.700 2178.955 3257.705 ;
        RECT 2178.625 3257.690 2179.210 3257.700 ;
        RECT 2178.625 3257.390 2179.410 3257.690 ;
        RECT 2178.625 3257.380 2179.210 3257.390 ;
        RECT 2178.625 3257.375 2178.955 3257.380 ;
        RECT 2178.830 3252.930 2179.210 3252.940 ;
        RECT 2677.725 3252.930 2678.055 3252.945 ;
        RECT 2178.830 3252.630 2678.055 3252.930 ;
        RECT 2178.830 3252.620 2179.210 3252.630 ;
        RECT 2677.725 3252.615 2678.055 3252.630 ;
        RECT 1448.605 246.650 1448.935 246.665 ;
        RECT 2677.725 246.650 2678.055 246.665 ;
        RECT 1448.605 246.350 2678.055 246.650 ;
        RECT 1448.605 246.335 1448.935 246.350 ;
        RECT 2677.725 246.335 2678.055 246.350 ;
      LAYER via3 ;
        RECT 2178.860 3257.380 2179.180 3257.700 ;
        RECT 2178.860 3252.620 2179.180 3252.940 ;
      LAYER met4 ;
        RECT 2178.855 3257.375 2179.185 3257.705 ;
        RECT 2178.870 3252.945 2179.170 3257.375 ;
        RECT 2178.855 3252.615 2179.185 3252.945 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 74.020 1469.630 74.080 ;
        RECT 2629.890 74.020 2630.210 74.080 ;
        RECT 1469.310 73.880 2630.210 74.020 ;
        RECT 1469.310 73.820 1469.630 73.880 ;
        RECT 2629.890 73.820 2630.210 73.880 ;
        RECT 1465.630 15.200 1465.950 15.260 ;
        RECT 1469.310 15.200 1469.630 15.260 ;
        RECT 1465.630 15.060 1469.630 15.200 ;
        RECT 1465.630 15.000 1465.950 15.060 ;
        RECT 1469.310 15.000 1469.630 15.060 ;
      LAYER via ;
        RECT 1469.340 73.820 1469.600 74.080 ;
        RECT 2629.920 73.820 2630.180 74.080 ;
        RECT 1465.660 15.000 1465.920 15.260 ;
        RECT 1469.340 15.000 1469.600 15.260 ;
      LAYER met2 ;
        RECT 2629.910 2367.915 2630.190 2368.285 ;
        RECT 2629.980 74.110 2630.120 2367.915 ;
        RECT 1469.340 73.790 1469.600 74.110 ;
        RECT 2629.920 73.790 2630.180 74.110 ;
        RECT 1469.400 15.290 1469.540 73.790 ;
        RECT 1465.660 14.970 1465.920 15.290 ;
        RECT 1469.340 14.970 1469.600 15.290 ;
        RECT 1465.720 2.400 1465.860 14.970 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
      LAYER via2 ;
        RECT 2629.910 2367.960 2630.190 2368.240 ;
      LAYER met3 ;
        RECT 2606.000 2368.250 2610.000 2368.640 ;
        RECT 2629.885 2368.250 2630.215 2368.265 ;
        RECT 2606.000 2368.040 2630.215 2368.250 ;
        RECT 2609.580 2367.950 2630.215 2368.040 ;
        RECT 2629.885 2367.935 2630.215 2367.950 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.570 20.640 1483.890 20.700 ;
        RECT 1489.550 20.640 1489.870 20.700 ;
        RECT 1483.570 20.500 1489.870 20.640 ;
        RECT 1483.570 20.440 1483.890 20.500 ;
        RECT 1489.550 20.440 1489.870 20.500 ;
      LAYER via ;
        RECT 1483.600 20.440 1483.860 20.700 ;
        RECT 1489.580 20.440 1489.840 20.700 ;
      LAYER met2 ;
        RECT 1489.570 106.235 1489.850 106.605 ;
        RECT 1489.640 20.730 1489.780 106.235 ;
        RECT 1483.600 20.410 1483.860 20.730 ;
        RECT 1489.580 20.410 1489.840 20.730 ;
        RECT 1483.660 2.400 1483.800 20.410 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
      LAYER via2 ;
        RECT 1489.570 106.280 1489.850 106.560 ;
      LAYER met3 ;
        RECT 2606.000 1458.200 2610.000 1458.800 ;
        RECT 2606.670 1457.060 2606.970 1458.200 ;
        RECT 2606.630 1456.740 2607.010 1457.060 ;
        RECT 1489.545 106.570 1489.875 106.585 ;
        RECT 2594.670 106.570 2595.050 106.580 ;
        RECT 1489.545 106.270 2595.050 106.570 ;
        RECT 1489.545 106.255 1489.875 106.270 ;
        RECT 2594.670 106.260 2595.050 106.270 ;
      LAYER via3 ;
        RECT 2606.660 1456.740 2606.980 1457.060 ;
        RECT 2594.700 106.260 2595.020 106.580 ;
      LAYER met4 ;
        RECT 2594.270 1456.310 2595.450 1457.490 ;
        RECT 2606.230 1456.310 2607.410 1457.490 ;
        RECT 2594.710 998.050 2595.010 1456.310 ;
        RECT 2593.790 997.750 2595.010 998.050 ;
        RECT 2593.790 984.450 2594.090 997.750 ;
        RECT 2593.790 984.150 2595.010 984.450 ;
        RECT 2594.710 736.250 2595.010 984.150 ;
        RECT 2591.950 735.950 2595.010 736.250 ;
        RECT 2591.950 702.250 2592.250 735.950 ;
        RECT 2591.950 701.950 2595.010 702.250 ;
        RECT 2594.710 106.585 2595.010 701.950 ;
        RECT 2594.695 106.255 2595.025 106.585 ;
      LAYER met5 ;
        RECT 2594.060 1456.100 2607.620 1457.700 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 302.750 3266.960 303.070 3267.020 ;
        RECT 1391.110 3266.960 1391.430 3267.020 ;
        RECT 302.750 3266.820 1391.430 3266.960 ;
        RECT 302.750 3266.760 303.070 3266.820 ;
        RECT 1391.110 3266.760 1391.430 3266.820 ;
        RECT 302.750 1014.120 303.070 1014.180 ;
        RECT 304.590 1014.120 304.910 1014.180 ;
        RECT 302.750 1013.980 304.910 1014.120 ;
        RECT 302.750 1013.920 303.070 1013.980 ;
        RECT 304.590 1013.920 304.910 1013.980 ;
        RECT 302.750 607.480 303.070 607.540 ;
        RECT 304.590 607.480 304.910 607.540 ;
        RECT 302.750 607.340 304.910 607.480 ;
        RECT 302.750 607.280 303.070 607.340 ;
        RECT 304.590 607.280 304.910 607.340 ;
        RECT 302.750 572.460 303.070 572.520 ;
        RECT 307.350 572.460 307.670 572.520 ;
        RECT 302.750 572.320 307.670 572.460 ;
        RECT 302.750 572.260 303.070 572.320 ;
        RECT 307.350 572.260 307.670 572.320 ;
        RECT 307.350 490.180 307.670 490.240 ;
        RECT 310.570 490.180 310.890 490.240 ;
        RECT 307.350 490.040 310.890 490.180 ;
        RECT 307.350 489.980 307.670 490.040 ;
        RECT 310.570 489.980 310.890 490.040 ;
        RECT 289.410 73.680 289.730 73.740 ;
        RECT 1497.370 73.680 1497.690 73.740 ;
        RECT 289.410 73.540 1497.690 73.680 ;
        RECT 289.410 73.480 289.730 73.540 ;
        RECT 1497.370 73.480 1497.690 73.540 ;
        RECT 1497.370 62.120 1497.690 62.180 ;
        RECT 1501.510 62.120 1501.830 62.180 ;
        RECT 1497.370 61.980 1501.830 62.120 ;
        RECT 1497.370 61.920 1497.690 61.980 ;
        RECT 1501.510 61.920 1501.830 61.980 ;
      LAYER via ;
        RECT 302.780 3266.760 303.040 3267.020 ;
        RECT 1391.140 3266.760 1391.400 3267.020 ;
        RECT 302.780 1013.920 303.040 1014.180 ;
        RECT 304.620 1013.920 304.880 1014.180 ;
        RECT 302.780 607.280 303.040 607.540 ;
        RECT 304.620 607.280 304.880 607.540 ;
        RECT 302.780 572.260 303.040 572.520 ;
        RECT 307.380 572.260 307.640 572.520 ;
        RECT 307.380 489.980 307.640 490.240 ;
        RECT 310.600 489.980 310.860 490.240 ;
        RECT 289.440 73.480 289.700 73.740 ;
        RECT 1497.400 73.480 1497.660 73.740 ;
        RECT 1497.400 61.920 1497.660 62.180 ;
        RECT 1501.540 61.920 1501.800 62.180 ;
      LAYER met2 ;
        RECT 302.780 3266.730 303.040 3267.050 ;
        RECT 1391.140 3266.730 1391.400 3267.050 ;
        RECT 302.840 1014.210 302.980 3266.730 ;
        RECT 1391.200 3260.000 1391.340 3266.730 ;
        RECT 1391.090 3256.000 1391.370 3260.000 ;
        RECT 302.780 1013.890 303.040 1014.210 ;
        RECT 304.620 1013.890 304.880 1014.210 ;
        RECT 304.680 607.570 304.820 1013.890 ;
        RECT 302.780 607.250 303.040 607.570 ;
        RECT 304.620 607.250 304.880 607.570 ;
        RECT 302.840 572.550 302.980 607.250 ;
        RECT 302.780 572.230 303.040 572.550 ;
        RECT 307.380 572.230 307.640 572.550 ;
        RECT 307.440 490.270 307.580 572.230 ;
        RECT 307.380 489.950 307.640 490.270 ;
        RECT 310.600 489.950 310.860 490.270 ;
        RECT 310.660 393.450 310.800 489.950 ;
        RECT 310.200 393.310 310.800 393.450 ;
        RECT 310.200 366.250 310.340 393.310 ;
        RECT 310.200 366.110 310.800 366.250 ;
        RECT 310.660 352.085 310.800 366.110 ;
        RECT 310.590 351.715 310.870 352.085 ;
        RECT 289.430 278.955 289.710 279.325 ;
        RECT 289.500 73.770 289.640 278.955 ;
        RECT 289.440 73.450 289.700 73.770 ;
        RECT 1497.400 73.450 1497.660 73.770 ;
        RECT 1497.460 62.210 1497.600 73.450 ;
        RECT 1497.400 61.890 1497.660 62.210 ;
        RECT 1501.540 61.890 1501.800 62.210 ;
        RECT 1501.600 2.400 1501.740 61.890 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
      LAYER via2 ;
        RECT 310.590 351.760 310.870 352.040 ;
        RECT 289.430 279.000 289.710 279.280 ;
      LAYER met3 ;
        RECT 299.270 352.050 299.650 352.060 ;
        RECT 310.565 352.050 310.895 352.065 ;
        RECT 299.270 351.750 310.895 352.050 ;
        RECT 299.270 351.740 299.650 351.750 ;
        RECT 310.565 351.735 310.895 351.750 ;
        RECT 289.405 279.290 289.735 279.305 ;
        RECT 299.270 279.290 299.650 279.300 ;
        RECT 289.405 278.990 299.650 279.290 ;
        RECT 289.405 278.975 289.735 278.990 ;
        RECT 299.270 278.980 299.650 278.990 ;
      LAYER via3 ;
        RECT 299.300 351.740 299.620 352.060 ;
        RECT 299.300 278.980 299.620 279.300 ;
      LAYER met4 ;
        RECT 299.295 351.735 299.625 352.065 ;
        RECT 299.310 279.305 299.610 351.735 ;
        RECT 299.295 278.975 299.625 279.305 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 218.860 1524.830 218.920 ;
        RECT 2611.950 218.860 2612.270 218.920 ;
        RECT 1524.510 218.720 2612.270 218.860 ;
        RECT 1524.510 218.660 1524.830 218.720 ;
        RECT 2611.950 218.660 2612.270 218.720 ;
        RECT 1518.990 20.640 1519.310 20.700 ;
        RECT 1524.510 20.640 1524.830 20.700 ;
        RECT 1518.990 20.500 1524.830 20.640 ;
        RECT 1518.990 20.440 1519.310 20.500 ;
        RECT 1524.510 20.440 1524.830 20.500 ;
      LAYER via ;
        RECT 1524.540 218.660 1524.800 218.920 ;
        RECT 2611.980 218.660 2612.240 218.920 ;
        RECT 1519.020 20.440 1519.280 20.700 ;
        RECT 1524.540 20.440 1524.800 20.700 ;
      LAYER met2 ;
        RECT 1563.170 3284.555 1563.450 3284.925 ;
        RECT 1563.240 3260.000 1563.380 3284.555 ;
        RECT 1563.130 3256.000 1563.410 3260.000 ;
        RECT 2606.910 2133.315 2607.190 2133.685 ;
        RECT 2606.980 2080.645 2607.120 2133.315 ;
        RECT 2606.910 2080.275 2607.190 2080.645 ;
        RECT 2607.830 1419.315 2608.110 1419.685 ;
        RECT 2607.900 1395.205 2608.040 1419.315 ;
        RECT 2607.830 1394.835 2608.110 1395.205 ;
        RECT 2607.830 1210.555 2608.110 1210.925 ;
        RECT 2607.900 1168.085 2608.040 1210.555 ;
        RECT 2607.830 1167.715 2608.110 1168.085 ;
        RECT 2608.290 498.595 2608.570 498.965 ;
        RECT 2608.360 379.965 2608.500 498.595 ;
        RECT 2608.290 379.595 2608.570 379.965 ;
        RECT 2611.970 278.955 2612.250 279.325 ;
        RECT 2612.040 218.950 2612.180 278.955 ;
        RECT 1524.540 218.630 1524.800 218.950 ;
        RECT 2611.980 218.630 2612.240 218.950 ;
        RECT 1524.600 20.730 1524.740 218.630 ;
        RECT 1519.020 20.410 1519.280 20.730 ;
        RECT 1524.540 20.410 1524.800 20.730 ;
        RECT 1519.080 2.400 1519.220 20.410 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
      LAYER via2 ;
        RECT 1563.170 3284.600 1563.450 3284.880 ;
        RECT 2606.910 2133.360 2607.190 2133.640 ;
        RECT 2606.910 2080.320 2607.190 2080.600 ;
        RECT 2607.830 1419.360 2608.110 1419.640 ;
        RECT 2607.830 1394.880 2608.110 1395.160 ;
        RECT 2607.830 1210.600 2608.110 1210.880 ;
        RECT 2607.830 1167.760 2608.110 1168.040 ;
        RECT 2608.290 498.640 2608.570 498.920 ;
        RECT 2608.290 379.640 2608.570 379.920 ;
        RECT 2611.970 279.000 2612.250 279.280 ;
      LAYER met3 ;
        RECT 1563.145 3284.890 1563.475 3284.905 ;
        RECT 2601.110 3284.890 2601.490 3284.900 ;
        RECT 1563.145 3284.590 2601.490 3284.890 ;
        RECT 1563.145 3284.575 1563.475 3284.590 ;
        RECT 2601.110 3284.580 2601.490 3284.590 ;
        RECT 2601.110 3263.810 2601.490 3263.820 ;
        RECT 2603.870 3263.810 2604.250 3263.820 ;
        RECT 2601.110 3263.510 2604.250 3263.810 ;
        RECT 2601.110 3263.500 2601.490 3263.510 ;
        RECT 2603.870 3263.500 2604.250 3263.510 ;
        RECT 2606.630 2329.490 2607.010 2329.500 ;
        RECT 2612.150 2329.490 2612.530 2329.500 ;
        RECT 2606.630 2329.190 2612.530 2329.490 ;
        RECT 2606.630 2329.180 2607.010 2329.190 ;
        RECT 2612.150 2329.180 2612.530 2329.190 ;
        RECT 2606.630 2283.250 2607.010 2283.260 ;
        RECT 2612.150 2283.250 2612.530 2283.260 ;
        RECT 2606.630 2282.950 2612.530 2283.250 ;
        RECT 2606.630 2282.940 2607.010 2282.950 ;
        RECT 2612.150 2282.940 2612.530 2282.950 ;
        RECT 2606.630 2175.130 2607.010 2175.140 ;
        RECT 2606.630 2174.830 2607.890 2175.130 ;
        RECT 2606.630 2174.820 2607.010 2174.830 ;
        RECT 2606.630 2173.770 2607.010 2173.780 ;
        RECT 2607.590 2173.770 2607.890 2174.830 ;
        RECT 2606.630 2173.470 2607.890 2173.770 ;
        RECT 2606.630 2173.460 2607.010 2173.470 ;
        RECT 2606.885 2133.660 2607.215 2133.665 ;
        RECT 2606.630 2133.650 2607.215 2133.660 ;
        RECT 2606.430 2133.350 2607.215 2133.650 ;
        RECT 2606.630 2133.340 2607.215 2133.350 ;
        RECT 2606.885 2133.335 2607.215 2133.340 ;
        RECT 2606.885 2080.610 2607.215 2080.625 ;
        RECT 2612.150 2080.610 2612.530 2080.620 ;
        RECT 2606.885 2080.310 2612.530 2080.610 ;
        RECT 2606.885 2080.295 2607.215 2080.310 ;
        RECT 2612.150 2080.300 2612.530 2080.310 ;
        RECT 2606.630 1419.650 2607.010 1419.660 ;
        RECT 2607.805 1419.650 2608.135 1419.665 ;
        RECT 2606.630 1419.350 2608.135 1419.650 ;
        RECT 2606.630 1419.340 2607.010 1419.350 ;
        RECT 2607.805 1419.335 2608.135 1419.350 ;
        RECT 2607.805 1395.170 2608.135 1395.185 ;
        RECT 2607.590 1394.855 2608.135 1395.170 ;
        RECT 2606.630 1393.980 2607.010 1393.990 ;
        RECT 2607.590 1393.980 2607.890 1394.855 ;
        RECT 2606.630 1393.680 2607.890 1393.980 ;
        RECT 2606.630 1393.670 2607.010 1393.680 ;
        RECT 2606.630 1342.130 2607.010 1342.140 ;
        RECT 2612.150 1342.130 2612.530 1342.140 ;
        RECT 2606.630 1341.830 2612.530 1342.130 ;
        RECT 2606.630 1341.820 2607.010 1341.830 ;
        RECT 2612.150 1341.820 2612.530 1341.830 ;
        RECT 2607.550 1307.450 2607.930 1307.460 ;
        RECT 2612.150 1307.450 2612.530 1307.460 ;
        RECT 2607.550 1307.150 2612.530 1307.450 ;
        RECT 2607.550 1307.140 2607.930 1307.150 ;
        RECT 2612.150 1307.140 2612.530 1307.150 ;
        RECT 2607.805 1210.900 2608.135 1210.905 ;
        RECT 2607.550 1210.890 2608.135 1210.900 ;
        RECT 2607.350 1210.590 2608.135 1210.890 ;
        RECT 2607.550 1210.580 2608.135 1210.590 ;
        RECT 2607.805 1210.575 2608.135 1210.580 ;
        RECT 2606.630 1168.050 2607.010 1168.060 ;
        RECT 2607.805 1168.050 2608.135 1168.065 ;
        RECT 2606.630 1167.750 2608.135 1168.050 ;
        RECT 2606.630 1167.740 2607.010 1167.750 ;
        RECT 2607.805 1167.735 2608.135 1167.750 ;
        RECT 2606.630 1103.820 2607.010 1104.140 ;
        RECT 2606.670 1102.780 2606.970 1103.820 ;
        RECT 2606.630 1102.460 2607.010 1102.780 ;
        RECT 2606.630 498.930 2607.010 498.940 ;
        RECT 2608.265 498.930 2608.595 498.945 ;
        RECT 2606.630 498.630 2608.595 498.930 ;
        RECT 2606.630 498.620 2607.010 498.630 ;
        RECT 2608.265 498.615 2608.595 498.630 ;
        RECT 2607.550 379.930 2607.930 379.940 ;
        RECT 2608.265 379.930 2608.595 379.945 ;
        RECT 2607.550 379.630 2608.595 379.930 ;
        RECT 2607.550 379.620 2607.930 379.630 ;
        RECT 2608.265 379.615 2608.595 379.630 ;
        RECT 2607.550 279.290 2607.930 279.300 ;
        RECT 2611.945 279.290 2612.275 279.305 ;
        RECT 2607.550 278.990 2612.275 279.290 ;
        RECT 2607.550 278.980 2607.930 278.990 ;
        RECT 2611.945 278.975 2612.275 278.990 ;
      LAYER via3 ;
        RECT 2601.140 3284.580 2601.460 3284.900 ;
        RECT 2601.140 3263.500 2601.460 3263.820 ;
        RECT 2603.900 3263.500 2604.220 3263.820 ;
        RECT 2606.660 2329.180 2606.980 2329.500 ;
        RECT 2612.180 2329.180 2612.500 2329.500 ;
        RECT 2606.660 2282.940 2606.980 2283.260 ;
        RECT 2612.180 2282.940 2612.500 2283.260 ;
        RECT 2606.660 2174.820 2606.980 2175.140 ;
        RECT 2606.660 2173.460 2606.980 2173.780 ;
        RECT 2606.660 2133.340 2606.980 2133.660 ;
        RECT 2612.180 2080.300 2612.500 2080.620 ;
        RECT 2606.660 1419.340 2606.980 1419.660 ;
        RECT 2606.660 1393.670 2606.980 1393.990 ;
        RECT 2606.660 1341.820 2606.980 1342.140 ;
        RECT 2612.180 1341.820 2612.500 1342.140 ;
        RECT 2607.580 1307.140 2607.900 1307.460 ;
        RECT 2612.180 1307.140 2612.500 1307.460 ;
        RECT 2607.580 1210.580 2607.900 1210.900 ;
        RECT 2606.660 1167.740 2606.980 1168.060 ;
        RECT 2606.660 1103.820 2606.980 1104.140 ;
        RECT 2606.660 1102.460 2606.980 1102.780 ;
        RECT 2606.660 498.620 2606.980 498.940 ;
        RECT 2607.580 379.620 2607.900 379.940 ;
        RECT 2607.580 278.980 2607.900 279.300 ;
      LAYER met4 ;
        RECT 2601.135 3284.575 2601.465 3284.905 ;
        RECT 2601.150 3263.825 2601.450 3284.575 ;
        RECT 2601.135 3263.495 2601.465 3263.825 ;
        RECT 2603.895 3263.495 2604.225 3263.825 ;
        RECT 2603.910 3191.050 2604.210 3263.495 ;
        RECT 2601.150 3190.750 2604.210 3191.050 ;
        RECT 2601.150 3129.850 2601.450 3190.750 ;
        RECT 2601.150 3129.550 2602.370 3129.850 ;
        RECT 2602.070 3061.850 2602.370 3129.550 ;
        RECT 2602.070 3061.550 2603.290 3061.850 ;
        RECT 2602.990 3027.850 2603.290 3061.550 ;
        RECT 2602.990 3027.550 2604.210 3027.850 ;
        RECT 2600.230 2966.350 2602.370 2966.650 ;
        RECT 2600.230 2898.650 2600.530 2966.350 ;
        RECT 2602.070 2963.250 2602.370 2966.350 ;
        RECT 2603.910 2963.250 2604.210 3027.550 ;
        RECT 2602.070 2962.950 2604.210 2963.250 ;
        RECT 2600.230 2898.350 2602.370 2898.650 ;
        RECT 2602.070 2874.850 2602.370 2898.350 ;
        RECT 2601.150 2874.550 2602.370 2874.850 ;
        RECT 2601.150 2862.610 2601.450 2874.550 ;
        RECT 2598.390 2862.310 2601.450 2862.610 ;
        RECT 2598.390 2815.690 2598.690 2862.310 ;
        RECT 2598.390 2815.390 2602.370 2815.690 ;
        RECT 2602.070 2694.650 2602.370 2815.390 ;
        RECT 2601.150 2694.350 2602.370 2694.650 ;
        RECT 2601.150 2691.250 2601.450 2694.350 ;
        RECT 2601.150 2690.950 2603.290 2691.250 ;
        RECT 2602.990 2684.450 2603.290 2690.950 ;
        RECT 2602.070 2684.150 2603.290 2684.450 ;
        RECT 2602.070 2613.490 2602.370 2684.150 ;
        RECT 2601.630 2612.310 2602.810 2613.490 ;
        RECT 2601.630 2602.110 2602.810 2603.290 ;
        RECT 2602.070 2572.250 2602.370 2602.110 ;
        RECT 2602.070 2571.950 2603.290 2572.250 ;
        RECT 2602.990 2558.650 2603.290 2571.950 ;
        RECT 2602.990 2558.350 2605.130 2558.650 ;
        RECT 2604.830 2551.850 2605.130 2558.350 ;
        RECT 2603.910 2551.550 2605.130 2551.850 ;
        RECT 2603.910 2497.450 2604.210 2551.550 ;
        RECT 2602.990 2497.150 2604.210 2497.450 ;
        RECT 2602.990 2466.850 2603.290 2497.150 ;
        RECT 2602.070 2466.550 2603.290 2466.850 ;
        RECT 2602.070 2419.690 2602.370 2466.550 ;
        RECT 2597.030 2418.510 2598.210 2419.690 ;
        RECT 2601.630 2418.510 2602.810 2419.690 ;
        RECT 2597.470 2361.890 2597.770 2418.510 ;
        RECT 2597.030 2360.710 2598.210 2361.890 ;
        RECT 2605.310 2360.710 2606.490 2361.890 ;
        RECT 2605.750 2329.490 2606.050 2360.710 ;
        RECT 2606.655 2329.490 2606.985 2329.505 ;
        RECT 2605.750 2329.190 2606.985 2329.490 ;
        RECT 2606.655 2329.175 2606.985 2329.190 ;
        RECT 2612.175 2329.175 2612.505 2329.505 ;
        RECT 2603.910 2286.350 2606.050 2286.650 ;
        RECT 2603.910 2232.250 2604.210 2286.350 ;
        RECT 2605.750 2283.250 2606.050 2286.350 ;
        RECT 2612.190 2283.265 2612.490 2329.175 ;
        RECT 2606.655 2283.250 2606.985 2283.265 ;
        RECT 2605.750 2282.950 2606.985 2283.250 ;
        RECT 2606.655 2282.935 2606.985 2282.950 ;
        RECT 2612.175 2282.935 2612.505 2283.265 ;
        RECT 2603.910 2231.950 2606.970 2232.250 ;
        RECT 2606.670 2175.145 2606.970 2231.950 ;
        RECT 2606.655 2174.815 2606.985 2175.145 ;
        RECT 2606.655 2173.455 2606.985 2173.785 ;
        RECT 2606.670 2171.050 2606.970 2173.455 ;
        RECT 2605.750 2170.750 2606.970 2171.050 ;
        RECT 2605.750 2133.650 2606.050 2170.750 ;
        RECT 2606.655 2133.650 2606.985 2133.665 ;
        RECT 2605.750 2133.350 2606.985 2133.650 ;
        RECT 2606.655 2133.335 2606.985 2133.350 ;
        RECT 2612.175 2080.295 2612.505 2080.625 ;
        RECT 2612.190 2062.690 2612.490 2080.295 ;
        RECT 2602.550 2061.510 2603.730 2062.690 ;
        RECT 2611.750 2061.510 2612.930 2062.690 ;
        RECT 2602.990 1997.650 2603.290 2061.510 ;
        RECT 2602.990 1997.350 2604.210 1997.650 ;
        RECT 2603.910 1943.250 2604.210 1997.350 ;
        RECT 2602.990 1942.950 2604.210 1943.250 ;
        RECT 2602.990 1916.050 2603.290 1942.950 ;
        RECT 2602.990 1915.750 2604.210 1916.050 ;
        RECT 2603.910 1905.850 2604.210 1915.750 ;
        RECT 2602.990 1905.550 2604.210 1905.850 ;
        RECT 2602.990 1746.050 2603.290 1905.550 ;
        RECT 2602.990 1745.750 2604.210 1746.050 ;
        RECT 2603.910 1739.250 2604.210 1745.750 ;
        RECT 2602.990 1738.950 2604.210 1739.250 ;
        RECT 2602.990 1705.250 2603.290 1738.950 ;
        RECT 2602.070 1704.950 2603.290 1705.250 ;
        RECT 2602.070 1698.450 2602.370 1704.950 ;
        RECT 2602.070 1698.150 2604.210 1698.450 ;
        RECT 2603.910 1624.090 2604.210 1698.150 ;
        RECT 2597.950 1622.910 2599.130 1624.090 ;
        RECT 2603.470 1622.910 2604.650 1624.090 ;
        RECT 2598.390 1607.090 2598.690 1622.910 ;
        RECT 2597.950 1605.910 2599.130 1607.090 ;
        RECT 2603.470 1605.910 2604.650 1607.090 ;
        RECT 2603.910 1542.050 2604.210 1605.910 ;
        RECT 2603.910 1541.750 2605.130 1542.050 ;
        RECT 2604.830 1497.850 2605.130 1541.750 ;
        RECT 2604.830 1497.550 2606.050 1497.850 ;
        RECT 2605.750 1460.450 2606.050 1497.550 ;
        RECT 2604.830 1460.150 2606.050 1460.450 ;
        RECT 2604.830 1419.650 2605.130 1460.150 ;
        RECT 2606.655 1419.650 2606.985 1419.665 ;
        RECT 2604.830 1419.350 2606.985 1419.650 ;
        RECT 2606.655 1419.335 2606.985 1419.350 ;
        RECT 2606.655 1393.665 2606.985 1393.995 ;
        RECT 2606.670 1342.145 2606.970 1393.665 ;
        RECT 2606.655 1341.815 2606.985 1342.145 ;
        RECT 2612.175 1341.815 2612.505 1342.145 ;
        RECT 2612.190 1307.465 2612.490 1341.815 ;
        RECT 2607.575 1307.135 2607.905 1307.465 ;
        RECT 2612.175 1307.135 2612.505 1307.465 ;
        RECT 2607.590 1210.905 2607.890 1307.135 ;
        RECT 2607.575 1210.575 2607.905 1210.905 ;
        RECT 2606.655 1168.050 2606.985 1168.065 ;
        RECT 2605.750 1167.750 2606.985 1168.050 ;
        RECT 2605.750 1161.250 2606.050 1167.750 ;
        RECT 2606.655 1167.735 2606.985 1167.750 ;
        RECT 2603.910 1160.950 2606.050 1161.250 ;
        RECT 2603.910 1104.130 2604.210 1160.950 ;
        RECT 2606.655 1104.130 2606.985 1104.145 ;
        RECT 2603.910 1103.830 2606.985 1104.130 ;
        RECT 2606.655 1103.815 2606.985 1103.830 ;
        RECT 2606.655 1102.455 2606.985 1102.785 ;
        RECT 2606.670 1028.650 2606.970 1102.455 ;
        RECT 2605.750 1028.350 2606.970 1028.650 ;
        RECT 2605.750 977.650 2606.050 1028.350 ;
        RECT 2603.910 977.350 2606.050 977.650 ;
        RECT 2603.910 879.050 2604.210 977.350 ;
        RECT 2603.910 878.750 2605.130 879.050 ;
        RECT 2604.830 787.250 2605.130 878.750 ;
        RECT 2604.830 786.950 2606.050 787.250 ;
        RECT 2605.750 770.250 2606.050 786.950 ;
        RECT 2604.830 769.950 2606.050 770.250 ;
        RECT 2604.830 766.850 2605.130 769.950 ;
        RECT 2603.910 766.550 2605.130 766.850 ;
        RECT 2603.910 739.650 2604.210 766.550 ;
        RECT 2603.910 739.350 2605.130 739.650 ;
        RECT 2604.830 664.850 2605.130 739.350 ;
        RECT 2604.830 664.550 2606.970 664.850 ;
        RECT 2606.670 603.650 2606.970 664.550 ;
        RECT 2605.750 603.350 2606.970 603.650 ;
        RECT 2605.750 573.050 2606.050 603.350 ;
        RECT 2602.070 572.750 2606.050 573.050 ;
        RECT 2602.070 501.650 2602.370 572.750 ;
        RECT 2602.070 501.350 2606.970 501.650 ;
        RECT 2606.670 498.945 2606.970 501.350 ;
        RECT 2606.655 498.615 2606.985 498.945 ;
        RECT 2607.575 379.615 2607.905 379.945 ;
        RECT 2607.590 279.305 2607.890 379.615 ;
        RECT 2607.575 278.975 2607.905 279.305 ;
      LAYER met5 ;
        RECT 2600.500 2612.100 2603.020 2613.700 ;
        RECT 2600.500 2603.500 2602.100 2612.100 ;
        RECT 2600.500 2601.900 2603.020 2603.500 ;
        RECT 2596.820 2418.300 2603.020 2419.900 ;
        RECT 2596.820 2360.500 2606.700 2362.100 ;
        RECT 2602.340 2061.300 2613.140 2062.900 ;
        RECT 2597.740 1622.700 2604.860 1624.300 ;
        RECT 2597.740 1605.700 2604.860 1607.300 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 289.945 3255.245 290.115 3256.095 ;
        RECT 303.285 3255.075 303.455 3255.415 ;
        RECT 303.285 3254.905 303.915 3255.075 ;
        RECT 337.785 3254.905 337.955 3256.435 ;
      LAYER mcon ;
        RECT 337.785 3256.265 337.955 3256.435 ;
        RECT 289.945 3255.925 290.115 3256.095 ;
        RECT 303.285 3255.245 303.455 3255.415 ;
        RECT 303.745 3254.905 303.915 3255.075 ;
      LAYER met1 ;
        RECT 337.725 3256.420 338.015 3256.465 ;
        RECT 989.070 3256.420 989.390 3256.480 ;
        RECT 337.725 3256.280 473.640 3256.420 ;
        RECT 337.725 3256.235 338.015 3256.280 ;
        RECT 279.290 3256.080 279.610 3256.140 ;
        RECT 289.885 3256.080 290.175 3256.125 ;
        RECT 279.290 3255.940 290.175 3256.080 ;
        RECT 279.290 3255.880 279.610 3255.940 ;
        RECT 289.885 3255.895 290.175 3255.940 ;
        RECT 473.500 3255.740 473.640 3256.280 ;
        RECT 497.420 3256.280 570.240 3256.420 ;
        RECT 497.420 3256.080 497.560 3256.280 ;
        RECT 496.960 3255.940 497.560 3256.080 ;
        RECT 496.960 3255.740 497.100 3255.940 ;
        RECT 473.500 3255.600 497.100 3255.740 ;
        RECT 570.100 3255.740 570.240 3256.280 ;
        RECT 809.760 3256.280 860.040 3256.420 ;
        RECT 592.640 3255.940 666.380 3256.080 ;
        RECT 592.640 3255.740 592.780 3255.940 ;
        RECT 570.100 3255.600 592.780 3255.740 ;
        RECT 666.240 3255.740 666.380 3255.940 ;
        RECT 713.620 3255.940 762.980 3256.080 ;
        RECT 666.240 3255.600 689.840 3255.740 ;
        RECT 289.885 3255.400 290.175 3255.445 ;
        RECT 303.225 3255.400 303.515 3255.445 ;
        RECT 289.885 3255.260 303.515 3255.400 ;
        RECT 689.700 3255.400 689.840 3255.600 ;
        RECT 713.620 3255.400 713.760 3255.940 ;
        RECT 762.840 3255.740 762.980 3255.940 ;
        RECT 762.840 3255.600 786.440 3255.740 ;
        RECT 689.700 3255.260 713.760 3255.400 ;
        RECT 786.300 3255.400 786.440 3255.600 ;
        RECT 809.760 3255.400 809.900 3256.280 ;
        RECT 859.900 3255.740 860.040 3256.280 ;
        RECT 931.660 3256.280 989.390 3256.420 ;
        RECT 931.660 3256.080 931.800 3256.280 ;
        RECT 989.070 3256.220 989.390 3256.280 ;
        RECT 883.360 3255.940 931.800 3256.080 ;
        RECT 859.900 3255.600 883.040 3255.740 ;
        RECT 786.300 3255.260 809.900 3255.400 ;
        RECT 882.900 3255.400 883.040 3255.600 ;
        RECT 883.360 3255.400 883.500 3255.940 ;
        RECT 882.900 3255.260 883.500 3255.400 ;
        RECT 289.885 3255.215 290.175 3255.260 ;
        RECT 303.225 3255.215 303.515 3255.260 ;
        RECT 303.685 3255.060 303.975 3255.105 ;
        RECT 337.725 3255.060 338.015 3255.105 ;
        RECT 303.685 3254.920 338.015 3255.060 ;
        RECT 303.685 3254.875 303.975 3254.920 ;
        RECT 337.725 3254.875 338.015 3254.920 ;
        RECT 264.570 676.500 264.890 676.560 ;
        RECT 279.290 676.500 279.610 676.560 ;
        RECT 264.570 676.360 279.610 676.500 ;
        RECT 264.570 676.300 264.890 676.360 ;
        RECT 279.290 676.300 279.610 676.360 ;
        RECT 310.570 263.060 310.890 263.120 ;
        RECT 351.510 263.060 351.830 263.120 ;
        RECT 310.570 262.920 351.830 263.060 ;
        RECT 310.570 262.860 310.890 262.920 ;
        RECT 351.510 262.860 351.830 262.920 ;
        RECT 711.230 20.640 711.550 20.700 ;
        RECT 716.290 20.640 716.610 20.700 ;
        RECT 711.230 20.500 716.610 20.640 ;
        RECT 711.230 20.440 711.550 20.500 ;
        RECT 716.290 20.440 716.610 20.500 ;
      LAYER via ;
        RECT 279.320 3255.880 279.580 3256.140 ;
        RECT 989.100 3256.220 989.360 3256.480 ;
        RECT 264.600 676.300 264.860 676.560 ;
        RECT 279.320 676.300 279.580 676.560 ;
        RECT 310.600 262.860 310.860 263.120 ;
        RECT 351.540 262.860 351.800 263.120 ;
        RECT 711.260 20.440 711.520 20.700 ;
        RECT 716.320 20.440 716.580 20.700 ;
      LAYER met2 ;
        RECT 990.890 3256.930 991.170 3260.000 ;
        RECT 989.160 3256.790 991.170 3256.930 ;
        RECT 989.160 3256.510 989.300 3256.790 ;
        RECT 989.100 3256.190 989.360 3256.510 ;
        RECT 279.320 3255.850 279.580 3256.170 ;
        RECT 990.890 3256.000 991.170 3256.790 ;
        RECT 279.380 676.590 279.520 3255.850 ;
        RECT 264.600 676.270 264.860 676.590 ;
        RECT 279.320 676.270 279.580 676.590 ;
        RECT 264.660 264.365 264.800 676.270 ;
        RECT 264.590 263.995 264.870 264.365 ;
        RECT 310.590 263.995 310.870 264.365 ;
        RECT 310.660 263.150 310.800 263.995 ;
        RECT 351.530 263.315 351.810 263.685 ;
        RECT 711.250 263.315 711.530 263.685 ;
        RECT 351.600 263.150 351.740 263.315 ;
        RECT 310.600 262.830 310.860 263.150 ;
        RECT 351.540 262.830 351.800 263.150 ;
        RECT 711.320 20.730 711.460 263.315 ;
        RECT 711.260 20.410 711.520 20.730 ;
        RECT 716.320 20.410 716.580 20.730 ;
        RECT 716.380 2.400 716.520 20.410 ;
        RECT 716.170 -4.800 716.730 2.400 ;
      LAYER via2 ;
        RECT 264.590 264.040 264.870 264.320 ;
        RECT 310.590 264.040 310.870 264.320 ;
        RECT 351.530 263.360 351.810 263.640 ;
        RECT 711.250 263.360 711.530 263.640 ;
      LAYER met3 ;
        RECT 264.565 264.330 264.895 264.345 ;
        RECT 310.565 264.330 310.895 264.345 ;
        RECT 264.565 264.030 310.895 264.330 ;
        RECT 264.565 264.015 264.895 264.030 ;
        RECT 310.565 264.015 310.895 264.030 ;
        RECT 351.505 263.650 351.835 263.665 ;
        RECT 711.225 263.650 711.555 263.665 ;
        RECT 351.505 263.350 711.555 263.650 ;
        RECT 351.505 263.335 351.835 263.350 ;
        RECT 711.225 263.335 711.555 263.350 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2122.050 3256.220 2122.370 3256.480 ;
        RECT 2122.140 3255.060 2122.280 3256.220 ;
        RECT 2637.250 3255.060 2637.570 3255.120 ;
        RECT 2122.140 3254.920 2637.570 3255.060 ;
        RECT 2637.250 3254.860 2637.570 3254.920 ;
        RECT 2637.250 345.340 2637.570 345.400 ;
        RECT 2629.520 345.200 2637.570 345.340 ;
        RECT 2629.520 345.060 2629.660 345.200 ;
        RECT 2637.250 345.140 2637.570 345.200 ;
        RECT 2629.430 344.800 2629.750 345.060 ;
        RECT 2563.190 263.060 2563.510 263.120 ;
        RECT 2629.430 263.060 2629.750 263.120 ;
        RECT 2563.190 262.920 2629.750 263.060 ;
        RECT 2563.190 262.860 2563.510 262.920 ;
        RECT 2629.430 262.860 2629.750 262.920 ;
        RECT 1536.930 19.960 1537.250 20.020 ;
        RECT 2563.190 19.960 2563.510 20.020 ;
        RECT 1536.930 19.820 2563.510 19.960 ;
        RECT 1536.930 19.760 1537.250 19.820 ;
        RECT 2563.190 19.760 2563.510 19.820 ;
      LAYER via ;
        RECT 2122.080 3256.220 2122.340 3256.480 ;
        RECT 2637.280 3254.860 2637.540 3255.120 ;
        RECT 2637.280 345.140 2637.540 345.400 ;
        RECT 2629.460 344.800 2629.720 345.060 ;
        RECT 2563.220 262.860 2563.480 263.120 ;
        RECT 2629.460 262.860 2629.720 263.120 ;
        RECT 1536.960 19.760 1537.220 20.020 ;
        RECT 2563.220 19.760 2563.480 20.020 ;
      LAYER met2 ;
        RECT 2120.650 3256.930 2120.930 3260.000 ;
        RECT 2120.650 3256.790 2122.280 3256.930 ;
        RECT 2120.650 3256.000 2120.930 3256.790 ;
        RECT 2122.140 3256.510 2122.280 3256.790 ;
        RECT 2122.080 3256.190 2122.340 3256.510 ;
        RECT 2637.280 3254.830 2637.540 3255.150 ;
        RECT 2637.340 345.430 2637.480 3254.830 ;
        RECT 2637.280 345.110 2637.540 345.430 ;
        RECT 2629.460 344.770 2629.720 345.090 ;
        RECT 2629.520 263.150 2629.660 344.770 ;
        RECT 2563.220 262.830 2563.480 263.150 ;
        RECT 2629.460 262.830 2629.720 263.150 ;
        RECT 2563.280 20.050 2563.420 262.830 ;
        RECT 1536.960 19.730 1537.220 20.050 ;
        RECT 2563.220 19.730 2563.480 20.050 ;
        RECT 1537.020 2.400 1537.160 19.730 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1499.670 244.020 1499.990 244.080 ;
        RECT 1503.810 244.020 1504.130 244.080 ;
        RECT 1499.670 243.880 1504.130 244.020 ;
        RECT 1499.670 243.820 1499.990 243.880 ;
        RECT 1503.810 243.820 1504.130 243.880 ;
        RECT 1503.810 169.220 1504.130 169.280 ;
        RECT 1552.570 169.220 1552.890 169.280 ;
        RECT 1503.810 169.080 1552.890 169.220 ;
        RECT 1503.810 169.020 1504.130 169.080 ;
        RECT 1552.570 169.020 1552.890 169.080 ;
        RECT 1552.570 14.180 1552.890 14.240 ;
        RECT 1552.570 14.040 1555.100 14.180 ;
        RECT 1552.570 13.980 1552.890 14.040 ;
        RECT 1554.960 13.900 1555.100 14.040 ;
        RECT 1554.870 13.640 1555.190 13.900 ;
      LAYER via ;
        RECT 1499.700 243.820 1499.960 244.080 ;
        RECT 1503.840 243.820 1504.100 244.080 ;
        RECT 1503.840 169.020 1504.100 169.280 ;
        RECT 1552.600 169.020 1552.860 169.280 ;
        RECT 1552.600 13.980 1552.860 14.240 ;
        RECT 1554.900 13.640 1555.160 13.900 ;
      LAYER met2 ;
        RECT 1499.650 260.000 1499.930 264.000 ;
        RECT 1499.760 244.110 1499.900 260.000 ;
        RECT 1499.700 243.790 1499.960 244.110 ;
        RECT 1503.840 243.790 1504.100 244.110 ;
        RECT 1503.900 169.310 1504.040 243.790 ;
        RECT 1503.840 168.990 1504.100 169.310 ;
        RECT 1552.600 168.990 1552.860 169.310 ;
        RECT 1552.660 14.270 1552.800 168.990 ;
        RECT 1552.600 13.950 1552.860 14.270 ;
        RECT 1554.900 13.610 1555.160 13.930 ;
        RECT 1554.960 2.400 1555.100 13.610 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2611.490 317.460 2611.810 317.520 ;
        RECT 2616.550 317.460 2616.870 317.520 ;
        RECT 2611.490 317.320 2616.870 317.460 ;
        RECT 2611.490 317.260 2611.810 317.320 ;
        RECT 2616.550 317.260 2616.870 317.320 ;
        RECT 1572.810 19.280 1573.130 19.340 ;
        RECT 2611.490 19.280 2611.810 19.340 ;
        RECT 1572.810 19.140 2611.810 19.280 ;
        RECT 1572.810 19.080 1573.130 19.140 ;
        RECT 2611.490 19.080 2611.810 19.140 ;
      LAYER via ;
        RECT 2611.520 317.260 2611.780 317.520 ;
        RECT 2616.580 317.260 2616.840 317.520 ;
        RECT 1572.840 19.080 1573.100 19.340 ;
        RECT 2611.520 19.080 2611.780 19.340 ;
      LAYER met2 ;
        RECT 2616.570 2219.675 2616.850 2220.045 ;
        RECT 2616.640 317.550 2616.780 2219.675 ;
        RECT 2611.520 317.230 2611.780 317.550 ;
        RECT 2616.580 317.230 2616.840 317.550 ;
        RECT 2611.580 19.370 2611.720 317.230 ;
        RECT 1572.840 19.050 1573.100 19.370 ;
        RECT 2611.520 19.050 2611.780 19.370 ;
        RECT 1572.900 2.400 1573.040 19.050 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 2616.570 2219.720 2616.850 2220.000 ;
      LAYER met3 ;
        RECT 2606.000 2220.010 2610.000 2220.400 ;
        RECT 2616.545 2220.010 2616.875 2220.025 ;
        RECT 2606.000 2219.800 2616.875 2220.010 ;
        RECT 2609.580 2219.710 2616.875 2219.800 ;
        RECT 2616.545 2219.695 2616.875 2219.710 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 3275.120 248.330 3275.180 ;
        RECT 547.470 3275.120 547.790 3275.180 ;
        RECT 248.010 3274.980 547.790 3275.120 ;
        RECT 248.010 3274.920 248.330 3274.980 ;
        RECT 547.470 3274.920 547.790 3274.980 ;
      LAYER via ;
        RECT 248.040 3274.920 248.300 3275.180 ;
        RECT 547.500 3274.920 547.760 3275.180 ;
      LAYER met2 ;
        RECT 248.040 3274.890 248.300 3275.210 ;
        RECT 547.500 3274.890 547.760 3275.210 ;
        RECT 248.100 18.205 248.240 3274.890 ;
        RECT 547.560 3260.000 547.700 3274.890 ;
        RECT 547.450 3256.000 547.730 3260.000 ;
        RECT 248.030 17.835 248.310 18.205 ;
        RECT 1590.310 17.835 1590.590 18.205 ;
        RECT 1590.380 2.400 1590.520 17.835 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
      LAYER via2 ;
        RECT 248.030 17.880 248.310 18.160 ;
        RECT 1590.310 17.880 1590.590 18.160 ;
      LAYER met3 ;
        RECT 248.005 18.170 248.335 18.185 ;
        RECT 1590.285 18.170 1590.615 18.185 ;
        RECT 248.005 17.870 1590.615 18.170 ;
        RECT 248.005 17.855 248.335 17.870 ;
        RECT 1590.285 17.855 1590.615 17.870 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1613.750 212.400 1614.070 212.460 ;
        RECT 2657.030 212.400 2657.350 212.460 ;
        RECT 1613.750 212.260 2657.350 212.400 ;
        RECT 1613.750 212.200 1614.070 212.260 ;
        RECT 2657.030 212.200 2657.350 212.260 ;
        RECT 1608.230 20.640 1608.550 20.700 ;
        RECT 1613.750 20.640 1614.070 20.700 ;
        RECT 1608.230 20.500 1614.070 20.640 ;
        RECT 1608.230 20.440 1608.550 20.500 ;
        RECT 1613.750 20.440 1614.070 20.500 ;
      LAYER via ;
        RECT 1613.780 212.200 1614.040 212.460 ;
        RECT 2657.060 212.200 2657.320 212.460 ;
        RECT 1608.260 20.440 1608.520 20.700 ;
        RECT 1613.780 20.440 1614.040 20.700 ;
      LAYER met2 ;
        RECT 2492.370 3272.315 2492.650 3272.685 ;
        RECT 2657.050 3272.315 2657.330 3272.685 ;
        RECT 2492.440 3260.000 2492.580 3272.315 ;
        RECT 2492.330 3256.000 2492.610 3260.000 ;
        RECT 2657.120 212.490 2657.260 3272.315 ;
        RECT 1613.780 212.170 1614.040 212.490 ;
        RECT 2657.060 212.170 2657.320 212.490 ;
        RECT 1613.840 20.730 1613.980 212.170 ;
        RECT 1608.260 20.410 1608.520 20.730 ;
        RECT 1613.780 20.410 1614.040 20.730 ;
        RECT 1608.320 2.400 1608.460 20.410 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
      LAYER via2 ;
        RECT 2492.370 3272.360 2492.650 3272.640 ;
        RECT 2657.050 3272.360 2657.330 3272.640 ;
      LAYER met3 ;
        RECT 2492.345 3272.650 2492.675 3272.665 ;
        RECT 2657.025 3272.650 2657.355 3272.665 ;
        RECT 2492.345 3272.350 2657.355 3272.650 ;
        RECT 2492.345 3272.335 2492.675 3272.350 ;
        RECT 2657.025 3272.335 2657.355 3272.350 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 505.170 3271.635 505.450 3272.005 ;
        RECT 505.240 3260.000 505.380 3271.635 ;
        RECT 505.130 3256.000 505.410 3260.000 ;
        RECT 1626.190 34.155 1626.470 34.525 ;
        RECT 1626.260 2.400 1626.400 34.155 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
      LAYER via2 ;
        RECT 505.170 3271.680 505.450 3271.960 ;
        RECT 1626.190 34.200 1626.470 34.480 ;
      LAYER met3 ;
        RECT 272.590 3271.970 272.970 3271.980 ;
        RECT 505.145 3271.970 505.475 3271.985 ;
        RECT 272.590 3271.670 505.475 3271.970 ;
        RECT 272.590 3271.660 272.970 3271.670 ;
        RECT 505.145 3271.655 505.475 3271.670 ;
        RECT 272.590 34.490 272.970 34.500 ;
        RECT 1626.165 34.490 1626.495 34.505 ;
        RECT 272.590 34.190 1626.495 34.490 ;
        RECT 272.590 34.180 272.970 34.190 ;
        RECT 1626.165 34.175 1626.495 34.190 ;
      LAYER via3 ;
        RECT 272.620 3271.660 272.940 3271.980 ;
        RECT 272.620 34.180 272.940 34.500 ;
      LAYER met4 ;
        RECT 272.615 3271.655 272.945 3271.985 ;
        RECT 272.630 34.505 272.930 3271.655 ;
        RECT 272.615 34.175 272.945 34.505 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.590 3266.280 1891.910 3266.340 ;
        RECT 2677.270 3266.280 2677.590 3266.340 ;
        RECT 1891.590 3266.140 2677.590 3266.280 ;
        RECT 1891.590 3266.080 1891.910 3266.140 ;
        RECT 2677.270 3266.080 2677.590 3266.140 ;
        RECT 1648.710 230.760 1649.030 230.820 ;
        RECT 2677.270 230.760 2677.590 230.820 ;
        RECT 1648.710 230.620 2677.590 230.760 ;
        RECT 1648.710 230.560 1649.030 230.620 ;
        RECT 2677.270 230.560 2677.590 230.620 ;
        RECT 1644.110 20.640 1644.430 20.700 ;
        RECT 1648.710 20.640 1649.030 20.700 ;
        RECT 1644.110 20.500 1649.030 20.640 ;
        RECT 1644.110 20.440 1644.430 20.500 ;
        RECT 1648.710 20.440 1649.030 20.500 ;
      LAYER via ;
        RECT 1891.620 3266.080 1891.880 3266.340 ;
        RECT 2677.300 3266.080 2677.560 3266.340 ;
        RECT 1648.740 230.560 1649.000 230.820 ;
        RECT 2677.300 230.560 2677.560 230.820 ;
        RECT 1644.140 20.440 1644.400 20.700 ;
        RECT 1648.740 20.440 1649.000 20.700 ;
      LAYER met2 ;
        RECT 1891.620 3266.050 1891.880 3266.370 ;
        RECT 2677.300 3266.050 2677.560 3266.370 ;
        RECT 1891.680 3260.000 1891.820 3266.050 ;
        RECT 1891.570 3256.000 1891.850 3260.000 ;
        RECT 2677.360 230.850 2677.500 3266.050 ;
        RECT 1648.740 230.530 1649.000 230.850 ;
        RECT 2677.300 230.530 2677.560 230.850 ;
        RECT 1648.800 20.730 1648.940 230.530 ;
        RECT 1644.140 20.410 1644.400 20.730 ;
        RECT 1648.740 20.410 1649.000 20.730 ;
        RECT 1644.200 2.400 1644.340 20.410 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 281.130 2480.200 281.450 2480.260 ;
        RECT 296.770 2480.200 297.090 2480.260 ;
        RECT 281.130 2480.060 297.090 2480.200 ;
        RECT 281.130 2480.000 281.450 2480.060 ;
        RECT 296.770 2480.000 297.090 2480.060 ;
        RECT 281.130 128.760 281.450 128.820 ;
        RECT 1656.070 128.760 1656.390 128.820 ;
        RECT 281.130 128.620 1656.390 128.760 ;
        RECT 281.130 128.560 281.450 128.620 ;
        RECT 1656.070 128.560 1656.390 128.620 ;
        RECT 1656.070 37.640 1656.390 37.700 ;
        RECT 1662.050 37.640 1662.370 37.700 ;
        RECT 1656.070 37.500 1662.370 37.640 ;
        RECT 1656.070 37.440 1656.390 37.500 ;
        RECT 1662.050 37.440 1662.370 37.500 ;
      LAYER via ;
        RECT 281.160 2480.000 281.420 2480.260 ;
        RECT 296.800 2480.000 297.060 2480.260 ;
        RECT 281.160 128.560 281.420 128.820 ;
        RECT 1656.100 128.560 1656.360 128.820 ;
        RECT 1656.100 37.440 1656.360 37.700 ;
        RECT 1662.080 37.440 1662.340 37.700 ;
      LAYER met2 ;
        RECT 296.790 2483.515 297.070 2483.885 ;
        RECT 296.860 2480.290 297.000 2483.515 ;
        RECT 281.160 2479.970 281.420 2480.290 ;
        RECT 296.800 2479.970 297.060 2480.290 ;
        RECT 281.220 128.850 281.360 2479.970 ;
        RECT 281.160 128.530 281.420 128.850 ;
        RECT 1656.100 128.530 1656.360 128.850 ;
        RECT 1656.160 37.730 1656.300 128.530 ;
        RECT 1656.100 37.410 1656.360 37.730 ;
        RECT 1662.080 37.410 1662.340 37.730 ;
        RECT 1662.140 2.400 1662.280 37.410 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
      LAYER via2 ;
        RECT 296.790 2483.560 297.070 2483.840 ;
      LAYER met3 ;
        RECT 296.765 2483.850 297.095 2483.865 ;
        RECT 310.000 2483.850 314.000 2484.240 ;
        RECT 296.765 2483.640 314.000 2483.850 ;
        RECT 296.765 2483.550 310.500 2483.640 ;
        RECT 296.765 2483.535 297.095 2483.550 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 217.500 294.330 217.560 ;
        RECT 1676.770 217.500 1677.090 217.560 ;
        RECT 294.010 217.360 1677.090 217.500 ;
        RECT 294.010 217.300 294.330 217.360 ;
        RECT 1676.770 217.300 1677.090 217.360 ;
      LAYER via ;
        RECT 294.040 217.300 294.300 217.560 ;
        RECT 1676.800 217.300 1677.060 217.560 ;
      LAYER met2 ;
        RECT 294.030 1383.275 294.310 1383.645 ;
        RECT 294.100 217.590 294.240 1383.275 ;
        RECT 294.040 217.270 294.300 217.590 ;
        RECT 1676.800 217.270 1677.060 217.590 ;
        RECT 1676.860 7.210 1677.000 217.270 ;
        RECT 1676.860 7.070 1679.760 7.210 ;
        RECT 1679.620 2.400 1679.760 7.070 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
      LAYER via2 ;
        RECT 294.030 1383.320 294.310 1383.600 ;
      LAYER met3 ;
        RECT 294.005 1383.610 294.335 1383.625 ;
        RECT 310.000 1383.610 314.000 1384.000 ;
        RECT 294.005 1383.400 314.000 1383.610 ;
        RECT 294.005 1383.310 310.500 1383.400 ;
        RECT 294.005 1383.295 294.335 1383.310 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 204.240 1704.230 204.300 ;
        RECT 2622.070 204.240 2622.390 204.300 ;
        RECT 1703.910 204.100 2622.390 204.240 ;
        RECT 1703.910 204.040 1704.230 204.100 ;
        RECT 2622.070 204.040 2622.390 204.100 ;
        RECT 1697.470 20.640 1697.790 20.700 ;
        RECT 1703.910 20.640 1704.230 20.700 ;
        RECT 1697.470 20.500 1704.230 20.640 ;
        RECT 1697.470 20.440 1697.790 20.500 ;
        RECT 1703.910 20.440 1704.230 20.500 ;
      LAYER via ;
        RECT 1703.940 204.040 1704.200 204.300 ;
        RECT 2622.100 204.040 2622.360 204.300 ;
        RECT 1697.500 20.440 1697.760 20.700 ;
        RECT 1703.940 20.440 1704.200 20.700 ;
      LAYER met2 ;
        RECT 2622.090 2790.875 2622.370 2791.245 ;
        RECT 2622.160 204.330 2622.300 2790.875 ;
        RECT 1703.940 204.010 1704.200 204.330 ;
        RECT 2622.100 204.010 2622.360 204.330 ;
        RECT 1704.000 20.730 1704.140 204.010 ;
        RECT 1697.500 20.410 1697.760 20.730 ;
        RECT 1703.940 20.410 1704.200 20.730 ;
        RECT 1697.560 2.400 1697.700 20.410 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
      LAYER via2 ;
        RECT 2622.090 2790.920 2622.370 2791.200 ;
      LAYER met3 ;
        RECT 2606.000 2791.210 2610.000 2791.600 ;
        RECT 2622.065 2791.210 2622.395 2791.225 ;
        RECT 2606.000 2791.000 2622.395 2791.210 ;
        RECT 2609.580 2790.910 2622.395 2791.000 ;
        RECT 2622.065 2790.895 2622.395 2790.910 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 372.745 263.245 372.915 264.095 ;
        RECT 394.825 263.245 394.995 264.095 ;
        RECT 448.645 263.245 448.815 264.095 ;
        RECT 593.085 263.585 593.715 263.755 ;
        RECT 628.045 262.565 628.215 263.415 ;
        RECT 675.885 262.565 676.055 263.755 ;
        RECT 689.685 263.585 690.315 263.755 ;
        RECT 731.545 48.365 731.715 96.475 ;
      LAYER mcon ;
        RECT 372.745 263.925 372.915 264.095 ;
        RECT 394.825 263.925 394.995 264.095 ;
        RECT 448.645 263.925 448.815 264.095 ;
        RECT 593.545 263.585 593.715 263.755 ;
        RECT 675.885 263.585 676.055 263.755 ;
        RECT 690.145 263.585 690.315 263.755 ;
        RECT 628.045 263.245 628.215 263.415 ;
        RECT 731.545 96.305 731.715 96.475 ;
      LAYER met1 ;
        RECT 299.990 3274.440 300.310 3274.500 ;
        RECT 590.710 3274.440 591.030 3274.500 ;
        RECT 299.990 3274.300 591.030 3274.440 ;
        RECT 299.990 3274.240 300.310 3274.300 ;
        RECT 590.710 3274.240 591.030 3274.300 ;
        RECT 279.290 628.220 279.610 628.280 ;
        RECT 299.990 628.220 300.310 628.280 ;
        RECT 279.290 628.080 300.310 628.220 ;
        RECT 279.290 628.020 279.610 628.080 ;
        RECT 299.990 628.020 300.310 628.080 ;
        RECT 279.290 264.080 279.610 264.140 ;
        RECT 372.685 264.080 372.975 264.125 ;
        RECT 279.290 263.940 372.975 264.080 ;
        RECT 279.290 263.880 279.610 263.940 ;
        RECT 372.685 263.895 372.975 263.940 ;
        RECT 394.765 264.080 395.055 264.125 ;
        RECT 448.585 264.080 448.875 264.125 ;
        RECT 394.765 263.940 448.875 264.080 ;
        RECT 394.765 263.895 395.055 263.940 ;
        RECT 448.585 263.895 448.875 263.940 ;
        RECT 696.140 263.940 731.240 264.080 ;
        RECT 593.025 263.740 593.315 263.785 ;
        RECT 545.260 263.600 593.315 263.740 ;
        RECT 372.685 263.400 372.975 263.445 ;
        RECT 394.765 263.400 395.055 263.445 ;
        RECT 372.685 263.260 395.055 263.400 ;
        RECT 372.685 263.215 372.975 263.260 ;
        RECT 394.765 263.215 395.055 263.260 ;
        RECT 448.585 263.400 448.875 263.445 ;
        RECT 545.260 263.400 545.400 263.600 ;
        RECT 593.025 263.555 593.315 263.600 ;
        RECT 593.485 263.740 593.775 263.785 ;
        RECT 675.825 263.740 676.115 263.785 ;
        RECT 689.625 263.740 689.915 263.785 ;
        RECT 593.485 263.600 594.620 263.740 ;
        RECT 593.485 263.555 593.775 263.600 ;
        RECT 448.585 263.260 545.400 263.400 ;
        RECT 594.480 263.400 594.620 263.600 ;
        RECT 675.825 263.600 689.915 263.740 ;
        RECT 675.825 263.555 676.115 263.600 ;
        RECT 689.625 263.555 689.915 263.600 ;
        RECT 690.085 263.740 690.375 263.785 ;
        RECT 696.140 263.740 696.280 263.940 ;
        RECT 731.100 263.800 731.240 263.940 ;
        RECT 690.085 263.600 696.280 263.740 ;
        RECT 690.085 263.555 690.375 263.600 ;
        RECT 731.010 263.540 731.330 263.800 ;
        RECT 627.985 263.400 628.275 263.445 ;
        RECT 594.480 263.260 628.275 263.400 ;
        RECT 448.585 263.215 448.875 263.260 ;
        RECT 627.985 263.215 628.275 263.260 ;
        RECT 627.985 262.720 628.275 262.765 ;
        RECT 675.825 262.720 676.115 262.765 ;
        RECT 627.985 262.580 676.115 262.720 ;
        RECT 627.985 262.535 628.275 262.580 ;
        RECT 675.825 262.535 676.115 262.580 ;
        RECT 731.470 96.460 731.790 96.520 ;
        RECT 731.275 96.320 731.790 96.460 ;
        RECT 731.470 96.260 731.790 96.320 ;
        RECT 731.485 48.520 731.775 48.565 ;
        RECT 734.230 48.520 734.550 48.580 ;
        RECT 731.485 48.380 734.550 48.520 ;
        RECT 731.485 48.335 731.775 48.380 ;
        RECT 734.230 48.320 734.550 48.380 ;
      LAYER via ;
        RECT 300.020 3274.240 300.280 3274.500 ;
        RECT 590.740 3274.240 591.000 3274.500 ;
        RECT 279.320 628.020 279.580 628.280 ;
        RECT 300.020 628.020 300.280 628.280 ;
        RECT 279.320 263.880 279.580 264.140 ;
        RECT 731.040 263.540 731.300 263.800 ;
        RECT 731.500 96.260 731.760 96.520 ;
        RECT 734.260 48.320 734.520 48.580 ;
      LAYER met2 ;
        RECT 300.020 3274.210 300.280 3274.530 ;
        RECT 590.740 3274.210 591.000 3274.530 ;
        RECT 300.080 628.310 300.220 3274.210 ;
        RECT 590.800 3260.000 590.940 3274.210 ;
        RECT 590.690 3256.000 590.970 3260.000 ;
        RECT 279.320 627.990 279.580 628.310 ;
        RECT 300.020 627.990 300.280 628.310 ;
        RECT 279.380 264.170 279.520 627.990 ;
        RECT 279.320 263.850 279.580 264.170 ;
        RECT 731.040 263.570 731.300 263.830 ;
        RECT 731.040 263.510 731.700 263.570 ;
        RECT 731.100 263.430 731.700 263.510 ;
        RECT 731.560 96.550 731.700 263.430 ;
        RECT 731.500 96.230 731.760 96.550 ;
        RECT 734.260 48.290 734.520 48.610 ;
        RECT 734.320 2.400 734.460 48.290 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 281.590 2497.880 281.910 2497.940 ;
        RECT 296.770 2497.880 297.090 2497.940 ;
        RECT 281.590 2497.740 297.090 2497.880 ;
        RECT 281.590 2497.680 281.910 2497.740 ;
        RECT 296.770 2497.680 297.090 2497.740 ;
        RECT 281.590 121.280 281.910 121.340 ;
        RECT 1711.270 121.280 1711.590 121.340 ;
        RECT 281.590 121.140 1711.590 121.280 ;
        RECT 281.590 121.080 281.910 121.140 ;
        RECT 1711.270 121.080 1711.590 121.140 ;
        RECT 1711.270 14.180 1711.590 14.240 ;
        RECT 1711.270 14.040 1715.640 14.180 ;
        RECT 1711.270 13.980 1711.590 14.040 ;
        RECT 1715.500 13.900 1715.640 14.040 ;
        RECT 1715.410 13.640 1715.730 13.900 ;
      LAYER via ;
        RECT 281.620 2497.680 281.880 2497.940 ;
        RECT 296.800 2497.680 297.060 2497.940 ;
        RECT 281.620 121.080 281.880 121.340 ;
        RECT 1711.300 121.080 1711.560 121.340 ;
        RECT 1711.300 13.980 1711.560 14.240 ;
        RECT 1715.440 13.640 1715.700 13.900 ;
      LAYER met2 ;
        RECT 296.790 2503.915 297.070 2504.285 ;
        RECT 296.860 2497.970 297.000 2503.915 ;
        RECT 281.620 2497.650 281.880 2497.970 ;
        RECT 296.800 2497.650 297.060 2497.970 ;
        RECT 281.680 121.370 281.820 2497.650 ;
        RECT 281.620 121.050 281.880 121.370 ;
        RECT 1711.300 121.050 1711.560 121.370 ;
        RECT 1711.360 54.810 1711.500 121.050 ;
        RECT 1711.360 54.670 1711.960 54.810 ;
        RECT 1711.820 48.690 1711.960 54.670 ;
        RECT 1711.360 48.550 1711.960 48.690 ;
        RECT 1711.360 14.270 1711.500 48.550 ;
        RECT 1711.300 13.950 1711.560 14.270 ;
        RECT 1715.440 13.610 1715.700 13.930 ;
        RECT 1715.500 2.400 1715.640 13.610 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
      LAYER via2 ;
        RECT 296.790 2503.960 297.070 2504.240 ;
      LAYER met3 ;
        RECT 296.765 2504.250 297.095 2504.265 ;
        RECT 310.000 2504.250 314.000 2504.640 ;
        RECT 296.765 2504.040 314.000 2504.250 ;
        RECT 296.765 2503.950 310.500 2504.040 ;
        RECT 296.765 2503.935 297.095 2503.950 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2657.565 447.865 2657.735 513.995 ;
        RECT 2657.565 399.925 2657.735 434.435 ;
        RECT 2658.025 144.925 2658.195 193.035 ;
        RECT 2658.485 33.745 2658.655 48.195 ;
      LAYER mcon ;
        RECT 2657.565 513.825 2657.735 513.995 ;
        RECT 2657.565 434.265 2657.735 434.435 ;
        RECT 2658.025 192.865 2658.195 193.035 ;
        RECT 2658.485 48.025 2658.655 48.195 ;
      LAYER met1 ;
        RECT 1277.030 3271.720 1277.350 3271.780 ;
        RECT 2497.870 3271.720 2498.190 3271.780 ;
        RECT 1277.030 3271.580 2498.190 3271.720 ;
        RECT 1277.030 3271.520 1277.350 3271.580 ;
        RECT 2497.870 3271.520 2498.190 3271.580 ;
        RECT 2497.870 3256.220 2498.190 3256.480 ;
        RECT 2497.960 3255.740 2498.100 3256.220 ;
        RECT 2611.490 3255.740 2611.810 3255.800 ;
        RECT 2497.960 3255.600 2611.810 3255.740 ;
        RECT 2611.490 3255.540 2611.810 3255.600 ;
        RECT 2611.490 513.980 2611.810 514.040 ;
        RECT 2657.505 513.980 2657.795 514.025 ;
        RECT 2611.490 513.840 2657.795 513.980 ;
        RECT 2611.490 513.780 2611.810 513.840 ;
        RECT 2657.505 513.795 2657.795 513.840 ;
        RECT 2657.505 448.020 2657.795 448.065 ;
        RECT 2657.950 448.020 2658.270 448.080 ;
        RECT 2657.505 447.880 2658.270 448.020 ;
        RECT 2657.505 447.835 2657.795 447.880 ;
        RECT 2657.950 447.820 2658.270 447.880 ;
        RECT 2657.505 434.420 2657.795 434.465 ;
        RECT 2657.950 434.420 2658.270 434.480 ;
        RECT 2657.505 434.280 2658.270 434.420 ;
        RECT 2657.505 434.235 2657.795 434.280 ;
        RECT 2657.950 434.220 2658.270 434.280 ;
        RECT 2657.490 400.080 2657.810 400.140 ;
        RECT 2657.295 399.940 2657.810 400.080 ;
        RECT 2657.490 399.880 2657.810 399.940 ;
        RECT 2657.490 351.800 2657.810 351.860 ;
        RECT 2659.790 351.800 2660.110 351.860 ;
        RECT 2657.490 351.660 2660.110 351.800 ;
        RECT 2657.490 351.600 2657.810 351.660 ;
        RECT 2659.790 351.600 2660.110 351.660 ;
        RECT 2657.950 303.520 2658.270 303.580 ;
        RECT 2659.790 303.520 2660.110 303.580 ;
        RECT 2657.950 303.380 2660.110 303.520 ;
        RECT 2657.950 303.320 2658.270 303.380 ;
        RECT 2659.790 303.320 2660.110 303.380 ;
        RECT 2657.950 255.580 2658.270 255.640 ;
        RECT 2659.790 255.580 2660.110 255.640 ;
        RECT 2657.950 255.440 2660.110 255.580 ;
        RECT 2657.950 255.380 2658.270 255.440 ;
        RECT 2659.790 255.380 2660.110 255.440 ;
        RECT 2657.950 207.300 2658.270 207.360 ;
        RECT 2659.790 207.300 2660.110 207.360 ;
        RECT 2657.950 207.160 2660.110 207.300 ;
        RECT 2657.950 207.100 2658.270 207.160 ;
        RECT 2659.790 207.100 2660.110 207.160 ;
        RECT 2657.950 193.020 2658.270 193.080 ;
        RECT 2657.755 192.880 2658.270 193.020 ;
        RECT 2657.950 192.820 2658.270 192.880 ;
        RECT 2657.965 145.080 2658.255 145.125 ;
        RECT 2658.410 145.080 2658.730 145.140 ;
        RECT 2657.965 144.940 2658.730 145.080 ;
        RECT 2657.965 144.895 2658.255 144.940 ;
        RECT 2658.410 144.880 2658.730 144.940 ;
        RECT 2658.410 48.180 2658.730 48.240 ;
        RECT 2658.215 48.040 2658.730 48.180 ;
        RECT 2658.410 47.980 2658.730 48.040 ;
        RECT 1733.350 33.900 1733.670 33.960 ;
        RECT 2658.425 33.900 2658.715 33.945 ;
        RECT 1733.350 33.760 2658.715 33.900 ;
        RECT 1733.350 33.700 1733.670 33.760 ;
        RECT 2658.425 33.715 2658.715 33.760 ;
      LAYER via ;
        RECT 1277.060 3271.520 1277.320 3271.780 ;
        RECT 2497.900 3271.520 2498.160 3271.780 ;
        RECT 2497.900 3256.220 2498.160 3256.480 ;
        RECT 2611.520 3255.540 2611.780 3255.800 ;
        RECT 2611.520 513.780 2611.780 514.040 ;
        RECT 2657.980 447.820 2658.240 448.080 ;
        RECT 2657.980 434.220 2658.240 434.480 ;
        RECT 2657.520 399.880 2657.780 400.140 ;
        RECT 2657.520 351.600 2657.780 351.860 ;
        RECT 2659.820 351.600 2660.080 351.860 ;
        RECT 2657.980 303.320 2658.240 303.580 ;
        RECT 2659.820 303.320 2660.080 303.580 ;
        RECT 2657.980 255.380 2658.240 255.640 ;
        RECT 2659.820 255.380 2660.080 255.640 ;
        RECT 2657.980 207.100 2658.240 207.360 ;
        RECT 2659.820 207.100 2660.080 207.360 ;
        RECT 2657.980 192.820 2658.240 193.080 ;
        RECT 2658.440 144.880 2658.700 145.140 ;
        RECT 2658.440 47.980 2658.700 48.240 ;
        RECT 1733.380 33.700 1733.640 33.960 ;
      LAYER met2 ;
        RECT 1277.060 3271.490 1277.320 3271.810 ;
        RECT 2497.900 3271.490 2498.160 3271.810 ;
        RECT 1277.120 3260.000 1277.260 3271.490 ;
        RECT 1277.010 3256.000 1277.290 3260.000 ;
        RECT 2497.960 3256.510 2498.100 3271.490 ;
        RECT 2497.900 3256.190 2498.160 3256.510 ;
        RECT 2611.520 3255.510 2611.780 3255.830 ;
        RECT 2611.580 514.070 2611.720 3255.510 ;
        RECT 2611.520 513.750 2611.780 514.070 ;
        RECT 2657.980 447.790 2658.240 448.110 ;
        RECT 2658.040 434.510 2658.180 447.790 ;
        RECT 2657.980 434.190 2658.240 434.510 ;
        RECT 2657.520 399.850 2657.780 400.170 ;
        RECT 2657.580 351.890 2657.720 399.850 ;
        RECT 2657.520 351.570 2657.780 351.890 ;
        RECT 2659.820 351.570 2660.080 351.890 ;
        RECT 2659.880 303.610 2660.020 351.570 ;
        RECT 2657.980 303.290 2658.240 303.610 ;
        RECT 2659.820 303.290 2660.080 303.610 ;
        RECT 2658.040 255.670 2658.180 303.290 ;
        RECT 2657.980 255.350 2658.240 255.670 ;
        RECT 2659.820 255.350 2660.080 255.670 ;
        RECT 2659.880 207.390 2660.020 255.350 ;
        RECT 2657.980 207.070 2658.240 207.390 ;
        RECT 2659.820 207.070 2660.080 207.390 ;
        RECT 2658.040 193.110 2658.180 207.070 ;
        RECT 2657.980 192.790 2658.240 193.110 ;
        RECT 2658.440 144.850 2658.700 145.170 ;
        RECT 2658.500 96.970 2658.640 144.850 ;
        RECT 2658.040 96.830 2658.640 96.970 ;
        RECT 2658.040 72.490 2658.180 96.830 ;
        RECT 2658.040 72.350 2658.640 72.490 ;
        RECT 2658.500 48.270 2658.640 72.350 ;
        RECT 2658.440 47.950 2658.700 48.270 ;
        RECT 1733.380 33.670 1733.640 33.990 ;
        RECT 1733.440 2.400 1733.580 33.670 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.510 241.640 1685.830 241.700 ;
        RECT 1689.650 241.640 1689.970 241.700 ;
        RECT 1685.510 241.500 1689.970 241.640 ;
        RECT 1685.510 241.440 1685.830 241.500 ;
        RECT 1689.650 241.440 1689.970 241.500 ;
        RECT 1689.650 24.380 1689.970 24.440 ;
        RECT 1751.290 24.380 1751.610 24.440 ;
        RECT 1689.650 24.240 1751.610 24.380 ;
        RECT 1689.650 24.180 1689.970 24.240 ;
        RECT 1751.290 24.180 1751.610 24.240 ;
      LAYER via ;
        RECT 1685.540 241.440 1685.800 241.700 ;
        RECT 1689.680 241.440 1689.940 241.700 ;
        RECT 1689.680 24.180 1689.940 24.440 ;
        RECT 1751.320 24.180 1751.580 24.440 ;
      LAYER met2 ;
        RECT 1685.490 260.000 1685.770 264.000 ;
        RECT 1685.600 241.730 1685.740 260.000 ;
        RECT 1685.540 241.410 1685.800 241.730 ;
        RECT 1689.680 241.410 1689.940 241.730 ;
        RECT 1689.740 24.470 1689.880 241.410 ;
        RECT 1689.680 24.150 1689.940 24.470 ;
        RECT 1751.320 24.150 1751.580 24.470 ;
        RECT 1751.380 2.400 1751.520 24.150 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1559.480 2615.490 1559.540 ;
        RECT 2638.630 1559.480 2638.950 1559.540 ;
        RECT 2615.170 1559.340 2638.950 1559.480 ;
        RECT 2615.170 1559.280 2615.490 1559.340 ;
        RECT 2638.630 1559.280 2638.950 1559.340 ;
        RECT 1768.770 51.580 1769.090 51.640 ;
        RECT 2638.630 51.580 2638.950 51.640 ;
        RECT 1768.770 51.440 2638.950 51.580 ;
        RECT 1768.770 51.380 1769.090 51.440 ;
        RECT 2638.630 51.380 2638.950 51.440 ;
      LAYER via ;
        RECT 2615.200 1559.280 2615.460 1559.540 ;
        RECT 2638.660 1559.280 2638.920 1559.540 ;
        RECT 1768.800 51.380 1769.060 51.640 ;
        RECT 2638.660 51.380 2638.920 51.640 ;
      LAYER met2 ;
        RECT 2615.190 1564.155 2615.470 1564.525 ;
        RECT 2615.260 1559.570 2615.400 1564.155 ;
        RECT 2615.200 1559.250 2615.460 1559.570 ;
        RECT 2638.660 1559.250 2638.920 1559.570 ;
        RECT 2638.720 51.670 2638.860 1559.250 ;
        RECT 1768.800 51.350 1769.060 51.670 ;
        RECT 2638.660 51.350 2638.920 51.670 ;
        RECT 1768.860 2.400 1769.000 51.350 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1564.200 2615.470 1564.480 ;
      LAYER met3 ;
        RECT 2606.000 1564.490 2610.000 1564.880 ;
        RECT 2615.165 1564.490 2615.495 1564.505 ;
        RECT 2606.000 1564.280 2615.495 1564.490 ;
        RECT 2609.580 1564.190 2615.495 1564.280 ;
        RECT 2615.165 1564.175 2615.495 1564.190 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 247.080 1787.030 247.140 ;
        RECT 2243.030 247.080 2243.350 247.140 ;
        RECT 1786.710 246.940 2243.350 247.080 ;
        RECT 1786.710 246.880 1787.030 246.940 ;
        RECT 2243.030 246.880 2243.350 246.940 ;
      LAYER via ;
        RECT 1786.740 246.880 1787.000 247.140 ;
        RECT 2243.060 246.880 2243.320 247.140 ;
      LAYER met2 ;
        RECT 2243.010 260.000 2243.290 264.000 ;
        RECT 2243.120 247.170 2243.260 260.000 ;
        RECT 1786.740 246.850 1787.000 247.170 ;
        RECT 2243.060 246.850 2243.320 247.170 ;
        RECT 1786.800 2.400 1786.940 246.850 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 898.910 244.020 899.230 244.080 ;
        RECT 903.510 244.020 903.830 244.080 ;
        RECT 898.910 243.880 903.830 244.020 ;
        RECT 898.910 243.820 899.230 243.880 ;
        RECT 903.510 243.820 903.830 243.880 ;
        RECT 903.510 135.220 903.830 135.280 ;
        RECT 1800.970 135.220 1801.290 135.280 ;
        RECT 903.510 135.080 1801.290 135.220 ;
        RECT 903.510 135.020 903.830 135.080 ;
        RECT 1800.970 135.020 1801.290 135.080 ;
        RECT 1800.970 62.120 1801.290 62.180 ;
        RECT 1804.650 62.120 1804.970 62.180 ;
        RECT 1800.970 61.980 1804.970 62.120 ;
        RECT 1800.970 61.920 1801.290 61.980 ;
        RECT 1804.650 61.920 1804.970 61.980 ;
      LAYER via ;
        RECT 898.940 243.820 899.200 244.080 ;
        RECT 903.540 243.820 903.800 244.080 ;
        RECT 903.540 135.020 903.800 135.280 ;
        RECT 1801.000 135.020 1801.260 135.280 ;
        RECT 1801.000 61.920 1801.260 62.180 ;
        RECT 1804.680 61.920 1804.940 62.180 ;
      LAYER met2 ;
        RECT 898.890 260.000 899.170 264.000 ;
        RECT 899.000 244.110 899.140 260.000 ;
        RECT 898.940 243.790 899.200 244.110 ;
        RECT 903.540 243.790 903.800 244.110 ;
        RECT 903.600 135.310 903.740 243.790 ;
        RECT 903.540 134.990 903.800 135.310 ;
        RECT 1801.000 134.990 1801.260 135.310 ;
        RECT 1801.060 62.210 1801.200 134.990 ;
        RECT 1801.000 61.890 1801.260 62.210 ;
        RECT 1804.680 61.890 1804.940 62.210 ;
        RECT 1804.740 2.400 1804.880 61.890 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2292.710 3260.840 2293.030 3260.900 ;
        RECT 2651.970 3260.840 2652.290 3260.900 ;
        RECT 2292.710 3260.700 2652.290 3260.840 ;
        RECT 2292.710 3260.640 2293.030 3260.700 ;
        RECT 2651.970 3260.640 2652.290 3260.700 ;
        RECT 1828.110 245.380 1828.430 245.440 ;
        RECT 2651.970 245.380 2652.290 245.440 ;
        RECT 1828.110 245.240 2652.290 245.380 ;
        RECT 1828.110 245.180 1828.430 245.240 ;
        RECT 2651.970 245.180 2652.290 245.240 ;
        RECT 1822.590 18.260 1822.910 18.320 ;
        RECT 1828.110 18.260 1828.430 18.320 ;
        RECT 1822.590 18.120 1828.430 18.260 ;
        RECT 1822.590 18.060 1822.910 18.120 ;
        RECT 1828.110 18.060 1828.430 18.120 ;
      LAYER via ;
        RECT 2292.740 3260.640 2293.000 3260.900 ;
        RECT 2652.000 3260.640 2652.260 3260.900 ;
        RECT 1828.140 245.180 1828.400 245.440 ;
        RECT 2652.000 245.180 2652.260 245.440 ;
        RECT 1822.620 18.060 1822.880 18.320 ;
        RECT 1828.140 18.060 1828.400 18.320 ;
      LAYER met2 ;
        RECT 2292.740 3260.610 2293.000 3260.930 ;
        RECT 2652.000 3260.610 2652.260 3260.930 ;
        RECT 2292.800 3260.000 2292.940 3260.610 ;
        RECT 2292.690 3256.000 2292.970 3260.000 ;
        RECT 2652.060 245.470 2652.200 3260.610 ;
        RECT 1828.140 245.150 1828.400 245.470 ;
        RECT 2652.000 245.150 2652.260 245.470 ;
        RECT 1828.200 18.350 1828.340 245.150 ;
        RECT 1822.620 18.030 1822.880 18.350 ;
        RECT 1828.140 18.030 1828.400 18.350 ;
        RECT 1822.680 2.400 1822.820 18.030 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 280.670 1911.380 280.990 1911.440 ;
        RECT 296.770 1911.380 297.090 1911.440 ;
        RECT 280.670 1911.240 297.090 1911.380 ;
        RECT 280.670 1911.180 280.990 1911.240 ;
        RECT 296.770 1911.180 297.090 1911.240 ;
        RECT 280.670 197.440 280.990 197.500 ;
        RECT 1835.470 197.440 1835.790 197.500 ;
        RECT 280.670 197.300 1835.790 197.440 ;
        RECT 280.670 197.240 280.990 197.300 ;
        RECT 1835.470 197.240 1835.790 197.300 ;
        RECT 1835.470 62.120 1835.790 62.180 ;
        RECT 1840.070 62.120 1840.390 62.180 ;
        RECT 1835.470 61.980 1840.390 62.120 ;
        RECT 1835.470 61.920 1835.790 61.980 ;
        RECT 1840.070 61.920 1840.390 61.980 ;
      LAYER via ;
        RECT 280.700 1911.180 280.960 1911.440 ;
        RECT 296.800 1911.180 297.060 1911.440 ;
        RECT 280.700 197.240 280.960 197.500 ;
        RECT 1835.500 197.240 1835.760 197.500 ;
        RECT 1835.500 61.920 1835.760 62.180 ;
        RECT 1840.100 61.920 1840.360 62.180 ;
      LAYER met2 ;
        RECT 296.790 1912.315 297.070 1912.685 ;
        RECT 296.860 1911.470 297.000 1912.315 ;
        RECT 280.700 1911.150 280.960 1911.470 ;
        RECT 296.800 1911.150 297.060 1911.470 ;
        RECT 280.760 197.530 280.900 1911.150 ;
        RECT 280.700 197.210 280.960 197.530 ;
        RECT 1835.500 197.210 1835.760 197.530 ;
        RECT 1835.560 62.210 1835.700 197.210 ;
        RECT 1835.500 61.890 1835.760 62.210 ;
        RECT 1840.100 61.890 1840.360 62.210 ;
        RECT 1840.160 2.400 1840.300 61.890 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
      LAYER via2 ;
        RECT 296.790 1912.360 297.070 1912.640 ;
      LAYER met3 ;
        RECT 296.765 1912.650 297.095 1912.665 ;
        RECT 310.000 1912.650 314.000 1913.040 ;
        RECT 296.765 1912.440 314.000 1912.650 ;
        RECT 296.765 1912.350 310.500 1912.440 ;
        RECT 296.765 1912.335 297.095 1912.350 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 313.405 1676.285 313.575 1690.395 ;
        RECT 312.485 1628.345 312.655 1676.115 ;
        RECT 312.945 1600.805 313.115 1628.515 ;
        RECT 312.945 1338.665 313.115 1386.775 ;
        RECT 312.945 1290.385 313.115 1304.495 ;
        RECT 312.945 1104.065 313.115 1200.455 ;
        RECT 313.405 628.065 313.575 676.175 ;
        RECT 313.405 485.265 313.575 517.395 ;
        RECT 312.945 324.445 313.115 372.555 ;
      LAYER mcon ;
        RECT 313.405 1690.225 313.575 1690.395 ;
        RECT 312.485 1675.945 312.655 1676.115 ;
        RECT 312.945 1628.345 313.115 1628.515 ;
        RECT 312.945 1386.605 313.115 1386.775 ;
        RECT 312.945 1304.325 313.115 1304.495 ;
        RECT 312.945 1200.285 313.115 1200.455 ;
        RECT 313.405 676.005 313.575 676.175 ;
        RECT 313.405 517.225 313.575 517.395 ;
        RECT 312.945 372.385 313.115 372.555 ;
      LAYER met1 ;
        RECT 313.330 1690.380 313.650 1690.440 ;
        RECT 313.135 1690.240 313.650 1690.380 ;
        RECT 313.330 1690.180 313.650 1690.240 ;
        RECT 313.345 1676.255 313.635 1676.485 ;
        RECT 312.425 1676.100 312.715 1676.145 ;
        RECT 313.420 1676.100 313.560 1676.255 ;
        RECT 312.425 1675.960 313.560 1676.100 ;
        RECT 312.425 1675.915 312.715 1675.960 ;
        RECT 312.425 1628.500 312.715 1628.545 ;
        RECT 312.885 1628.500 313.175 1628.545 ;
        RECT 312.425 1628.360 313.175 1628.500 ;
        RECT 312.425 1628.315 312.715 1628.360 ;
        RECT 312.885 1628.315 313.175 1628.360 ;
        RECT 312.870 1600.960 313.190 1601.020 ;
        RECT 312.675 1600.820 313.190 1600.960 ;
        RECT 312.870 1600.760 313.190 1600.820 ;
        RECT 311.950 1531.940 312.270 1532.000 ;
        RECT 312.870 1531.940 313.190 1532.000 ;
        RECT 311.950 1531.800 313.190 1531.940 ;
        RECT 311.950 1531.740 312.270 1531.800 ;
        RECT 312.870 1531.740 313.190 1531.800 ;
        RECT 311.490 1448.980 311.810 1449.040 ;
        RECT 312.410 1448.980 312.730 1449.040 ;
        RECT 311.490 1448.840 312.730 1448.980 ;
        RECT 311.490 1448.780 311.810 1448.840 ;
        RECT 312.410 1448.780 312.730 1448.840 ;
        RECT 312.870 1386.760 313.190 1386.820 ;
        RECT 312.675 1386.620 313.190 1386.760 ;
        RECT 312.870 1386.560 313.190 1386.620 ;
        RECT 312.885 1338.820 313.175 1338.865 ;
        RECT 313.330 1338.820 313.650 1338.880 ;
        RECT 312.885 1338.680 313.650 1338.820 ;
        RECT 312.885 1338.635 313.175 1338.680 ;
        RECT 313.330 1338.620 313.650 1338.680 ;
        RECT 312.870 1304.480 313.190 1304.540 ;
        RECT 312.675 1304.340 313.190 1304.480 ;
        RECT 312.870 1304.280 313.190 1304.340 ;
        RECT 312.870 1290.540 313.190 1290.600 ;
        RECT 312.675 1290.400 313.190 1290.540 ;
        RECT 312.870 1290.340 313.190 1290.400 ;
        RECT 312.870 1255.860 313.190 1255.920 ;
        RECT 313.330 1255.860 313.650 1255.920 ;
        RECT 312.870 1255.720 313.650 1255.860 ;
        RECT 312.870 1255.660 313.190 1255.720 ;
        RECT 313.330 1255.660 313.650 1255.720 ;
        RECT 312.885 1200.440 313.175 1200.485 ;
        RECT 313.330 1200.440 313.650 1200.500 ;
        RECT 312.885 1200.300 313.650 1200.440 ;
        RECT 312.885 1200.255 313.175 1200.300 ;
        RECT 313.330 1200.240 313.650 1200.300 ;
        RECT 312.870 1104.220 313.190 1104.280 ;
        RECT 312.675 1104.080 313.190 1104.220 ;
        RECT 312.870 1104.020 313.190 1104.080 ;
        RECT 312.870 1062.400 313.190 1062.460 ;
        RECT 313.330 1062.400 313.650 1062.460 ;
        RECT 312.870 1062.260 313.650 1062.400 ;
        RECT 312.870 1062.200 313.190 1062.260 ;
        RECT 313.330 1062.200 313.650 1062.260 ;
        RECT 312.870 724.440 313.190 724.500 ;
        RECT 313.330 724.440 313.650 724.500 ;
        RECT 312.870 724.300 313.650 724.440 ;
        RECT 312.870 724.240 313.190 724.300 ;
        RECT 313.330 724.240 313.650 724.300 ;
        RECT 313.330 676.160 313.650 676.220 ;
        RECT 313.135 676.020 313.650 676.160 ;
        RECT 313.330 675.960 313.650 676.020 ;
        RECT 313.330 628.220 313.650 628.280 ;
        RECT 313.135 628.080 313.650 628.220 ;
        RECT 313.330 628.020 313.650 628.080 ;
        RECT 313.330 593.680 313.650 593.940 ;
        RECT 313.420 593.260 313.560 593.680 ;
        RECT 313.330 593.000 313.650 593.260 ;
        RECT 313.330 517.380 313.650 517.440 ;
        RECT 313.135 517.240 313.650 517.380 ;
        RECT 313.330 517.180 313.650 517.240 ;
        RECT 313.345 485.420 313.635 485.465 ;
        RECT 313.790 485.420 314.110 485.480 ;
        RECT 313.345 485.280 314.110 485.420 ;
        RECT 313.345 485.235 313.635 485.280 ;
        RECT 313.790 485.220 314.110 485.280 ;
        RECT 312.870 386.480 313.190 386.540 ;
        RECT 314.250 386.480 314.570 386.540 ;
        RECT 312.870 386.340 314.570 386.480 ;
        RECT 312.870 386.280 313.190 386.340 ;
        RECT 314.250 386.280 314.570 386.340 ;
        RECT 312.870 372.540 313.190 372.600 ;
        RECT 312.675 372.400 313.190 372.540 ;
        RECT 312.870 372.340 313.190 372.400 ;
        RECT 312.885 324.600 313.175 324.645 ;
        RECT 313.330 324.600 313.650 324.660 ;
        RECT 312.885 324.460 313.650 324.600 ;
        RECT 312.885 324.415 313.175 324.460 ;
        RECT 313.330 324.400 313.650 324.460 ;
        RECT 311.030 300.120 311.350 300.180 ;
        RECT 313.330 300.120 313.650 300.180 ;
        RECT 311.030 299.980 313.650 300.120 ;
        RECT 311.030 299.920 311.350 299.980 ;
        RECT 313.330 299.920 313.650 299.980 ;
        RECT 311.030 211.720 311.350 211.780 ;
        RECT 1856.170 211.720 1856.490 211.780 ;
        RECT 311.030 211.580 1856.490 211.720 ;
        RECT 311.030 211.520 311.350 211.580 ;
        RECT 1856.170 211.520 1856.490 211.580 ;
        RECT 1856.170 96.460 1856.490 96.520 ;
        RECT 1857.550 96.460 1857.870 96.520 ;
        RECT 1856.170 96.320 1857.870 96.460 ;
        RECT 1856.170 96.260 1856.490 96.320 ;
        RECT 1857.550 96.260 1857.870 96.320 ;
      LAYER via ;
        RECT 313.360 1690.180 313.620 1690.440 ;
        RECT 312.900 1600.760 313.160 1601.020 ;
        RECT 311.980 1531.740 312.240 1532.000 ;
        RECT 312.900 1531.740 313.160 1532.000 ;
        RECT 311.520 1448.780 311.780 1449.040 ;
        RECT 312.440 1448.780 312.700 1449.040 ;
        RECT 312.900 1386.560 313.160 1386.820 ;
        RECT 313.360 1338.620 313.620 1338.880 ;
        RECT 312.900 1304.280 313.160 1304.540 ;
        RECT 312.900 1290.340 313.160 1290.600 ;
        RECT 312.900 1255.660 313.160 1255.920 ;
        RECT 313.360 1255.660 313.620 1255.920 ;
        RECT 313.360 1200.240 313.620 1200.500 ;
        RECT 312.900 1104.020 313.160 1104.280 ;
        RECT 312.900 1062.200 313.160 1062.460 ;
        RECT 313.360 1062.200 313.620 1062.460 ;
        RECT 312.900 724.240 313.160 724.500 ;
        RECT 313.360 724.240 313.620 724.500 ;
        RECT 313.360 675.960 313.620 676.220 ;
        RECT 313.360 628.020 313.620 628.280 ;
        RECT 313.360 593.680 313.620 593.940 ;
        RECT 313.360 593.000 313.620 593.260 ;
        RECT 313.360 517.180 313.620 517.440 ;
        RECT 313.820 485.220 314.080 485.480 ;
        RECT 312.900 386.280 313.160 386.540 ;
        RECT 314.280 386.280 314.540 386.540 ;
        RECT 312.900 372.340 313.160 372.600 ;
        RECT 313.360 324.400 313.620 324.660 ;
        RECT 311.060 299.920 311.320 300.180 ;
        RECT 313.360 299.920 313.620 300.180 ;
        RECT 311.060 211.520 311.320 211.780 ;
        RECT 1856.200 211.520 1856.460 211.780 ;
        RECT 1856.200 96.260 1856.460 96.520 ;
        RECT 1857.580 96.260 1857.840 96.520 ;
      LAYER met2 ;
        RECT 312.890 1740.955 313.170 1741.325 ;
        RECT 312.960 1704.490 313.100 1740.955 ;
        RECT 312.960 1704.350 313.560 1704.490 ;
        RECT 313.420 1690.470 313.560 1704.350 ;
        RECT 313.360 1690.150 313.620 1690.470 ;
        RECT 312.900 1600.730 313.160 1601.050 ;
        RECT 312.960 1580.165 313.100 1600.730 ;
        RECT 311.970 1579.795 312.250 1580.165 ;
        RECT 312.890 1579.795 313.170 1580.165 ;
        RECT 312.040 1532.030 312.180 1579.795 ;
        RECT 311.980 1531.710 312.240 1532.030 ;
        RECT 312.900 1531.710 313.160 1532.030 ;
        RECT 312.960 1514.770 313.100 1531.710 ;
        RECT 312.500 1514.630 313.100 1514.770 ;
        RECT 312.500 1449.070 312.640 1514.630 ;
        RECT 311.520 1448.750 311.780 1449.070 ;
        RECT 312.440 1448.750 312.700 1449.070 ;
        RECT 311.580 1435.210 311.720 1448.750 ;
        RECT 311.580 1435.070 313.100 1435.210 ;
        RECT 312.960 1386.850 313.100 1435.070 ;
        RECT 312.900 1386.530 313.160 1386.850 ;
        RECT 313.360 1338.650 313.620 1338.910 ;
        RECT 312.960 1338.590 313.620 1338.650 ;
        RECT 312.960 1338.510 313.560 1338.590 ;
        RECT 312.960 1304.570 313.100 1338.510 ;
        RECT 312.900 1304.250 313.160 1304.570 ;
        RECT 312.900 1290.310 313.160 1290.630 ;
        RECT 312.960 1255.950 313.100 1290.310 ;
        RECT 312.900 1255.630 313.160 1255.950 ;
        RECT 313.360 1255.630 313.620 1255.950 ;
        RECT 313.420 1200.530 313.560 1255.630 ;
        RECT 313.360 1200.210 313.620 1200.530 ;
        RECT 312.900 1103.990 313.160 1104.310 ;
        RECT 312.960 1062.490 313.100 1103.990 ;
        RECT 312.900 1062.170 313.160 1062.490 ;
        RECT 313.360 1062.170 313.620 1062.490 ;
        RECT 313.420 870.130 313.560 1062.170 ;
        RECT 312.960 869.990 313.560 870.130 ;
        RECT 312.960 869.620 313.100 869.990 ;
        RECT 312.960 869.480 313.560 869.620 ;
        RECT 313.420 724.530 313.560 869.480 ;
        RECT 312.900 724.210 313.160 724.530 ;
        RECT 313.360 724.210 313.620 724.530 ;
        RECT 312.960 677.125 313.100 724.210 ;
        RECT 312.890 676.755 313.170 677.125 ;
        RECT 313.350 676.075 313.630 676.445 ;
        RECT 313.360 675.930 313.620 676.075 ;
        RECT 313.360 627.990 313.620 628.310 ;
        RECT 313.420 593.970 313.560 627.990 ;
        RECT 313.360 593.650 313.620 593.970 ;
        RECT 313.360 592.970 313.620 593.290 ;
        RECT 313.420 517.470 313.560 592.970 ;
        RECT 313.360 517.150 313.620 517.470 ;
        RECT 313.820 485.190 314.080 485.510 ;
        RECT 313.880 483.210 314.020 485.190 ;
        RECT 313.880 483.070 314.480 483.210 ;
        RECT 314.340 386.570 314.480 483.070 ;
        RECT 312.900 386.250 313.160 386.570 ;
        RECT 314.280 386.250 314.540 386.570 ;
        RECT 312.960 372.630 313.100 386.250 ;
        RECT 312.900 372.310 313.160 372.630 ;
        RECT 313.360 324.370 313.620 324.690 ;
        RECT 313.420 300.210 313.560 324.370 ;
        RECT 311.060 299.890 311.320 300.210 ;
        RECT 313.360 299.890 313.620 300.210 ;
        RECT 311.120 211.810 311.260 299.890 ;
        RECT 311.060 211.490 311.320 211.810 ;
        RECT 1856.200 211.490 1856.460 211.810 ;
        RECT 1856.260 96.550 1856.400 211.490 ;
        RECT 1856.200 96.230 1856.460 96.550 ;
        RECT 1857.580 96.230 1857.840 96.550 ;
        RECT 1857.640 61.610 1857.780 96.230 ;
        RECT 1857.640 61.470 1858.240 61.610 ;
        RECT 1858.100 2.400 1858.240 61.470 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
      LAYER via2 ;
        RECT 312.890 1741.000 313.170 1741.280 ;
        RECT 311.970 1579.840 312.250 1580.120 ;
        RECT 312.890 1579.840 313.170 1580.120 ;
        RECT 312.890 676.800 313.170 677.080 ;
        RECT 313.350 676.120 313.630 676.400 ;
      LAYER met3 ;
        RECT 310.000 1743.800 314.000 1744.400 ;
        RECT 313.110 1741.305 313.410 1743.800 ;
        RECT 312.865 1740.990 313.410 1741.305 ;
        RECT 312.865 1740.975 313.195 1740.990 ;
        RECT 311.945 1580.130 312.275 1580.145 ;
        RECT 312.865 1580.130 313.195 1580.145 ;
        RECT 311.945 1579.830 313.195 1580.130 ;
        RECT 311.945 1579.815 312.275 1579.830 ;
        RECT 312.865 1579.815 313.195 1579.830 ;
        RECT 312.865 677.090 313.195 677.105 ;
        RECT 312.865 676.775 313.410 677.090 ;
        RECT 313.110 676.425 313.410 676.775 ;
        RECT 313.110 676.110 313.655 676.425 ;
        RECT 313.325 676.095 313.655 676.110 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2935.120 2615.490 2935.180 ;
        RECT 2637.710 2935.120 2638.030 2935.180 ;
        RECT 2615.170 2934.980 2638.030 2935.120 ;
        RECT 2615.170 2934.920 2615.490 2934.980 ;
        RECT 2637.710 2934.920 2638.030 2934.980 ;
        RECT 1876.410 246.400 1876.730 246.460 ;
        RECT 2637.710 246.400 2638.030 246.460 ;
        RECT 1876.410 246.260 2638.030 246.400 ;
        RECT 1876.410 246.200 1876.730 246.260 ;
        RECT 2637.710 246.200 2638.030 246.260 ;
      LAYER via ;
        RECT 2615.200 2934.920 2615.460 2935.180 ;
        RECT 2637.740 2934.920 2638.000 2935.180 ;
        RECT 1876.440 246.200 1876.700 246.460 ;
        RECT 2637.740 246.200 2638.000 246.460 ;
      LAYER met2 ;
        RECT 2615.190 2937.755 2615.470 2938.125 ;
        RECT 2615.260 2935.210 2615.400 2937.755 ;
        RECT 2615.200 2934.890 2615.460 2935.210 ;
        RECT 2637.740 2934.890 2638.000 2935.210 ;
        RECT 2637.800 246.490 2637.940 2934.890 ;
        RECT 1876.440 246.170 1876.700 246.490 ;
        RECT 2637.740 246.170 2638.000 246.490 ;
        RECT 1876.500 17.410 1876.640 246.170 ;
        RECT 1876.040 17.270 1876.640 17.410 ;
        RECT 1876.040 2.400 1876.180 17.270 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2937.800 2615.470 2938.080 ;
      LAYER met3 ;
        RECT 2606.000 2938.090 2610.000 2938.480 ;
        RECT 2615.165 2938.090 2615.495 2938.105 ;
        RECT 2606.000 2937.880 2615.495 2938.090 ;
        RECT 2609.580 2937.790 2615.495 2937.880 ;
        RECT 2615.165 2937.775 2615.495 2937.790 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 244.330 869.620 244.650 869.680 ;
        RECT 296.770 869.620 297.090 869.680 ;
        RECT 244.330 869.480 297.090 869.620 ;
        RECT 244.330 869.420 244.650 869.480 ;
        RECT 296.770 869.420 297.090 869.480 ;
        RECT 244.330 30.500 244.650 30.560 ;
        RECT 752.170 30.500 752.490 30.560 ;
        RECT 244.330 30.360 752.490 30.500 ;
        RECT 244.330 30.300 244.650 30.360 ;
        RECT 752.170 30.300 752.490 30.360 ;
      LAYER via ;
        RECT 244.360 869.420 244.620 869.680 ;
        RECT 296.800 869.420 297.060 869.680 ;
        RECT 244.360 30.300 244.620 30.560 ;
        RECT 752.200 30.300 752.460 30.560 ;
      LAYER met2 ;
        RECT 296.790 875.995 297.070 876.365 ;
        RECT 296.860 869.710 297.000 875.995 ;
        RECT 244.360 869.390 244.620 869.710 ;
        RECT 296.800 869.390 297.060 869.710 ;
        RECT 244.420 30.590 244.560 869.390 ;
        RECT 244.360 30.270 244.620 30.590 ;
        RECT 752.200 30.270 752.460 30.590 ;
        RECT 752.260 2.400 752.400 30.270 ;
        RECT 752.050 -4.800 752.610 2.400 ;
      LAYER via2 ;
        RECT 296.790 876.040 297.070 876.320 ;
      LAYER met3 ;
        RECT 296.765 876.330 297.095 876.345 ;
        RECT 310.000 876.330 314.000 876.720 ;
        RECT 296.765 876.120 314.000 876.330 ;
        RECT 296.765 876.030 310.500 876.120 ;
        RECT 296.765 876.015 297.095 876.030 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1890.745 48.365 1890.915 96.475 ;
      LAYER mcon ;
        RECT 1890.745 96.305 1890.915 96.475 ;
      LAYER met1 ;
        RECT 1890.670 96.460 1890.990 96.520 ;
        RECT 1890.475 96.320 1890.990 96.460 ;
        RECT 1890.670 96.260 1890.990 96.320 ;
        RECT 1890.685 48.520 1890.975 48.565 ;
        RECT 1893.890 48.520 1894.210 48.580 ;
        RECT 1890.685 48.380 1894.210 48.520 ;
        RECT 1890.685 48.335 1890.975 48.380 ;
        RECT 1893.890 48.320 1894.210 48.380 ;
      LAYER via ;
        RECT 1890.700 96.260 1890.960 96.520 ;
        RECT 1893.920 48.320 1894.180 48.580 ;
      LAYER met2 ;
        RECT 1891.150 113.715 1891.430 114.085 ;
        RECT 1891.220 96.970 1891.360 113.715 ;
        RECT 1890.760 96.830 1891.360 96.970 ;
        RECT 1890.760 96.550 1890.900 96.830 ;
        RECT 1890.700 96.230 1890.960 96.550 ;
        RECT 1893.920 48.290 1894.180 48.610 ;
        RECT 1893.980 2.400 1894.120 48.290 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
      LAYER via2 ;
        RECT 1891.150 113.760 1891.430 114.040 ;
      LAYER met3 ;
        RECT 279.950 2546.410 280.330 2546.420 ;
        RECT 310.000 2546.410 314.000 2546.800 ;
        RECT 279.950 2546.200 314.000 2546.410 ;
        RECT 279.950 2546.110 310.500 2546.200 ;
        RECT 279.950 2546.100 280.330 2546.110 ;
        RECT 279.950 114.050 280.330 114.060 ;
        RECT 1891.125 114.050 1891.455 114.065 ;
        RECT 279.950 113.750 1891.455 114.050 ;
        RECT 279.950 113.740 280.330 113.750 ;
        RECT 1891.125 113.735 1891.455 113.750 ;
      LAYER via3 ;
        RECT 279.980 2546.100 280.300 2546.420 ;
        RECT 279.980 113.740 280.300 114.060 ;
      LAYER met4 ;
        RECT 279.975 2546.095 280.305 2546.425 ;
        RECT 279.990 114.065 280.290 2546.095 ;
        RECT 279.975 113.735 280.305 114.065 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1806.030 3279.200 1806.350 3279.260 ;
        RECT 2697.970 3279.200 2698.290 3279.260 ;
        RECT 1806.030 3279.060 2698.290 3279.200 ;
        RECT 1806.030 3279.000 1806.350 3279.060 ;
        RECT 2697.970 3279.000 2698.290 3279.060 ;
        RECT 1911.830 30.500 1912.150 30.560 ;
        RECT 2697.970 30.500 2698.290 30.560 ;
        RECT 1911.830 30.360 2698.290 30.500 ;
        RECT 1911.830 30.300 1912.150 30.360 ;
        RECT 2697.970 30.300 2698.290 30.360 ;
      LAYER via ;
        RECT 1806.060 3279.000 1806.320 3279.260 ;
        RECT 2698.000 3279.000 2698.260 3279.260 ;
        RECT 1911.860 30.300 1912.120 30.560 ;
        RECT 2698.000 30.300 2698.260 30.560 ;
      LAYER met2 ;
        RECT 1806.060 3278.970 1806.320 3279.290 ;
        RECT 2698.000 3278.970 2698.260 3279.290 ;
        RECT 1806.120 3260.000 1806.260 3278.970 ;
        RECT 1806.010 3256.000 1806.290 3260.000 ;
        RECT 2698.060 30.590 2698.200 3278.970 ;
        RECT 1911.860 30.270 1912.120 30.590 ;
        RECT 2698.000 30.270 2698.260 30.590 ;
        RECT 1911.920 2.400 1912.060 30.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2221.410 3256.220 2221.730 3256.480 ;
        RECT 2221.500 3255.400 2221.640 3256.220 ;
        RECT 2656.570 3255.400 2656.890 3255.460 ;
        RECT 2221.500 3255.260 2656.890 3255.400 ;
        RECT 2656.570 3255.200 2656.890 3255.260 ;
        RECT 1929.310 18.260 1929.630 18.320 ;
        RECT 2656.570 18.260 2656.890 18.320 ;
        RECT 1929.310 18.120 2656.890 18.260 ;
        RECT 1929.310 18.060 1929.630 18.120 ;
        RECT 2656.570 18.060 2656.890 18.120 ;
      LAYER via ;
        RECT 2221.440 3256.220 2221.700 3256.480 ;
        RECT 2656.600 3255.200 2656.860 3255.460 ;
        RECT 1929.340 18.060 1929.600 18.320 ;
        RECT 2656.600 18.060 2656.860 18.320 ;
      LAYER met2 ;
        RECT 2220.930 3256.930 2221.210 3260.000 ;
        RECT 2220.930 3256.790 2221.640 3256.930 ;
        RECT 2220.930 3256.000 2221.210 3256.790 ;
        RECT 2221.500 3256.510 2221.640 3256.790 ;
        RECT 2221.440 3256.190 2221.700 3256.510 ;
        RECT 2656.600 3255.170 2656.860 3255.490 ;
        RECT 2656.660 18.350 2656.800 3255.170 ;
        RECT 1929.340 18.030 1929.600 18.350 ;
        RECT 2656.600 18.030 2656.860 18.350 ;
        RECT 1929.400 2.400 1929.540 18.030 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1945.870 71.980 1946.190 72.040 ;
        RECT 1946.790 71.980 1947.110 72.040 ;
        RECT 1945.870 71.840 1947.110 71.980 ;
        RECT 1945.870 71.780 1946.190 71.840 ;
        RECT 1946.790 71.780 1947.110 71.840 ;
      LAYER via ;
        RECT 1945.900 71.780 1946.160 72.040 ;
        RECT 1946.820 71.780 1947.080 72.040 ;
      LAYER met2 ;
        RECT 1945.890 203.475 1946.170 203.845 ;
        RECT 1945.960 72.070 1946.100 203.475 ;
        RECT 1945.900 71.750 1946.160 72.070 ;
        RECT 1946.820 71.750 1947.080 72.070 ;
        RECT 1946.880 61.610 1947.020 71.750 ;
        RECT 1946.880 61.470 1947.480 61.610 ;
        RECT 1947.340 2.400 1947.480 61.470 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1945.890 203.520 1946.170 203.800 ;
      LAYER met3 ;
        RECT 280.870 2652.490 281.250 2652.500 ;
        RECT 310.000 2652.490 314.000 2652.880 ;
        RECT 280.870 2652.280 314.000 2652.490 ;
        RECT 280.870 2652.190 310.500 2652.280 ;
        RECT 280.870 2652.180 281.250 2652.190 ;
        RECT 280.870 203.810 281.250 203.820 ;
        RECT 1945.865 203.810 1946.195 203.825 ;
        RECT 280.870 203.510 1946.195 203.810 ;
        RECT 280.870 203.500 281.250 203.510 ;
        RECT 1945.865 203.495 1946.195 203.510 ;
      LAYER via3 ;
        RECT 280.900 2652.180 281.220 2652.500 ;
        RECT 280.900 203.500 281.220 203.820 ;
      LAYER met4 ;
        RECT 280.895 2652.175 281.225 2652.505 ;
        RECT 280.910 203.825 281.210 2652.175 ;
        RECT 280.895 203.495 281.225 203.825 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1332.020 2615.490 1332.080 ;
        RECT 2680.490 1332.020 2680.810 1332.080 ;
        RECT 2615.170 1331.880 2680.810 1332.020 ;
        RECT 2615.170 1331.820 2615.490 1331.880 ;
        RECT 2680.490 1331.820 2680.810 1331.880 ;
        RECT 1966.110 227.700 1966.430 227.760 ;
        RECT 2680.490 227.700 2680.810 227.760 ;
        RECT 1966.110 227.560 2680.810 227.700 ;
        RECT 1966.110 227.500 1966.430 227.560 ;
        RECT 2680.490 227.500 2680.810 227.560 ;
        RECT 1966.110 14.180 1966.430 14.240 ;
        RECT 1965.280 14.040 1966.430 14.180 ;
        RECT 1965.280 13.900 1965.420 14.040 ;
        RECT 1966.110 13.980 1966.430 14.040 ;
        RECT 1965.190 13.640 1965.510 13.900 ;
      LAYER via ;
        RECT 2615.200 1331.820 2615.460 1332.080 ;
        RECT 2680.520 1331.820 2680.780 1332.080 ;
        RECT 1966.140 227.500 1966.400 227.760 ;
        RECT 2680.520 227.500 2680.780 227.760 ;
        RECT 1966.140 13.980 1966.400 14.240 ;
        RECT 1965.220 13.640 1965.480 13.900 ;
      LAYER met2 ;
        RECT 2615.200 1331.965 2615.460 1332.110 ;
        RECT 2615.190 1331.595 2615.470 1331.965 ;
        RECT 2680.520 1331.790 2680.780 1332.110 ;
        RECT 2680.580 227.790 2680.720 1331.790 ;
        RECT 1966.140 227.470 1966.400 227.790 ;
        RECT 2680.520 227.470 2680.780 227.790 ;
        RECT 1966.200 14.270 1966.340 227.470 ;
        RECT 1966.140 13.950 1966.400 14.270 ;
        RECT 1965.220 13.610 1965.480 13.930 ;
        RECT 1965.280 2.400 1965.420 13.610 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1331.640 2615.470 1331.920 ;
      LAYER met3 ;
        RECT 2606.000 1331.930 2610.000 1332.320 ;
        RECT 2615.165 1331.930 2615.495 1331.945 ;
        RECT 2606.000 1331.720 2615.495 1331.930 ;
        RECT 2609.580 1331.630 2615.495 1331.720 ;
        RECT 2615.165 1331.615 2615.495 1331.630 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1056.230 244.020 1056.550 244.080 ;
        RECT 1061.750 244.020 1062.070 244.080 ;
        RECT 1056.230 243.880 1062.070 244.020 ;
        RECT 1056.230 243.820 1056.550 243.880 ;
        RECT 1061.750 243.820 1062.070 243.880 ;
        RECT 1061.750 79.800 1062.070 79.860 ;
        RECT 1980.370 79.800 1980.690 79.860 ;
        RECT 1061.750 79.660 1980.690 79.800 ;
        RECT 1061.750 79.600 1062.070 79.660 ;
        RECT 1980.370 79.600 1980.690 79.660 ;
        RECT 1980.370 62.120 1980.690 62.180 ;
        RECT 1983.130 62.120 1983.450 62.180 ;
        RECT 1980.370 61.980 1983.450 62.120 ;
        RECT 1980.370 61.920 1980.690 61.980 ;
        RECT 1983.130 61.920 1983.450 61.980 ;
      LAYER via ;
        RECT 1056.260 243.820 1056.520 244.080 ;
        RECT 1061.780 243.820 1062.040 244.080 ;
        RECT 1061.780 79.600 1062.040 79.860 ;
        RECT 1980.400 79.600 1980.660 79.860 ;
        RECT 1980.400 61.920 1980.660 62.180 ;
        RECT 1983.160 61.920 1983.420 62.180 ;
      LAYER met2 ;
        RECT 1056.210 260.000 1056.490 264.000 ;
        RECT 1056.320 244.110 1056.460 260.000 ;
        RECT 1056.260 243.790 1056.520 244.110 ;
        RECT 1061.780 243.790 1062.040 244.110 ;
        RECT 1061.840 79.890 1061.980 243.790 ;
        RECT 1061.780 79.570 1062.040 79.890 ;
        RECT 1980.400 79.570 1980.660 79.890 ;
        RECT 1980.460 62.210 1980.600 79.570 ;
        RECT 1980.400 61.890 1980.660 62.210 ;
        RECT 1983.160 61.890 1983.420 62.210 ;
        RECT 1983.220 2.400 1983.360 61.890 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1384.670 246.400 1384.990 246.460 ;
        RECT 1618.350 246.400 1618.670 246.460 ;
        RECT 1384.670 246.260 1618.670 246.400 ;
        RECT 1384.670 246.200 1384.990 246.260 ;
        RECT 1618.350 246.200 1618.670 246.260 ;
        RECT 1618.350 107.340 1618.670 107.400 ;
        RECT 2001.070 107.340 2001.390 107.400 ;
        RECT 1618.350 107.200 2001.390 107.340 ;
        RECT 1618.350 107.140 1618.670 107.200 ;
        RECT 2001.070 107.140 2001.390 107.200 ;
      LAYER via ;
        RECT 1384.700 246.200 1384.960 246.460 ;
        RECT 1618.380 246.200 1618.640 246.460 ;
        RECT 1618.380 107.140 1618.640 107.400 ;
        RECT 2001.100 107.140 2001.360 107.400 ;
      LAYER met2 ;
        RECT 1384.650 260.000 1384.930 264.000 ;
        RECT 1384.760 246.490 1384.900 260.000 ;
        RECT 1384.700 246.170 1384.960 246.490 ;
        RECT 1618.380 246.170 1618.640 246.490 ;
        RECT 1618.440 107.430 1618.580 246.170 ;
        RECT 1618.380 107.110 1618.640 107.430 ;
        RECT 2001.100 107.110 2001.360 107.430 ;
        RECT 2001.160 2.400 2001.300 107.110 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 220.410 73.340 220.730 73.400 ;
        RECT 2014.870 73.340 2015.190 73.400 ;
        RECT 220.410 73.200 2015.190 73.340 ;
        RECT 220.410 73.140 220.730 73.200 ;
        RECT 2014.870 73.140 2015.190 73.200 ;
        RECT 2014.870 14.180 2015.190 14.240 ;
        RECT 2014.870 14.040 2018.780 14.180 ;
        RECT 2014.870 13.980 2015.190 14.040 ;
        RECT 2018.640 13.900 2018.780 14.040 ;
        RECT 2018.550 13.640 2018.870 13.900 ;
      LAYER via ;
        RECT 220.440 73.140 220.700 73.400 ;
        RECT 2014.900 73.140 2015.160 73.400 ;
        RECT 2014.900 13.980 2015.160 14.240 ;
        RECT 2018.580 13.640 2018.840 13.900 ;
      LAYER met2 ;
        RECT 220.430 3258.035 220.710 3258.405 ;
        RECT 662.030 3258.290 662.310 3258.405 ;
        RECT 662.450 3258.290 662.730 3260.000 ;
        RECT 662.030 3258.150 662.730 3258.290 ;
        RECT 662.030 3258.035 662.310 3258.150 ;
        RECT 220.500 73.430 220.640 3258.035 ;
        RECT 662.450 3256.000 662.730 3258.150 ;
        RECT 220.440 73.110 220.700 73.430 ;
        RECT 2014.900 73.110 2015.160 73.430 ;
        RECT 2014.960 14.270 2015.100 73.110 ;
        RECT 2014.900 13.950 2015.160 14.270 ;
        RECT 2018.580 13.610 2018.840 13.930 ;
        RECT 2018.640 2.400 2018.780 13.610 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
      LAYER via2 ;
        RECT 220.430 3258.080 220.710 3258.360 ;
        RECT 662.030 3258.080 662.310 3258.360 ;
      LAYER met3 ;
        RECT 220.405 3258.370 220.735 3258.385 ;
        RECT 662.005 3258.370 662.335 3258.385 ;
        RECT 220.405 3258.070 662.335 3258.370 ;
        RECT 220.405 3258.055 220.735 3258.070 ;
        RECT 662.005 3258.055 662.335 3258.070 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2035.645 144.925 2035.815 192.695 ;
        RECT 2035.645 48.365 2035.815 96.475 ;
      LAYER mcon ;
        RECT 2035.645 192.525 2035.815 192.695 ;
        RECT 2035.645 96.305 2035.815 96.475 ;
      LAYER met1 ;
        RECT 1377.310 3265.940 1377.630 3266.000 ;
        RECT 2621.150 3265.940 2621.470 3266.000 ;
        RECT 1377.310 3265.800 2621.470 3265.940 ;
        RECT 1377.310 3265.740 1377.630 3265.800 ;
        RECT 2621.150 3265.740 2621.470 3265.800 ;
        RECT 2614.710 372.540 2615.030 372.600 ;
        RECT 2621.150 372.540 2621.470 372.600 ;
        RECT 2614.710 372.400 2621.470 372.540 ;
        RECT 2614.710 372.340 2615.030 372.400 ;
        RECT 2621.150 372.340 2621.470 372.400 ;
        RECT 2615.170 264.080 2615.490 264.140 ;
        RECT 2035.660 263.940 2615.490 264.080 ;
        RECT 2035.660 263.800 2035.800 263.940 ;
        RECT 2615.170 263.880 2615.490 263.940 ;
        RECT 2035.570 263.540 2035.890 263.800 ;
        RECT 2035.570 193.840 2035.890 194.100 ;
        RECT 2035.660 193.420 2035.800 193.840 ;
        RECT 2035.570 193.160 2035.890 193.420 ;
        RECT 2035.570 192.680 2035.890 192.740 ;
        RECT 2035.375 192.540 2035.890 192.680 ;
        RECT 2035.570 192.480 2035.890 192.540 ;
        RECT 2035.570 145.080 2035.890 145.140 ;
        RECT 2035.375 144.940 2035.890 145.080 ;
        RECT 2035.570 144.880 2035.890 144.940 ;
        RECT 2035.570 96.460 2035.890 96.520 ;
        RECT 2035.375 96.320 2035.890 96.460 ;
        RECT 2035.570 96.260 2035.890 96.320 ;
        RECT 2035.570 48.520 2035.890 48.580 ;
        RECT 2035.375 48.380 2035.890 48.520 ;
        RECT 2035.570 48.320 2035.890 48.380 ;
        RECT 2035.570 14.180 2035.890 14.240 ;
        RECT 2035.570 14.040 2036.720 14.180 ;
        RECT 2035.570 13.980 2035.890 14.040 ;
        RECT 2036.580 13.900 2036.720 14.040 ;
        RECT 2036.490 13.640 2036.810 13.900 ;
      LAYER via ;
        RECT 1377.340 3265.740 1377.600 3266.000 ;
        RECT 2621.180 3265.740 2621.440 3266.000 ;
        RECT 2614.740 372.340 2615.000 372.600 ;
        RECT 2621.180 372.340 2621.440 372.600 ;
        RECT 2615.200 263.880 2615.460 264.140 ;
        RECT 2035.600 263.540 2035.860 263.800 ;
        RECT 2035.600 193.840 2035.860 194.100 ;
        RECT 2035.600 193.160 2035.860 193.420 ;
        RECT 2035.600 192.480 2035.860 192.740 ;
        RECT 2035.600 144.880 2035.860 145.140 ;
        RECT 2035.600 96.260 2035.860 96.520 ;
        RECT 2035.600 48.320 2035.860 48.580 ;
        RECT 2035.600 13.980 2035.860 14.240 ;
        RECT 2036.520 13.640 2036.780 13.900 ;
      LAYER met2 ;
        RECT 1377.340 3265.710 1377.600 3266.030 ;
        RECT 2621.180 3265.710 2621.440 3266.030 ;
        RECT 1377.400 3260.000 1377.540 3265.710 ;
        RECT 1377.290 3256.000 1377.570 3260.000 ;
        RECT 2621.240 372.630 2621.380 3265.710 ;
        RECT 2614.740 372.310 2615.000 372.630 ;
        RECT 2621.180 372.310 2621.440 372.630 ;
        RECT 2614.800 291.450 2614.940 372.310 ;
        RECT 2614.800 291.310 2615.400 291.450 ;
        RECT 2615.260 264.170 2615.400 291.310 ;
        RECT 2615.200 263.850 2615.460 264.170 ;
        RECT 2035.600 263.510 2035.860 263.830 ;
        RECT 2035.660 194.130 2035.800 263.510 ;
        RECT 2035.600 193.810 2035.860 194.130 ;
        RECT 2035.600 193.130 2035.860 193.450 ;
        RECT 2035.660 192.770 2035.800 193.130 ;
        RECT 2035.600 192.450 2035.860 192.770 ;
        RECT 2035.600 144.850 2035.860 145.170 ;
        RECT 2035.660 96.550 2035.800 144.850 ;
        RECT 2035.600 96.230 2035.860 96.550 ;
        RECT 2035.600 48.290 2035.860 48.610 ;
        RECT 2035.660 14.270 2035.800 48.290 ;
        RECT 2035.600 13.950 2035.860 14.270 ;
        RECT 2036.520 13.610 2036.780 13.930 ;
        RECT 2036.580 2.400 2036.720 13.610 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2055.885 48.365 2056.055 96.475 ;
      LAYER mcon ;
        RECT 2055.885 96.305 2056.055 96.475 ;
      LAYER met1 ;
        RECT 2620.690 2346.240 2621.010 2346.300 ;
        RECT 2638.170 2346.240 2638.490 2346.300 ;
        RECT 2620.690 2346.100 2638.490 2346.240 ;
        RECT 2620.690 2346.040 2621.010 2346.100 ;
        RECT 2638.170 2346.040 2638.490 2346.100 ;
        RECT 2055.350 135.220 2055.670 135.280 ;
        RECT 2638.170 135.220 2638.490 135.280 ;
        RECT 2055.350 135.080 2638.490 135.220 ;
        RECT 2055.350 135.020 2055.670 135.080 ;
        RECT 2638.170 135.020 2638.490 135.080 ;
        RECT 2055.810 96.460 2056.130 96.520 ;
        RECT 2055.615 96.320 2056.130 96.460 ;
        RECT 2055.810 96.260 2056.130 96.320 ;
        RECT 2055.810 48.520 2056.130 48.580 ;
        RECT 2055.615 48.380 2056.130 48.520 ;
        RECT 2055.810 48.320 2056.130 48.380 ;
      LAYER via ;
        RECT 2620.720 2346.040 2620.980 2346.300 ;
        RECT 2638.200 2346.040 2638.460 2346.300 ;
        RECT 2055.380 135.020 2055.640 135.280 ;
        RECT 2638.200 135.020 2638.460 135.280 ;
        RECT 2055.840 96.260 2056.100 96.520 ;
        RECT 2055.840 48.320 2056.100 48.580 ;
      LAYER met2 ;
        RECT 2620.710 2346.155 2620.990 2346.525 ;
        RECT 2620.720 2346.010 2620.980 2346.155 ;
        RECT 2638.200 2346.010 2638.460 2346.330 ;
        RECT 2638.260 135.310 2638.400 2346.010 ;
        RECT 2055.380 134.990 2055.640 135.310 ;
        RECT 2638.200 134.990 2638.460 135.310 ;
        RECT 2055.440 96.970 2055.580 134.990 ;
        RECT 2055.440 96.830 2056.040 96.970 ;
        RECT 2055.900 96.550 2056.040 96.830 ;
        RECT 2055.840 96.230 2056.100 96.550 ;
        RECT 2055.840 48.290 2056.100 48.610 ;
        RECT 2055.900 14.010 2056.040 48.290 ;
        RECT 2054.980 13.870 2056.040 14.010 ;
        RECT 2054.980 13.330 2055.120 13.870 ;
        RECT 2054.520 13.190 2055.120 13.330 ;
        RECT 2054.520 2.400 2054.660 13.190 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
      LAYER via2 ;
        RECT 2620.710 2346.200 2620.990 2346.480 ;
      LAYER met3 ;
        RECT 2606.000 2346.490 2610.000 2346.880 ;
        RECT 2620.685 2346.490 2621.015 2346.505 ;
        RECT 2606.000 2346.280 2621.015 2346.490 ;
        RECT 2609.580 2346.190 2621.015 2346.280 ;
        RECT 2620.685 2346.175 2621.015 2346.190 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 261.810 3275.800 262.130 3275.860 ;
        RECT 490.430 3275.800 490.750 3275.860 ;
        RECT 261.810 3275.660 490.750 3275.800 ;
        RECT 261.810 3275.600 262.130 3275.660 ;
        RECT 490.430 3275.600 490.750 3275.660 ;
      LAYER via ;
        RECT 261.840 3275.600 262.100 3275.860 ;
        RECT 490.460 3275.600 490.720 3275.860 ;
      LAYER met2 ;
        RECT 261.840 3275.570 262.100 3275.890 ;
        RECT 490.460 3275.570 490.720 3275.890 ;
        RECT 261.900 20.245 262.040 3275.570 ;
        RECT 490.520 3260.000 490.660 3275.570 ;
        RECT 490.410 3256.000 490.690 3260.000 ;
        RECT 261.830 19.875 262.110 20.245 ;
        RECT 769.670 19.875 769.950 20.245 ;
        RECT 769.740 2.400 769.880 19.875 ;
        RECT 769.530 -4.800 770.090 2.400 ;
      LAYER via2 ;
        RECT 261.830 19.920 262.110 20.200 ;
        RECT 769.670 19.920 769.950 20.200 ;
      LAYER met3 ;
        RECT 261.805 20.210 262.135 20.225 ;
        RECT 769.645 20.210 769.975 20.225 ;
        RECT 261.805 19.910 769.975 20.210 ;
        RECT 261.805 19.895 262.135 19.910 ;
        RECT 769.645 19.895 769.975 19.910 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 232.370 2629.120 232.690 2629.180 ;
        RECT 296.770 2629.120 297.090 2629.180 ;
        RECT 232.370 2628.980 297.090 2629.120 ;
        RECT 232.370 2628.920 232.690 2628.980 ;
        RECT 296.770 2628.920 297.090 2628.980 ;
        RECT 232.370 47.160 232.690 47.220 ;
        RECT 2072.370 47.160 2072.690 47.220 ;
        RECT 232.370 47.020 2072.690 47.160 ;
        RECT 232.370 46.960 232.690 47.020 ;
        RECT 2072.370 46.960 2072.690 47.020 ;
      LAYER via ;
        RECT 232.400 2628.920 232.660 2629.180 ;
        RECT 296.800 2628.920 297.060 2629.180 ;
        RECT 232.400 46.960 232.660 47.220 ;
        RECT 2072.400 46.960 2072.660 47.220 ;
      LAYER met2 ;
        RECT 296.790 2630.395 297.070 2630.765 ;
        RECT 296.860 2629.210 297.000 2630.395 ;
        RECT 232.400 2628.890 232.660 2629.210 ;
        RECT 296.800 2628.890 297.060 2629.210 ;
        RECT 232.460 47.250 232.600 2628.890 ;
        RECT 232.400 46.930 232.660 47.250 ;
        RECT 2072.400 46.930 2072.660 47.250 ;
        RECT 2072.460 2.400 2072.600 46.930 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
      LAYER via2 ;
        RECT 296.790 2630.440 297.070 2630.720 ;
      LAYER met3 ;
        RECT 296.765 2630.730 297.095 2630.745 ;
        RECT 310.000 2630.730 314.000 2631.120 ;
        RECT 296.765 2630.520 314.000 2630.730 ;
        RECT 296.765 2630.430 310.500 2630.520 ;
        RECT 296.765 2630.415 297.095 2630.430 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 219.950 3112.260 220.270 3112.320 ;
        RECT 296.770 3112.260 297.090 3112.320 ;
        RECT 219.950 3112.120 297.090 3112.260 ;
        RECT 219.950 3112.060 220.270 3112.120 ;
        RECT 296.770 3112.060 297.090 3112.120 ;
        RECT 219.950 72.660 220.270 72.720 ;
        RECT 2084.330 72.660 2084.650 72.720 ;
        RECT 219.950 72.520 2084.650 72.660 ;
        RECT 219.950 72.460 220.270 72.520 ;
        RECT 2084.330 72.460 2084.650 72.520 ;
        RECT 2084.790 2.960 2085.110 3.020 ;
        RECT 2089.850 2.960 2090.170 3.020 ;
        RECT 2084.790 2.820 2090.170 2.960 ;
        RECT 2084.790 2.760 2085.110 2.820 ;
        RECT 2089.850 2.760 2090.170 2.820 ;
      LAYER via ;
        RECT 219.980 3112.060 220.240 3112.320 ;
        RECT 296.800 3112.060 297.060 3112.320 ;
        RECT 219.980 72.460 220.240 72.720 ;
        RECT 2084.360 72.460 2084.620 72.720 ;
        RECT 2084.820 2.760 2085.080 3.020 ;
        RECT 2089.880 2.760 2090.140 3.020 ;
      LAYER met2 ;
        RECT 296.790 3117.275 297.070 3117.645 ;
        RECT 296.860 3112.350 297.000 3117.275 ;
        RECT 219.980 3112.030 220.240 3112.350 ;
        RECT 296.800 3112.030 297.060 3112.350 ;
        RECT 220.040 72.750 220.180 3112.030 ;
        RECT 219.980 72.430 220.240 72.750 ;
        RECT 2084.360 72.430 2084.620 72.750 ;
        RECT 2084.420 38.490 2084.560 72.430 ;
        RECT 2084.420 38.350 2085.020 38.490 ;
        RECT 2084.880 3.050 2085.020 38.350 ;
        RECT 2084.820 2.730 2085.080 3.050 ;
        RECT 2089.880 2.730 2090.140 3.050 ;
        RECT 2089.940 2.400 2090.080 2.730 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
      LAYER via2 ;
        RECT 296.790 3117.320 297.070 3117.600 ;
      LAYER met3 ;
        RECT 296.765 3117.610 297.095 3117.625 ;
        RECT 310.000 3117.610 314.000 3118.000 ;
        RECT 296.765 3117.400 314.000 3117.610 ;
        RECT 296.765 3117.310 310.500 3117.400 ;
        RECT 296.765 3117.295 297.095 3117.310 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1014.460 2615.490 1014.520 ;
        RECT 2631.730 1014.460 2632.050 1014.520 ;
        RECT 2615.170 1014.320 2632.050 1014.460 ;
        RECT 2615.170 1014.260 2615.490 1014.320 ;
        RECT 2631.730 1014.260 2632.050 1014.320 ;
        RECT 2111.010 246.060 2111.330 246.120 ;
        RECT 2631.730 246.060 2632.050 246.120 ;
        RECT 2111.010 245.920 2632.050 246.060 ;
        RECT 2111.010 245.860 2111.330 245.920 ;
        RECT 2631.730 245.860 2632.050 245.920 ;
        RECT 2107.790 17.920 2108.110 17.980 ;
        RECT 2111.010 17.920 2111.330 17.980 ;
        RECT 2107.790 17.780 2111.330 17.920 ;
        RECT 2107.790 17.720 2108.110 17.780 ;
        RECT 2111.010 17.720 2111.330 17.780 ;
      LAYER via ;
        RECT 2615.200 1014.260 2615.460 1014.520 ;
        RECT 2631.760 1014.260 2632.020 1014.520 ;
        RECT 2111.040 245.860 2111.300 246.120 ;
        RECT 2631.760 245.860 2632.020 246.120 ;
        RECT 2107.820 17.720 2108.080 17.980 ;
        RECT 2111.040 17.720 2111.300 17.980 ;
      LAYER met2 ;
        RECT 2615.190 1014.715 2615.470 1015.085 ;
        RECT 2615.260 1014.550 2615.400 1014.715 ;
        RECT 2615.200 1014.230 2615.460 1014.550 ;
        RECT 2631.760 1014.230 2632.020 1014.550 ;
        RECT 2631.820 246.150 2631.960 1014.230 ;
        RECT 2111.040 245.830 2111.300 246.150 ;
        RECT 2631.760 245.830 2632.020 246.150 ;
        RECT 2111.100 18.010 2111.240 245.830 ;
        RECT 2107.820 17.690 2108.080 18.010 ;
        RECT 2111.040 17.690 2111.300 18.010 ;
        RECT 2107.880 2.400 2108.020 17.690 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1014.760 2615.470 1015.040 ;
      LAYER met3 ;
        RECT 2606.000 1015.050 2610.000 1015.440 ;
        RECT 2615.165 1015.050 2615.495 1015.065 ;
        RECT 2606.000 1014.840 2615.495 1015.050 ;
        RECT 2609.580 1014.750 2615.495 1014.840 ;
        RECT 2615.165 1014.735 2615.495 1014.750 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1591.670 3272.060 1591.990 3272.120 ;
        RECT 2539.270 3272.060 2539.590 3272.120 ;
        RECT 1591.670 3271.920 2539.590 3272.060 ;
        RECT 1591.670 3271.860 1591.990 3271.920 ;
        RECT 2539.270 3271.860 2539.590 3271.920 ;
        RECT 2539.270 3268.320 2539.590 3268.380 ;
        RECT 2643.690 3268.320 2644.010 3268.380 ;
        RECT 2539.270 3268.180 2644.010 3268.320 ;
        RECT 2539.270 3268.120 2539.590 3268.180 ;
        RECT 2643.690 3268.120 2644.010 3268.180 ;
        RECT 2125.270 263.400 2125.590 263.460 ;
        RECT 2643.690 263.400 2644.010 263.460 ;
        RECT 2125.270 263.260 2644.010 263.400 ;
        RECT 2125.270 263.200 2125.590 263.260 ;
        RECT 2643.690 263.200 2644.010 263.260 ;
      LAYER via ;
        RECT 1591.700 3271.860 1591.960 3272.120 ;
        RECT 2539.300 3271.860 2539.560 3272.120 ;
        RECT 2539.300 3268.120 2539.560 3268.380 ;
        RECT 2643.720 3268.120 2643.980 3268.380 ;
        RECT 2125.300 263.200 2125.560 263.460 ;
        RECT 2643.720 263.200 2643.980 263.460 ;
      LAYER met2 ;
        RECT 1591.700 3271.830 1591.960 3272.150 ;
        RECT 2539.300 3271.830 2539.560 3272.150 ;
        RECT 1591.760 3260.000 1591.900 3271.830 ;
        RECT 2539.360 3268.410 2539.500 3271.830 ;
        RECT 2539.300 3268.090 2539.560 3268.410 ;
        RECT 2643.720 3268.090 2643.980 3268.410 ;
        RECT 1591.650 3256.000 1591.930 3260.000 ;
        RECT 2643.780 263.490 2643.920 3268.090 ;
        RECT 2125.300 263.170 2125.560 263.490 ;
        RECT 2643.720 263.170 2643.980 263.490 ;
        RECT 2125.360 37.130 2125.500 263.170 ;
        RECT 2125.360 36.990 2125.960 37.130 ;
        RECT 2125.820 2.400 2125.960 36.990 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2102.345 16.745 2102.515 17.935 ;
      LAYER mcon ;
        RECT 2102.345 17.765 2102.515 17.935 ;
      LAYER met1 ;
        RECT 279.750 704.040 280.070 704.100 ;
        RECT 296.770 704.040 297.090 704.100 ;
        RECT 279.750 703.900 297.090 704.040 ;
        RECT 279.750 703.840 280.070 703.900 ;
        RECT 296.770 703.840 297.090 703.900 ;
        RECT 279.750 17.920 280.070 17.980 ;
        RECT 2102.285 17.920 2102.575 17.965 ;
        RECT 279.750 17.780 2102.575 17.920 ;
        RECT 279.750 17.720 280.070 17.780 ;
        RECT 2102.285 17.735 2102.575 17.780 ;
        RECT 2102.285 16.900 2102.575 16.945 ;
        RECT 2143.670 16.900 2143.990 16.960 ;
        RECT 2102.285 16.760 2143.990 16.900 ;
        RECT 2102.285 16.715 2102.575 16.760 ;
        RECT 2143.670 16.700 2143.990 16.760 ;
      LAYER via ;
        RECT 279.780 703.840 280.040 704.100 ;
        RECT 296.800 703.840 297.060 704.100 ;
        RECT 279.780 17.720 280.040 17.980 ;
        RECT 2143.700 16.700 2143.960 16.960 ;
      LAYER met2 ;
        RECT 296.790 707.355 297.070 707.725 ;
        RECT 296.860 704.130 297.000 707.355 ;
        RECT 279.780 703.810 280.040 704.130 ;
        RECT 296.800 703.810 297.060 704.130 ;
        RECT 279.840 18.010 279.980 703.810 ;
        RECT 279.780 17.690 280.040 18.010 ;
        RECT 2143.700 16.670 2143.960 16.990 ;
        RECT 2143.760 2.400 2143.900 16.670 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
      LAYER via2 ;
        RECT 296.790 707.400 297.070 707.680 ;
      LAYER met3 ;
        RECT 296.765 707.690 297.095 707.705 ;
        RECT 310.000 707.690 314.000 708.080 ;
        RECT 296.765 707.480 314.000 707.690 ;
        RECT 296.765 707.390 310.500 707.480 ;
        RECT 296.765 707.375 297.095 707.390 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.210 247.420 2166.530 247.480 ;
        RECT 2609.650 247.420 2609.970 247.480 ;
        RECT 2166.210 247.280 2609.970 247.420 ;
        RECT 2166.210 247.220 2166.530 247.280 ;
        RECT 2609.650 247.220 2609.970 247.280 ;
        RECT 2161.610 14.520 2161.930 14.580 ;
        RECT 2166.210 14.520 2166.530 14.580 ;
        RECT 2161.610 14.380 2166.530 14.520 ;
        RECT 2161.610 14.320 2161.930 14.380 ;
        RECT 2166.210 14.320 2166.530 14.380 ;
      LAYER via ;
        RECT 2166.240 247.220 2166.500 247.480 ;
        RECT 2609.680 247.220 2609.940 247.480 ;
        RECT 2161.640 14.320 2161.900 14.580 ;
        RECT 2166.240 14.320 2166.500 14.580 ;
      LAYER met2 ;
        RECT 2609.670 1373.075 2609.950 1373.445 ;
        RECT 2609.740 247.510 2609.880 1373.075 ;
        RECT 2166.240 247.190 2166.500 247.510 ;
        RECT 2609.680 247.190 2609.940 247.510 ;
        RECT 2166.300 14.610 2166.440 247.190 ;
        RECT 2161.640 14.290 2161.900 14.610 ;
        RECT 2166.240 14.290 2166.500 14.610 ;
        RECT 2161.700 2.400 2161.840 14.290 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 2609.670 1373.120 2609.950 1373.400 ;
      LAYER met3 ;
        RECT 2606.000 1373.880 2610.000 1374.480 ;
        RECT 2609.430 1373.425 2609.730 1373.880 ;
        RECT 2609.430 1373.110 2609.975 1373.425 ;
        RECT 2609.645 1373.095 2609.975 1373.110 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 14.180 2180.330 14.240 ;
        RECT 2179.180 14.040 2180.330 14.180 ;
        RECT 2179.180 13.900 2179.320 14.040 ;
        RECT 2180.010 13.980 2180.330 14.040 ;
        RECT 2179.090 13.640 2179.410 13.900 ;
      LAYER via ;
        RECT 2180.040 13.980 2180.300 14.240 ;
        RECT 2179.120 13.640 2179.380 13.900 ;
      LAYER met2 ;
        RECT 2180.030 155.195 2180.310 155.565 ;
        RECT 2180.100 14.270 2180.240 155.195 ;
        RECT 2180.040 13.950 2180.300 14.270 ;
        RECT 2179.120 13.610 2179.380 13.930 ;
        RECT 2179.180 2.400 2179.320 13.610 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
      LAYER via2 ;
        RECT 2180.030 155.240 2180.310 155.520 ;
      LAYER met3 ;
        RECT 2606.000 2747.480 2610.000 2748.080 ;
        RECT 2606.670 2744.300 2606.970 2747.480 ;
        RECT 2606.630 2743.980 2607.010 2744.300 ;
        RECT 2180.005 155.530 2180.335 155.545 ;
        RECT 2600.190 155.530 2600.570 155.540 ;
        RECT 2180.005 155.230 2600.570 155.530 ;
        RECT 2180.005 155.215 2180.335 155.230 ;
        RECT 2600.190 155.220 2600.570 155.230 ;
      LAYER via3 ;
        RECT 2606.660 2743.980 2606.980 2744.300 ;
        RECT 2600.220 155.220 2600.540 155.540 ;
      LAYER met4 ;
        RECT 2606.655 2743.975 2606.985 2744.305 ;
        RECT 2606.670 2715.490 2606.970 2743.975 ;
        RECT 2597.950 2714.310 2599.130 2715.490 ;
        RECT 2606.230 2714.310 2607.410 2715.490 ;
        RECT 2598.390 2677.650 2598.690 2714.310 ;
        RECT 2598.390 2677.350 2600.530 2677.650 ;
        RECT 2600.230 2415.850 2600.530 2677.350 ;
        RECT 2598.390 2415.550 2600.530 2415.850 ;
        RECT 2598.390 2405.650 2598.690 2415.550 ;
        RECT 2598.390 2405.350 2600.530 2405.650 ;
        RECT 2600.230 2358.050 2600.530 2405.350 ;
        RECT 2597.470 2357.750 2600.530 2358.050 ;
        RECT 2597.470 2324.050 2597.770 2357.750 ;
        RECT 2597.470 2323.750 2600.530 2324.050 ;
        RECT 2600.230 2001.050 2600.530 2323.750 ;
        RECT 2598.390 2000.750 2600.530 2001.050 ;
        RECT 2598.390 1939.850 2598.690 2000.750 ;
        RECT 2598.390 1939.550 2600.530 1939.850 ;
        RECT 2600.230 1875.250 2600.530 1939.550 ;
        RECT 2598.390 1874.950 2600.530 1875.250 ;
        RECT 2598.390 1851.450 2598.690 1874.950 ;
        RECT 2598.390 1851.150 2599.610 1851.450 ;
        RECT 2599.310 1810.650 2599.610 1851.150 ;
        RECT 2599.310 1810.350 2600.530 1810.650 ;
        RECT 2600.230 1752.850 2600.530 1810.350 ;
        RECT 2598.390 1752.550 2600.530 1752.850 ;
        RECT 2598.390 1742.650 2598.690 1752.550 ;
        RECT 2598.390 1742.350 2599.610 1742.650 ;
        RECT 2599.310 1739.250 2599.610 1742.350 ;
        RECT 2599.310 1738.950 2600.530 1739.250 ;
        RECT 2600.230 1718.850 2600.530 1738.950 ;
        RECT 2597.470 1718.550 2600.530 1718.850 ;
        RECT 2597.470 1661.050 2597.770 1718.550 ;
        RECT 2597.470 1660.750 2600.530 1661.050 ;
        RECT 2600.230 1559.050 2600.530 1660.750 ;
        RECT 2599.310 1558.750 2600.530 1559.050 ;
        RECT 2599.310 1535.250 2599.610 1558.750 ;
        RECT 2598.390 1534.950 2599.610 1535.250 ;
        RECT 2598.390 1474.050 2598.690 1534.950 ;
        RECT 2598.390 1473.750 2600.530 1474.050 ;
        RECT 2600.230 1242.850 2600.530 1473.750 ;
        RECT 2600.230 1242.550 2601.450 1242.850 ;
        RECT 2601.150 1236.050 2601.450 1242.550 ;
        RECT 2600.230 1235.750 2601.450 1236.050 ;
        RECT 2600.230 1191.850 2600.530 1235.750 ;
        RECT 2600.230 1191.550 2604.210 1191.850 ;
        RECT 2603.910 1174.850 2604.210 1191.550 ;
        RECT 2602.990 1174.550 2604.210 1174.850 ;
        RECT 2602.990 1103.450 2603.290 1174.550 ;
        RECT 2600.230 1103.150 2603.290 1103.450 ;
        RECT 2600.230 1038.850 2600.530 1103.150 ;
        RECT 2600.230 1038.550 2601.450 1038.850 ;
        RECT 2601.150 1032.050 2601.450 1038.550 ;
        RECT 2600.230 1031.750 2601.450 1032.050 ;
        RECT 2600.230 749.850 2600.530 1031.750 ;
        RECT 2600.230 749.550 2602.370 749.850 ;
        RECT 2602.070 736.250 2602.370 749.550 ;
        RECT 2600.230 735.950 2602.370 736.250 ;
        RECT 2600.230 719.250 2600.530 735.950 ;
        RECT 2598.390 718.950 2600.530 719.250 ;
        RECT 2598.390 692.050 2598.690 718.950 ;
        RECT 2598.390 691.750 2600.530 692.050 ;
        RECT 2600.230 634.250 2600.530 691.750 ;
        RECT 2599.310 633.950 2600.530 634.250 ;
        RECT 2599.310 610.450 2599.610 633.950 ;
        RECT 2598.390 610.150 2599.610 610.450 ;
        RECT 2598.390 607.050 2598.690 610.150 ;
        RECT 2598.390 606.750 2599.610 607.050 ;
        RECT 2599.310 559.450 2599.610 606.750 ;
        RECT 2599.310 559.150 2600.530 559.450 ;
        RECT 2600.230 505.050 2600.530 559.150 ;
        RECT 2599.310 504.750 2600.530 505.050 ;
        RECT 2599.310 501.650 2599.610 504.750 ;
        RECT 2599.310 501.350 2600.530 501.650 ;
        RECT 2600.230 426.850 2600.530 501.350 ;
        RECT 2599.310 426.550 2600.530 426.850 ;
        RECT 2599.310 352.050 2599.610 426.550 ;
        RECT 2599.310 351.750 2600.530 352.050 ;
        RECT 2600.230 155.545 2600.530 351.750 ;
        RECT 2600.215 155.215 2600.545 155.545 ;
      LAYER met5 ;
        RECT 2597.740 2714.100 2607.620 2715.700 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2507.070 3275.800 2507.390 3275.860 ;
        RECT 2646.910 3275.800 2647.230 3275.860 ;
        RECT 2507.070 3275.660 2647.230 3275.800 ;
        RECT 2507.070 3275.600 2507.390 3275.660 ;
        RECT 2646.910 3275.600 2647.230 3275.660 ;
        RECT 2197.030 18.940 2197.350 19.000 ;
        RECT 2200.710 18.940 2201.030 19.000 ;
        RECT 2197.030 18.800 2201.030 18.940 ;
        RECT 2197.030 18.740 2197.350 18.800 ;
        RECT 2200.710 18.740 2201.030 18.800 ;
      LAYER via ;
        RECT 2507.100 3275.600 2507.360 3275.860 ;
        RECT 2646.940 3275.600 2647.200 3275.860 ;
        RECT 2197.060 18.740 2197.320 19.000 ;
        RECT 2200.740 18.740 2201.000 19.000 ;
      LAYER met2 ;
        RECT 2507.100 3275.570 2507.360 3275.890 ;
        RECT 2646.940 3275.570 2647.200 3275.890 ;
        RECT 2507.160 3260.000 2507.300 3275.570 ;
        RECT 2507.050 3256.000 2507.330 3260.000 ;
        RECT 2647.000 260.285 2647.140 3275.570 ;
        RECT 2201.190 260.170 2201.470 260.285 ;
        RECT 2200.800 260.030 2201.470 260.170 ;
        RECT 2200.800 19.030 2200.940 260.030 ;
        RECT 2201.190 259.915 2201.470 260.030 ;
        RECT 2646.930 259.915 2647.210 260.285 ;
        RECT 2197.060 18.710 2197.320 19.030 ;
        RECT 2200.740 18.710 2201.000 19.030 ;
        RECT 2197.120 2.400 2197.260 18.710 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
      LAYER via2 ;
        RECT 2201.190 259.960 2201.470 260.240 ;
        RECT 2646.930 259.960 2647.210 260.240 ;
      LAYER met3 ;
        RECT 2201.165 260.250 2201.495 260.265 ;
        RECT 2646.905 260.250 2647.235 260.265 ;
        RECT 2201.165 259.950 2647.235 260.250 ;
        RECT 2201.165 259.935 2201.495 259.950 ;
        RECT 2646.905 259.935 2647.235 259.950 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.990 19.195 2215.270 19.565 ;
        RECT 2585.290 19.195 2585.570 19.565 ;
        RECT 2215.060 2.400 2215.200 19.195 ;
        RECT 2585.360 15.485 2585.500 19.195 ;
        RECT 2585.290 15.115 2585.570 15.485 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
      LAYER via2 ;
        RECT 2214.990 19.240 2215.270 19.520 ;
        RECT 2585.290 19.240 2585.570 19.520 ;
        RECT 2585.290 15.160 2585.570 15.440 ;
      LAYER met3 ;
        RECT 2606.000 804.250 2610.000 804.640 ;
        RECT 2620.430 804.250 2620.810 804.260 ;
        RECT 2606.000 804.040 2620.810 804.250 ;
        RECT 2609.580 803.950 2620.810 804.040 ;
        RECT 2620.430 803.940 2620.810 803.950 ;
        RECT 2214.965 19.530 2215.295 19.545 ;
        RECT 2585.265 19.530 2585.595 19.545 ;
        RECT 2214.965 19.230 2585.595 19.530 ;
        RECT 2214.965 19.215 2215.295 19.230 ;
        RECT 2585.265 19.215 2585.595 19.230 ;
        RECT 2585.265 15.450 2585.595 15.465 ;
        RECT 2598.350 15.450 2598.730 15.460 ;
        RECT 2585.265 15.150 2598.730 15.450 ;
        RECT 2585.265 15.135 2585.595 15.150 ;
        RECT 2598.350 15.140 2598.730 15.150 ;
      LAYER via3 ;
        RECT 2620.460 803.940 2620.780 804.260 ;
        RECT 2598.380 15.140 2598.700 15.460 ;
      LAYER met4 ;
        RECT 2620.455 803.935 2620.785 804.265 ;
        RECT 2620.470 536.090 2620.770 803.935 ;
        RECT 2597.950 534.910 2599.130 536.090 ;
        RECT 2620.030 534.910 2621.210 536.090 ;
        RECT 2598.390 15.465 2598.690 534.910 ;
        RECT 2598.375 15.135 2598.705 15.465 ;
      LAYER met5 ;
        RECT 2597.740 534.700 2621.420 536.300 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2228.770 62.120 2229.090 62.180 ;
        RECT 2232.910 62.120 2233.230 62.180 ;
        RECT 2228.770 61.980 2233.230 62.120 ;
        RECT 2228.770 61.920 2229.090 61.980 ;
        RECT 2232.910 61.920 2233.230 61.980 ;
      LAYER via ;
        RECT 2228.800 61.920 2229.060 62.180 ;
        RECT 2232.940 61.920 2233.200 62.180 ;
      LAYER met2 ;
        RECT 2228.790 189.195 2229.070 189.565 ;
        RECT 2228.860 62.210 2229.000 189.195 ;
        RECT 2228.800 61.890 2229.060 62.210 ;
        RECT 2232.940 61.890 2233.200 62.210 ;
        RECT 2233.000 2.400 2233.140 61.890 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
      LAYER via2 ;
        RECT 2228.790 189.240 2229.070 189.520 ;
      LAYER met3 ;
        RECT 279.030 2103.050 279.410 2103.060 ;
        RECT 310.000 2103.050 314.000 2103.440 ;
        RECT 279.030 2102.840 314.000 2103.050 ;
        RECT 279.030 2102.750 310.500 2102.840 ;
        RECT 279.030 2102.740 279.410 2102.750 ;
        RECT 279.030 189.530 279.410 189.540 ;
        RECT 2228.765 189.530 2229.095 189.545 ;
        RECT 279.030 189.230 2229.095 189.530 ;
        RECT 279.030 189.220 279.410 189.230 ;
        RECT 2228.765 189.215 2229.095 189.230 ;
      LAYER via3 ;
        RECT 279.060 2102.740 279.380 2103.060 ;
        RECT 279.060 189.220 279.380 189.540 ;
      LAYER met4 ;
        RECT 279.055 2102.735 279.385 2103.065 ;
        RECT 279.070 189.545 279.370 2102.735 ;
        RECT 279.055 189.215 279.385 189.545 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 73.000 793.430 73.060 ;
        RECT 2620.690 73.000 2621.010 73.060 ;
        RECT 793.110 72.860 2621.010 73.000 ;
        RECT 793.110 72.800 793.430 72.860 ;
        RECT 2620.690 72.800 2621.010 72.860 ;
        RECT 787.590 20.640 787.910 20.700 ;
        RECT 793.110 20.640 793.430 20.700 ;
        RECT 787.590 20.500 793.430 20.640 ;
        RECT 787.590 20.440 787.910 20.500 ;
        RECT 793.110 20.440 793.430 20.500 ;
      LAYER via ;
        RECT 793.140 72.800 793.400 73.060 ;
        RECT 2620.720 72.800 2620.980 73.060 ;
        RECT 787.620 20.440 787.880 20.700 ;
        RECT 793.140 20.440 793.400 20.700 ;
      LAYER met2 ;
        RECT 2620.710 718.235 2620.990 718.605 ;
        RECT 2620.780 73.090 2620.920 718.235 ;
        RECT 793.140 72.770 793.400 73.090 ;
        RECT 2620.720 72.770 2620.980 73.090 ;
        RECT 793.200 20.730 793.340 72.770 ;
        RECT 787.620 20.410 787.880 20.730 ;
        RECT 793.140 20.410 793.400 20.730 ;
        RECT 787.680 2.400 787.820 20.410 ;
        RECT 787.470 -4.800 788.030 2.400 ;
      LAYER via2 ;
        RECT 2620.710 718.280 2620.990 718.560 ;
      LAYER met3 ;
        RECT 2606.000 718.570 2610.000 718.960 ;
        RECT 2620.685 718.570 2621.015 718.585 ;
        RECT 2606.000 718.360 2621.015 718.570 ;
        RECT 2609.580 718.270 2621.015 718.360 ;
        RECT 2620.685 718.255 2621.015 718.270 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1092.570 3258.120 1092.890 3258.180 ;
        RECT 2616.090 3258.120 2616.410 3258.180 ;
        RECT 1092.570 3257.980 2616.410 3258.120 ;
        RECT 1092.570 3257.920 1092.890 3257.980 ;
        RECT 2616.090 3257.920 2616.410 3257.980 ;
        RECT 2614.710 665.960 2615.030 666.020 ;
        RECT 2616.090 665.960 2616.410 666.020 ;
        RECT 2614.710 665.820 2616.410 665.960 ;
        RECT 2614.710 665.760 2615.030 665.820 ;
        RECT 2616.090 665.760 2616.410 665.820 ;
        RECT 2614.710 393.280 2615.030 393.340 ;
        RECT 2634.030 393.280 2634.350 393.340 ;
        RECT 2614.710 393.140 2634.350 393.280 ;
        RECT 2614.710 393.080 2615.030 393.140 ;
        RECT 2634.030 393.080 2634.350 393.140 ;
      LAYER via ;
        RECT 1092.600 3257.920 1092.860 3258.180 ;
        RECT 2616.120 3257.920 2616.380 3258.180 ;
        RECT 2614.740 665.760 2615.000 666.020 ;
        RECT 2616.120 665.760 2616.380 666.020 ;
        RECT 2614.740 393.080 2615.000 393.340 ;
        RECT 2634.060 393.080 2634.320 393.340 ;
      LAYER met2 ;
        RECT 1091.170 3258.290 1091.450 3260.000 ;
        RECT 1091.170 3258.210 1092.800 3258.290 ;
        RECT 1091.170 3258.150 1092.860 3258.210 ;
        RECT 1091.170 3256.000 1091.450 3258.150 ;
        RECT 1092.600 3257.890 1092.860 3258.150 ;
        RECT 2616.120 3257.890 2616.380 3258.210 ;
        RECT 2616.180 666.050 2616.320 3257.890 ;
        RECT 2614.740 665.730 2615.000 666.050 ;
        RECT 2616.120 665.730 2616.380 666.050 ;
        RECT 2614.800 393.370 2614.940 665.730 ;
        RECT 2614.740 393.050 2615.000 393.370 ;
        RECT 2634.060 393.050 2634.320 393.370 ;
        RECT 2634.120 270.485 2634.260 393.050 ;
        RECT 2634.050 270.115 2634.330 270.485 ;
        RECT 2250.870 33.475 2251.150 33.845 ;
        RECT 2250.940 2.400 2251.080 33.475 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
      LAYER via2 ;
        RECT 2634.050 270.160 2634.330 270.440 ;
        RECT 2250.870 33.520 2251.150 33.800 ;
      LAYER met3 ;
        RECT 2626.870 270.450 2627.250 270.460 ;
        RECT 2634.025 270.450 2634.355 270.465 ;
        RECT 2626.870 270.150 2634.355 270.450 ;
        RECT 2626.870 270.140 2627.250 270.150 ;
        RECT 2634.025 270.135 2634.355 270.150 ;
        RECT 2250.845 33.810 2251.175 33.825 ;
        RECT 2589.150 33.810 2589.530 33.820 ;
        RECT 2250.845 33.510 2589.530 33.810 ;
        RECT 2250.845 33.495 2251.175 33.510 ;
        RECT 2589.150 33.500 2589.530 33.510 ;
      LAYER via3 ;
        RECT 2626.900 270.140 2627.220 270.460 ;
        RECT 2589.180 33.500 2589.500 33.820 ;
      LAYER met4 ;
        RECT 2626.470 269.710 2627.650 270.890 ;
        RECT 2588.750 266.310 2589.930 267.490 ;
        RECT 2589.190 33.825 2589.490 266.310 ;
        RECT 2589.175 33.495 2589.505 33.825 ;
      LAYER met5 ;
        RECT 2588.540 269.500 2627.860 271.100 ;
        RECT 2588.540 266.100 2590.140 269.500 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 546.280 2619.170 546.340 ;
        RECT 2626.210 546.280 2626.530 546.340 ;
        RECT 2618.850 546.140 2626.530 546.280 ;
        RECT 2618.850 546.080 2619.170 546.140 ;
        RECT 2626.210 546.080 2626.530 546.140 ;
        RECT 2268.330 18.940 2268.650 19.000 ;
        RECT 2626.210 18.940 2626.530 19.000 ;
        RECT 2268.330 18.800 2626.530 18.940 ;
        RECT 2268.330 18.740 2268.650 18.800 ;
        RECT 2626.210 18.740 2626.530 18.800 ;
      LAYER via ;
        RECT 2618.880 546.080 2619.140 546.340 ;
        RECT 2626.240 546.080 2626.500 546.340 ;
        RECT 2268.360 18.740 2268.620 19.000 ;
        RECT 2626.240 18.740 2626.500 19.000 ;
      LAYER met2 ;
        RECT 2618.870 908.635 2619.150 909.005 ;
        RECT 2618.940 546.370 2619.080 908.635 ;
        RECT 2618.880 546.050 2619.140 546.370 ;
        RECT 2626.240 546.050 2626.500 546.370 ;
        RECT 2626.300 19.030 2626.440 546.050 ;
        RECT 2268.360 18.710 2268.620 19.030 ;
        RECT 2626.240 18.710 2626.500 19.030 ;
        RECT 2268.420 2.400 2268.560 18.710 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
      LAYER via2 ;
        RECT 2618.870 908.680 2619.150 908.960 ;
      LAYER met3 ;
        RECT 2606.000 908.970 2610.000 909.360 ;
        RECT 2618.845 908.970 2619.175 908.985 ;
        RECT 2606.000 908.760 2619.175 908.970 ;
        RECT 2609.580 908.670 2619.175 908.760 ;
        RECT 2618.845 908.655 2619.175 908.670 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.870 243.340 842.190 243.400 ;
        RECT 847.850 243.340 848.170 243.400 ;
        RECT 841.870 243.200 848.170 243.340 ;
        RECT 841.870 243.140 842.190 243.200 ;
        RECT 847.850 243.140 848.170 243.200 ;
        RECT 847.850 38.660 848.170 38.720 ;
        RECT 2286.270 38.660 2286.590 38.720 ;
        RECT 847.850 38.520 2286.590 38.660 ;
        RECT 847.850 38.460 848.170 38.520 ;
        RECT 2286.270 38.460 2286.590 38.520 ;
      LAYER via ;
        RECT 841.900 243.140 842.160 243.400 ;
        RECT 847.880 243.140 848.140 243.400 ;
        RECT 847.880 38.460 848.140 38.720 ;
        RECT 2286.300 38.460 2286.560 38.720 ;
      LAYER met2 ;
        RECT 841.850 260.000 842.130 264.000 ;
        RECT 841.960 243.430 842.100 260.000 ;
        RECT 841.900 243.110 842.160 243.430 ;
        RECT 847.880 243.110 848.140 243.430 ;
        RECT 847.940 38.750 848.080 243.110 ;
        RECT 847.880 38.430 848.140 38.750 ;
        RECT 2286.300 38.430 2286.560 38.750 ;
        RECT 2286.360 2.400 2286.500 38.430 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 287.110 1442.180 287.430 1442.240 ;
        RECT 296.770 1442.180 297.090 1442.240 ;
        RECT 287.110 1442.040 297.090 1442.180 ;
        RECT 287.110 1441.980 287.430 1442.040 ;
        RECT 296.770 1441.980 297.090 1442.040 ;
        RECT 287.110 141.340 287.430 141.400 ;
        RECT 2297.770 141.340 2298.090 141.400 ;
        RECT 287.110 141.200 2298.090 141.340 ;
        RECT 287.110 141.140 287.430 141.200 ;
        RECT 2297.770 141.140 2298.090 141.200 ;
        RECT 2297.770 37.640 2298.090 37.700 ;
        RECT 2304.210 37.640 2304.530 37.700 ;
        RECT 2297.770 37.500 2304.530 37.640 ;
        RECT 2297.770 37.440 2298.090 37.500 ;
        RECT 2304.210 37.440 2304.530 37.500 ;
      LAYER via ;
        RECT 287.140 1441.980 287.400 1442.240 ;
        RECT 296.800 1441.980 297.060 1442.240 ;
        RECT 287.140 141.140 287.400 141.400 ;
        RECT 2297.800 141.140 2298.060 141.400 ;
        RECT 2297.800 37.440 2298.060 37.700 ;
        RECT 2304.240 37.440 2304.500 37.700 ;
      LAYER met2 ;
        RECT 296.790 1447.195 297.070 1447.565 ;
        RECT 296.860 1442.270 297.000 1447.195 ;
        RECT 287.140 1441.950 287.400 1442.270 ;
        RECT 296.800 1441.950 297.060 1442.270 ;
        RECT 287.200 141.430 287.340 1441.950 ;
        RECT 287.140 141.110 287.400 141.430 ;
        RECT 2297.800 141.110 2298.060 141.430 ;
        RECT 2297.860 37.730 2298.000 141.110 ;
        RECT 2297.800 37.410 2298.060 37.730 ;
        RECT 2304.240 37.410 2304.500 37.730 ;
        RECT 2304.300 2.400 2304.440 37.410 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
      LAYER via2 ;
        RECT 296.790 1447.240 297.070 1447.520 ;
      LAYER met3 ;
        RECT 296.765 1447.530 297.095 1447.545 ;
        RECT 310.000 1447.530 314.000 1447.920 ;
        RECT 296.765 1447.320 314.000 1447.530 ;
        RECT 296.765 1447.230 310.500 1447.320 ;
        RECT 296.765 1447.215 297.095 1447.230 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.910 3271.380 2049.230 3271.440 ;
        RECT 2671.750 3271.380 2672.070 3271.440 ;
        RECT 2048.910 3271.240 2672.070 3271.380 ;
        RECT 2048.910 3271.180 2049.230 3271.240 ;
        RECT 2671.750 3271.180 2672.070 3271.240 ;
        RECT 2322.150 32.540 2322.470 32.600 ;
        RECT 2671.750 32.540 2672.070 32.600 ;
        RECT 2322.150 32.400 2672.070 32.540 ;
        RECT 2322.150 32.340 2322.470 32.400 ;
        RECT 2671.750 32.340 2672.070 32.400 ;
      LAYER via ;
        RECT 2048.940 3271.180 2049.200 3271.440 ;
        RECT 2671.780 3271.180 2672.040 3271.440 ;
        RECT 2322.180 32.340 2322.440 32.600 ;
        RECT 2671.780 32.340 2672.040 32.600 ;
      LAYER met2 ;
        RECT 2048.940 3271.150 2049.200 3271.470 ;
        RECT 2671.780 3271.150 2672.040 3271.470 ;
        RECT 2049.000 3260.000 2049.140 3271.150 ;
        RECT 2048.890 3256.000 2049.170 3260.000 ;
        RECT 2671.840 32.630 2671.980 3271.150 ;
        RECT 2322.180 32.310 2322.440 32.630 ;
        RECT 2671.780 32.310 2672.040 32.630 ;
        RECT 2322.240 2.400 2322.380 32.310 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 244.360 2345.930 244.420 ;
        RECT 2472.110 244.360 2472.430 244.420 ;
        RECT 2345.610 244.220 2472.430 244.360 ;
        RECT 2345.610 244.160 2345.930 244.220 ;
        RECT 2472.110 244.160 2472.430 244.220 ;
        RECT 2339.630 14.860 2339.950 14.920 ;
        RECT 2345.610 14.860 2345.930 14.920 ;
        RECT 2339.630 14.720 2345.930 14.860 ;
        RECT 2339.630 14.660 2339.950 14.720 ;
        RECT 2345.610 14.660 2345.930 14.720 ;
      LAYER via ;
        RECT 2345.640 244.160 2345.900 244.420 ;
        RECT 2472.140 244.160 2472.400 244.420 ;
        RECT 2339.660 14.660 2339.920 14.920 ;
        RECT 2345.640 14.660 2345.900 14.920 ;
      LAYER met2 ;
        RECT 2472.090 260.000 2472.370 264.000 ;
        RECT 2472.200 244.450 2472.340 260.000 ;
        RECT 2345.640 244.130 2345.900 244.450 ;
        RECT 2472.140 244.130 2472.400 244.450 ;
        RECT 2345.700 14.950 2345.840 244.130 ;
        RECT 2339.660 14.630 2339.920 14.950 ;
        RECT 2345.640 14.630 2345.900 14.950 ;
        RECT 2339.720 2.400 2339.860 14.630 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1720.470 3272.740 1720.790 3272.800 ;
        RECT 2650.130 3272.740 2650.450 3272.800 ;
        RECT 1720.470 3272.600 2650.450 3272.740 ;
        RECT 1720.470 3272.540 1720.790 3272.600 ;
        RECT 2650.130 3272.540 2650.450 3272.600 ;
        RECT 2650.130 16.560 2650.450 16.620 ;
        RECT 2404.580 16.420 2650.450 16.560 ;
        RECT 2357.570 16.220 2357.890 16.280 ;
        RECT 2404.580 16.220 2404.720 16.420 ;
        RECT 2650.130 16.360 2650.450 16.420 ;
        RECT 2357.570 16.080 2404.720 16.220 ;
        RECT 2357.570 16.020 2357.890 16.080 ;
      LAYER via ;
        RECT 1720.500 3272.540 1720.760 3272.800 ;
        RECT 2650.160 3272.540 2650.420 3272.800 ;
        RECT 2357.600 16.020 2357.860 16.280 ;
        RECT 2650.160 16.360 2650.420 16.620 ;
      LAYER met2 ;
        RECT 1720.500 3272.510 1720.760 3272.830 ;
        RECT 2650.160 3272.510 2650.420 3272.830 ;
        RECT 1720.560 3260.000 1720.700 3272.510 ;
        RECT 1720.450 3256.000 1720.730 3260.000 ;
        RECT 2650.220 16.650 2650.360 3272.510 ;
        RECT 2650.160 16.330 2650.420 16.650 ;
        RECT 2357.600 15.990 2357.860 16.310 ;
        RECT 2357.660 2.400 2357.800 15.990 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2380.110 244.700 2380.430 244.760 ;
        RECT 2414.150 244.700 2414.470 244.760 ;
        RECT 2380.110 244.560 2414.470 244.700 ;
        RECT 2380.110 244.500 2380.430 244.560 ;
        RECT 2414.150 244.500 2414.470 244.560 ;
        RECT 2375.510 16.560 2375.830 16.620 ;
        RECT 2380.110 16.560 2380.430 16.620 ;
        RECT 2375.510 16.420 2380.430 16.560 ;
        RECT 2375.510 16.360 2375.830 16.420 ;
        RECT 2380.110 16.360 2380.430 16.420 ;
      LAYER via ;
        RECT 2380.140 244.500 2380.400 244.760 ;
        RECT 2414.180 244.500 2414.440 244.760 ;
        RECT 2375.540 16.360 2375.800 16.620 ;
        RECT 2380.140 16.360 2380.400 16.620 ;
      LAYER met2 ;
        RECT 2414.130 260.000 2414.410 264.000 ;
        RECT 2414.240 244.790 2414.380 260.000 ;
        RECT 2380.140 244.470 2380.400 244.790 ;
        RECT 2414.180 244.470 2414.440 244.790 ;
        RECT 2380.200 16.650 2380.340 244.470 ;
        RECT 2375.540 16.330 2375.800 16.650 ;
        RECT 2380.140 16.330 2380.400 16.650 ;
        RECT 2375.600 2.400 2375.740 16.330 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 607.480 2615.490 607.540 ;
        RECT 2667.610 607.480 2667.930 607.540 ;
        RECT 2615.170 607.340 2667.930 607.480 ;
        RECT 2615.170 607.280 2615.490 607.340 ;
        RECT 2667.610 607.280 2667.930 607.340 ;
        RECT 2393.450 247.080 2393.770 247.140 ;
        RECT 2667.610 247.080 2667.930 247.140 ;
        RECT 2393.450 246.940 2667.930 247.080 ;
        RECT 2393.450 246.880 2393.770 246.940 ;
        RECT 2667.610 246.880 2667.930 246.940 ;
      LAYER via ;
        RECT 2615.200 607.280 2615.460 607.540 ;
        RECT 2667.640 607.280 2667.900 607.540 ;
        RECT 2393.480 246.880 2393.740 247.140 ;
        RECT 2667.640 246.880 2667.900 247.140 ;
      LAYER met2 ;
        RECT 2615.190 613.515 2615.470 613.885 ;
        RECT 2615.260 607.570 2615.400 613.515 ;
        RECT 2615.200 607.250 2615.460 607.570 ;
        RECT 2667.640 607.250 2667.900 607.570 ;
        RECT 2667.700 247.170 2667.840 607.250 ;
        RECT 2393.480 246.850 2393.740 247.170 ;
        RECT 2667.640 246.850 2667.900 247.170 ;
        RECT 2393.540 2.400 2393.680 246.850 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
      LAYER via2 ;
        RECT 2615.190 613.560 2615.470 613.840 ;
      LAYER met3 ;
        RECT 2606.000 613.850 2610.000 614.240 ;
        RECT 2615.165 613.850 2615.495 613.865 ;
        RECT 2606.000 613.640 2615.495 613.850 ;
        RECT 2609.580 613.550 2615.495 613.640 ;
        RECT 2615.165 613.535 2615.495 613.550 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 273.770 1952.860 274.090 1952.920 ;
        RECT 296.770 1952.860 297.090 1952.920 ;
        RECT 273.770 1952.720 297.090 1952.860 ;
        RECT 273.770 1952.660 274.090 1952.720 ;
        RECT 296.770 1952.660 297.090 1952.720 ;
        RECT 273.770 99.860 274.090 99.920 ;
        RECT 2408.170 99.860 2408.490 99.920 ;
        RECT 273.770 99.720 2408.490 99.860 ;
        RECT 273.770 99.660 274.090 99.720 ;
        RECT 2408.170 99.660 2408.490 99.720 ;
        RECT 2408.170 62.120 2408.490 62.180 ;
        RECT 2411.390 62.120 2411.710 62.180 ;
        RECT 2408.170 61.980 2411.710 62.120 ;
        RECT 2408.170 61.920 2408.490 61.980 ;
        RECT 2411.390 61.920 2411.710 61.980 ;
      LAYER via ;
        RECT 273.800 1952.660 274.060 1952.920 ;
        RECT 296.800 1952.660 297.060 1952.920 ;
        RECT 273.800 99.660 274.060 99.920 ;
        RECT 2408.200 99.660 2408.460 99.920 ;
        RECT 2408.200 61.920 2408.460 62.180 ;
        RECT 2411.420 61.920 2411.680 62.180 ;
      LAYER met2 ;
        RECT 296.790 1954.475 297.070 1954.845 ;
        RECT 296.860 1952.950 297.000 1954.475 ;
        RECT 273.800 1952.630 274.060 1952.950 ;
        RECT 296.800 1952.630 297.060 1952.950 ;
        RECT 273.860 99.950 274.000 1952.630 ;
        RECT 273.800 99.630 274.060 99.950 ;
        RECT 2408.200 99.630 2408.460 99.950 ;
        RECT 2408.260 62.210 2408.400 99.630 ;
        RECT 2408.200 61.890 2408.460 62.210 ;
        RECT 2411.420 61.890 2411.680 62.210 ;
        RECT 2411.480 2.400 2411.620 61.890 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 296.790 1954.520 297.070 1954.800 ;
      LAYER met3 ;
        RECT 296.765 1954.810 297.095 1954.825 ;
        RECT 310.000 1954.810 314.000 1955.200 ;
        RECT 296.765 1954.600 314.000 1954.810 ;
        RECT 296.765 1954.510 310.500 1954.600 ;
        RECT 296.765 1954.495 297.095 1954.510 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1897.645 246.585 1897.815 247.775 ;
        RECT 1945.485 246.585 1945.655 248.115 ;
      LAYER mcon ;
        RECT 1945.485 247.945 1945.655 248.115 ;
        RECT 1897.645 247.605 1897.815 247.775 ;
      LAYER met1 ;
        RECT 1945.425 248.100 1945.715 248.145 ;
        RECT 2013.950 248.100 2014.270 248.160 ;
        RECT 1801.060 247.960 1849.500 248.100 ;
        RECT 1797.290 247.760 1797.610 247.820 ;
        RECT 1801.060 247.760 1801.200 247.960 ;
        RECT 1797.290 247.620 1801.200 247.760 ;
        RECT 1849.360 247.760 1849.500 247.960 ;
        RECT 1945.425 247.960 2014.270 248.100 ;
        RECT 1945.425 247.915 1945.715 247.960 ;
        RECT 2013.950 247.900 2014.270 247.960 ;
        RECT 1897.585 247.760 1897.875 247.805 ;
        RECT 1849.360 247.620 1897.875 247.760 ;
        RECT 1797.290 247.560 1797.610 247.620 ;
        RECT 1897.585 247.575 1897.875 247.620 ;
        RECT 1897.585 246.740 1897.875 246.785 ;
        RECT 1945.425 246.740 1945.715 246.785 ;
        RECT 1897.585 246.600 1945.715 246.740 ;
        RECT 1897.585 246.555 1897.875 246.600 ;
        RECT 1945.425 246.555 1945.715 246.600 ;
        RECT 806.910 155.620 807.230 155.680 ;
        RECT 1797.290 155.620 1797.610 155.680 ;
        RECT 806.910 155.480 1797.610 155.620 ;
        RECT 806.910 155.420 807.230 155.480 ;
        RECT 1797.290 155.420 1797.610 155.480 ;
        RECT 805.530 14.180 805.850 14.240 ;
        RECT 806.910 14.180 807.230 14.240 ;
        RECT 805.530 14.040 807.230 14.180 ;
        RECT 805.530 13.980 805.850 14.040 ;
        RECT 806.910 13.980 807.230 14.040 ;
      LAYER via ;
        RECT 1797.320 247.560 1797.580 247.820 ;
        RECT 2013.980 247.900 2014.240 248.160 ;
        RECT 806.940 155.420 807.200 155.680 ;
        RECT 1797.320 155.420 1797.580 155.680 ;
        RECT 805.560 13.980 805.820 14.240 ;
        RECT 806.940 13.980 807.200 14.240 ;
      LAYER met2 ;
        RECT 2013.930 260.000 2014.210 264.000 ;
        RECT 2014.040 248.190 2014.180 260.000 ;
        RECT 2013.980 247.870 2014.240 248.190 ;
        RECT 1797.320 247.530 1797.580 247.850 ;
        RECT 1797.380 155.710 1797.520 247.530 ;
        RECT 806.940 155.390 807.200 155.710 ;
        RECT 1797.320 155.390 1797.580 155.710 ;
        RECT 807.000 14.270 807.140 155.390 ;
        RECT 805.560 13.950 805.820 14.270 ;
        RECT 806.940 13.950 807.200 14.270 ;
        RECT 805.620 2.400 805.760 13.950 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 10.190 51.580 10.510 51.640 ;
        RECT 1242.070 51.580 1242.390 51.640 ;
        RECT 10.190 51.440 1242.390 51.580 ;
        RECT 10.190 51.380 10.510 51.440 ;
        RECT 1242.070 51.380 1242.390 51.440 ;
        RECT 2.830 16.900 3.150 16.960 ;
        RECT 10.190 16.900 10.510 16.960 ;
        RECT 2.830 16.760 10.510 16.900 ;
        RECT 2.830 16.700 3.150 16.760 ;
        RECT 10.190 16.700 10.510 16.760 ;
      LAYER via ;
        RECT 10.220 51.380 10.480 51.640 ;
        RECT 1242.100 51.380 1242.360 51.640 ;
        RECT 2.860 16.700 3.120 16.960 ;
        RECT 10.220 16.700 10.480 16.960 ;
      LAYER met2 ;
        RECT 1242.050 260.000 1242.330 264.000 ;
        RECT 1242.160 51.670 1242.300 260.000 ;
        RECT 10.220 51.350 10.480 51.670 ;
        RECT 1242.100 51.350 1242.360 51.670 ;
        RECT 10.280 16.990 10.420 51.350 ;
        RECT 2.860 16.670 3.120 16.990 ;
        RECT 10.220 16.670 10.480 16.990 ;
        RECT 2.920 2.400 3.060 16.670 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 99.890 2884.460 100.210 2884.520 ;
        RECT 296.770 2884.460 297.090 2884.520 ;
        RECT 99.890 2884.320 297.090 2884.460 ;
        RECT 99.890 2884.260 100.210 2884.320 ;
        RECT 296.770 2884.260 297.090 2884.320 ;
        RECT 8.350 18.600 8.670 18.660 ;
        RECT 99.890 18.600 100.210 18.660 ;
        RECT 8.350 18.460 100.210 18.600 ;
        RECT 8.350 18.400 8.670 18.460 ;
        RECT 99.890 18.400 100.210 18.460 ;
      LAYER via ;
        RECT 99.920 2884.260 100.180 2884.520 ;
        RECT 296.800 2884.260 297.060 2884.520 ;
        RECT 8.380 18.400 8.640 18.660 ;
        RECT 99.920 18.400 100.180 18.660 ;
      LAYER met2 ;
        RECT 296.790 2884.715 297.070 2885.085 ;
        RECT 296.860 2884.550 297.000 2884.715 ;
        RECT 99.920 2884.230 100.180 2884.550 ;
        RECT 296.800 2884.230 297.060 2884.550 ;
        RECT 99.980 18.690 100.120 2884.230 ;
        RECT 8.380 18.370 8.640 18.690 ;
        RECT 99.920 18.370 100.180 18.690 ;
        RECT 8.440 2.400 8.580 18.370 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 296.790 2884.760 297.070 2885.040 ;
      LAYER met3 ;
        RECT 296.765 2885.050 297.095 2885.065 ;
        RECT 310.000 2885.050 314.000 2885.440 ;
        RECT 296.765 2884.840 314.000 2885.050 ;
        RECT 296.765 2884.750 310.500 2884.840 ;
        RECT 296.765 2884.735 297.095 2884.750 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.290 3258.460 72.610 3258.520 ;
        RECT 1104.070 3258.460 1104.390 3258.520 ;
        RECT 72.290 3258.320 1104.390 3258.460 ;
        RECT 72.290 3258.260 72.610 3258.320 ;
        RECT 1104.070 3258.260 1104.390 3258.320 ;
        RECT 14.330 18.940 14.650 19.000 ;
        RECT 72.290 18.940 72.610 19.000 ;
        RECT 14.330 18.800 72.610 18.940 ;
        RECT 14.330 18.740 14.650 18.800 ;
        RECT 72.290 18.740 72.610 18.800 ;
      LAYER via ;
        RECT 72.320 3258.260 72.580 3258.520 ;
        RECT 1104.100 3258.260 1104.360 3258.520 ;
        RECT 14.360 18.740 14.620 19.000 ;
        RECT 72.320 18.740 72.580 19.000 ;
      LAYER met2 ;
        RECT 72.320 3258.230 72.580 3258.550 ;
        RECT 1104.100 3258.290 1104.360 3258.550 ;
        RECT 1104.970 3258.290 1105.250 3260.000 ;
        RECT 1104.100 3258.230 1105.250 3258.290 ;
        RECT 72.380 19.030 72.520 3258.230 ;
        RECT 1104.160 3258.150 1105.250 3258.230 ;
        RECT 1104.970 3256.000 1105.250 3258.150 ;
        RECT 14.360 18.710 14.620 19.030 ;
        RECT 72.320 18.710 72.580 19.030 ;
        RECT 14.420 2.400 14.560 18.710 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.750 1552.680 142.070 1552.740 ;
        RECT 296.770 1552.680 297.090 1552.740 ;
        RECT 141.750 1552.540 297.090 1552.680 ;
        RECT 141.750 1552.480 142.070 1552.540 ;
        RECT 296.770 1552.480 297.090 1552.540 ;
        RECT 141.750 17.920 142.070 17.980 ;
        RECT 136.320 17.780 142.070 17.920 ;
        RECT 38.250 17.580 38.570 17.640 ;
        RECT 136.320 17.580 136.460 17.780 ;
        RECT 141.750 17.720 142.070 17.780 ;
        RECT 38.250 17.440 136.460 17.580 ;
        RECT 38.250 17.380 38.570 17.440 ;
      LAYER via ;
        RECT 141.780 1552.480 142.040 1552.740 ;
        RECT 296.800 1552.480 297.060 1552.740 ;
        RECT 38.280 17.380 38.540 17.640 ;
        RECT 141.780 17.720 142.040 17.980 ;
      LAYER met2 ;
        RECT 296.790 1553.275 297.070 1553.645 ;
        RECT 296.860 1552.770 297.000 1553.275 ;
        RECT 141.780 1552.450 142.040 1552.770 ;
        RECT 296.800 1552.450 297.060 1552.770 ;
        RECT 141.840 18.010 141.980 1552.450 ;
        RECT 141.780 17.690 142.040 18.010 ;
        RECT 38.280 17.350 38.540 17.670 ;
        RECT 38.340 2.400 38.480 17.350 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 296.790 1553.320 297.070 1553.600 ;
      LAYER met3 ;
        RECT 296.765 1553.610 297.095 1553.625 ;
        RECT 310.000 1553.610 314.000 1554.000 ;
        RECT 296.765 1553.400 314.000 1553.610 ;
        RECT 296.765 1553.310 310.500 1553.400 ;
        RECT 296.765 1553.295 297.095 1553.310 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.750 175.595 240.030 175.965 ;
        RECT 239.820 3.130 239.960 175.595 ;
        RECT 239.820 2.990 240.880 3.130 ;
        RECT 240.740 2.400 240.880 2.990 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 239.750 175.640 240.030 175.920 ;
      LAYER met3 ;
        RECT 2606.000 2917.690 2610.000 2918.080 ;
        RECT 2636.990 2917.690 2637.370 2917.700 ;
        RECT 2606.000 2917.480 2637.370 2917.690 ;
        RECT 2609.580 2917.390 2637.370 2917.480 ;
        RECT 2636.990 2917.380 2637.370 2917.390 ;
        RECT 239.725 175.930 240.055 175.945 ;
        RECT 2636.990 175.930 2637.370 175.940 ;
        RECT 239.725 175.630 2637.370 175.930 ;
        RECT 239.725 175.615 240.055 175.630 ;
        RECT 2636.990 175.620 2637.370 175.630 ;
      LAYER via3 ;
        RECT 2637.020 2917.380 2637.340 2917.700 ;
        RECT 2637.020 175.620 2637.340 175.940 ;
      LAYER met4 ;
        RECT 2637.015 2917.375 2637.345 2917.705 ;
        RECT 2637.030 175.945 2637.330 2917.375 ;
        RECT 2637.015 175.615 2637.345 175.945 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1107.290 246.740 1107.610 246.800 ;
        RECT 1756.350 246.740 1756.670 246.800 ;
        RECT 1107.290 246.600 1756.670 246.740 ;
        RECT 1107.290 246.540 1107.610 246.600 ;
        RECT 1756.350 246.540 1756.670 246.600 ;
        RECT 258.130 34.240 258.450 34.300 ;
        RECT 1107.290 34.240 1107.610 34.300 ;
        RECT 258.130 34.100 1107.610 34.240 ;
        RECT 258.130 34.040 258.450 34.100 ;
        RECT 1107.290 34.040 1107.610 34.100 ;
      LAYER via ;
        RECT 1107.320 246.540 1107.580 246.800 ;
        RECT 1756.380 246.540 1756.640 246.800 ;
        RECT 258.160 34.040 258.420 34.300 ;
        RECT 1107.320 34.040 1107.580 34.300 ;
      LAYER met2 ;
        RECT 1756.330 260.000 1756.610 264.000 ;
        RECT 1756.440 246.830 1756.580 260.000 ;
        RECT 1107.320 246.510 1107.580 246.830 ;
        RECT 1756.380 246.510 1756.640 246.830 ;
        RECT 1107.380 34.330 1107.520 246.510 ;
        RECT 258.160 34.010 258.420 34.330 ;
        RECT 1107.320 34.010 1107.580 34.330 ;
        RECT 258.220 2.400 258.360 34.010 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 87.280 282.830 87.340 ;
        RECT 883.270 87.280 883.590 87.340 ;
        RECT 282.510 87.140 883.590 87.280 ;
        RECT 282.510 87.080 282.830 87.140 ;
        RECT 883.270 87.080 883.590 87.140 ;
        RECT 276.070 20.640 276.390 20.700 ;
        RECT 282.510 20.640 282.830 20.700 ;
        RECT 276.070 20.500 282.830 20.640 ;
        RECT 276.070 20.440 276.390 20.500 ;
        RECT 282.510 20.440 282.830 20.500 ;
      LAYER via ;
        RECT 282.540 87.080 282.800 87.340 ;
        RECT 883.300 87.080 883.560 87.340 ;
        RECT 276.100 20.440 276.360 20.700 ;
        RECT 282.540 20.440 282.800 20.700 ;
      LAYER met2 ;
        RECT 884.170 260.170 884.450 264.000 ;
        RECT 883.360 260.030 884.450 260.170 ;
        RECT 883.360 87.370 883.500 260.030 ;
        RECT 884.170 260.000 884.450 260.030 ;
        RECT 282.540 87.050 282.800 87.370 ;
        RECT 883.300 87.050 883.560 87.370 ;
        RECT 282.600 20.730 282.740 87.050 ;
        RECT 276.100 20.410 276.360 20.730 ;
        RECT 282.540 20.410 282.800 20.730 ;
        RECT 276.160 2.400 276.300 20.410 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1852.490 241.640 1852.810 241.700 ;
        RECT 1856.630 241.640 1856.950 241.700 ;
        RECT 1852.490 241.500 1856.950 241.640 ;
        RECT 1852.490 241.440 1852.810 241.500 ;
        RECT 1856.630 241.440 1856.950 241.500 ;
        RECT 296.310 93.740 296.630 93.800 ;
        RECT 1852.490 93.740 1852.810 93.800 ;
        RECT 296.310 93.600 1852.810 93.740 ;
        RECT 296.310 93.540 296.630 93.600 ;
        RECT 1852.490 93.540 1852.810 93.600 ;
        RECT 294.010 20.640 294.330 20.700 ;
        RECT 296.310 20.640 296.630 20.700 ;
        RECT 294.010 20.500 296.630 20.640 ;
        RECT 294.010 20.440 294.330 20.500 ;
        RECT 296.310 20.440 296.630 20.500 ;
      LAYER via ;
        RECT 1852.520 241.440 1852.780 241.700 ;
        RECT 1856.660 241.440 1856.920 241.700 ;
        RECT 296.340 93.540 296.600 93.800 ;
        RECT 1852.520 93.540 1852.780 93.800 ;
        RECT 294.040 20.440 294.300 20.700 ;
        RECT 296.340 20.440 296.600 20.700 ;
      LAYER met2 ;
        RECT 1856.610 260.000 1856.890 264.000 ;
        RECT 1856.720 241.730 1856.860 260.000 ;
        RECT 1852.520 241.410 1852.780 241.730 ;
        RECT 1856.660 241.410 1856.920 241.730 ;
        RECT 1852.580 93.830 1852.720 241.410 ;
        RECT 296.340 93.510 296.600 93.830 ;
        RECT 1852.520 93.510 1852.780 93.830 ;
        RECT 296.400 20.730 296.540 93.510 ;
        RECT 294.040 20.410 294.300 20.730 ;
        RECT 296.340 20.410 296.600 20.730 ;
        RECT 294.100 2.400 294.240 20.410 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 226.390 3271.040 226.710 3271.100 ;
        RECT 347.830 3271.040 348.150 3271.100 ;
        RECT 226.390 3270.900 348.150 3271.040 ;
        RECT 226.390 3270.840 226.710 3270.900 ;
        RECT 347.830 3270.840 348.150 3270.900 ;
        RECT 226.390 238.920 226.710 238.980 ;
        RECT 310.570 238.920 310.890 238.980 ;
        RECT 226.390 238.780 310.890 238.920 ;
        RECT 226.390 238.720 226.710 238.780 ;
        RECT 310.570 238.720 310.890 238.780 ;
        RECT 310.570 2.960 310.890 3.020 ;
        RECT 311.950 2.960 312.270 3.020 ;
        RECT 310.570 2.820 312.270 2.960 ;
        RECT 310.570 2.760 310.890 2.820 ;
        RECT 311.950 2.760 312.270 2.820 ;
      LAYER via ;
        RECT 226.420 3270.840 226.680 3271.100 ;
        RECT 347.860 3270.840 348.120 3271.100 ;
        RECT 226.420 238.720 226.680 238.980 ;
        RECT 310.600 238.720 310.860 238.980 ;
        RECT 310.600 2.760 310.860 3.020 ;
        RECT 311.980 2.760 312.240 3.020 ;
      LAYER met2 ;
        RECT 226.420 3270.810 226.680 3271.130 ;
        RECT 347.860 3270.810 348.120 3271.130 ;
        RECT 226.480 239.010 226.620 3270.810 ;
        RECT 347.920 3260.000 348.060 3270.810 ;
        RECT 347.810 3256.000 348.090 3260.000 ;
        RECT 226.420 238.690 226.680 239.010 ;
        RECT 310.600 238.690 310.860 239.010 ;
        RECT 310.660 3.050 310.800 238.690 ;
        RECT 310.600 2.730 310.860 3.050 ;
        RECT 311.980 2.730 312.240 3.050 ;
        RECT 312.040 2.400 312.180 2.730 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 233.290 2987.820 233.610 2987.880 ;
        RECT 296.770 2987.820 297.090 2987.880 ;
        RECT 233.290 2987.680 297.090 2987.820 ;
        RECT 233.290 2987.620 233.610 2987.680 ;
        RECT 296.770 2987.620 297.090 2987.680 ;
        RECT 233.290 18.600 233.610 18.660 ;
        RECT 329.890 18.600 330.210 18.660 ;
        RECT 233.290 18.460 330.210 18.600 ;
        RECT 233.290 18.400 233.610 18.460 ;
        RECT 329.890 18.400 330.210 18.460 ;
      LAYER via ;
        RECT 233.320 2987.620 233.580 2987.880 ;
        RECT 296.800 2987.620 297.060 2987.880 ;
        RECT 233.320 18.400 233.580 18.660 ;
        RECT 329.920 18.400 330.180 18.660 ;
      LAYER met2 ;
        RECT 296.790 2990.795 297.070 2991.165 ;
        RECT 296.860 2987.910 297.000 2990.795 ;
        RECT 233.320 2987.590 233.580 2987.910 ;
        RECT 296.800 2987.590 297.060 2987.910 ;
        RECT 233.380 18.690 233.520 2987.590 ;
        RECT 233.320 18.370 233.580 18.690 ;
        RECT 329.920 18.370 330.180 18.690 ;
        RECT 329.980 2.400 330.120 18.370 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 296.790 2990.840 297.070 2991.120 ;
      LAYER met3 ;
        RECT 296.765 2991.130 297.095 2991.145 ;
        RECT 310.000 2991.130 314.000 2991.520 ;
        RECT 296.765 2990.920 314.000 2991.130 ;
        RECT 296.765 2990.830 310.500 2990.920 ;
        RECT 296.765 2990.815 297.095 2990.830 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.170 3266.280 246.490 3266.340 ;
        RECT 1419.630 3266.280 1419.950 3266.340 ;
        RECT 246.170 3266.140 1419.950 3266.280 ;
        RECT 246.170 3266.080 246.490 3266.140 ;
        RECT 1419.630 3266.080 1419.950 3266.140 ;
        RECT 246.170 261.360 246.490 261.420 ;
        RECT 345.070 261.360 345.390 261.420 ;
        RECT 246.170 261.220 345.390 261.360 ;
        RECT 246.170 261.160 246.490 261.220 ;
        RECT 345.070 261.160 345.390 261.220 ;
        RECT 345.070 18.600 345.390 18.660 ;
        RECT 347.370 18.600 347.690 18.660 ;
        RECT 345.070 18.460 347.690 18.600 ;
        RECT 345.070 18.400 345.390 18.460 ;
        RECT 347.370 18.400 347.690 18.460 ;
      LAYER via ;
        RECT 246.200 3266.080 246.460 3266.340 ;
        RECT 1419.660 3266.080 1419.920 3266.340 ;
        RECT 246.200 261.160 246.460 261.420 ;
        RECT 345.100 261.160 345.360 261.420 ;
        RECT 345.100 18.400 345.360 18.660 ;
        RECT 347.400 18.400 347.660 18.660 ;
      LAYER met2 ;
        RECT 246.200 3266.050 246.460 3266.370 ;
        RECT 1419.660 3266.050 1419.920 3266.370 ;
        RECT 246.260 261.450 246.400 3266.050 ;
        RECT 1419.720 3260.000 1419.860 3266.050 ;
        RECT 1419.610 3256.000 1419.890 3260.000 ;
        RECT 246.200 261.130 246.460 261.450 ;
        RECT 345.100 261.130 345.360 261.450 ;
        RECT 345.160 18.690 345.300 261.130 ;
        RECT 345.100 18.370 345.360 18.690 ;
        RECT 347.400 18.370 347.660 18.690 ;
        RECT 347.460 2.400 347.600 18.370 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 274.690 3174.140 275.010 3174.200 ;
        RECT 296.770 3174.140 297.090 3174.200 ;
        RECT 274.690 3174.000 297.090 3174.140 ;
        RECT 274.690 3173.940 275.010 3174.000 ;
        RECT 296.770 3173.940 297.090 3174.000 ;
        RECT 274.690 38.320 275.010 38.380 ;
        RECT 365.310 38.320 365.630 38.380 ;
        RECT 274.690 38.180 365.630 38.320 ;
        RECT 274.690 38.120 275.010 38.180 ;
        RECT 365.310 38.120 365.630 38.180 ;
      LAYER via ;
        RECT 274.720 3173.940 274.980 3174.200 ;
        RECT 296.800 3173.940 297.060 3174.200 ;
        RECT 274.720 38.120 274.980 38.380 ;
        RECT 365.340 38.120 365.600 38.380 ;
      LAYER met2 ;
        RECT 296.790 3179.835 297.070 3180.205 ;
        RECT 296.860 3174.230 297.000 3179.835 ;
        RECT 274.720 3173.910 274.980 3174.230 ;
        RECT 296.800 3173.910 297.060 3174.230 ;
        RECT 274.780 38.410 274.920 3173.910 ;
        RECT 274.720 38.090 274.980 38.410 ;
        RECT 365.340 38.090 365.600 38.410 ;
        RECT 365.400 2.400 365.540 38.090 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 296.790 3179.880 297.070 3180.160 ;
      LAYER met3 ;
        RECT 296.765 3180.170 297.095 3180.185 ;
        RECT 310.000 3180.170 314.000 3180.560 ;
        RECT 296.765 3179.960 314.000 3180.170 ;
        RECT 296.765 3179.870 310.500 3179.960 ;
        RECT 296.765 3179.855 297.095 3179.870 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 233.750 255.920 234.070 255.980 ;
        RECT 380.030 255.920 380.350 255.980 ;
        RECT 233.750 255.780 380.350 255.920 ;
        RECT 233.750 255.720 234.070 255.780 ;
        RECT 380.030 255.720 380.350 255.780 ;
        RECT 380.030 19.620 380.350 19.680 ;
        RECT 383.250 19.620 383.570 19.680 ;
        RECT 380.030 19.480 383.570 19.620 ;
        RECT 380.030 19.420 380.350 19.480 ;
        RECT 383.250 19.420 383.570 19.480 ;
      LAYER via ;
        RECT 233.780 255.720 234.040 255.980 ;
        RECT 380.060 255.720 380.320 255.980 ;
        RECT 380.060 19.420 380.320 19.680 ;
        RECT 383.280 19.420 383.540 19.680 ;
      LAYER met2 ;
        RECT 2335.050 3264.155 2335.330 3264.525 ;
        RECT 2335.120 3260.000 2335.260 3264.155 ;
        RECT 2335.010 3256.000 2335.290 3260.000 ;
        RECT 233.770 261.955 234.050 262.325 ;
        RECT 233.840 256.010 233.980 261.955 ;
        RECT 233.780 255.690 234.040 256.010 ;
        RECT 380.060 255.690 380.320 256.010 ;
        RECT 380.120 19.710 380.260 255.690 ;
        RECT 380.060 19.390 380.320 19.710 ;
        RECT 383.280 19.390 383.540 19.710 ;
        RECT 383.340 2.400 383.480 19.390 ;
        RECT 383.130 -4.800 383.690 2.400 ;
      LAYER via2 ;
        RECT 2335.050 3264.200 2335.330 3264.480 ;
        RECT 233.770 262.000 234.050 262.280 ;
      LAYER met3 ;
        RECT 233.950 3264.490 234.330 3264.500 ;
        RECT 2335.025 3264.490 2335.355 3264.505 ;
        RECT 233.950 3264.190 2335.355 3264.490 ;
        RECT 233.950 3264.180 234.330 3264.190 ;
        RECT 2335.025 3264.175 2335.355 3264.190 ;
        RECT 233.745 262.300 234.075 262.305 ;
        RECT 233.745 262.290 234.330 262.300 ;
        RECT 233.745 261.990 234.530 262.290 ;
        RECT 233.745 261.980 234.330 261.990 ;
        RECT 233.745 261.975 234.075 261.980 ;
      LAYER via3 ;
        RECT 233.980 3264.180 234.300 3264.500 ;
        RECT 233.980 261.980 234.300 262.300 ;
      LAYER met4 ;
        RECT 233.975 3264.175 234.305 3264.505 ;
        RECT 233.990 262.305 234.290 3264.175 ;
        RECT 233.975 261.975 234.305 262.305 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 400.345 48.365 400.515 137.955 ;
      LAYER mcon ;
        RECT 400.345 137.785 400.515 137.955 ;
      LAYER met1 ;
        RECT 238.810 3264.920 239.130 3264.980 ;
        RECT 1777.510 3264.920 1777.830 3264.980 ;
        RECT 238.810 3264.780 1777.830 3264.920 ;
        RECT 238.810 3264.720 239.130 3264.780 ;
        RECT 1777.510 3264.720 1777.830 3264.780 ;
        RECT 238.810 260.340 239.130 260.400 ;
        RECT 400.270 260.340 400.590 260.400 ;
        RECT 238.810 260.200 400.590 260.340 ;
        RECT 238.810 260.140 239.130 260.200 ;
        RECT 400.270 260.140 400.590 260.200 ;
        RECT 400.270 193.020 400.590 193.080 ;
        RECT 400.730 193.020 401.050 193.080 ;
        RECT 400.270 192.880 401.050 193.020 ;
        RECT 400.270 192.820 400.590 192.880 ;
        RECT 400.730 192.820 401.050 192.880 ;
        RECT 400.270 137.940 400.590 138.000 ;
        RECT 400.075 137.800 400.590 137.940 ;
        RECT 400.270 137.740 400.590 137.800 ;
        RECT 400.285 48.520 400.575 48.565 ;
        RECT 401.190 48.520 401.510 48.580 ;
        RECT 400.285 48.380 401.510 48.520 ;
        RECT 400.285 48.335 400.575 48.380 ;
        RECT 401.190 48.320 401.510 48.380 ;
      LAYER via ;
        RECT 238.840 3264.720 239.100 3264.980 ;
        RECT 1777.540 3264.720 1777.800 3264.980 ;
        RECT 238.840 260.140 239.100 260.400 ;
        RECT 400.300 260.140 400.560 260.400 ;
        RECT 400.300 192.820 400.560 193.080 ;
        RECT 400.760 192.820 401.020 193.080 ;
        RECT 400.300 137.740 400.560 138.000 ;
        RECT 401.220 48.320 401.480 48.580 ;
      LAYER met2 ;
        RECT 238.840 3264.690 239.100 3265.010 ;
        RECT 1777.540 3264.690 1777.800 3265.010 ;
        RECT 238.900 260.430 239.040 3264.690 ;
        RECT 1777.600 3260.000 1777.740 3264.690 ;
        RECT 1777.490 3256.000 1777.770 3260.000 ;
        RECT 238.840 260.110 239.100 260.430 ;
        RECT 400.300 260.110 400.560 260.430 ;
        RECT 400.360 193.110 400.500 260.110 ;
        RECT 400.300 192.790 400.560 193.110 ;
        RECT 400.760 192.790 401.020 193.110 ;
        RECT 400.820 145.250 400.960 192.790 ;
        RECT 400.360 145.110 400.960 145.250 ;
        RECT 400.360 138.030 400.500 145.110 ;
        RECT 400.300 137.710 400.560 138.030 ;
        RECT 401.220 48.290 401.480 48.610 ;
        RECT 401.280 2.400 401.420 48.290 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2617.930 1243.620 2618.250 1243.680 ;
        RECT 2639.550 1243.620 2639.870 1243.680 ;
        RECT 2617.930 1243.480 2639.870 1243.620 ;
        RECT 2617.930 1243.420 2618.250 1243.480 ;
        RECT 2639.550 1243.420 2639.870 1243.480 ;
        RECT 62.170 37.980 62.490 38.040 ;
        RECT 2639.550 37.980 2639.870 38.040 ;
        RECT 62.170 37.840 2639.870 37.980 ;
        RECT 62.170 37.780 62.490 37.840 ;
        RECT 2639.550 37.780 2639.870 37.840 ;
      LAYER via ;
        RECT 2617.960 1243.420 2618.220 1243.680 ;
        RECT 2639.580 1243.420 2639.840 1243.680 ;
        RECT 62.200 37.780 62.460 38.040 ;
        RECT 2639.580 37.780 2639.840 38.040 ;
      LAYER met2 ;
        RECT 2617.950 1247.275 2618.230 1247.645 ;
        RECT 2618.020 1243.710 2618.160 1247.275 ;
        RECT 2617.960 1243.390 2618.220 1243.710 ;
        RECT 2639.580 1243.390 2639.840 1243.710 ;
        RECT 2639.640 38.070 2639.780 1243.390 ;
        RECT 62.200 37.750 62.460 38.070 ;
        RECT 2639.580 37.750 2639.840 38.070 ;
        RECT 62.260 2.400 62.400 37.750 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 2617.950 1247.320 2618.230 1247.600 ;
      LAYER met3 ;
        RECT 2606.000 1247.610 2610.000 1248.000 ;
        RECT 2617.925 1247.610 2618.255 1247.625 ;
        RECT 2606.000 1247.400 2618.255 1247.610 ;
        RECT 2609.580 1247.310 2618.255 1247.400 ;
        RECT 2617.925 1247.295 2618.255 1247.310 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.510 246.060 420.830 246.120 ;
        RECT 1185.030 246.060 1185.350 246.120 ;
        RECT 420.510 245.920 1185.350 246.060 ;
        RECT 420.510 245.860 420.830 245.920 ;
        RECT 1185.030 245.860 1185.350 245.920 ;
        RECT 419.130 14.180 419.450 14.240 ;
        RECT 420.510 14.180 420.830 14.240 ;
        RECT 419.130 14.040 420.830 14.180 ;
        RECT 419.130 13.980 419.450 14.040 ;
        RECT 420.510 13.980 420.830 14.040 ;
      LAYER via ;
        RECT 420.540 245.860 420.800 246.120 ;
        RECT 1185.060 245.860 1185.320 246.120 ;
        RECT 419.160 13.980 419.420 14.240 ;
        RECT 420.540 13.980 420.800 14.240 ;
      LAYER met2 ;
        RECT 1185.010 260.000 1185.290 264.000 ;
        RECT 1185.120 246.150 1185.260 260.000 ;
        RECT 420.540 245.830 420.800 246.150 ;
        RECT 1185.060 245.830 1185.320 246.150 ;
        RECT 420.600 14.270 420.740 245.830 ;
        RECT 419.160 13.950 419.420 14.270 ;
        RECT 420.540 13.950 420.800 14.270 ;
        RECT 419.220 2.400 419.360 13.950 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 271.930 1421.780 272.250 1421.840 ;
        RECT 296.770 1421.780 297.090 1421.840 ;
        RECT 271.930 1421.640 297.090 1421.780 ;
        RECT 271.930 1421.580 272.250 1421.640 ;
        RECT 296.770 1421.580 297.090 1421.640 ;
        RECT 271.930 24.380 272.250 24.440 ;
        RECT 436.610 24.380 436.930 24.440 ;
        RECT 271.930 24.240 436.930 24.380 ;
        RECT 271.930 24.180 272.250 24.240 ;
        RECT 436.610 24.180 436.930 24.240 ;
      LAYER via ;
        RECT 271.960 1421.580 272.220 1421.840 ;
        RECT 296.800 1421.580 297.060 1421.840 ;
        RECT 271.960 24.180 272.220 24.440 ;
        RECT 436.640 24.180 436.900 24.440 ;
      LAYER met2 ;
        RECT 296.790 1425.435 297.070 1425.805 ;
        RECT 296.860 1421.870 297.000 1425.435 ;
        RECT 271.960 1421.550 272.220 1421.870 ;
        RECT 296.800 1421.550 297.060 1421.870 ;
        RECT 272.020 24.470 272.160 1421.550 ;
        RECT 271.960 24.150 272.220 24.470 ;
        RECT 436.640 24.150 436.900 24.470 ;
        RECT 436.700 2.400 436.840 24.150 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 296.790 1425.480 297.070 1425.760 ;
      LAYER met3 ;
        RECT 296.765 1425.770 297.095 1425.785 ;
        RECT 310.000 1425.770 314.000 1426.160 ;
        RECT 296.765 1425.560 314.000 1425.770 ;
        RECT 296.765 1425.470 310.500 1425.560 ;
        RECT 296.765 1425.455 297.095 1425.470 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 272.850 1718.260 273.170 1718.320 ;
        RECT 296.770 1718.260 297.090 1718.320 ;
        RECT 272.850 1718.120 297.090 1718.260 ;
        RECT 272.850 1718.060 273.170 1718.120 ;
        RECT 296.770 1718.060 297.090 1718.120 ;
        RECT 272.850 168.880 273.170 168.940 ;
        RECT 448.570 168.880 448.890 168.940 ;
        RECT 272.850 168.740 448.890 168.880 ;
        RECT 272.850 168.680 273.170 168.740 ;
        RECT 448.570 168.680 448.890 168.740 ;
        RECT 448.570 38.320 448.890 38.380 ;
        RECT 454.550 38.320 454.870 38.380 ;
        RECT 448.570 38.180 454.870 38.320 ;
        RECT 448.570 38.120 448.890 38.180 ;
        RECT 454.550 38.120 454.870 38.180 ;
      LAYER via ;
        RECT 272.880 1718.060 273.140 1718.320 ;
        RECT 296.800 1718.060 297.060 1718.320 ;
        RECT 272.880 168.680 273.140 168.940 ;
        RECT 448.600 168.680 448.860 168.940 ;
        RECT 448.600 38.120 448.860 38.380 ;
        RECT 454.580 38.120 454.840 38.380 ;
      LAYER met2 ;
        RECT 296.790 1721.915 297.070 1722.285 ;
        RECT 296.860 1718.350 297.000 1721.915 ;
        RECT 272.880 1718.030 273.140 1718.350 ;
        RECT 296.800 1718.030 297.060 1718.350 ;
        RECT 272.940 168.970 273.080 1718.030 ;
        RECT 272.880 168.650 273.140 168.970 ;
        RECT 448.600 168.650 448.860 168.970 ;
        RECT 448.660 38.410 448.800 168.650 ;
        RECT 448.600 38.090 448.860 38.410 ;
        RECT 454.580 38.090 454.840 38.410 ;
        RECT 454.640 2.400 454.780 38.090 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 296.790 1721.960 297.070 1722.240 ;
      LAYER met3 ;
        RECT 296.765 1722.250 297.095 1722.265 ;
        RECT 310.000 1722.250 314.000 1722.640 ;
        RECT 296.765 1722.040 314.000 1722.250 ;
        RECT 296.765 1721.950 310.500 1722.040 ;
        RECT 296.765 1721.935 297.095 1721.950 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 244.790 1214.720 245.110 1214.780 ;
        RECT 296.770 1214.720 297.090 1214.780 ;
        RECT 244.790 1214.580 297.090 1214.720 ;
        RECT 244.790 1214.520 245.110 1214.580 ;
        RECT 296.770 1214.520 297.090 1214.580 ;
        RECT 244.790 16.560 245.110 16.620 ;
        RECT 472.490 16.560 472.810 16.620 ;
        RECT 244.790 16.420 472.810 16.560 ;
        RECT 244.790 16.360 245.110 16.420 ;
        RECT 472.490 16.360 472.810 16.420 ;
      LAYER via ;
        RECT 244.820 1214.520 245.080 1214.780 ;
        RECT 296.800 1214.520 297.060 1214.780 ;
        RECT 244.820 16.360 245.080 16.620 ;
        RECT 472.520 16.360 472.780 16.620 ;
      LAYER met2 ;
        RECT 244.820 1214.490 245.080 1214.810 ;
        RECT 296.790 1214.635 297.070 1215.005 ;
        RECT 296.800 1214.490 297.060 1214.635 ;
        RECT 244.880 16.650 245.020 1214.490 ;
        RECT 244.820 16.330 245.080 16.650 ;
        RECT 472.520 16.330 472.780 16.650 ;
        RECT 472.580 2.400 472.720 16.330 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 296.790 1214.680 297.070 1214.960 ;
      LAYER met3 ;
        RECT 296.765 1214.970 297.095 1214.985 ;
        RECT 310.000 1214.970 314.000 1215.360 ;
        RECT 296.765 1214.760 314.000 1214.970 ;
        RECT 296.765 1214.670 310.500 1214.760 ;
        RECT 296.765 1214.655 297.095 1214.670 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1305.570 3274.355 1305.850 3274.725 ;
        RECT 1305.640 3260.000 1305.780 3274.355 ;
        RECT 1305.530 3256.000 1305.810 3260.000 ;
        RECT 490.450 260.595 490.730 260.965 ;
        RECT 490.520 2.400 490.660 260.595 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 1305.570 3274.400 1305.850 3274.680 ;
        RECT 490.450 260.640 490.730 260.920 ;
      LAYER met3 ;
        RECT 281.790 3274.690 282.170 3274.700 ;
        RECT 1305.545 3274.690 1305.875 3274.705 ;
        RECT 281.790 3274.390 1305.875 3274.690 ;
        RECT 281.790 3274.380 282.170 3274.390 ;
        RECT 1305.545 3274.375 1305.875 3274.390 ;
        RECT 281.790 260.930 282.170 260.940 ;
        RECT 490.425 260.930 490.755 260.945 ;
        RECT 281.790 260.630 490.755 260.930 ;
        RECT 281.790 260.620 282.170 260.630 ;
        RECT 490.425 260.615 490.755 260.630 ;
      LAYER via3 ;
        RECT 281.820 3274.380 282.140 3274.700 ;
        RECT 281.820 260.620 282.140 260.940 ;
      LAYER met4 ;
        RECT 281.815 3274.375 282.145 3274.705 ;
        RECT 281.830 260.945 282.130 3274.375 ;
        RECT 281.815 260.615 282.145 260.945 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 476.170 3271.040 476.490 3271.100 ;
        RECT 2406.790 3271.040 2407.110 3271.100 ;
        RECT 476.170 3270.900 2407.110 3271.040 ;
        RECT 476.170 3270.840 476.490 3270.900 ;
        RECT 2406.790 3270.840 2407.110 3270.900 ;
        RECT 503.770 16.560 504.090 16.620 ;
        RECT 507.910 16.560 508.230 16.620 ;
        RECT 503.770 16.420 508.230 16.560 ;
        RECT 503.770 16.360 504.090 16.420 ;
        RECT 507.910 16.360 508.230 16.420 ;
      LAYER via ;
        RECT 476.200 3270.840 476.460 3271.100 ;
        RECT 2406.820 3270.840 2407.080 3271.100 ;
        RECT 503.800 16.360 504.060 16.620 ;
        RECT 507.940 16.360 508.200 16.620 ;
      LAYER met2 ;
        RECT 476.190 3272.995 476.470 3273.365 ;
        RECT 476.260 3271.130 476.400 3272.995 ;
        RECT 476.200 3270.810 476.460 3271.130 ;
        RECT 2406.820 3270.810 2407.080 3271.130 ;
        RECT 2406.880 3260.000 2407.020 3270.810 ;
        RECT 2406.770 3256.000 2407.050 3260.000 ;
        RECT 503.790 258.555 504.070 258.925 ;
        RECT 503.860 16.650 504.000 258.555 ;
        RECT 503.800 16.330 504.060 16.650 ;
        RECT 507.940 16.330 508.200 16.650 ;
        RECT 508.000 2.400 508.140 16.330 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 476.190 3273.040 476.470 3273.320 ;
        RECT 503.790 258.600 504.070 258.880 ;
      LAYER met3 ;
        RECT 266.150 3273.330 266.530 3273.340 ;
        RECT 476.165 3273.330 476.495 3273.345 ;
        RECT 266.150 3273.030 476.495 3273.330 ;
        RECT 266.150 3273.020 266.530 3273.030 ;
        RECT 476.165 3273.015 476.495 3273.030 ;
        RECT 266.150 258.890 266.530 258.900 ;
        RECT 503.765 258.890 504.095 258.905 ;
        RECT 266.150 258.590 504.095 258.890 ;
        RECT 266.150 258.580 266.530 258.590 ;
        RECT 503.765 258.575 504.095 258.590 ;
      LAYER via3 ;
        RECT 266.180 3273.020 266.500 3273.340 ;
        RECT 266.180 258.580 266.500 258.900 ;
      LAYER met4 ;
        RECT 266.175 3273.015 266.505 3273.345 ;
        RECT 266.190 258.905 266.490 3273.015 ;
        RECT 266.175 258.575 266.505 258.905 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 273.310 1821.960 273.630 1822.020 ;
        RECT 296.770 1821.960 297.090 1822.020 ;
        RECT 273.310 1821.820 297.090 1821.960 ;
        RECT 273.310 1821.760 273.630 1821.820 ;
        RECT 296.770 1821.760 297.090 1821.820 ;
        RECT 273.310 162.080 273.630 162.140 ;
        RECT 524.470 162.080 524.790 162.140 ;
        RECT 273.310 161.940 524.790 162.080 ;
        RECT 273.310 161.880 273.630 161.940 ;
        RECT 524.470 161.880 524.790 161.940 ;
      LAYER via ;
        RECT 273.340 1821.760 273.600 1822.020 ;
        RECT 296.800 1821.760 297.060 1822.020 ;
        RECT 273.340 161.880 273.600 162.140 ;
        RECT 524.500 161.880 524.760 162.140 ;
      LAYER met2 ;
        RECT 296.790 1827.995 297.070 1828.365 ;
        RECT 296.860 1822.050 297.000 1827.995 ;
        RECT 273.340 1821.730 273.600 1822.050 ;
        RECT 296.800 1821.730 297.060 1822.050 ;
        RECT 273.400 162.170 273.540 1821.730 ;
        RECT 273.340 161.850 273.600 162.170 ;
        RECT 524.500 161.850 524.760 162.170 ;
        RECT 524.560 3.130 524.700 161.850 ;
        RECT 524.560 2.990 526.080 3.130 ;
        RECT 525.940 2.400 526.080 2.990 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 296.790 1828.040 297.070 1828.320 ;
      LAYER met3 ;
        RECT 296.765 1828.330 297.095 1828.345 ;
        RECT 310.000 1828.330 314.000 1828.720 ;
        RECT 296.765 1828.120 314.000 1828.330 ;
        RECT 296.765 1828.030 310.500 1828.120 ;
        RECT 296.765 1828.015 297.095 1828.030 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.210 260.000 303.530 260.060 ;
        RECT 538.270 260.000 538.590 260.060 ;
        RECT 303.210 259.860 538.590 260.000 ;
        RECT 303.210 259.800 303.530 259.860 ;
        RECT 538.270 259.800 538.590 259.860 ;
        RECT 538.270 2.960 538.590 3.020 ;
        RECT 543.790 2.960 544.110 3.020 ;
        RECT 538.270 2.820 544.110 2.960 ;
        RECT 538.270 2.760 538.590 2.820 ;
        RECT 543.790 2.760 544.110 2.820 ;
      LAYER via ;
        RECT 303.240 259.800 303.500 260.060 ;
        RECT 538.300 259.800 538.560 260.060 ;
        RECT 538.300 2.760 538.560 3.020 ;
        RECT 543.820 2.760 544.080 3.020 ;
      LAYER met2 ;
        RECT 303.230 348.315 303.510 348.685 ;
        RECT 303.300 260.090 303.440 348.315 ;
        RECT 303.240 259.770 303.500 260.090 ;
        RECT 538.300 259.770 538.560 260.090 ;
        RECT 538.360 3.050 538.500 259.770 ;
        RECT 538.300 2.730 538.560 3.050 ;
        RECT 543.820 2.730 544.080 3.050 ;
        RECT 543.880 2.400 544.020 2.730 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 303.230 348.360 303.510 348.640 ;
      LAYER met3 ;
        RECT 303.205 348.650 303.535 348.665 ;
        RECT 310.000 348.650 314.000 349.040 ;
        RECT 303.205 348.440 314.000 348.650 ;
        RECT 303.205 348.350 310.500 348.440 ;
        RECT 303.205 348.335 303.535 348.350 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 38.320 562.050 38.380 ;
        RECT 2617.010 38.320 2617.330 38.380 ;
        RECT 561.730 38.180 2617.330 38.320 ;
        RECT 561.730 38.120 562.050 38.180 ;
        RECT 2617.010 38.120 2617.330 38.180 ;
      LAYER via ;
        RECT 561.760 38.120 562.020 38.380 ;
        RECT 2617.040 38.120 2617.300 38.380 ;
      LAYER met2 ;
        RECT 2617.030 760.395 2617.310 760.765 ;
        RECT 2617.100 38.410 2617.240 760.395 ;
        RECT 561.760 38.090 562.020 38.410 ;
        RECT 2617.040 38.090 2617.300 38.410 ;
        RECT 561.820 2.400 561.960 38.090 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 2617.030 760.440 2617.310 760.720 ;
      LAYER met3 ;
        RECT 2606.000 760.730 2610.000 761.120 ;
        RECT 2617.005 760.730 2617.335 760.745 ;
        RECT 2606.000 760.520 2617.335 760.730 ;
        RECT 2609.580 760.430 2617.335 760.520 ;
        RECT 2617.005 760.415 2617.335 760.430 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.690 51.155 579.970 51.525 ;
        RECT 579.760 2.400 579.900 51.155 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 579.690 51.200 579.970 51.480 ;
      LAYER met3 ;
        RECT 2606.000 2430.810 2610.000 2431.200 ;
        RECT 2637.910 2430.810 2638.290 2430.820 ;
        RECT 2606.000 2430.600 2638.290 2430.810 ;
        RECT 2609.580 2430.510 2638.290 2430.600 ;
        RECT 2637.910 2430.500 2638.290 2430.510 ;
        RECT 579.665 51.490 579.995 51.505 ;
        RECT 2637.910 51.490 2638.290 51.500 ;
        RECT 579.665 51.190 2638.290 51.490 ;
        RECT 579.665 51.175 579.995 51.190 ;
        RECT 2637.910 51.180 2638.290 51.190 ;
      LAYER via3 ;
        RECT 2637.940 2430.500 2638.260 2430.820 ;
        RECT 2637.940 51.180 2638.260 51.500 ;
      LAYER met4 ;
        RECT 2637.935 2430.495 2638.265 2430.825 ;
        RECT 2637.950 51.505 2638.250 2430.495 ;
        RECT 2637.935 51.175 2638.265 51.505 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 89.310 3258.800 89.630 3258.860 ;
        RECT 1260.470 3258.800 1260.790 3258.860 ;
        RECT 89.310 3258.660 1260.790 3258.800 ;
        RECT 89.310 3258.600 89.630 3258.660 ;
        RECT 1260.470 3258.600 1260.790 3258.660 ;
        RECT 86.090 16.900 86.410 16.960 ;
        RECT 89.310 16.900 89.630 16.960 ;
        RECT 86.090 16.760 89.630 16.900 ;
        RECT 86.090 16.700 86.410 16.760 ;
        RECT 89.310 16.700 89.630 16.760 ;
      LAYER via ;
        RECT 89.340 3258.600 89.600 3258.860 ;
        RECT 1260.500 3258.600 1260.760 3258.860 ;
        RECT 86.120 16.700 86.380 16.960 ;
        RECT 89.340 16.700 89.600 16.960 ;
      LAYER met2 ;
        RECT 1262.290 3258.970 1262.570 3260.000 ;
        RECT 1260.560 3258.890 1262.570 3258.970 ;
        RECT 89.340 3258.570 89.600 3258.890 ;
        RECT 1260.500 3258.830 1262.570 3258.890 ;
        RECT 1260.500 3258.570 1260.760 3258.830 ;
        RECT 89.400 16.990 89.540 3258.570 ;
        RECT 1262.290 3256.000 1262.570 3258.830 ;
        RECT 86.120 16.670 86.380 16.990 ;
        RECT 89.340 16.670 89.600 16.990 ;
        RECT 86.180 2.400 86.320 16.670 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 239.730 3257.440 240.050 3257.500 ;
        RECT 817.950 3257.440 818.270 3257.500 ;
        RECT 239.730 3257.300 818.270 3257.440 ;
        RECT 239.730 3257.240 240.050 3257.300 ;
        RECT 817.950 3257.240 818.270 3257.300 ;
        RECT 239.730 245.040 240.050 245.100 ;
        RECT 593.470 245.040 593.790 245.100 ;
        RECT 239.730 244.900 593.790 245.040 ;
        RECT 239.730 244.840 240.050 244.900 ;
        RECT 593.470 244.840 593.790 244.900 ;
        RECT 593.470 18.940 593.790 19.000 ;
        RECT 597.150 18.940 597.470 19.000 ;
        RECT 593.470 18.800 597.470 18.940 ;
        RECT 593.470 18.740 593.790 18.800 ;
        RECT 597.150 18.740 597.470 18.800 ;
      LAYER via ;
        RECT 239.760 3257.240 240.020 3257.500 ;
        RECT 817.980 3257.240 818.240 3257.500 ;
        RECT 239.760 244.840 240.020 245.100 ;
        RECT 593.500 244.840 593.760 245.100 ;
        RECT 593.500 18.740 593.760 19.000 ;
        RECT 597.180 18.740 597.440 19.000 ;
      LAYER met2 ;
        RECT 819.770 3257.610 820.050 3260.000 ;
        RECT 818.040 3257.530 820.050 3257.610 ;
        RECT 239.760 3257.210 240.020 3257.530 ;
        RECT 817.980 3257.470 820.050 3257.530 ;
        RECT 817.980 3257.210 818.240 3257.470 ;
        RECT 239.820 245.130 239.960 3257.210 ;
        RECT 819.770 3256.000 820.050 3257.470 ;
        RECT 239.760 244.810 240.020 245.130 ;
        RECT 593.500 244.810 593.760 245.130 ;
        RECT 593.560 19.030 593.700 244.810 ;
        RECT 593.500 18.710 593.760 19.030 ;
        RECT 597.180 18.710 597.440 19.030 ;
        RECT 597.240 2.400 597.380 18.710 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 20.640 615.410 20.700 ;
        RECT 620.610 20.640 620.930 20.700 ;
        RECT 615.090 20.500 620.930 20.640 ;
        RECT 615.090 20.440 615.410 20.500 ;
        RECT 620.610 20.440 620.930 20.500 ;
      LAYER via ;
        RECT 615.120 20.440 615.380 20.700 ;
        RECT 620.640 20.440 620.900 20.700 ;
      LAYER met2 ;
        RECT 620.630 85.835 620.910 86.205 ;
        RECT 620.700 20.730 620.840 85.835 ;
        RECT 615.120 20.410 615.380 20.730 ;
        RECT 620.640 20.410 620.900 20.730 ;
        RECT 615.180 2.400 615.320 20.410 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 620.630 85.880 620.910 86.160 ;
      LAYER met3 ;
        RECT 2606.000 2410.410 2610.000 2410.800 ;
        RECT 2638.830 2410.410 2639.210 2410.420 ;
        RECT 2606.000 2410.200 2639.210 2410.410 ;
        RECT 2609.580 2410.110 2639.210 2410.200 ;
        RECT 2638.830 2410.100 2639.210 2410.110 ;
        RECT 620.605 86.170 620.935 86.185 ;
        RECT 2638.830 86.170 2639.210 86.180 ;
        RECT 620.605 85.870 2639.210 86.170 ;
        RECT 620.605 85.855 620.935 85.870 ;
        RECT 2638.830 85.860 2639.210 85.870 ;
      LAYER via3 ;
        RECT 2638.860 2410.100 2639.180 2410.420 ;
        RECT 2638.860 85.860 2639.180 86.180 ;
      LAYER met4 ;
        RECT 2638.855 2410.095 2639.185 2410.425 ;
        RECT 2638.870 86.185 2639.170 2410.095 ;
        RECT 2638.855 85.855 2639.185 86.185 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 46.480 109.870 46.540 ;
        RECT 2111.470 46.480 2111.790 46.540 ;
        RECT 109.550 46.340 2111.790 46.480 ;
        RECT 109.550 46.280 109.870 46.340 ;
        RECT 2111.470 46.280 2111.790 46.340 ;
      LAYER via ;
        RECT 109.580 46.280 109.840 46.540 ;
        RECT 2111.500 46.280 2111.760 46.540 ;
      LAYER met2 ;
        RECT 2114.210 260.170 2114.490 264.000 ;
        RECT 2111.560 260.030 2114.490 260.170 ;
        RECT 2111.560 46.570 2111.700 260.030 ;
        RECT 2114.210 260.000 2114.490 260.030 ;
        RECT 109.580 46.250 109.840 46.570 ;
        RECT 2111.500 46.250 2111.760 46.570 ;
        RECT 109.640 2.400 109.780 46.250 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1035.070 251.160 1035.390 251.220 ;
        RECT 1041.510 251.160 1041.830 251.220 ;
        RECT 1035.070 251.020 1041.830 251.160 ;
        RECT 1035.070 250.960 1035.390 251.020 ;
        RECT 1041.510 250.960 1041.830 251.020 ;
        RECT 133.470 32.880 133.790 32.940 ;
        RECT 1035.070 32.880 1035.390 32.940 ;
        RECT 133.470 32.740 1035.390 32.880 ;
        RECT 133.470 32.680 133.790 32.740 ;
        RECT 1035.070 32.680 1035.390 32.740 ;
      LAYER via ;
        RECT 1035.100 250.960 1035.360 251.220 ;
        RECT 1041.540 250.960 1041.800 251.220 ;
        RECT 133.500 32.680 133.760 32.940 ;
        RECT 1035.100 32.680 1035.360 32.940 ;
      LAYER met2 ;
        RECT 1041.490 260.000 1041.770 264.000 ;
        RECT 1041.600 251.250 1041.740 260.000 ;
        RECT 1035.100 250.930 1035.360 251.250 ;
        RECT 1041.540 250.930 1041.800 251.250 ;
        RECT 1035.160 32.970 1035.300 250.930 ;
        RECT 133.500 32.650 133.760 32.970 ;
        RECT 1035.100 32.650 1035.360 32.970 ;
        RECT 133.560 2.400 133.700 32.650 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 303.860 169.670 303.920 ;
        RECT 296.770 303.860 297.090 303.920 ;
        RECT 169.350 303.720 297.090 303.860 ;
        RECT 169.350 303.660 169.670 303.720 ;
        RECT 296.770 303.660 297.090 303.720 ;
        RECT 151.410 20.980 151.730 21.040 ;
        RECT 169.350 20.980 169.670 21.040 ;
        RECT 151.410 20.840 169.670 20.980 ;
        RECT 151.410 20.780 151.730 20.840 ;
        RECT 169.350 20.780 169.670 20.840 ;
      LAYER via ;
        RECT 169.380 303.660 169.640 303.920 ;
        RECT 296.800 303.660 297.060 303.920 ;
        RECT 151.440 20.780 151.700 21.040 ;
        RECT 169.380 20.780 169.640 21.040 ;
      LAYER met2 ;
        RECT 296.790 306.155 297.070 306.525 ;
        RECT 296.860 303.950 297.000 306.155 ;
        RECT 169.380 303.630 169.640 303.950 ;
        RECT 296.800 303.630 297.060 303.950 ;
        RECT 169.440 21.070 169.580 303.630 ;
        RECT 151.440 20.750 151.700 21.070 ;
        RECT 169.380 20.750 169.640 21.070 ;
        RECT 151.500 2.400 151.640 20.750 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 296.790 306.200 297.070 306.480 ;
      LAYER met3 ;
        RECT 296.765 306.490 297.095 306.505 ;
        RECT 310.000 306.490 314.000 306.880 ;
        RECT 296.765 306.280 314.000 306.490 ;
        RECT 296.765 306.190 310.500 306.280 ;
        RECT 296.765 306.175 297.095 306.190 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1003.790 247.080 1004.110 247.140 ;
        RECT 1213.550 247.080 1213.870 247.140 ;
        RECT 1003.790 246.940 1213.870 247.080 ;
        RECT 1003.790 246.880 1004.110 246.940 ;
        RECT 1213.550 246.880 1213.870 246.940 ;
        RECT 172.110 169.220 172.430 169.280 ;
        RECT 1003.790 169.220 1004.110 169.280 ;
        RECT 172.110 169.080 1004.110 169.220 ;
        RECT 172.110 169.020 172.430 169.080 ;
        RECT 1003.790 169.020 1004.110 169.080 ;
        RECT 169.350 17.580 169.670 17.640 ;
        RECT 172.110 17.580 172.430 17.640 ;
        RECT 169.350 17.440 172.430 17.580 ;
        RECT 169.350 17.380 169.670 17.440 ;
        RECT 172.110 17.380 172.430 17.440 ;
      LAYER via ;
        RECT 1003.820 246.880 1004.080 247.140 ;
        RECT 1213.580 246.880 1213.840 247.140 ;
        RECT 172.140 169.020 172.400 169.280 ;
        RECT 1003.820 169.020 1004.080 169.280 ;
        RECT 169.380 17.380 169.640 17.640 ;
        RECT 172.140 17.380 172.400 17.640 ;
      LAYER met2 ;
        RECT 1213.530 260.000 1213.810 264.000 ;
        RECT 1213.640 247.170 1213.780 260.000 ;
        RECT 1003.820 246.850 1004.080 247.170 ;
        RECT 1213.580 246.850 1213.840 247.170 ;
        RECT 1003.880 169.310 1004.020 246.850 ;
        RECT 172.140 168.990 172.400 169.310 ;
        RECT 1003.820 168.990 1004.080 169.310 ;
        RECT 172.200 17.670 172.340 168.990 ;
        RECT 169.380 17.350 169.640 17.670 ;
        RECT 172.140 17.350 172.400 17.670 ;
        RECT 169.440 2.400 169.580 17.350 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 3259.480 193.130 3259.540 ;
        RECT 1360.750 3259.480 1361.070 3259.540 ;
        RECT 192.810 3259.340 1361.070 3259.480 ;
        RECT 192.810 3259.280 193.130 3259.340 ;
        RECT 1360.750 3259.280 1361.070 3259.340 ;
        RECT 186.830 17.580 187.150 17.640 ;
        RECT 192.810 17.580 193.130 17.640 ;
        RECT 186.830 17.440 193.130 17.580 ;
        RECT 186.830 17.380 187.150 17.440 ;
        RECT 192.810 17.380 193.130 17.440 ;
      LAYER via ;
        RECT 192.840 3259.280 193.100 3259.540 ;
        RECT 1360.780 3259.280 1361.040 3259.540 ;
        RECT 186.860 17.380 187.120 17.640 ;
        RECT 192.840 17.380 193.100 17.640 ;
      LAYER met2 ;
        RECT 1362.570 3259.650 1362.850 3260.000 ;
        RECT 1360.840 3259.570 1362.850 3259.650 ;
        RECT 192.840 3259.250 193.100 3259.570 ;
        RECT 1360.780 3259.510 1362.850 3259.570 ;
        RECT 1360.780 3259.250 1361.040 3259.510 ;
        RECT 192.900 17.670 193.040 3259.250 ;
        RECT 1362.570 3256.000 1362.850 3259.510 ;
        RECT 186.860 17.350 187.120 17.670 ;
        RECT 192.840 17.350 193.100 17.670 ;
        RECT 186.920 2.400 187.060 17.350 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 45.120 205.090 45.180 ;
        RECT 2366.770 45.120 2367.090 45.180 ;
        RECT 204.770 44.980 2367.090 45.120 ;
        RECT 204.770 44.920 205.090 44.980 ;
        RECT 2366.770 44.920 2367.090 44.980 ;
      LAYER via ;
        RECT 204.800 44.920 205.060 45.180 ;
        RECT 2366.800 44.920 2367.060 45.180 ;
      LAYER met2 ;
        RECT 2371.810 260.170 2372.090 264.000 ;
        RECT 2366.860 260.030 2372.090 260.170 ;
        RECT 2366.860 45.210 2367.000 260.030 ;
        RECT 2371.810 260.000 2372.090 260.030 ;
        RECT 204.800 44.890 205.060 45.210 ;
        RECT 2366.800 44.890 2367.060 45.210 ;
        RECT 204.860 2.400 205.000 44.890 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 1539.080 2615.490 1539.140 ;
        RECT 2639.090 1539.080 2639.410 1539.140 ;
        RECT 2615.170 1538.940 2639.410 1539.080 ;
        RECT 2615.170 1538.880 2615.490 1538.940 ;
        RECT 2639.090 1538.880 2639.410 1538.940 ;
        RECT 226.390 120.600 226.710 120.660 ;
        RECT 2639.090 120.600 2639.410 120.660 ;
        RECT 226.390 120.460 2639.410 120.600 ;
        RECT 226.390 120.400 226.710 120.460 ;
        RECT 2639.090 120.400 2639.410 120.460 ;
        RECT 222.710 17.580 223.030 17.640 ;
        RECT 226.390 17.580 226.710 17.640 ;
        RECT 222.710 17.440 226.710 17.580 ;
        RECT 222.710 17.380 223.030 17.440 ;
        RECT 226.390 17.380 226.710 17.440 ;
      LAYER via ;
        RECT 2615.200 1538.880 2615.460 1539.140 ;
        RECT 2639.120 1538.880 2639.380 1539.140 ;
        RECT 226.420 120.400 226.680 120.660 ;
        RECT 2639.120 120.400 2639.380 120.660 ;
        RECT 222.740 17.380 223.000 17.640 ;
        RECT 226.420 17.380 226.680 17.640 ;
      LAYER met2 ;
        RECT 2615.190 1543.755 2615.470 1544.125 ;
        RECT 2615.260 1539.170 2615.400 1543.755 ;
        RECT 2615.200 1538.850 2615.460 1539.170 ;
        RECT 2639.120 1538.850 2639.380 1539.170 ;
        RECT 2639.180 120.690 2639.320 1538.850 ;
        RECT 226.420 120.370 226.680 120.690 ;
        RECT 2639.120 120.370 2639.380 120.690 ;
        RECT 226.480 17.670 226.620 120.370 ;
        RECT 222.740 17.350 223.000 17.670 ;
        RECT 226.420 17.350 226.680 17.670 ;
        RECT 222.800 2.400 222.940 17.350 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 2615.190 1543.800 2615.470 1544.080 ;
      LAYER met3 ;
        RECT 2606.000 1544.090 2610.000 1544.480 ;
        RECT 2615.165 1544.090 2615.495 1544.105 ;
        RECT 2606.000 1543.880 2615.495 1544.090 ;
        RECT 2609.580 1543.790 2615.495 1543.880 ;
        RECT 2615.165 1543.775 2615.495 1543.790 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.150 510.920 45.470 510.980 ;
        RECT 296.770 510.920 297.090 510.980 ;
        RECT 45.150 510.780 297.090 510.920 ;
        RECT 45.150 510.720 45.470 510.780 ;
        RECT 296.770 510.720 297.090 510.780 ;
        RECT 20.310 15.200 20.630 15.260 ;
        RECT 45.150 15.200 45.470 15.260 ;
        RECT 20.310 15.060 45.470 15.200 ;
        RECT 20.310 15.000 20.630 15.060 ;
        RECT 45.150 15.000 45.470 15.060 ;
      LAYER via ;
        RECT 45.180 510.720 45.440 510.980 ;
        RECT 296.800 510.720 297.060 510.980 ;
        RECT 20.340 15.000 20.600 15.260 ;
        RECT 45.180 15.000 45.440 15.260 ;
      LAYER met2 ;
        RECT 296.790 516.955 297.070 517.325 ;
        RECT 296.860 511.010 297.000 516.955 ;
        RECT 45.180 510.690 45.440 511.010 ;
        RECT 296.800 510.690 297.060 511.010 ;
        RECT 45.240 15.290 45.380 510.690 ;
        RECT 20.340 14.970 20.600 15.290 ;
        RECT 45.180 14.970 45.440 15.290 ;
        RECT 20.400 2.400 20.540 14.970 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 296.790 517.000 297.070 517.280 ;
      LAYER met3 ;
        RECT 296.765 517.290 297.095 517.305 ;
        RECT 310.000 517.290 314.000 517.680 ;
        RECT 296.765 517.080 314.000 517.290 ;
        RECT 296.765 516.990 310.500 517.080 ;
        RECT 296.765 516.975 297.095 516.990 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 983.090 245.720 983.410 245.780 ;
        RECT 1899.870 245.720 1900.190 245.780 ;
        RECT 983.090 245.580 1900.190 245.720 ;
        RECT 983.090 245.520 983.410 245.580 ;
        RECT 1899.870 245.520 1900.190 245.580 ;
        RECT 47.910 134.880 48.230 134.940 ;
        RECT 983.090 134.880 983.410 134.940 ;
        RECT 47.910 134.740 983.410 134.880 ;
        RECT 47.910 134.680 48.230 134.740 ;
        RECT 983.090 134.680 983.410 134.740 ;
        RECT 44.230 15.540 44.550 15.600 ;
        RECT 47.910 15.540 48.230 15.600 ;
        RECT 44.230 15.400 48.230 15.540 ;
        RECT 44.230 15.340 44.550 15.400 ;
        RECT 47.910 15.340 48.230 15.400 ;
      LAYER via ;
        RECT 983.120 245.520 983.380 245.780 ;
        RECT 1899.900 245.520 1900.160 245.780 ;
        RECT 47.940 134.680 48.200 134.940 ;
        RECT 983.120 134.680 983.380 134.940 ;
        RECT 44.260 15.340 44.520 15.600 ;
        RECT 47.940 15.340 48.200 15.600 ;
      LAYER met2 ;
        RECT 1899.850 260.000 1900.130 264.000 ;
        RECT 1899.960 245.810 1900.100 260.000 ;
        RECT 983.120 245.490 983.380 245.810 ;
        RECT 1899.900 245.490 1900.160 245.810 ;
        RECT 983.180 134.970 983.320 245.490 ;
        RECT 47.940 134.650 48.200 134.970 ;
        RECT 983.120 134.650 983.380 134.970 ;
        RECT 48.000 15.630 48.140 134.650 ;
        RECT 44.260 15.310 44.520 15.630 ;
        RECT 47.940 15.310 48.200 15.630 ;
        RECT 44.320 2.400 44.460 15.310 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 247.550 3260.160 247.870 3260.220 ;
        RECT 1174.910 3260.160 1175.230 3260.220 ;
        RECT 247.550 3260.020 1175.230 3260.160 ;
        RECT 247.550 3259.960 247.870 3260.020 ;
        RECT 1174.910 3259.960 1175.230 3260.020 ;
      LAYER via ;
        RECT 247.580 3259.960 247.840 3260.220 ;
        RECT 1174.940 3259.960 1175.200 3260.220 ;
      LAYER met2 ;
        RECT 247.580 3259.930 247.840 3260.250 ;
        RECT 1174.940 3259.930 1175.200 3260.250 ;
        RECT 247.640 3.130 247.780 3259.930 ;
        RECT 1175.000 3259.650 1175.140 3259.930 ;
        RECT 1176.730 3259.650 1177.010 3260.000 ;
        RECT 1175.000 3259.510 1177.010 3259.650 ;
        RECT 1176.730 3256.000 1177.010 3259.510 ;
        RECT 246.720 2.990 247.780 3.130 ;
        RECT 246.720 2.400 246.860 2.990 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1252.190 247.080 1252.510 247.140 ;
        RECT 1656.990 247.080 1657.310 247.140 ;
        RECT 1252.190 246.940 1657.310 247.080 ;
        RECT 1252.190 246.880 1252.510 246.940 ;
        RECT 1656.990 246.880 1657.310 246.940 ;
        RECT 268.710 66.200 269.030 66.260 ;
        RECT 1252.190 66.200 1252.510 66.260 ;
        RECT 268.710 66.060 1252.510 66.200 ;
        RECT 268.710 66.000 269.030 66.060 ;
        RECT 1252.190 66.000 1252.510 66.060 ;
        RECT 264.110 17.920 264.430 17.980 ;
        RECT 268.710 17.920 269.030 17.980 ;
        RECT 264.110 17.780 269.030 17.920 ;
        RECT 264.110 17.720 264.430 17.780 ;
        RECT 268.710 17.720 269.030 17.780 ;
      LAYER via ;
        RECT 1252.220 246.880 1252.480 247.140 ;
        RECT 1657.020 246.880 1657.280 247.140 ;
        RECT 268.740 66.000 269.000 66.260 ;
        RECT 1252.220 66.000 1252.480 66.260 ;
        RECT 264.140 17.720 264.400 17.980 ;
        RECT 268.740 17.720 269.000 17.980 ;
      LAYER met2 ;
        RECT 1656.970 260.000 1657.250 264.000 ;
        RECT 1657.080 247.170 1657.220 260.000 ;
        RECT 1252.220 246.850 1252.480 247.170 ;
        RECT 1657.020 246.850 1657.280 247.170 ;
        RECT 1252.280 66.290 1252.420 246.850 ;
        RECT 268.740 65.970 269.000 66.290 ;
        RECT 1252.220 65.970 1252.480 66.290 ;
        RECT 268.800 18.010 268.940 65.970 ;
        RECT 264.140 17.690 264.400 18.010 ;
        RECT 268.740 17.690 269.000 18.010 ;
        RECT 264.200 2.400 264.340 17.690 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1814.845 245.225 1815.015 246.415 ;
      LAYER mcon ;
        RECT 1814.845 246.245 1815.015 246.415 ;
      LAYER met1 ;
        RECT 1814.785 246.400 1815.075 246.445 ;
        RECT 1871.350 246.400 1871.670 246.460 ;
        RECT 1814.785 246.260 1871.670 246.400 ;
        RECT 1814.785 246.215 1815.075 246.260 ;
        RECT 1871.350 246.200 1871.670 246.260 ;
        RECT 1811.090 245.380 1811.410 245.440 ;
        RECT 1814.785 245.380 1815.075 245.425 ;
        RECT 1811.090 245.240 1815.075 245.380 ;
        RECT 1811.090 245.180 1811.410 245.240 ;
        RECT 1814.785 245.195 1815.075 245.240 ;
        RECT 280.670 128.420 280.990 128.480 ;
        RECT 1811.090 128.420 1811.410 128.480 ;
        RECT 280.670 128.280 1811.410 128.420 ;
        RECT 280.670 128.220 280.990 128.280 ;
        RECT 1811.090 128.220 1811.410 128.280 ;
      LAYER via ;
        RECT 1871.380 246.200 1871.640 246.460 ;
        RECT 1811.120 245.180 1811.380 245.440 ;
        RECT 280.700 128.220 280.960 128.480 ;
        RECT 1811.120 128.220 1811.380 128.480 ;
      LAYER met2 ;
        RECT 1871.330 260.000 1871.610 264.000 ;
        RECT 1871.440 246.490 1871.580 260.000 ;
        RECT 1871.380 246.170 1871.640 246.490 ;
        RECT 1811.120 245.150 1811.380 245.470 ;
        RECT 1811.180 128.510 1811.320 245.150 ;
        RECT 280.700 128.190 280.960 128.510 ;
        RECT 1811.120 128.190 1811.380 128.510 ;
        RECT 280.760 3.130 280.900 128.190 ;
        RECT 280.760 2.990 282.280 3.130 ;
        RECT 282.140 2.400 282.280 2.990 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 38.660 300.310 38.720 ;
        RECT 724.570 38.660 724.890 38.720 ;
        RECT 299.990 38.520 724.890 38.660 ;
        RECT 299.990 38.460 300.310 38.520 ;
        RECT 724.570 38.460 724.890 38.520 ;
      LAYER via ;
        RECT 300.020 38.460 300.280 38.720 ;
        RECT 724.600 38.460 724.860 38.720 ;
      LAYER met2 ;
        RECT 726.850 260.170 727.130 264.000 ;
        RECT 724.660 260.030 727.130 260.170 ;
        RECT 724.660 38.750 724.800 260.030 ;
        RECT 726.850 260.000 727.130 260.030 ;
        RECT 300.020 38.430 300.280 38.750 ;
        RECT 724.600 38.430 724.860 38.750 ;
        RECT 300.080 2.400 300.220 38.430 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 250.770 855.680 251.090 855.740 ;
        RECT 296.770 855.680 297.090 855.740 ;
        RECT 250.770 855.540 297.090 855.680 ;
        RECT 250.770 855.480 251.090 855.540 ;
        RECT 296.770 855.480 297.090 855.540 ;
        RECT 250.770 16.900 251.090 16.960 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 250.770 16.760 318.250 16.900 ;
        RECT 250.770 16.700 251.090 16.760 ;
        RECT 317.930 16.700 318.250 16.760 ;
      LAYER via ;
        RECT 250.800 855.480 251.060 855.740 ;
        RECT 296.800 855.480 297.060 855.740 ;
        RECT 250.800 16.700 251.060 16.960 ;
        RECT 317.960 16.700 318.220 16.960 ;
      LAYER met2 ;
        RECT 250.800 855.450 251.060 855.770 ;
        RECT 296.790 855.595 297.070 855.965 ;
        RECT 296.800 855.450 297.060 855.595 ;
        RECT 250.860 16.990 251.000 855.450 ;
        RECT 250.800 16.670 251.060 16.990 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 296.790 855.640 297.070 855.920 ;
      LAYER met3 ;
        RECT 296.765 855.930 297.095 855.945 ;
        RECT 310.000 855.930 314.000 856.320 ;
        RECT 296.765 855.720 314.000 855.930 ;
        RECT 296.765 855.630 310.500 855.720 ;
        RECT 296.765 855.615 297.095 855.630 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2063.245 247.265 2063.415 248.115 ;
        RECT 400.805 23.885 401.435 24.055 ;
        RECT 400.805 23.545 400.975 23.885 ;
        RECT 448.185 23.545 448.815 23.715 ;
        RECT 462.445 22.525 462.615 23.715 ;
        RECT 510.285 22.525 510.455 23.715 ;
        RECT 518.105 23.375 518.275 23.715 ;
        RECT 517.645 23.205 518.275 23.375 ;
        RECT 651.505 23.205 651.675 24.055 ;
        RECT 662.545 22.525 662.715 24.055 ;
        RECT 800.545 22.865 800.715 24.055 ;
        RECT 848.385 22.865 848.555 23.715 ;
        RECT 848.845 22.525 849.015 23.375 ;
        RECT 1000.645 22.525 1000.815 23.375 ;
        RECT 1038.825 22.525 1038.995 23.715 ;
        RECT 1200.285 22.865 1200.455 23.715 ;
        RECT 1242.145 22.525 1242.315 23.375 ;
        RECT 1289.985 22.525 1290.155 23.375 ;
        RECT 1297.345 22.525 1297.515 23.375 ;
        RECT 1345.645 22.525 1345.815 24.055 ;
        RECT 1393.945 22.525 1394.115 24.055 ;
        RECT 1441.785 22.525 1441.955 23.715 ;
        RECT 1607.385 23.205 1608.015 23.375 ;
        RECT 1628.545 23.205 1628.715 24.395 ;
        RECT 1676.385 23.545 1676.555 24.395 ;
        RECT 1676.845 22.525 1677.015 23.375 ;
        RECT 1724.685 22.525 1724.855 23.715 ;
        RECT 1731.585 23.545 1732.215 23.715 ;
        RECT 1786.785 23.545 1787.415 23.715 ;
        RECT 1787.245 23.205 1787.415 23.545 ;
        RECT 1821.745 23.205 1821.915 24.055 ;
        RECT 1869.585 23.205 1869.755 24.055 ;
        RECT 1918.345 22.525 1918.515 23.375 ;
        RECT 1966.185 22.525 1966.355 24.055 ;
        RECT 2028.745 23.885 2028.915 27.455 ;
      LAYER mcon ;
        RECT 2063.245 247.945 2063.415 248.115 ;
        RECT 2028.745 27.285 2028.915 27.455 ;
        RECT 1628.545 24.225 1628.715 24.395 ;
        RECT 401.265 23.885 401.435 24.055 ;
        RECT 651.505 23.885 651.675 24.055 ;
        RECT 448.645 23.545 448.815 23.715 ;
        RECT 462.445 23.545 462.615 23.715 ;
        RECT 510.285 23.545 510.455 23.715 ;
        RECT 518.105 23.545 518.275 23.715 ;
        RECT 662.545 23.885 662.715 24.055 ;
        RECT 800.545 23.885 800.715 24.055 ;
        RECT 1345.645 23.885 1345.815 24.055 ;
        RECT 848.385 23.545 848.555 23.715 ;
        RECT 1038.825 23.545 1038.995 23.715 ;
        RECT 848.845 23.205 849.015 23.375 ;
        RECT 1000.645 23.205 1000.815 23.375 ;
        RECT 1200.285 23.545 1200.455 23.715 ;
        RECT 1242.145 23.205 1242.315 23.375 ;
        RECT 1289.985 23.205 1290.155 23.375 ;
        RECT 1297.345 23.205 1297.515 23.375 ;
        RECT 1393.945 23.885 1394.115 24.055 ;
        RECT 1441.785 23.545 1441.955 23.715 ;
        RECT 1676.385 24.225 1676.555 24.395 ;
        RECT 1821.745 23.885 1821.915 24.055 ;
        RECT 1724.685 23.545 1724.855 23.715 ;
        RECT 1732.045 23.545 1732.215 23.715 ;
        RECT 1607.845 23.205 1608.015 23.375 ;
        RECT 1676.845 23.205 1677.015 23.375 ;
        RECT 1869.585 23.885 1869.755 24.055 ;
        RECT 1966.185 23.885 1966.355 24.055 ;
        RECT 1918.345 23.205 1918.515 23.375 ;
      LAYER met1 ;
        RECT 2063.185 248.100 2063.475 248.145 ;
        RECT 2199.790 248.100 2200.110 248.160 ;
        RECT 2063.185 247.960 2200.110 248.100 ;
        RECT 2063.185 247.915 2063.475 247.960 ;
        RECT 2199.790 247.900 2200.110 247.960 ;
        RECT 2059.490 247.420 2059.810 247.480 ;
        RECT 2063.185 247.420 2063.475 247.465 ;
        RECT 2059.490 247.280 2063.475 247.420 ;
        RECT 2059.490 247.220 2059.810 247.280 ;
        RECT 2063.185 247.235 2063.475 247.280 ;
        RECT 2028.685 27.440 2028.975 27.485 ;
        RECT 2059.490 27.440 2059.810 27.500 ;
        RECT 2028.685 27.300 2059.810 27.440 ;
        RECT 2028.685 27.255 2028.975 27.300 ;
        RECT 2059.490 27.240 2059.810 27.300 ;
        RECT 1628.485 24.380 1628.775 24.425 ;
        RECT 1676.325 24.380 1676.615 24.425 ;
        RECT 1628.485 24.240 1676.615 24.380 ;
        RECT 1628.485 24.195 1628.775 24.240 ;
        RECT 1676.325 24.195 1676.615 24.240 ;
        RECT 401.205 24.040 401.495 24.085 ;
        RECT 651.445 24.040 651.735 24.085 ;
        RECT 662.485 24.040 662.775 24.085 ;
        RECT 800.485 24.040 800.775 24.085 ;
        RECT 401.205 23.900 420.740 24.040 ;
        RECT 401.205 23.855 401.495 23.900 ;
        RECT 335.870 23.700 336.190 23.760 ;
        RECT 400.745 23.700 401.035 23.745 ;
        RECT 335.870 23.560 401.035 23.700 ;
        RECT 420.600 23.700 420.740 23.900 ;
        RECT 651.445 23.900 662.775 24.040 ;
        RECT 651.445 23.855 651.735 23.900 ;
        RECT 662.485 23.855 662.775 23.900 ;
        RECT 758.700 23.900 800.775 24.040 ;
        RECT 448.125 23.700 448.415 23.745 ;
        RECT 420.600 23.560 448.415 23.700 ;
        RECT 335.870 23.500 336.190 23.560 ;
        RECT 400.745 23.515 401.035 23.560 ;
        RECT 448.125 23.515 448.415 23.560 ;
        RECT 448.585 23.700 448.875 23.745 ;
        RECT 462.385 23.700 462.675 23.745 ;
        RECT 448.585 23.560 462.675 23.700 ;
        RECT 448.585 23.515 448.875 23.560 ;
        RECT 462.385 23.515 462.675 23.560 ;
        RECT 510.225 23.700 510.515 23.745 ;
        RECT 518.045 23.700 518.335 23.745 ;
        RECT 565.410 23.700 565.730 23.760 ;
        RECT 758.700 23.700 758.840 23.900 ;
        RECT 800.485 23.855 800.775 23.900 ;
        RECT 1345.585 24.040 1345.875 24.085 ;
        RECT 1393.885 24.040 1394.175 24.085 ;
        RECT 1345.585 23.900 1394.175 24.040 ;
        RECT 1345.585 23.855 1345.875 23.900 ;
        RECT 1393.885 23.855 1394.175 23.900 ;
        RECT 1821.685 24.040 1821.975 24.085 ;
        RECT 1869.525 24.040 1869.815 24.085 ;
        RECT 1821.685 23.900 1869.815 24.040 ;
        RECT 1821.685 23.855 1821.975 23.900 ;
        RECT 1869.525 23.855 1869.815 23.900 ;
        RECT 1966.125 24.040 1966.415 24.085 ;
        RECT 2028.685 24.040 2028.975 24.085 ;
        RECT 1966.125 23.900 2028.975 24.040 ;
        RECT 1966.125 23.855 1966.415 23.900 ;
        RECT 2028.685 23.855 2028.975 23.900 ;
        RECT 510.225 23.560 517.800 23.700 ;
        RECT 510.225 23.515 510.515 23.560 ;
        RECT 517.660 23.405 517.800 23.560 ;
        RECT 518.045 23.560 565.730 23.700 ;
        RECT 518.045 23.515 518.335 23.560 ;
        RECT 565.410 23.500 565.730 23.560 ;
        RECT 734.780 23.560 758.840 23.700 ;
        RECT 848.325 23.700 848.615 23.745 ;
        RECT 1038.765 23.700 1039.055 23.745 ;
        RECT 1200.225 23.700 1200.515 23.745 ;
        RECT 848.325 23.560 849.000 23.700 ;
        RECT 517.585 23.175 517.875 23.405 ;
        RECT 566.330 23.360 566.650 23.420 ;
        RECT 651.445 23.360 651.735 23.405 ;
        RECT 734.780 23.360 734.920 23.560 ;
        RECT 848.325 23.515 848.615 23.560 ;
        RECT 848.860 23.405 849.000 23.560 ;
        RECT 1038.765 23.560 1061.980 23.700 ;
        RECT 1038.765 23.515 1039.055 23.560 ;
        RECT 566.330 23.220 651.735 23.360 ;
        RECT 566.330 23.160 566.650 23.220 ;
        RECT 651.445 23.175 651.735 23.220 ;
        RECT 710.400 23.220 734.920 23.360 ;
        RECT 710.400 23.020 710.540 23.220 ;
        RECT 848.785 23.175 849.075 23.405 ;
        RECT 1000.585 23.360 1000.875 23.405 ;
        RECT 934.880 23.220 952.500 23.360 ;
        RECT 693.840 22.880 710.540 23.020 ;
        RECT 800.485 23.020 800.775 23.065 ;
        RECT 848.325 23.020 848.615 23.065 ;
        RECT 800.485 22.880 848.615 23.020 ;
        RECT 462.385 22.680 462.675 22.725 ;
        RECT 510.225 22.680 510.515 22.725 ;
        RECT 462.385 22.540 510.515 22.680 ;
        RECT 462.385 22.495 462.675 22.540 ;
        RECT 510.225 22.495 510.515 22.540 ;
        RECT 662.485 22.680 662.775 22.725 ;
        RECT 693.840 22.680 693.980 22.880 ;
        RECT 800.485 22.835 800.775 22.880 ;
        RECT 848.325 22.835 848.615 22.880 ;
        RECT 662.485 22.540 693.980 22.680 ;
        RECT 848.785 22.680 849.075 22.725 ;
        RECT 934.880 22.680 935.020 23.220 ;
        RECT 952.360 23.020 952.500 23.220 ;
        RECT 1000.200 23.220 1000.875 23.360 ;
        RECT 1061.840 23.360 1061.980 23.560 ;
        RECT 1077.020 23.560 1111.200 23.700 ;
        RECT 1077.020 23.360 1077.160 23.560 ;
        RECT 1061.840 23.220 1077.160 23.360 ;
        RECT 1111.060 23.360 1111.200 23.560 ;
        RECT 1135.900 23.560 1200.515 23.700 ;
        RECT 1135.900 23.360 1136.040 23.560 ;
        RECT 1200.225 23.515 1200.515 23.560 ;
        RECT 1441.725 23.700 1442.015 23.745 ;
        RECT 1442.170 23.700 1442.490 23.760 ;
        RECT 1441.725 23.560 1442.490 23.700 ;
        RECT 1441.725 23.515 1442.015 23.560 ;
        RECT 1442.170 23.500 1442.490 23.560 ;
        RECT 1497.460 23.560 1545.440 23.700 ;
        RECT 1242.085 23.360 1242.375 23.405 ;
        RECT 1111.060 23.220 1136.040 23.360 ;
        RECT 1200.300 23.220 1242.375 23.360 ;
        RECT 1000.200 23.020 1000.340 23.220 ;
        RECT 1000.585 23.175 1000.875 23.220 ;
        RECT 1200.300 23.065 1200.440 23.220 ;
        RECT 1242.085 23.175 1242.375 23.220 ;
        RECT 1289.925 23.360 1290.215 23.405 ;
        RECT 1297.285 23.360 1297.575 23.405 ;
        RECT 1289.925 23.220 1297.575 23.360 ;
        RECT 1289.925 23.175 1290.215 23.220 ;
        RECT 1297.285 23.175 1297.575 23.220 ;
        RECT 1442.630 23.360 1442.950 23.420 ;
        RECT 1497.460 23.360 1497.600 23.560 ;
        RECT 1442.630 23.220 1497.600 23.360 ;
        RECT 1545.300 23.360 1545.440 23.560 ;
        RECT 1676.325 23.515 1676.615 23.745 ;
        RECT 1724.625 23.700 1724.915 23.745 ;
        RECT 1731.525 23.700 1731.815 23.745 ;
        RECT 1724.625 23.560 1731.815 23.700 ;
        RECT 1724.625 23.515 1724.915 23.560 ;
        RECT 1731.525 23.515 1731.815 23.560 ;
        RECT 1731.985 23.700 1732.275 23.745 ;
        RECT 1786.725 23.700 1787.015 23.745 ;
        RECT 1731.985 23.560 1787.015 23.700 ;
        RECT 1731.985 23.515 1732.275 23.560 ;
        RECT 1786.725 23.515 1787.015 23.560 ;
        RECT 1607.325 23.360 1607.615 23.405 ;
        RECT 1545.300 23.220 1607.615 23.360 ;
        RECT 1442.630 23.160 1442.950 23.220 ;
        RECT 1607.325 23.175 1607.615 23.220 ;
        RECT 1607.785 23.360 1608.075 23.405 ;
        RECT 1628.485 23.360 1628.775 23.405 ;
        RECT 1607.785 23.220 1628.775 23.360 ;
        RECT 1676.400 23.360 1676.540 23.515 ;
        RECT 1676.785 23.360 1677.075 23.405 ;
        RECT 1676.400 23.220 1677.075 23.360 ;
        RECT 1607.785 23.175 1608.075 23.220 ;
        RECT 1628.485 23.175 1628.775 23.220 ;
        RECT 1676.785 23.175 1677.075 23.220 ;
        RECT 1787.185 23.360 1787.475 23.405 ;
        RECT 1821.685 23.360 1821.975 23.405 ;
        RECT 1787.185 23.220 1821.975 23.360 ;
        RECT 1787.185 23.175 1787.475 23.220 ;
        RECT 1821.685 23.175 1821.975 23.220 ;
        RECT 1869.525 23.360 1869.815 23.405 ;
        RECT 1918.285 23.360 1918.575 23.405 ;
        RECT 1869.525 23.220 1918.575 23.360 ;
        RECT 1869.525 23.175 1869.815 23.220 ;
        RECT 1918.285 23.175 1918.575 23.220 ;
        RECT 952.360 22.880 1000.340 23.020 ;
        RECT 1200.225 22.835 1200.515 23.065 ;
        RECT 1313.000 22.880 1345.800 23.020 ;
        RECT 848.785 22.540 935.020 22.680 ;
        RECT 1000.585 22.680 1000.875 22.725 ;
        RECT 1038.765 22.680 1039.055 22.725 ;
        RECT 1000.585 22.540 1039.055 22.680 ;
        RECT 662.485 22.495 662.775 22.540 ;
        RECT 848.785 22.495 849.075 22.540 ;
        RECT 1000.585 22.495 1000.875 22.540 ;
        RECT 1038.765 22.495 1039.055 22.540 ;
        RECT 1242.085 22.680 1242.375 22.725 ;
        RECT 1289.925 22.680 1290.215 22.725 ;
        RECT 1242.085 22.540 1290.215 22.680 ;
        RECT 1242.085 22.495 1242.375 22.540 ;
        RECT 1289.925 22.495 1290.215 22.540 ;
        RECT 1297.285 22.680 1297.575 22.725 ;
        RECT 1313.000 22.680 1313.140 22.880 ;
        RECT 1345.660 22.725 1345.800 22.880 ;
        RECT 1297.285 22.540 1313.140 22.680 ;
        RECT 1297.285 22.495 1297.575 22.540 ;
        RECT 1345.585 22.495 1345.875 22.725 ;
        RECT 1393.885 22.680 1394.175 22.725 ;
        RECT 1441.725 22.680 1442.015 22.725 ;
        RECT 1393.885 22.540 1442.015 22.680 ;
        RECT 1393.885 22.495 1394.175 22.540 ;
        RECT 1441.725 22.495 1442.015 22.540 ;
        RECT 1676.785 22.680 1677.075 22.725 ;
        RECT 1724.625 22.680 1724.915 22.725 ;
        RECT 1676.785 22.540 1724.915 22.680 ;
        RECT 1676.785 22.495 1677.075 22.540 ;
        RECT 1724.625 22.495 1724.915 22.540 ;
        RECT 1918.285 22.680 1918.575 22.725 ;
        RECT 1966.125 22.680 1966.415 22.725 ;
        RECT 1918.285 22.540 1966.415 22.680 ;
        RECT 1918.285 22.495 1918.575 22.540 ;
        RECT 1966.125 22.495 1966.415 22.540 ;
      LAYER via ;
        RECT 2199.820 247.900 2200.080 248.160 ;
        RECT 2059.520 247.220 2059.780 247.480 ;
        RECT 2059.520 27.240 2059.780 27.500 ;
        RECT 335.900 23.500 336.160 23.760 ;
        RECT 565.440 23.500 565.700 23.760 ;
        RECT 566.360 23.160 566.620 23.420 ;
        RECT 1442.200 23.500 1442.460 23.760 ;
        RECT 1442.660 23.160 1442.920 23.420 ;
      LAYER met2 ;
        RECT 2199.770 260.000 2200.050 264.000 ;
        RECT 2199.880 248.190 2200.020 260.000 ;
        RECT 2199.820 247.870 2200.080 248.190 ;
        RECT 2059.520 247.190 2059.780 247.510 ;
        RECT 2059.580 27.530 2059.720 247.190 ;
        RECT 2059.520 27.210 2059.780 27.530 ;
        RECT 565.500 24.070 566.560 24.210 ;
        RECT 565.500 23.790 565.640 24.070 ;
        RECT 335.900 23.470 336.160 23.790 ;
        RECT 565.440 23.470 565.700 23.790 ;
        RECT 335.960 2.400 336.100 23.470 ;
        RECT 566.420 23.450 566.560 24.070 ;
        RECT 1442.200 23.530 1442.460 23.790 ;
        RECT 1442.200 23.470 1442.860 23.530 ;
        RECT 1442.260 23.450 1442.860 23.470 ;
        RECT 566.360 23.130 566.620 23.450 ;
        RECT 1442.260 23.390 1442.920 23.450 ;
        RECT 1442.660 23.130 1442.920 23.390 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 352.505 186.405 352.675 234.515 ;
        RECT 352.505 48.365 352.675 137.955 ;
      LAYER mcon ;
        RECT 352.505 234.345 352.675 234.515 ;
        RECT 352.505 137.785 352.675 137.955 ;
      LAYER met1 ;
        RECT 219.490 3270.700 219.810 3270.760 ;
        RECT 418.670 3270.700 418.990 3270.760 ;
        RECT 219.490 3270.560 418.990 3270.700 ;
        RECT 219.490 3270.500 219.810 3270.560 ;
        RECT 418.670 3270.500 418.990 3270.560 ;
        RECT 219.490 260.680 219.810 260.740 ;
        RECT 352.430 260.680 352.750 260.740 ;
        RECT 219.490 260.540 352.750 260.680 ;
        RECT 219.490 260.480 219.810 260.540 ;
        RECT 352.430 260.480 352.750 260.540 ;
        RECT 352.430 234.500 352.750 234.560 ;
        RECT 352.235 234.360 352.750 234.500 ;
        RECT 352.430 234.300 352.750 234.360 ;
        RECT 352.430 186.560 352.750 186.620 ;
        RECT 352.235 186.420 352.750 186.560 ;
        RECT 352.430 186.360 352.750 186.420 ;
        RECT 352.430 137.940 352.750 138.000 ;
        RECT 352.235 137.800 352.750 137.940 ;
        RECT 352.430 137.740 352.750 137.800 ;
        RECT 352.445 48.520 352.735 48.565 ;
        RECT 353.350 48.520 353.670 48.580 ;
        RECT 352.445 48.380 353.670 48.520 ;
        RECT 352.445 48.335 352.735 48.380 ;
        RECT 353.350 48.320 353.670 48.380 ;
      LAYER via ;
        RECT 219.520 3270.500 219.780 3270.760 ;
        RECT 418.700 3270.500 418.960 3270.760 ;
        RECT 219.520 260.480 219.780 260.740 ;
        RECT 352.460 260.480 352.720 260.740 ;
        RECT 352.460 234.300 352.720 234.560 ;
        RECT 352.460 186.360 352.720 186.620 ;
        RECT 352.460 137.740 352.720 138.000 ;
        RECT 353.380 48.320 353.640 48.580 ;
      LAYER met2 ;
        RECT 219.520 3270.470 219.780 3270.790 ;
        RECT 418.700 3270.470 418.960 3270.790 ;
        RECT 219.580 260.770 219.720 3270.470 ;
        RECT 418.760 3260.000 418.900 3270.470 ;
        RECT 418.650 3256.000 418.930 3260.000 ;
        RECT 219.520 260.450 219.780 260.770 ;
        RECT 352.460 260.450 352.720 260.770 ;
        RECT 352.520 234.590 352.660 260.450 ;
        RECT 352.460 234.270 352.720 234.590 ;
        RECT 352.460 186.330 352.720 186.650 ;
        RECT 352.520 138.030 352.660 186.330 ;
        RECT 352.460 137.710 352.720 138.030 ;
        RECT 353.380 48.290 353.640 48.610 ;
        RECT 353.440 2.400 353.580 48.290 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 371.290 39.000 371.610 39.060 ;
        RECT 1435.730 39.000 1436.050 39.060 ;
        RECT 371.290 38.860 1436.050 39.000 ;
        RECT 371.290 38.800 371.610 38.860 ;
        RECT 1435.730 38.800 1436.050 38.860 ;
      LAYER via ;
        RECT 371.320 38.800 371.580 39.060 ;
        RECT 1435.760 38.800 1436.020 39.060 ;
      LAYER met2 ;
        RECT 1441.690 260.170 1441.970 264.000 ;
        RECT 1435.820 260.030 1441.970 260.170 ;
        RECT 1435.820 39.090 1435.960 260.030 ;
        RECT 1441.690 260.000 1441.970 260.030 ;
        RECT 371.320 38.770 371.580 39.090 ;
        RECT 1435.760 38.770 1436.020 39.090 ;
        RECT 371.380 2.400 371.520 38.770 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 370.445 16.065 370.615 19.635 ;
      LAYER mcon ;
        RECT 370.445 19.465 370.615 19.635 ;
      LAYER met1 ;
        RECT 224.090 1635.640 224.410 1635.700 ;
        RECT 296.770 1635.640 297.090 1635.700 ;
        RECT 224.090 1635.500 297.090 1635.640 ;
        RECT 224.090 1635.440 224.410 1635.500 ;
        RECT 296.770 1635.440 297.090 1635.500 ;
        RECT 224.090 19.620 224.410 19.680 ;
        RECT 370.385 19.620 370.675 19.665 ;
        RECT 224.090 19.480 370.675 19.620 ;
        RECT 224.090 19.420 224.410 19.480 ;
        RECT 370.385 19.435 370.675 19.480 ;
        RECT 370.385 16.220 370.675 16.265 ;
        RECT 389.230 16.220 389.550 16.280 ;
        RECT 370.385 16.080 389.550 16.220 ;
        RECT 370.385 16.035 370.675 16.080 ;
        RECT 389.230 16.020 389.550 16.080 ;
      LAYER via ;
        RECT 224.120 1635.440 224.380 1635.700 ;
        RECT 296.800 1635.440 297.060 1635.700 ;
        RECT 224.120 19.420 224.380 19.680 ;
        RECT 389.260 16.020 389.520 16.280 ;
      LAYER met2 ;
        RECT 296.790 1637.595 297.070 1637.965 ;
        RECT 296.860 1635.730 297.000 1637.595 ;
        RECT 224.120 1635.410 224.380 1635.730 ;
        RECT 296.800 1635.410 297.060 1635.730 ;
        RECT 224.180 19.710 224.320 1635.410 ;
        RECT 224.120 19.390 224.380 19.710 ;
        RECT 389.260 15.990 389.520 16.310 ;
        RECT 389.320 2.400 389.460 15.990 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 296.790 1637.640 297.070 1637.920 ;
      LAYER met3 ;
        RECT 296.765 1637.930 297.095 1637.945 ;
        RECT 310.000 1637.930 314.000 1638.320 ;
        RECT 296.765 1637.720 314.000 1637.930 ;
        RECT 296.765 1637.630 310.500 1637.720 ;
        RECT 296.765 1637.615 297.095 1637.630 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1791.310 3273.760 1791.630 3273.820 ;
        RECT 2363.550 3273.760 2363.870 3273.820 ;
        RECT 1791.310 3273.620 2363.870 3273.760 ;
        RECT 1791.310 3273.560 1791.630 3273.620 ;
        RECT 2363.550 3273.560 2363.870 3273.620 ;
      LAYER via ;
        RECT 1791.340 3273.560 1791.600 3273.820 ;
        RECT 2363.580 3273.560 2363.840 3273.820 ;
      LAYER met2 ;
        RECT 1791.340 3273.530 1791.600 3273.850 ;
        RECT 2363.580 3273.530 2363.840 3273.850 ;
        RECT 1791.400 3261.125 1791.540 3273.530 ;
        RECT 1791.330 3260.755 1791.610 3261.125 ;
        RECT 2363.640 3260.000 2363.780 3273.530 ;
        RECT 2363.530 3256.000 2363.810 3260.000 ;
        RECT 411.790 96.035 412.070 96.405 ;
        RECT 411.860 48.805 412.000 96.035 ;
        RECT 411.790 48.435 412.070 48.805 ;
        RECT 407.190 17.155 407.470 17.525 ;
        RECT 407.260 2.400 407.400 17.155 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 1791.330 3260.800 1791.610 3261.080 ;
        RECT 411.790 96.080 412.070 96.360 ;
        RECT 411.790 48.480 412.070 48.760 ;
        RECT 407.190 17.200 407.470 17.480 ;
      LAYER met3 ;
        RECT 425.310 3261.090 425.690 3261.100 ;
        RECT 1791.305 3261.090 1791.635 3261.105 ;
        RECT 425.310 3260.790 1791.635 3261.090 ;
        RECT 425.310 3260.780 425.690 3260.790 ;
        RECT 1791.305 3260.775 1791.635 3260.790 ;
        RECT 411.765 96.370 412.095 96.385 ;
        RECT 412.430 96.370 412.810 96.380 ;
        RECT 411.765 96.070 412.810 96.370 ;
        RECT 411.765 96.055 412.095 96.070 ;
        RECT 412.430 96.060 412.810 96.070 ;
        RECT 411.765 48.780 412.095 48.785 ;
        RECT 411.510 48.770 412.095 48.780 ;
        RECT 411.310 48.470 412.095 48.770 ;
        RECT 411.510 48.460 412.095 48.470 ;
        RECT 411.765 48.455 412.095 48.460 ;
        RECT 407.165 17.490 407.495 17.505 ;
        RECT 411.510 17.490 411.890 17.500 ;
        RECT 407.165 17.190 411.890 17.490 ;
        RECT 407.165 17.175 407.495 17.190 ;
        RECT 411.510 17.180 411.890 17.190 ;
      LAYER via3 ;
        RECT 425.340 3260.780 425.660 3261.100 ;
        RECT 412.460 96.060 412.780 96.380 ;
        RECT 411.540 48.460 411.860 48.780 ;
        RECT 411.540 17.180 411.860 17.500 ;
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 3260.000 367.020 3528.900 ;
        RECT 425.335 3260.775 425.665 3261.105 ;
        RECT 425.350 3249.290 425.650 3260.775 ;
        RECT 544.020 3260.000 547.020 3528.900 ;
        RECT 724.020 3260.000 727.020 3528.900 ;
        RECT 904.020 3260.000 907.020 3528.900 ;
        RECT 1084.020 3260.000 1087.020 3528.900 ;
        RECT 1264.020 3260.000 1267.020 3528.900 ;
        RECT 1444.020 3260.000 1447.020 3528.900 ;
        RECT 1624.020 3260.000 1627.020 3528.900 ;
        RECT 1804.020 3260.000 1807.020 3528.900 ;
        RECT 1984.020 3260.000 1987.020 3528.900 ;
        RECT 2164.020 3260.000 2167.020 3528.900 ;
        RECT 2344.020 3260.000 2347.020 3528.900 ;
        RECT 2524.020 3260.000 2527.020 3528.900 ;
        RECT 424.910 3248.110 426.090 3249.290 ;
        RECT 407.840 3228.890 409.440 3246.800 ;
        RECT 407.840 3227.710 409.530 3228.890 ;
        RECT 407.840 2970.490 409.440 3227.710 ;
        RECT 407.430 2969.310 409.440 2970.490 ;
        RECT 407.840 2960.290 409.440 2969.310 ;
        RECT 407.840 2959.110 409.530 2960.290 ;
        RECT 407.840 2797.090 409.440 2959.110 ;
        RECT 407.430 2795.910 409.440 2797.090 ;
        RECT 407.840 2776.690 409.440 2795.910 ;
        RECT 407.840 2775.510 409.530 2776.690 ;
        RECT 407.840 2606.690 409.440 2775.510 ;
        RECT 407.840 2605.510 409.530 2606.690 ;
        RECT 407.840 2599.890 409.440 2605.510 ;
        RECT 407.430 2598.710 409.440 2599.890 ;
        RECT 407.840 2525.090 409.440 2598.710 ;
        RECT 407.840 2523.910 409.530 2525.090 ;
        RECT 407.840 2498.390 409.440 2523.910 ;
        RECT 407.840 2497.210 409.530 2498.390 ;
        RECT 407.840 2256.490 409.440 2497.210 ;
        RECT 407.840 2255.310 409.530 2256.490 ;
        RECT 407.840 2236.090 409.440 2255.310 ;
        RECT 407.430 2234.910 409.440 2236.090 ;
        RECT 407.840 2168.090 409.440 2234.910 ;
        RECT 407.430 2166.910 409.440 2168.090 ;
        RECT 407.840 2146.490 409.440 2166.910 ;
        RECT 407.840 2145.310 409.530 2146.490 ;
        RECT 407.840 2072.890 409.440 2145.310 ;
        RECT 407.430 2071.710 409.440 2072.890 ;
        RECT 407.840 2059.290 409.440 2071.710 ;
        RECT 407.430 2058.110 409.440 2059.290 ;
        RECT 407.840 1797.490 409.440 2058.110 ;
        RECT 407.430 1796.310 409.440 1797.490 ;
        RECT 407.840 1787.290 409.440 1796.310 ;
        RECT 407.430 1786.110 409.440 1787.290 ;
        RECT 407.840 1256.890 409.440 1786.110 ;
        RECT 407.840 1255.710 409.530 1256.890 ;
        RECT 407.840 1250.090 409.440 1255.710 ;
        RECT 407.430 1248.910 409.440 1250.090 ;
        RECT 407.840 988.290 409.440 1248.910 ;
        RECT 407.840 987.110 409.530 988.290 ;
        RECT 407.840 971.290 409.440 987.110 ;
        RECT 407.430 970.110 409.440 971.290 ;
        RECT 407.840 631.290 409.440 970.110 ;
        RECT 407.430 630.110 409.440 631.290 ;
        RECT 407.840 621.090 409.440 630.110 ;
        RECT 407.430 619.910 409.440 621.090 ;
        RECT 407.840 539.490 409.440 619.910 ;
        RECT 407.840 538.310 409.530 539.490 ;
        RECT 407.840 529.290 409.440 538.310 ;
        RECT 407.430 528.110 409.440 529.290 ;
        RECT 407.840 359.290 409.440 528.110 ;
        RECT 407.840 358.110 409.530 359.290 ;
        RECT 407.840 338.890 409.440 358.110 ;
        RECT 407.840 337.710 409.530 338.890 ;
        RECT 407.840 270.640 409.440 337.710 ;
        RECT 364.020 -9.220 367.020 260.000 ;
        RECT 408.790 256.850 409.090 270.640 ;
        RECT 408.790 256.550 410.930 256.850 ;
        RECT 410.630 158.250 410.930 256.550 ;
        RECT 410.630 157.950 411.850 158.250 ;
        RECT 411.550 110.650 411.850 157.950 ;
        RECT 411.550 110.350 412.770 110.650 ;
        RECT 412.470 96.385 412.770 110.350 ;
        RECT 412.455 96.055 412.785 96.385 ;
        RECT 411.535 48.455 411.865 48.785 ;
        RECT 411.550 17.505 411.850 48.455 ;
        RECT 411.535 17.175 411.865 17.505 ;
        RECT 544.020 -9.220 547.020 260.000 ;
        RECT 724.020 -9.220 727.020 260.000 ;
        RECT 904.020 -9.220 907.020 260.000 ;
        RECT 1084.020 -9.220 1087.020 260.000 ;
        RECT 1264.020 -9.220 1267.020 260.000 ;
        RECT 1444.020 -9.220 1447.020 260.000 ;
        RECT 1624.020 -9.220 1627.020 260.000 ;
        RECT 1804.020 -9.220 1807.020 260.000 ;
        RECT 1984.020 -9.220 1987.020 260.000 ;
        RECT 2164.020 -9.220 2167.020 260.000 ;
        RECT 2344.020 -9.220 2347.020 260.000 ;
        RECT 2524.020 -9.220 2527.020 260.000 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 408.350 3227.710 409.530 3228.890 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 408.350 2959.110 409.530 2960.290 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 408.350 2775.510 409.530 2776.690 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 408.350 2605.510 409.530 2606.690 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 408.350 2523.910 409.530 2525.090 ;
        RECT 408.350 2497.210 409.530 2498.390 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 408.350 2255.310 409.530 2256.490 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 408.350 2145.310 409.530 2146.490 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 408.350 1255.710 409.530 1256.890 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 408.350 987.110 409.530 988.290 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 408.350 538.310 409.530 539.490 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 408.350 358.110 409.530 359.290 ;
        RECT 408.350 337.710 409.530 338.890 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 424.700 3246.100 426.300 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT 409.980 3244.500 426.300 3246.100 ;
        RECT 409.980 3229.100 411.580 3244.500 ;
        RECT 408.140 3227.500 411.580 3229.100 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT 407.220 2969.100 409.740 2970.700 ;
        RECT 408.140 2958.900 409.740 2969.100 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT 407.220 2776.900 408.820 2797.300 ;
        RECT 407.220 2775.300 409.740 2776.900 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT 408.140 2605.300 411.580 2606.900 ;
        RECT 409.980 2600.100 411.580 2605.300 ;
        RECT 407.220 2598.500 411.580 2600.100 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT 408.140 2523.700 411.580 2525.300 ;
        RECT 409.980 2508.300 411.580 2523.700 ;
        RECT 408.140 2506.700 411.580 2508.300 ;
        RECT 408.140 2497.000 409.740 2506.700 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT 406.300 2255.100 409.740 2256.700 ;
        RECT 406.300 2236.300 407.900 2255.100 ;
        RECT 406.300 2234.700 408.820 2236.300 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT 407.220 2167.400 408.820 2168.300 ;
        RECT 406.300 2165.800 408.820 2167.400 ;
        RECT 406.300 2161.500 407.900 2165.800 ;
        RECT 403.540 2159.900 407.900 2161.500 ;
        RECT 403.540 2147.900 405.140 2159.900 ;
        RECT 403.540 2146.300 407.900 2147.900 ;
        RECT 406.300 2144.500 407.900 2146.300 ;
        RECT 408.140 2144.500 409.740 2146.700 ;
        RECT 406.300 2142.900 409.740 2144.500 ;
        RECT 407.220 2057.900 408.820 2073.100 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT 407.220 1796.100 409.740 1797.700 ;
        RECT 408.140 1787.500 409.740 1796.100 ;
        RECT 407.220 1785.900 409.740 1787.500 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT 406.300 1255.500 409.740 1257.100 ;
        RECT 406.300 1250.300 407.900 1255.500 ;
        RECT 406.300 1248.700 408.820 1250.300 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT 408.140 986.900 411.580 988.500 ;
        RECT 409.980 985.100 411.580 986.900 ;
        RECT 407.220 983.500 411.580 985.100 ;
        RECT 407.220 969.900 408.820 983.500 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT 407.220 629.900 410.660 631.500 ;
        RECT 409.060 621.300 410.660 629.900 ;
        RECT 407.220 619.700 410.660 621.300 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT 407.220 538.100 409.740 539.700 ;
        RECT 407.220 527.900 408.820 538.100 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT 406.300 357.900 409.740 359.500 ;
        RECT 406.300 345.900 407.900 357.900 ;
        RECT 406.300 344.300 409.740 345.900 ;
        RECT 408.140 337.500 409.740 344.300 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.610 107.000 68.930 107.060 ;
        RECT 1669.870 107.000 1670.190 107.060 ;
        RECT 68.610 106.860 1670.190 107.000 ;
        RECT 68.610 106.800 68.930 106.860 ;
        RECT 1669.870 106.800 1670.190 106.860 ;
      LAYER via ;
        RECT 68.640 106.800 68.900 107.060 ;
        RECT 1669.900 106.800 1670.160 107.060 ;
      LAYER met2 ;
        RECT 1670.770 260.170 1671.050 264.000 ;
        RECT 1669.960 260.030 1671.050 260.170 ;
        RECT 1669.960 107.090 1670.100 260.030 ;
        RECT 1670.770 260.000 1671.050 260.030 ;
        RECT 68.640 106.770 68.900 107.090 ;
        RECT 1669.900 106.770 1670.160 107.090 ;
        RECT 68.700 17.410 68.840 106.770 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2349.770 3264.835 2350.050 3265.205 ;
        RECT 2349.840 3260.000 2349.980 3264.835 ;
        RECT 2349.730 3256.000 2350.010 3260.000 ;
        RECT 421.910 240.195 422.190 240.565 ;
        RECT 421.980 194.325 422.120 240.195 ;
        RECT 421.910 193.955 422.190 194.325 ;
        RECT 424.670 17.155 424.950 17.525 ;
        RECT 424.740 2.400 424.880 17.155 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 2349.770 3264.880 2350.050 3265.160 ;
        RECT 421.910 240.240 422.190 240.520 ;
        RECT 421.910 194.000 422.190 194.280 ;
        RECT 424.670 17.200 424.950 17.480 ;
      LAYER met3 ;
        RECT 259.710 3265.170 260.090 3265.180 ;
        RECT 2349.745 3265.170 2350.075 3265.185 ;
        RECT 259.710 3264.870 2350.075 3265.170 ;
        RECT 259.710 3264.860 260.090 3264.870 ;
        RECT 2349.745 3264.855 2350.075 3264.870 ;
        RECT 259.710 1800.820 260.090 1801.140 ;
        RECT 259.750 1799.780 260.050 1800.820 ;
        RECT 259.710 1799.460 260.090 1799.780 ;
        RECT 259.710 290.540 260.090 290.860 ;
        RECT 259.750 290.180 260.050 290.540 ;
        RECT 259.710 289.860 260.090 290.180 ;
        RECT 421.885 240.530 422.215 240.545 ;
        RECT 422.550 240.530 422.930 240.540 ;
        RECT 421.885 240.230 422.930 240.530 ;
        RECT 421.885 240.215 422.215 240.230 ;
        RECT 422.550 240.220 422.930 240.230 ;
        RECT 421.885 194.290 422.215 194.305 ;
        RECT 421.670 193.975 422.215 194.290 ;
        RECT 421.670 193.620 421.970 193.975 ;
        RECT 421.630 193.300 422.010 193.620 ;
        RECT 421.630 17.490 422.010 17.500 ;
        RECT 424.645 17.490 424.975 17.505 ;
        RECT 421.630 17.190 424.975 17.490 ;
        RECT 421.630 17.180 422.010 17.190 ;
        RECT 424.645 17.175 424.975 17.190 ;
      LAYER via3 ;
        RECT 259.740 3264.860 260.060 3265.180 ;
        RECT 259.740 1800.820 260.060 1801.140 ;
        RECT 259.740 1799.460 260.060 1799.780 ;
        RECT 259.740 290.540 260.060 290.860 ;
        RECT 259.740 289.860 260.060 290.180 ;
        RECT 422.580 240.220 422.900 240.540 ;
        RECT 421.660 193.300 421.980 193.620 ;
        RECT 421.660 17.180 421.980 17.500 ;
      LAYER met4 ;
        RECT 259.735 3264.855 260.065 3265.185 ;
        RECT 259.750 1801.145 260.050 3264.855 ;
        RECT 259.735 1800.815 260.065 1801.145 ;
        RECT 259.735 1799.455 260.065 1799.785 ;
        RECT 259.750 290.865 260.050 1799.455 ;
        RECT 259.735 290.535 260.065 290.865 ;
        RECT 259.735 289.855 260.065 290.185 ;
        RECT 259.750 257.290 260.050 289.855 ;
        RECT 259.310 256.110 260.490 257.290 ;
        RECT 422.150 256.110 423.330 257.290 ;
        RECT 422.590 240.545 422.890 256.110 ;
        RECT 422.575 240.215 422.905 240.545 ;
        RECT 421.655 193.295 421.985 193.625 ;
        RECT 421.670 17.505 421.970 193.295 ;
        RECT 421.655 17.175 421.985 17.505 ;
      LAYER met5 ;
        RECT 259.100 255.900 423.540 257.500 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 210.360 448.430 210.420 ;
        RECT 2698.430 210.360 2698.750 210.420 ;
        RECT 448.110 210.220 2698.750 210.360 ;
        RECT 448.110 210.160 448.430 210.220 ;
        RECT 2698.430 210.160 2698.750 210.220 ;
        RECT 442.590 19.620 442.910 19.680 ;
        RECT 448.110 19.620 448.430 19.680 ;
        RECT 442.590 19.480 448.430 19.620 ;
        RECT 442.590 19.420 442.910 19.480 ;
        RECT 448.110 19.420 448.430 19.480 ;
      LAYER via ;
        RECT 448.140 210.160 448.400 210.420 ;
        RECT 2698.460 210.160 2698.720 210.420 ;
        RECT 442.620 19.420 442.880 19.680 ;
        RECT 448.140 19.420 448.400 19.680 ;
      LAYER met2 ;
        RECT 2592.650 3270.955 2592.930 3271.325 ;
        RECT 2698.450 3270.955 2698.730 3271.325 ;
        RECT 2592.720 3260.000 2592.860 3270.955 ;
        RECT 2592.610 3256.000 2592.890 3260.000 ;
        RECT 2698.520 210.450 2698.660 3270.955 ;
        RECT 448.140 210.130 448.400 210.450 ;
        RECT 2698.460 210.130 2698.720 210.450 ;
        RECT 448.200 19.710 448.340 210.130 ;
        RECT 442.620 19.390 442.880 19.710 ;
        RECT 448.140 19.390 448.400 19.710 ;
        RECT 442.680 2.400 442.820 19.390 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 2592.650 3271.000 2592.930 3271.280 ;
        RECT 2698.450 3271.000 2698.730 3271.280 ;
      LAYER met3 ;
        RECT 2592.625 3271.290 2592.955 3271.305 ;
        RECT 2698.425 3271.290 2698.755 3271.305 ;
        RECT 2592.625 3270.990 2698.755 3271.290 ;
        RECT 2592.625 3270.975 2592.955 3270.990 ;
        RECT 2698.425 3270.975 2698.755 3270.990 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 456.925 144.925 457.095 234.515 ;
        RECT 456.465 48.365 456.635 96.475 ;
      LAYER mcon ;
        RECT 456.925 234.345 457.095 234.515 ;
        RECT 456.465 96.305 456.635 96.475 ;
      LAYER met1 ;
        RECT 456.390 240.960 456.710 241.020 ;
        RECT 457.310 240.960 457.630 241.020 ;
        RECT 456.390 240.820 457.630 240.960 ;
        RECT 456.390 240.760 456.710 240.820 ;
        RECT 457.310 240.760 457.630 240.820 ;
        RECT 456.865 234.500 457.155 234.545 ;
        RECT 457.310 234.500 457.630 234.560 ;
        RECT 456.865 234.360 457.630 234.500 ;
        RECT 456.865 234.315 457.155 234.360 ;
        RECT 457.310 234.300 457.630 234.360 ;
        RECT 456.850 145.080 457.170 145.140 ;
        RECT 456.655 144.940 457.170 145.080 ;
        RECT 456.850 144.880 457.170 144.940 ;
        RECT 456.390 96.460 456.710 96.520 ;
        RECT 456.195 96.320 456.710 96.460 ;
        RECT 456.390 96.260 456.710 96.320 ;
        RECT 456.405 48.520 456.695 48.565 ;
        RECT 456.850 48.520 457.170 48.580 ;
        RECT 456.405 48.380 457.170 48.520 ;
        RECT 456.405 48.335 456.695 48.380 ;
        RECT 456.850 48.320 457.170 48.380 ;
        RECT 456.850 19.620 457.170 19.680 ;
        RECT 460.530 19.620 460.850 19.680 ;
        RECT 456.850 19.480 460.850 19.620 ;
        RECT 456.850 19.420 457.170 19.480 ;
        RECT 460.530 19.420 460.850 19.480 ;
      LAYER via ;
        RECT 456.420 240.760 456.680 241.020 ;
        RECT 457.340 240.760 457.600 241.020 ;
        RECT 457.340 234.300 457.600 234.560 ;
        RECT 456.880 144.880 457.140 145.140 ;
        RECT 456.420 96.260 456.680 96.520 ;
        RECT 456.880 48.320 457.140 48.580 ;
        RECT 456.880 19.420 457.140 19.680 ;
        RECT 460.560 19.420 460.820 19.680 ;
      LAYER met2 ;
        RECT 2063.650 3275.715 2063.930 3276.085 ;
        RECT 2063.720 3260.000 2063.860 3275.715 ;
        RECT 2063.610 3256.000 2063.890 3260.000 ;
        RECT 258.150 2719.475 258.430 2719.845 ;
        RECT 258.220 2698.085 258.360 2719.475 ;
        RECT 258.150 2697.715 258.430 2698.085 ;
        RECT 258.150 2641.275 258.430 2641.645 ;
        RECT 258.220 2594.725 258.360 2641.275 ;
        RECT 258.150 2594.355 258.430 2594.725 ;
        RECT 258.150 2524.995 258.430 2525.365 ;
        RECT 258.220 2478.445 258.360 2524.995 ;
        RECT 258.150 2478.075 258.430 2478.445 ;
        RECT 258.150 2380.155 258.430 2380.525 ;
        RECT 258.220 2375.085 258.360 2380.155 ;
        RECT 258.150 2374.715 258.430 2375.085 ;
        RECT 259.530 2325.075 259.810 2325.445 ;
        RECT 259.600 2283.285 259.740 2325.075 ;
        RECT 259.530 2282.915 259.810 2283.285 ;
        RECT 258.150 2187.035 258.430 2187.405 ;
        RECT 258.220 2180.605 258.360 2187.035 ;
        RECT 258.150 2180.235 258.430 2180.605 ;
        RECT 259.530 2131.275 259.810 2131.645 ;
        RECT 259.600 2090.165 259.740 2131.275 ;
        RECT 259.530 2089.795 259.810 2090.165 ;
        RECT 257.690 1946.315 257.970 1946.685 ;
        RECT 257.760 1910.645 257.900 1946.315 ;
        RECT 257.690 1910.275 257.970 1910.645 ;
        RECT 258.150 1621.275 258.430 1621.645 ;
        RECT 258.220 1574.725 258.360 1621.275 ;
        RECT 258.150 1574.355 258.430 1574.725 ;
        RECT 259.990 1572.315 260.270 1572.685 ;
        RECT 260.060 1535.285 260.200 1572.315 ;
        RECT 259.990 1534.915 260.270 1535.285 ;
        RECT 258.150 1455.355 258.430 1455.725 ;
        RECT 258.220 1414.245 258.360 1455.355 ;
        RECT 258.150 1413.875 258.430 1414.245 ;
        RECT 258.150 1317.315 258.430 1317.685 ;
        RECT 258.220 1270.765 258.360 1317.315 ;
        RECT 258.150 1270.395 258.430 1270.765 ;
        RECT 257.690 1142.555 257.970 1142.925 ;
        RECT 257.760 1124.565 257.900 1142.555 ;
        RECT 257.690 1124.195 257.970 1124.565 ;
        RECT 256.310 854.915 256.590 855.285 ;
        RECT 256.380 807.685 256.520 854.915 ;
        RECT 256.310 807.315 256.590 807.685 ;
        RECT 256.310 751.555 256.590 751.925 ;
        RECT 256.380 705.005 256.520 751.555 ;
        RECT 256.310 704.635 256.590 705.005 ;
        RECT 256.310 703.275 256.590 703.645 ;
        RECT 256.380 656.725 256.520 703.275 ;
        RECT 256.310 656.355 256.590 656.725 ;
        RECT 261.370 613.515 261.650 613.885 ;
        RECT 261.440 532.285 261.580 613.515 ;
        RECT 261.370 531.915 261.650 532.285 ;
        RECT 256.310 516.955 256.590 517.325 ;
        RECT 256.380 470.405 256.520 516.955 ;
        RECT 256.310 470.035 256.590 470.405 ;
        RECT 456.410 261.275 456.690 261.645 ;
        RECT 456.480 241.050 456.620 261.275 ;
        RECT 456.420 240.730 456.680 241.050 ;
        RECT 457.340 240.730 457.600 241.050 ;
        RECT 457.400 234.590 457.540 240.730 ;
        RECT 457.340 234.270 457.600 234.590 ;
        RECT 456.880 144.850 457.140 145.170 ;
        RECT 456.940 110.570 457.080 144.850 ;
        RECT 456.480 110.430 457.080 110.570 ;
        RECT 456.480 96.550 456.620 110.430 ;
        RECT 456.420 96.230 456.680 96.550 ;
        RECT 456.880 48.290 457.140 48.610 ;
        RECT 456.940 19.710 457.080 48.290 ;
        RECT 456.880 19.390 457.140 19.710 ;
        RECT 460.560 19.390 460.820 19.710 ;
        RECT 460.620 2.400 460.760 19.390 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 2063.650 3275.760 2063.930 3276.040 ;
        RECT 258.150 2719.520 258.430 2719.800 ;
        RECT 258.150 2697.760 258.430 2698.040 ;
        RECT 258.150 2641.320 258.430 2641.600 ;
        RECT 258.150 2594.400 258.430 2594.680 ;
        RECT 258.150 2525.040 258.430 2525.320 ;
        RECT 258.150 2478.120 258.430 2478.400 ;
        RECT 258.150 2380.200 258.430 2380.480 ;
        RECT 258.150 2374.760 258.430 2375.040 ;
        RECT 259.530 2325.120 259.810 2325.400 ;
        RECT 259.530 2282.960 259.810 2283.240 ;
        RECT 258.150 2187.080 258.430 2187.360 ;
        RECT 258.150 2180.280 258.430 2180.560 ;
        RECT 259.530 2131.320 259.810 2131.600 ;
        RECT 259.530 2089.840 259.810 2090.120 ;
        RECT 257.690 1946.360 257.970 1946.640 ;
        RECT 257.690 1910.320 257.970 1910.600 ;
        RECT 258.150 1621.320 258.430 1621.600 ;
        RECT 258.150 1574.400 258.430 1574.680 ;
        RECT 259.990 1572.360 260.270 1572.640 ;
        RECT 259.990 1534.960 260.270 1535.240 ;
        RECT 258.150 1455.400 258.430 1455.680 ;
        RECT 258.150 1413.920 258.430 1414.200 ;
        RECT 258.150 1317.360 258.430 1317.640 ;
        RECT 258.150 1270.440 258.430 1270.720 ;
        RECT 257.690 1142.600 257.970 1142.880 ;
        RECT 257.690 1124.240 257.970 1124.520 ;
        RECT 256.310 854.960 256.590 855.240 ;
        RECT 256.310 807.360 256.590 807.640 ;
        RECT 256.310 751.600 256.590 751.880 ;
        RECT 256.310 704.680 256.590 704.960 ;
        RECT 256.310 703.320 256.590 703.600 ;
        RECT 256.310 656.400 256.590 656.680 ;
        RECT 261.370 613.560 261.650 613.840 ;
        RECT 261.370 531.960 261.650 532.240 ;
        RECT 256.310 517.000 256.590 517.280 ;
        RECT 256.310 470.080 256.590 470.360 ;
        RECT 456.410 261.320 456.690 261.600 ;
      LAYER met3 ;
        RECT 542.150 3276.050 542.530 3276.060 ;
        RECT 548.590 3276.050 548.970 3276.060 ;
        RECT 542.150 3275.750 548.970 3276.050 ;
        RECT 542.150 3275.740 542.530 3275.750 ;
        RECT 548.590 3275.740 548.970 3275.750 ;
        RECT 2063.625 3276.050 2063.955 3276.065 ;
        RECT 2064.750 3276.050 2065.130 3276.060 ;
        RECT 2063.625 3275.750 2065.130 3276.050 ;
        RECT 2063.625 3275.735 2063.955 3275.750 ;
        RECT 2064.750 3275.740 2065.130 3275.750 ;
        RECT 260.630 2747.690 261.010 2747.700 ;
        RECT 257.910 2747.390 261.010 2747.690 ;
        RECT 257.910 2747.020 258.210 2747.390 ;
        RECT 260.630 2747.380 261.010 2747.390 ;
        RECT 257.870 2746.700 258.250 2747.020 ;
        RECT 258.125 2719.820 258.455 2719.825 ;
        RECT 257.870 2719.810 258.455 2719.820 ;
        RECT 257.870 2719.510 258.680 2719.810 ;
        RECT 257.870 2719.500 258.455 2719.510 ;
        RECT 258.125 2719.495 258.455 2719.500 ;
        RECT 258.125 2698.060 258.455 2698.065 ;
        RECT 257.870 2698.050 258.455 2698.060 ;
        RECT 257.670 2697.750 258.455 2698.050 ;
        RECT 257.870 2697.740 258.455 2697.750 ;
        RECT 258.125 2697.735 258.455 2697.740 ;
        RECT 257.870 2641.980 258.250 2642.300 ;
        RECT 257.910 2641.625 258.210 2641.980 ;
        RECT 257.910 2641.310 258.455 2641.625 ;
        RECT 258.125 2641.295 258.455 2641.310 ;
        RECT 258.125 2594.700 258.455 2594.705 ;
        RECT 257.870 2594.690 258.455 2594.700 ;
        RECT 257.870 2594.390 258.680 2594.690 ;
        RECT 257.870 2594.380 258.455 2594.390 ;
        RECT 258.125 2594.375 258.455 2594.380 ;
        RECT 258.125 2525.340 258.455 2525.345 ;
        RECT 257.870 2525.330 258.455 2525.340 ;
        RECT 257.870 2525.030 258.680 2525.330 ;
        RECT 257.870 2525.020 258.455 2525.030 ;
        RECT 258.125 2525.015 258.455 2525.020 ;
        RECT 258.125 2478.410 258.455 2478.425 ;
        RECT 258.125 2478.110 259.130 2478.410 ;
        RECT 258.125 2478.095 258.455 2478.110 ;
        RECT 258.830 2477.060 259.130 2478.110 ;
        RECT 258.790 2476.740 259.170 2477.060 ;
        RECT 258.125 2380.490 258.455 2380.505 ;
        RECT 258.790 2380.490 259.170 2380.500 ;
        RECT 258.125 2380.190 259.170 2380.490 ;
        RECT 258.125 2380.175 258.455 2380.190 ;
        RECT 258.790 2380.180 259.170 2380.190 ;
        RECT 258.125 2375.050 258.455 2375.065 ;
        RECT 258.125 2374.750 259.130 2375.050 ;
        RECT 258.125 2374.735 258.455 2374.750 ;
        RECT 258.830 2374.380 259.130 2374.750 ;
        RECT 258.790 2374.060 259.170 2374.380 ;
        RECT 258.790 2325.410 259.170 2325.420 ;
        RECT 259.505 2325.410 259.835 2325.425 ;
        RECT 258.790 2325.110 259.835 2325.410 ;
        RECT 258.790 2325.100 259.170 2325.110 ;
        RECT 259.505 2325.095 259.835 2325.110 ;
        RECT 258.790 2283.250 259.170 2283.260 ;
        RECT 259.505 2283.250 259.835 2283.265 ;
        RECT 258.790 2282.950 259.835 2283.250 ;
        RECT 258.790 2282.940 259.170 2282.950 ;
        RECT 259.505 2282.935 259.835 2282.950 ;
        RECT 258.125 2187.370 258.455 2187.385 ;
        RECT 258.790 2187.370 259.170 2187.380 ;
        RECT 258.125 2187.070 259.170 2187.370 ;
        RECT 258.125 2187.055 258.455 2187.070 ;
        RECT 258.790 2187.060 259.170 2187.070 ;
        RECT 258.125 2180.570 258.455 2180.585 ;
        RECT 258.790 2180.570 259.170 2180.580 ;
        RECT 258.125 2180.270 259.170 2180.570 ;
        RECT 258.125 2180.255 258.455 2180.270 ;
        RECT 258.790 2180.260 259.170 2180.270 ;
        RECT 258.790 2131.610 259.170 2131.620 ;
        RECT 259.505 2131.610 259.835 2131.625 ;
        RECT 258.790 2131.310 259.835 2131.610 ;
        RECT 258.790 2131.300 259.170 2131.310 ;
        RECT 259.505 2131.295 259.835 2131.310 ;
        RECT 258.790 2090.130 259.170 2090.140 ;
        RECT 259.505 2090.130 259.835 2090.145 ;
        RECT 258.790 2089.830 259.835 2090.130 ;
        RECT 258.790 2089.820 259.170 2089.830 ;
        RECT 259.505 2089.815 259.835 2089.830 ;
        RECT 258.790 2043.890 259.170 2043.900 ;
        RECT 257.910 2043.590 259.170 2043.890 ;
        RECT 257.910 2043.220 258.210 2043.590 ;
        RECT 258.790 2043.580 259.170 2043.590 ;
        RECT 257.870 2042.900 258.250 2043.220 ;
        RECT 258.790 2001.730 259.170 2001.740 ;
        RECT 257.910 2001.430 259.170 2001.730 ;
        RECT 257.910 2000.380 258.210 2001.430 ;
        RECT 258.790 2001.420 259.170 2001.430 ;
        RECT 257.870 2000.060 258.250 2000.380 ;
        RECT 257.665 1946.660 257.995 1946.665 ;
        RECT 257.665 1946.650 258.250 1946.660 ;
        RECT 257.440 1946.350 258.250 1946.650 ;
        RECT 257.665 1946.340 258.250 1946.350 ;
        RECT 257.665 1946.335 257.995 1946.340 ;
        RECT 256.950 1910.610 257.330 1910.620 ;
        RECT 257.665 1910.610 257.995 1910.625 ;
        RECT 256.950 1910.310 257.995 1910.610 ;
        RECT 256.950 1910.300 257.330 1910.310 ;
        RECT 257.665 1910.295 257.995 1910.310 ;
        RECT 258.790 1790.930 259.170 1790.940 ;
        RECT 260.630 1790.930 261.010 1790.940 ;
        RECT 258.790 1790.630 261.010 1790.930 ;
        RECT 258.790 1790.620 259.170 1790.630 ;
        RECT 260.630 1790.620 261.010 1790.630 ;
        RECT 257.870 1703.890 258.250 1703.900 ;
        RECT 260.630 1703.890 261.010 1703.900 ;
        RECT 257.870 1703.590 261.010 1703.890 ;
        RECT 257.870 1703.580 258.250 1703.590 ;
        RECT 260.630 1703.580 261.010 1703.590 ;
        RECT 256.950 1622.970 257.330 1622.980 ;
        RECT 258.790 1622.970 259.170 1622.980 ;
        RECT 256.950 1622.670 259.170 1622.970 ;
        RECT 256.950 1622.660 257.330 1622.670 ;
        RECT 258.790 1622.660 259.170 1622.670 ;
        RECT 258.125 1621.610 258.455 1621.625 ;
        RECT 258.790 1621.610 259.170 1621.620 ;
        RECT 258.125 1621.310 259.170 1621.610 ;
        RECT 258.125 1621.295 258.455 1621.310 ;
        RECT 258.790 1621.300 259.170 1621.310 ;
        RECT 258.125 1574.690 258.455 1574.705 ;
        RECT 257.910 1574.375 258.455 1574.690 ;
        RECT 257.910 1574.020 258.210 1574.375 ;
        RECT 257.870 1573.700 258.250 1574.020 ;
        RECT 258.790 1572.650 259.170 1572.660 ;
        RECT 259.965 1572.650 260.295 1572.665 ;
        RECT 258.790 1572.350 260.295 1572.650 ;
        RECT 258.790 1572.340 259.170 1572.350 ;
        RECT 259.965 1572.335 260.295 1572.350 ;
        RECT 257.870 1535.250 258.250 1535.260 ;
        RECT 259.965 1535.250 260.295 1535.265 ;
        RECT 257.870 1534.950 260.295 1535.250 ;
        RECT 257.870 1534.940 258.250 1534.950 ;
        RECT 259.965 1534.935 260.295 1534.950 ;
        RECT 258.125 1455.690 258.455 1455.705 ;
        RECT 258.790 1455.690 259.170 1455.700 ;
        RECT 258.125 1455.390 259.170 1455.690 ;
        RECT 258.125 1455.375 258.455 1455.390 ;
        RECT 258.790 1455.380 259.170 1455.390 ;
        RECT 258.125 1414.210 258.455 1414.225 ;
        RECT 258.790 1414.210 259.170 1414.220 ;
        RECT 258.125 1413.910 259.170 1414.210 ;
        RECT 258.125 1413.895 258.455 1413.910 ;
        RECT 258.790 1413.900 259.170 1413.910 ;
        RECT 258.790 1367.290 259.170 1367.300 ;
        RECT 257.910 1366.990 259.170 1367.290 ;
        RECT 257.910 1366.620 258.210 1366.990 ;
        RECT 258.790 1366.980 259.170 1366.990 ;
        RECT 257.870 1366.300 258.250 1366.620 ;
        RECT 258.125 1317.650 258.455 1317.665 ;
        RECT 258.790 1317.650 259.170 1317.660 ;
        RECT 258.125 1317.350 259.170 1317.650 ;
        RECT 258.125 1317.335 258.455 1317.350 ;
        RECT 258.790 1317.340 259.170 1317.350 ;
        RECT 258.125 1270.730 258.455 1270.745 ;
        RECT 257.910 1270.415 258.455 1270.730 ;
        RECT 257.910 1270.060 258.210 1270.415 ;
        RECT 257.870 1269.740 258.250 1270.060 ;
        RECT 257.665 1142.900 257.995 1142.905 ;
        RECT 257.665 1142.890 258.250 1142.900 ;
        RECT 257.440 1142.590 258.250 1142.890 ;
        RECT 257.665 1142.580 258.250 1142.590 ;
        RECT 257.665 1142.575 257.995 1142.580 ;
        RECT 257.665 1124.530 257.995 1124.545 ;
        RECT 258.790 1124.530 259.170 1124.540 ;
        RECT 257.665 1124.230 259.170 1124.530 ;
        RECT 257.665 1124.215 257.995 1124.230 ;
        RECT 258.790 1124.220 259.170 1124.230 ;
        RECT 258.790 1027.970 259.170 1027.980 ;
        RECT 260.630 1027.970 261.010 1027.980 ;
        RECT 258.790 1027.670 261.010 1027.970 ;
        RECT 258.790 1027.660 259.170 1027.670 ;
        RECT 260.630 1027.660 261.010 1027.670 ;
        RECT 257.870 917.130 258.250 917.140 ;
        RECT 260.630 917.130 261.010 917.140 ;
        RECT 257.870 916.830 261.010 917.130 ;
        RECT 257.870 916.820 258.250 916.830 ;
        RECT 260.630 916.820 261.010 916.830 ;
        RECT 256.950 857.290 257.330 857.300 ;
        RECT 256.950 856.990 259.130 857.290 ;
        RECT 256.950 856.980 257.330 856.990 ;
        RECT 258.830 856.620 259.130 856.990 ;
        RECT 258.790 856.300 259.170 856.620 ;
        RECT 256.285 855.250 256.615 855.265 ;
        RECT 258.790 855.250 259.170 855.260 ;
        RECT 256.285 854.950 259.170 855.250 ;
        RECT 256.285 854.935 256.615 854.950 ;
        RECT 258.790 854.940 259.170 854.950 ;
        RECT 256.285 807.650 256.615 807.665 ;
        RECT 256.950 807.650 257.330 807.660 ;
        RECT 256.285 807.350 257.330 807.650 ;
        RECT 256.285 807.335 256.615 807.350 ;
        RECT 256.950 807.340 257.330 807.350 ;
        RECT 256.950 799.860 257.330 800.180 ;
        RECT 256.990 799.490 257.290 799.860 ;
        RECT 257.870 799.490 258.250 799.500 ;
        RECT 256.990 799.190 258.250 799.490 ;
        RECT 257.870 799.180 258.250 799.190 ;
        RECT 256.285 751.890 256.615 751.905 ;
        RECT 257.870 751.890 258.250 751.900 ;
        RECT 256.285 751.590 258.250 751.890 ;
        RECT 256.285 751.575 256.615 751.590 ;
        RECT 257.870 751.580 258.250 751.590 ;
        RECT 256.285 704.970 256.615 704.985 ;
        RECT 257.870 704.970 258.250 704.980 ;
        RECT 256.285 704.670 258.250 704.970 ;
        RECT 256.285 704.655 256.615 704.670 ;
        RECT 257.870 704.660 258.250 704.670 ;
        RECT 256.285 703.610 256.615 703.625 ;
        RECT 257.870 703.610 258.250 703.620 ;
        RECT 256.285 703.310 258.250 703.610 ;
        RECT 256.285 703.295 256.615 703.310 ;
        RECT 257.870 703.300 258.250 703.310 ;
        RECT 256.285 656.690 256.615 656.705 ;
        RECT 256.285 656.390 257.290 656.690 ;
        RECT 256.285 656.375 256.615 656.390 ;
        RECT 256.990 656.020 257.290 656.390 ;
        RECT 256.950 655.700 257.330 656.020 ;
        RECT 258.790 613.850 259.170 613.860 ;
        RECT 261.345 613.850 261.675 613.865 ;
        RECT 258.790 613.550 261.675 613.850 ;
        RECT 258.790 613.540 259.170 613.550 ;
        RECT 261.345 613.535 261.675 613.550 ;
        RECT 257.870 532.250 258.250 532.260 ;
        RECT 261.345 532.250 261.675 532.265 ;
        RECT 257.870 531.950 261.675 532.250 ;
        RECT 257.870 531.940 258.250 531.950 ;
        RECT 261.345 531.935 261.675 531.950 ;
        RECT 256.285 517.290 256.615 517.305 ;
        RECT 257.870 517.290 258.250 517.300 ;
        RECT 256.285 516.990 258.250 517.290 ;
        RECT 256.285 516.975 256.615 516.990 ;
        RECT 257.870 516.980 258.250 516.990 ;
        RECT 256.285 470.370 256.615 470.385 ;
        RECT 256.285 470.070 257.290 470.370 ;
        RECT 256.285 470.055 256.615 470.070 ;
        RECT 256.990 469.700 257.290 470.070 ;
        RECT 256.950 469.380 257.330 469.700 ;
        RECT 258.790 261.610 259.170 261.620 ;
        RECT 456.385 261.610 456.715 261.625 ;
        RECT 258.790 261.310 456.715 261.610 ;
        RECT 258.790 261.300 259.170 261.310 ;
        RECT 456.385 261.295 456.715 261.310 ;
      LAYER via3 ;
        RECT 542.180 3275.740 542.500 3276.060 ;
        RECT 548.620 3275.740 548.940 3276.060 ;
        RECT 2064.780 3275.740 2065.100 3276.060 ;
        RECT 260.660 2747.380 260.980 2747.700 ;
        RECT 257.900 2746.700 258.220 2747.020 ;
        RECT 257.900 2719.500 258.220 2719.820 ;
        RECT 257.900 2697.740 258.220 2698.060 ;
        RECT 257.900 2641.980 258.220 2642.300 ;
        RECT 257.900 2594.380 258.220 2594.700 ;
        RECT 257.900 2525.020 258.220 2525.340 ;
        RECT 258.820 2476.740 259.140 2477.060 ;
        RECT 258.820 2380.180 259.140 2380.500 ;
        RECT 258.820 2374.060 259.140 2374.380 ;
        RECT 258.820 2325.100 259.140 2325.420 ;
        RECT 258.820 2282.940 259.140 2283.260 ;
        RECT 258.820 2187.060 259.140 2187.380 ;
        RECT 258.820 2180.260 259.140 2180.580 ;
        RECT 258.820 2131.300 259.140 2131.620 ;
        RECT 258.820 2089.820 259.140 2090.140 ;
        RECT 258.820 2043.580 259.140 2043.900 ;
        RECT 257.900 2042.900 258.220 2043.220 ;
        RECT 258.820 2001.420 259.140 2001.740 ;
        RECT 257.900 2000.060 258.220 2000.380 ;
        RECT 257.900 1946.340 258.220 1946.660 ;
        RECT 256.980 1910.300 257.300 1910.620 ;
        RECT 258.820 1790.620 259.140 1790.940 ;
        RECT 260.660 1790.620 260.980 1790.940 ;
        RECT 257.900 1703.580 258.220 1703.900 ;
        RECT 260.660 1703.580 260.980 1703.900 ;
        RECT 256.980 1622.660 257.300 1622.980 ;
        RECT 258.820 1622.660 259.140 1622.980 ;
        RECT 258.820 1621.300 259.140 1621.620 ;
        RECT 257.900 1573.700 258.220 1574.020 ;
        RECT 258.820 1572.340 259.140 1572.660 ;
        RECT 257.900 1534.940 258.220 1535.260 ;
        RECT 258.820 1455.380 259.140 1455.700 ;
        RECT 258.820 1413.900 259.140 1414.220 ;
        RECT 258.820 1366.980 259.140 1367.300 ;
        RECT 257.900 1366.300 258.220 1366.620 ;
        RECT 258.820 1317.340 259.140 1317.660 ;
        RECT 257.900 1269.740 258.220 1270.060 ;
        RECT 257.900 1142.580 258.220 1142.900 ;
        RECT 258.820 1124.220 259.140 1124.540 ;
        RECT 258.820 1027.660 259.140 1027.980 ;
        RECT 260.660 1027.660 260.980 1027.980 ;
        RECT 257.900 916.820 258.220 917.140 ;
        RECT 260.660 916.820 260.980 917.140 ;
        RECT 256.980 856.980 257.300 857.300 ;
        RECT 258.820 856.300 259.140 856.620 ;
        RECT 258.820 854.940 259.140 855.260 ;
        RECT 256.980 807.340 257.300 807.660 ;
        RECT 256.980 799.860 257.300 800.180 ;
        RECT 257.900 799.180 258.220 799.500 ;
        RECT 257.900 751.580 258.220 751.900 ;
        RECT 257.900 704.660 258.220 704.980 ;
        RECT 257.900 703.300 258.220 703.620 ;
        RECT 256.980 655.700 257.300 656.020 ;
        RECT 258.820 613.540 259.140 613.860 ;
        RECT 257.900 531.940 258.220 532.260 ;
        RECT 257.900 516.980 258.220 517.300 ;
        RECT 256.980 469.380 257.300 469.700 ;
        RECT 258.820 261.300 259.140 261.620 ;
      LAYER met4 ;
        RECT 260.230 3275.310 261.410 3276.490 ;
        RECT 541.750 3275.310 542.930 3276.490 ;
        RECT 548.190 3275.310 549.370 3276.490 ;
        RECT 2064.350 3275.310 2065.530 3276.490 ;
        RECT 260.670 2747.705 260.970 3275.310 ;
        RECT 260.655 2747.375 260.985 2747.705 ;
        RECT 257.895 2746.695 258.225 2747.025 ;
        RECT 257.910 2719.825 258.210 2746.695 ;
        RECT 257.895 2719.495 258.225 2719.825 ;
        RECT 257.895 2698.050 258.225 2698.065 ;
        RECT 256.990 2697.750 258.225 2698.050 ;
        RECT 256.990 2657.250 257.290 2697.750 ;
        RECT 257.895 2697.735 258.225 2697.750 ;
        RECT 256.990 2656.950 258.440 2657.250 ;
        RECT 258.140 2653.850 258.440 2656.950 ;
        RECT 257.910 2653.550 258.440 2653.850 ;
        RECT 257.910 2642.305 258.210 2653.550 ;
        RECT 257.895 2641.975 258.225 2642.305 ;
        RECT 257.895 2594.375 258.225 2594.705 ;
        RECT 257.910 2525.345 258.210 2594.375 ;
        RECT 257.895 2525.015 258.225 2525.345 ;
        RECT 258.815 2476.735 259.145 2477.065 ;
        RECT 258.830 2380.505 259.130 2476.735 ;
        RECT 258.815 2380.175 259.145 2380.505 ;
        RECT 258.815 2374.055 259.145 2374.385 ;
        RECT 258.830 2325.425 259.130 2374.055 ;
        RECT 258.815 2325.095 259.145 2325.425 ;
        RECT 258.815 2282.935 259.145 2283.265 ;
        RECT 258.830 2259.450 259.130 2282.935 ;
        RECT 257.910 2259.150 259.130 2259.450 ;
        RECT 257.910 2235.650 258.210 2259.150 ;
        RECT 257.910 2235.350 259.130 2235.650 ;
        RECT 258.830 2187.385 259.130 2235.350 ;
        RECT 258.815 2187.055 259.145 2187.385 ;
        RECT 258.815 2180.255 259.145 2180.585 ;
        RECT 258.830 2131.625 259.130 2180.255 ;
        RECT 258.815 2131.295 259.145 2131.625 ;
        RECT 258.815 2089.815 259.145 2090.145 ;
        RECT 258.830 2043.905 259.130 2089.815 ;
        RECT 258.815 2043.575 259.145 2043.905 ;
        RECT 257.895 2042.895 258.225 2043.225 ;
        RECT 257.910 2041.850 258.210 2042.895 ;
        RECT 257.910 2041.550 259.130 2041.850 ;
        RECT 258.830 2001.745 259.130 2041.550 ;
        RECT 258.815 2001.415 259.145 2001.745 ;
        RECT 257.895 2000.055 258.225 2000.385 ;
        RECT 257.910 1946.665 258.210 2000.055 ;
        RECT 257.895 1946.335 258.225 1946.665 ;
        RECT 256.975 1910.295 257.305 1910.625 ;
        RECT 256.990 1899.050 257.290 1910.295 ;
        RECT 256.070 1898.750 257.290 1899.050 ;
        RECT 256.070 1837.850 256.370 1898.750 ;
        RECT 256.070 1837.550 259.130 1837.850 ;
        RECT 258.830 1790.945 259.130 1837.550 ;
        RECT 258.815 1790.615 259.145 1790.945 ;
        RECT 260.655 1790.615 260.985 1790.945 ;
        RECT 260.670 1703.905 260.970 1790.615 ;
        RECT 257.895 1703.575 258.225 1703.905 ;
        RECT 260.655 1703.575 260.985 1703.905 ;
        RECT 257.910 1657.650 258.210 1703.575 ;
        RECT 256.990 1657.350 258.210 1657.650 ;
        RECT 256.990 1622.985 257.290 1657.350 ;
        RECT 256.975 1622.655 257.305 1622.985 ;
        RECT 258.815 1622.655 259.145 1622.985 ;
        RECT 258.830 1621.625 259.130 1622.655 ;
        RECT 258.815 1621.295 259.145 1621.625 ;
        RECT 257.895 1573.695 258.225 1574.025 ;
        RECT 257.910 1572.650 258.210 1573.695 ;
        RECT 258.815 1572.650 259.145 1572.665 ;
        RECT 257.910 1572.350 259.145 1572.650 ;
        RECT 258.815 1572.335 259.145 1572.350 ;
        RECT 257.895 1534.935 258.225 1535.265 ;
        RECT 257.910 1487.650 258.210 1534.935 ;
        RECT 257.910 1487.350 259.130 1487.650 ;
        RECT 258.830 1455.705 259.130 1487.350 ;
        RECT 258.815 1455.375 259.145 1455.705 ;
        RECT 258.815 1413.895 259.145 1414.225 ;
        RECT 258.830 1367.305 259.130 1413.895 ;
        RECT 258.815 1366.975 259.145 1367.305 ;
        RECT 257.895 1366.295 258.225 1366.625 ;
        RECT 257.910 1365.250 258.210 1366.295 ;
        RECT 257.910 1364.950 259.130 1365.250 ;
        RECT 258.830 1317.665 259.130 1364.950 ;
        RECT 258.815 1317.335 259.145 1317.665 ;
        RECT 257.895 1269.735 258.225 1270.065 ;
        RECT 257.910 1142.905 258.210 1269.735 ;
        RECT 257.895 1142.575 258.225 1142.905 ;
        RECT 258.815 1124.215 259.145 1124.545 ;
        RECT 258.830 1027.985 259.130 1124.215 ;
        RECT 258.815 1027.655 259.145 1027.985 ;
        RECT 260.655 1027.655 260.985 1027.985 ;
        RECT 260.670 917.145 260.970 1027.655 ;
        RECT 257.895 916.815 258.225 917.145 ;
        RECT 260.655 916.815 260.985 917.145 ;
        RECT 257.910 885.850 258.210 916.815 ;
        RECT 256.990 885.550 258.210 885.850 ;
        RECT 256.990 857.305 257.290 885.550 ;
        RECT 256.975 856.975 257.305 857.305 ;
        RECT 258.815 856.295 259.145 856.625 ;
        RECT 258.830 855.265 259.130 856.295 ;
        RECT 258.815 854.935 259.145 855.265 ;
        RECT 256.975 807.335 257.305 807.665 ;
        RECT 256.990 800.185 257.290 807.335 ;
        RECT 256.975 799.855 257.305 800.185 ;
        RECT 257.895 799.175 258.225 799.505 ;
        RECT 257.910 751.905 258.210 799.175 ;
        RECT 257.895 751.575 258.225 751.905 ;
        RECT 257.895 704.655 258.225 704.985 ;
        RECT 257.910 703.625 258.210 704.655 ;
        RECT 257.895 703.295 258.225 703.625 ;
        RECT 256.975 655.695 257.305 656.025 ;
        RECT 256.990 637.650 257.290 655.695 ;
        RECT 256.990 637.350 258.210 637.650 ;
        RECT 257.910 613.850 258.210 637.350 ;
        RECT 258.815 613.850 259.145 613.865 ;
        RECT 257.910 613.550 259.145 613.850 ;
        RECT 258.815 613.535 259.145 613.550 ;
        RECT 257.895 531.935 258.225 532.265 ;
        RECT 257.910 517.305 258.210 531.935 ;
        RECT 257.895 516.975 258.225 517.305 ;
        RECT 256.975 469.375 257.305 469.705 ;
        RECT 256.990 447.250 257.290 469.375 ;
        RECT 256.990 446.950 258.210 447.250 ;
        RECT 257.910 403.050 258.210 446.950 ;
        RECT 256.990 402.750 258.210 403.050 ;
        RECT 256.990 386.050 257.290 402.750 ;
        RECT 256.990 385.750 258.210 386.050 ;
        RECT 257.910 362.250 258.210 385.750 ;
        RECT 256.990 361.950 258.210 362.250 ;
        RECT 256.990 301.050 257.290 361.950 ;
        RECT 256.990 300.750 259.130 301.050 ;
        RECT 258.830 261.625 259.130 300.750 ;
        RECT 258.815 261.295 259.145 261.625 ;
      LAYER met5 ;
        RECT 639.980 3280.100 642.500 3283.500 ;
        RECT 736.580 3280.100 739.100 3283.500 ;
        RECT 929.780 3280.100 932.300 3283.500 ;
        RECT 1026.380 3280.100 1028.900 3283.500 ;
        RECT 1219.580 3281.900 1242.340 3283.500 ;
        RECT 1219.580 3280.100 1221.180 3281.900 ;
        RECT 299.580 3278.500 304.860 3280.100 ;
        RECT 299.580 3276.700 301.180 3278.500 ;
        RECT 260.020 3275.100 301.180 3276.700 ;
        RECT 303.260 3276.700 304.860 3278.500 ;
        RECT 398.940 3278.500 449.300 3280.100 ;
        RECT 398.940 3276.700 400.540 3278.500 ;
        RECT 303.260 3275.100 400.540 3276.700 ;
        RECT 447.700 3276.700 449.300 3278.500 ;
        RECT 592.140 3278.500 597.420 3280.100 ;
        RECT 592.140 3276.700 593.740 3278.500 ;
        RECT 447.700 3275.100 543.140 3276.700 ;
        RECT 547.980 3275.100 593.740 3276.700 ;
        RECT 595.820 3276.700 597.420 3278.500 ;
        RECT 638.140 3278.500 645.260 3280.100 ;
        RECT 638.140 3276.700 639.740 3278.500 ;
        RECT 595.820 3275.100 639.740 3276.700 ;
        RECT 643.660 3276.700 645.260 3278.500 ;
        RECT 685.980 3278.500 691.260 3280.100 ;
        RECT 685.980 3276.700 687.580 3278.500 ;
        RECT 643.660 3275.100 687.580 3276.700 ;
        RECT 689.660 3276.700 691.260 3278.500 ;
        RECT 736.580 3278.500 741.860 3280.100 ;
        RECT 736.580 3276.700 738.180 3278.500 ;
        RECT 689.660 3275.100 738.180 3276.700 ;
        RECT 740.260 3276.700 741.860 3278.500 ;
        RECT 782.580 3278.500 835.700 3280.100 ;
        RECT 782.580 3276.700 784.180 3278.500 ;
        RECT 740.260 3275.100 784.180 3276.700 ;
        RECT 834.100 3276.700 835.700 3278.500 ;
        RECT 881.940 3276.700 884.460 3280.100 ;
        RECT 929.780 3278.500 935.060 3280.100 ;
        RECT 929.780 3276.700 931.380 3278.500 ;
        RECT 834.100 3275.100 931.380 3276.700 ;
        RECT 933.460 3276.700 935.060 3278.500 ;
        RECT 975.780 3278.500 983.820 3280.100 ;
        RECT 975.780 3276.700 977.380 3278.500 ;
        RECT 933.460 3275.100 977.380 3276.700 ;
        RECT 982.220 3276.700 983.820 3278.500 ;
        RECT 1024.540 3278.500 1031.660 3280.100 ;
        RECT 1024.540 3276.700 1026.140 3278.500 ;
        RECT 982.220 3275.100 1026.140 3276.700 ;
        RECT 1030.060 3276.700 1031.660 3278.500 ;
        RECT 1171.740 3278.500 1177.020 3280.100 ;
        RECT 1171.740 3276.700 1173.340 3278.500 ;
        RECT 1030.060 3275.100 1173.340 3276.700 ;
        RECT 1175.420 3276.700 1177.020 3278.500 ;
        RECT 1217.740 3278.500 1221.180 3280.100 ;
        RECT 1217.740 3276.700 1219.340 3278.500 ;
        RECT 1175.420 3275.100 1219.340 3276.700 ;
        RECT 1240.740 3276.700 1242.340 3281.900 ;
        RECT 1412.780 3280.100 1415.300 3283.500 ;
        RECT 1509.380 3280.100 1511.900 3283.500 ;
        RECT 1702.580 3281.900 1725.340 3283.500 ;
        RECT 1702.580 3280.100 1704.180 3281.900 ;
        RECT 1313.420 3278.500 1318.700 3280.100 ;
        RECT 1313.420 3276.700 1315.020 3278.500 ;
        RECT 1240.740 3275.100 1315.020 3276.700 ;
        RECT 1317.100 3276.700 1318.700 3278.500 ;
        RECT 1365.860 3278.500 1463.140 3280.100 ;
        RECT 1365.860 3276.700 1367.460 3278.500 ;
        RECT 1317.100 3275.100 1367.460 3276.700 ;
        RECT 1461.540 3276.700 1463.140 3278.500 ;
        RECT 1507.540 3278.500 1559.740 3280.100 ;
        RECT 1507.540 3276.700 1509.140 3278.500 ;
        RECT 1461.540 3275.100 1509.140 3276.700 ;
        RECT 1558.140 3276.700 1559.740 3278.500 ;
        RECT 1655.660 3278.500 1704.180 3280.100 ;
        RECT 1655.660 3276.700 1657.260 3278.500 ;
        RECT 1558.140 3275.100 1657.260 3276.700 ;
        RECT 1723.740 3276.700 1725.340 3281.900 ;
        RECT 1772.500 3281.900 1821.940 3283.500 ;
        RECT 1772.500 3276.700 1774.100 3281.900 ;
        RECT 1723.740 3275.100 1774.100 3276.700 ;
        RECT 1820.340 3276.700 1821.940 3281.900 ;
        RECT 1869.100 3281.900 1898.300 3283.500 ;
        RECT 1869.100 3276.700 1870.700 3281.900 ;
        RECT 1896.700 3280.100 1898.300 3281.900 ;
        RECT 1965.700 3281.900 1994.900 3283.500 ;
        RECT 1896.700 3278.500 1946.140 3280.100 ;
        RECT 1820.340 3275.100 1870.700 3276.700 ;
        RECT 1944.540 3276.700 1946.140 3278.500 ;
        RECT 1965.700 3276.700 1967.300 3281.900 ;
        RECT 1993.300 3280.100 1994.900 3281.900 ;
        RECT 1993.300 3278.500 2042.740 3280.100 ;
        RECT 1944.540 3275.100 1967.300 3276.700 ;
        RECT 2041.140 3276.700 2042.740 3278.500 ;
        RECT 2041.140 3275.100 2065.740 3276.700 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1072.790 247.420 1073.110 247.480 ;
        RECT 1227.350 247.420 1227.670 247.480 ;
        RECT 1072.790 247.280 1227.670 247.420 ;
        RECT 1072.790 247.220 1073.110 247.280 ;
        RECT 1227.350 247.220 1227.670 247.280 ;
        RECT 482.610 142.360 482.930 142.420 ;
        RECT 1072.790 142.360 1073.110 142.420 ;
        RECT 482.610 142.220 1073.110 142.360 ;
        RECT 482.610 142.160 482.930 142.220 ;
        RECT 1072.790 142.160 1073.110 142.220 ;
        RECT 478.470 19.620 478.790 19.680 ;
        RECT 482.610 19.620 482.930 19.680 ;
        RECT 478.470 19.480 482.930 19.620 ;
        RECT 478.470 19.420 478.790 19.480 ;
        RECT 482.610 19.420 482.930 19.480 ;
      LAYER via ;
        RECT 1072.820 247.220 1073.080 247.480 ;
        RECT 1227.380 247.220 1227.640 247.480 ;
        RECT 482.640 142.160 482.900 142.420 ;
        RECT 1072.820 142.160 1073.080 142.420 ;
        RECT 478.500 19.420 478.760 19.680 ;
        RECT 482.640 19.420 482.900 19.680 ;
      LAYER met2 ;
        RECT 1227.330 260.000 1227.610 264.000 ;
        RECT 1227.440 247.510 1227.580 260.000 ;
        RECT 1072.820 247.190 1073.080 247.510 ;
        RECT 1227.380 247.190 1227.640 247.510 ;
        RECT 1072.880 142.450 1073.020 247.190 ;
        RECT 482.640 142.130 482.900 142.450 ;
        RECT 1072.820 142.130 1073.080 142.450 ;
        RECT 482.700 19.710 482.840 142.130 ;
        RECT 478.500 19.390 478.760 19.710 ;
        RECT 482.640 19.390 482.900 19.710 ;
        RECT 478.560 2.400 478.700 19.390 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 3273.760 227.630 3273.820 ;
        RECT 361.630 3273.760 361.950 3273.820 ;
        RECT 227.310 3273.620 361.950 3273.760 ;
        RECT 227.310 3273.560 227.630 3273.620 ;
        RECT 361.630 3273.560 361.950 3273.620 ;
        RECT 227.310 29.820 227.630 29.880 ;
        RECT 496.410 29.820 496.730 29.880 ;
        RECT 227.310 29.680 496.730 29.820 ;
        RECT 227.310 29.620 227.630 29.680 ;
        RECT 496.410 29.620 496.730 29.680 ;
      LAYER via ;
        RECT 227.340 3273.560 227.600 3273.820 ;
        RECT 361.660 3273.560 361.920 3273.820 ;
        RECT 227.340 29.620 227.600 29.880 ;
        RECT 496.440 29.620 496.700 29.880 ;
      LAYER met2 ;
        RECT 227.340 3273.530 227.600 3273.850 ;
        RECT 361.660 3273.530 361.920 3273.850 ;
        RECT 227.400 29.910 227.540 3273.530 ;
        RECT 361.720 3260.000 361.860 3273.530 ;
        RECT 361.610 3256.000 361.890 3260.000 ;
        RECT 227.340 29.590 227.600 29.910 ;
        RECT 496.440 29.590 496.700 29.910 ;
        RECT 496.500 2.400 496.640 29.590 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 511.205 186.405 511.375 234.515 ;
        RECT 511.205 48.365 511.375 137.955 ;
      LAYER mcon ;
        RECT 511.205 234.345 511.375 234.515 ;
        RECT 511.205 137.785 511.375 137.955 ;
      LAYER met1 ;
        RECT 274.230 2353.040 274.550 2353.100 ;
        RECT 296.770 2353.040 297.090 2353.100 ;
        RECT 274.230 2352.900 297.090 2353.040 ;
        RECT 274.230 2352.840 274.550 2352.900 ;
        RECT 296.770 2352.840 297.090 2352.900 ;
        RECT 274.230 246.740 274.550 246.800 ;
        RECT 511.130 246.740 511.450 246.800 ;
        RECT 274.230 246.600 511.450 246.740 ;
        RECT 274.230 246.540 274.550 246.600 ;
        RECT 511.130 246.540 511.450 246.600 ;
        RECT 511.130 234.500 511.450 234.560 ;
        RECT 510.935 234.360 511.450 234.500 ;
        RECT 511.130 234.300 511.450 234.360 ;
        RECT 511.130 186.560 511.450 186.620 ;
        RECT 510.935 186.420 511.450 186.560 ;
        RECT 511.130 186.360 511.450 186.420 ;
        RECT 511.130 137.940 511.450 138.000 ;
        RECT 510.935 137.800 511.450 137.940 ;
        RECT 511.130 137.740 511.450 137.800 ;
        RECT 511.145 48.520 511.435 48.565 ;
        RECT 513.890 48.520 514.210 48.580 ;
        RECT 511.145 48.380 514.210 48.520 ;
        RECT 511.145 48.335 511.435 48.380 ;
        RECT 513.890 48.320 514.210 48.380 ;
      LAYER via ;
        RECT 274.260 2352.840 274.520 2353.100 ;
        RECT 296.800 2352.840 297.060 2353.100 ;
        RECT 274.260 246.540 274.520 246.800 ;
        RECT 511.160 246.540 511.420 246.800 ;
        RECT 511.160 234.300 511.420 234.560 ;
        RECT 511.160 186.360 511.420 186.620 ;
        RECT 511.160 137.740 511.420 138.000 ;
        RECT 513.920 48.320 514.180 48.580 ;
      LAYER met2 ;
        RECT 296.790 2355.675 297.070 2356.045 ;
        RECT 296.860 2353.130 297.000 2355.675 ;
        RECT 274.260 2352.810 274.520 2353.130 ;
        RECT 296.800 2352.810 297.060 2353.130 ;
        RECT 274.320 246.830 274.460 2352.810 ;
        RECT 274.260 246.510 274.520 246.830 ;
        RECT 511.160 246.510 511.420 246.830 ;
        RECT 511.220 234.590 511.360 246.510 ;
        RECT 511.160 234.270 511.420 234.590 ;
        RECT 511.160 186.330 511.420 186.650 ;
        RECT 511.220 138.030 511.360 186.330 ;
        RECT 511.160 137.710 511.420 138.030 ;
        RECT 513.920 48.290 514.180 48.610 ;
        RECT 513.980 2.400 514.120 48.290 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 296.790 2355.720 297.070 2356.000 ;
      LAYER met3 ;
        RECT 296.765 2356.010 297.095 2356.025 ;
        RECT 310.000 2356.010 314.000 2356.400 ;
        RECT 296.765 2355.800 314.000 2356.010 ;
        RECT 296.765 2355.710 310.500 2355.800 ;
        RECT 296.765 2355.695 297.095 2355.710 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 3259.140 246.950 3259.200 ;
        RECT 1462.410 3259.140 1462.730 3259.200 ;
        RECT 246.630 3259.000 1462.730 3259.140 ;
        RECT 246.630 3258.940 246.950 3259.000 ;
        RECT 1462.410 3258.940 1462.730 3259.000 ;
      LAYER via ;
        RECT 246.660 3258.940 246.920 3259.200 ;
        RECT 1462.440 3258.940 1462.700 3259.200 ;
      LAYER met2 ;
        RECT 246.660 3258.910 246.920 3259.230 ;
        RECT 1462.440 3258.970 1462.700 3259.230 ;
        RECT 1462.850 3258.970 1463.130 3260.000 ;
        RECT 1462.440 3258.910 1463.130 3258.970 ;
        RECT 246.720 244.645 246.860 3258.910 ;
        RECT 1462.500 3258.830 1463.130 3258.910 ;
        RECT 1462.850 3256.000 1463.130 3258.830 ;
        RECT 246.650 244.275 246.930 244.645 ;
        RECT 531.390 244.275 531.670 244.645 ;
        RECT 531.460 7.890 531.600 244.275 ;
        RECT 531.460 7.750 532.060 7.890 ;
        RECT 531.920 2.400 532.060 7.750 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 246.650 244.320 246.930 244.600 ;
        RECT 531.390 244.320 531.670 244.600 ;
      LAYER met3 ;
        RECT 246.625 244.610 246.955 244.625 ;
        RECT 531.365 244.610 531.695 244.625 ;
        RECT 246.625 244.310 531.695 244.610 ;
        RECT 246.625 244.295 246.955 244.310 ;
        RECT 531.365 244.295 531.695 244.310 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 2277.220 2615.490 2277.280 ;
        RECT 2673.130 2277.220 2673.450 2277.280 ;
        RECT 2615.170 2277.080 2673.450 2277.220 ;
        RECT 2615.170 2277.020 2615.490 2277.080 ;
        RECT 2673.130 2277.020 2673.450 2277.080 ;
        RECT 549.770 2.960 550.090 3.020 ;
        RECT 551.610 2.960 551.930 3.020 ;
        RECT 549.770 2.820 551.930 2.960 ;
        RECT 549.770 2.760 550.090 2.820 ;
        RECT 551.610 2.760 551.930 2.820 ;
      LAYER via ;
        RECT 2615.200 2277.020 2615.460 2277.280 ;
        RECT 2673.160 2277.020 2673.420 2277.280 ;
        RECT 549.800 2.760 550.060 3.020 ;
        RECT 551.640 2.760 551.900 3.020 ;
      LAYER met2 ;
        RECT 2615.190 2283.595 2615.470 2283.965 ;
        RECT 2615.260 2277.310 2615.400 2283.595 ;
        RECT 2615.200 2276.990 2615.460 2277.310 ;
        RECT 2673.160 2276.990 2673.420 2277.310 ;
        RECT 2673.220 244.645 2673.360 2276.990 ;
        RECT 551.630 244.275 551.910 244.645 ;
        RECT 2673.150 244.275 2673.430 244.645 ;
        RECT 551.700 3.050 551.840 244.275 ;
        RECT 549.800 2.730 550.060 3.050 ;
        RECT 551.640 2.730 551.900 3.050 ;
        RECT 549.860 2.400 550.000 2.730 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 2615.190 2283.640 2615.470 2283.920 ;
        RECT 551.630 244.320 551.910 244.600 ;
        RECT 2673.150 244.320 2673.430 244.600 ;
      LAYER met3 ;
        RECT 2606.000 2283.930 2610.000 2284.320 ;
        RECT 2615.165 2283.930 2615.495 2283.945 ;
        RECT 2606.000 2283.720 2615.495 2283.930 ;
        RECT 2609.580 2283.630 2615.495 2283.720 ;
        RECT 2615.165 2283.615 2615.495 2283.630 ;
        RECT 551.605 244.610 551.935 244.625 ;
        RECT 2673.125 244.610 2673.455 244.625 ;
        RECT 551.605 244.310 2673.455 244.610 ;
        RECT 551.605 244.295 551.935 244.310 ;
        RECT 2673.125 244.295 2673.455 244.310 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.730 58.635 568.010 59.005 ;
        RECT 567.800 2.400 567.940 58.635 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 567.730 58.680 568.010 58.960 ;
      LAYER met3 ;
        RECT 2606.000 2326.090 2610.000 2326.480 ;
        RECT 2643.430 2326.090 2643.810 2326.100 ;
        RECT 2606.000 2325.880 2643.810 2326.090 ;
        RECT 2609.580 2325.790 2643.810 2325.880 ;
        RECT 2643.430 2325.780 2643.810 2325.790 ;
        RECT 567.705 58.970 568.035 58.985 ;
        RECT 2643.430 58.970 2643.810 58.980 ;
        RECT 567.705 58.670 2643.810 58.970 ;
        RECT 567.705 58.655 568.035 58.670 ;
        RECT 2643.430 58.660 2643.810 58.670 ;
      LAYER via3 ;
        RECT 2643.460 2325.780 2643.780 2326.100 ;
        RECT 2643.460 58.660 2643.780 58.980 ;
      LAYER met4 ;
        RECT 2643.455 2325.775 2643.785 2326.105 ;
        RECT 2643.470 58.985 2643.770 2325.775 ;
        RECT 2643.455 58.655 2643.785 58.985 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 293.090 917.900 293.410 917.960 ;
        RECT 300.450 917.900 300.770 917.960 ;
        RECT 293.090 917.760 300.770 917.900 ;
        RECT 293.090 917.700 293.410 917.760 ;
        RECT 300.450 917.700 300.770 917.760 ;
      LAYER via ;
        RECT 293.120 917.700 293.380 917.960 ;
        RECT 300.480 917.700 300.740 917.960 ;
      LAYER met2 ;
        RECT 300.470 3223.355 300.750 3223.725 ;
        RECT 300.540 917.990 300.680 3223.355 ;
        RECT 293.120 917.670 293.380 917.990 ;
        RECT 300.480 917.670 300.740 917.990 ;
        RECT 293.180 16.165 293.320 917.670 ;
        RECT 293.110 15.795 293.390 16.165 ;
        RECT 585.670 15.795 585.950 16.165 ;
        RECT 585.740 2.400 585.880 15.795 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 300.470 3223.400 300.750 3223.680 ;
        RECT 293.110 15.840 293.390 16.120 ;
        RECT 585.670 15.840 585.950 16.120 ;
      LAYER met3 ;
        RECT 300.445 3223.690 300.775 3223.705 ;
        RECT 310.000 3223.690 314.000 3224.080 ;
        RECT 300.445 3223.480 314.000 3223.690 ;
        RECT 300.445 3223.390 310.500 3223.480 ;
        RECT 300.445 3223.375 300.775 3223.390 ;
        RECT 293.085 16.130 293.415 16.145 ;
        RECT 585.645 16.130 585.975 16.145 ;
        RECT 293.085 15.830 585.975 16.130 ;
        RECT 293.085 15.815 293.415 15.830 ;
        RECT 585.645 15.815 585.975 15.830 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.590 247.420 948.910 247.480 ;
        RECT 1070.030 247.420 1070.350 247.480 ;
        RECT 948.590 247.280 1070.350 247.420 ;
        RECT 948.590 247.220 948.910 247.280 ;
        RECT 1070.030 247.220 1070.350 247.280 ;
        RECT 96.210 182.820 96.530 182.880 ;
        RECT 948.590 182.820 948.910 182.880 ;
        RECT 96.210 182.680 948.910 182.820 ;
        RECT 96.210 182.620 96.530 182.680 ;
        RECT 948.590 182.620 948.910 182.680 ;
        RECT 91.610 16.900 91.930 16.960 ;
        RECT 96.210 16.900 96.530 16.960 ;
        RECT 91.610 16.760 96.530 16.900 ;
        RECT 91.610 16.700 91.930 16.760 ;
        RECT 96.210 16.700 96.530 16.760 ;
      LAYER via ;
        RECT 948.620 247.220 948.880 247.480 ;
        RECT 1070.060 247.220 1070.320 247.480 ;
        RECT 96.240 182.620 96.500 182.880 ;
        RECT 948.620 182.620 948.880 182.880 ;
        RECT 91.640 16.700 91.900 16.960 ;
        RECT 96.240 16.700 96.500 16.960 ;
      LAYER met2 ;
        RECT 1070.010 260.000 1070.290 264.000 ;
        RECT 1070.120 247.510 1070.260 260.000 ;
        RECT 948.620 247.190 948.880 247.510 ;
        RECT 1070.060 247.190 1070.320 247.510 ;
        RECT 948.680 182.910 948.820 247.190 ;
        RECT 96.240 182.590 96.500 182.910 ;
        RECT 948.620 182.590 948.880 182.910 ;
        RECT 96.300 16.990 96.440 182.590 ;
        RECT 91.640 16.670 91.900 16.990 ;
        RECT 96.240 16.670 96.500 16.990 ;
        RECT 91.700 2.400 91.840 16.670 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 862.820 2615.490 862.880 ;
        RECT 2681.410 862.820 2681.730 862.880 ;
        RECT 2615.170 862.680 2681.730 862.820 ;
        RECT 2615.170 862.620 2615.490 862.680 ;
        RECT 2681.410 862.620 2681.730 862.680 ;
        RECT 606.810 245.040 607.130 245.100 ;
        RECT 2681.410 245.040 2681.730 245.100 ;
        RECT 606.810 244.900 2681.730 245.040 ;
        RECT 606.810 244.840 607.130 244.900 ;
        RECT 2681.410 244.840 2681.730 244.900 ;
        RECT 603.130 20.640 603.450 20.700 ;
        RECT 606.810 20.640 607.130 20.700 ;
        RECT 603.130 20.500 607.130 20.640 ;
        RECT 603.130 20.440 603.450 20.500 ;
        RECT 606.810 20.440 607.130 20.500 ;
      LAYER via ;
        RECT 2615.200 862.620 2615.460 862.880 ;
        RECT 2681.440 862.620 2681.700 862.880 ;
        RECT 606.840 244.840 607.100 245.100 ;
        RECT 2681.440 244.840 2681.700 245.100 ;
        RECT 603.160 20.440 603.420 20.700 ;
        RECT 606.840 20.440 607.100 20.700 ;
      LAYER met2 ;
        RECT 2615.190 866.475 2615.470 866.845 ;
        RECT 2615.260 862.910 2615.400 866.475 ;
        RECT 2615.200 862.590 2615.460 862.910 ;
        RECT 2681.440 862.590 2681.700 862.910 ;
        RECT 2681.500 245.130 2681.640 862.590 ;
        RECT 606.840 244.810 607.100 245.130 ;
        RECT 2681.440 244.810 2681.700 245.130 ;
        RECT 606.900 20.730 607.040 244.810 ;
        RECT 603.160 20.410 603.420 20.730 ;
        RECT 606.840 20.410 607.100 20.730 ;
        RECT 603.220 2.400 603.360 20.410 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 2615.190 866.520 2615.470 866.800 ;
      LAYER met3 ;
        RECT 2606.000 866.810 2610.000 867.200 ;
        RECT 2615.165 866.810 2615.495 866.825 ;
        RECT 2606.000 866.600 2615.495 866.810 ;
        RECT 2609.580 866.510 2615.495 866.600 ;
        RECT 2615.165 866.495 2615.495 866.510 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2615.170 966.180 2615.490 966.240 ;
        RECT 2674.050 966.180 2674.370 966.240 ;
        RECT 2615.170 966.040 2674.370 966.180 ;
        RECT 2615.170 965.980 2615.490 966.040 ;
        RECT 2674.050 965.980 2674.370 966.040 ;
        RECT 627.510 211.040 627.830 211.100 ;
        RECT 2674.050 211.040 2674.370 211.100 ;
        RECT 627.510 210.900 2674.370 211.040 ;
        RECT 627.510 210.840 627.830 210.900 ;
        RECT 2674.050 210.840 2674.370 210.900 ;
        RECT 621.070 20.640 621.390 20.700 ;
        RECT 627.510 20.640 627.830 20.700 ;
        RECT 621.070 20.500 627.830 20.640 ;
        RECT 621.070 20.440 621.390 20.500 ;
        RECT 627.510 20.440 627.830 20.500 ;
      LAYER via ;
        RECT 2615.200 965.980 2615.460 966.240 ;
        RECT 2674.080 965.980 2674.340 966.240 ;
        RECT 627.540 210.840 627.800 211.100 ;
        RECT 2674.080 210.840 2674.340 211.100 ;
        RECT 621.100 20.440 621.360 20.700 ;
        RECT 627.540 20.440 627.800 20.700 ;
      LAYER met2 ;
        RECT 2615.190 972.555 2615.470 972.925 ;
        RECT 2615.260 966.270 2615.400 972.555 ;
        RECT 2615.200 965.950 2615.460 966.270 ;
        RECT 2674.080 965.950 2674.340 966.270 ;
        RECT 2674.140 211.130 2674.280 965.950 ;
        RECT 627.540 210.810 627.800 211.130 ;
        RECT 2674.080 210.810 2674.340 211.130 ;
        RECT 627.600 20.730 627.740 210.810 ;
        RECT 621.100 20.410 621.360 20.730 ;
        RECT 627.540 20.410 627.800 20.730 ;
        RECT 621.160 2.400 621.300 20.410 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 2615.190 972.600 2615.470 972.880 ;
      LAYER met3 ;
        RECT 2606.000 972.890 2610.000 973.280 ;
        RECT 2615.165 972.890 2615.495 972.905 ;
        RECT 2606.000 972.680 2615.495 972.890 ;
        RECT 2609.580 972.590 2615.495 972.680 ;
        RECT 2615.165 972.575 2615.495 972.590 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2266.490 241.640 2266.810 241.700 ;
        RECT 2271.550 241.640 2271.870 241.700 ;
        RECT 2266.490 241.500 2271.870 241.640 ;
        RECT 2266.490 241.440 2266.810 241.500 ;
        RECT 2271.550 241.440 2271.870 241.500 ;
        RECT 115.530 45.800 115.850 45.860 ;
        RECT 2266.490 45.800 2266.810 45.860 ;
        RECT 115.530 45.660 2266.810 45.800 ;
        RECT 115.530 45.600 115.850 45.660 ;
        RECT 2266.490 45.600 2266.810 45.660 ;
      LAYER via ;
        RECT 2266.520 241.440 2266.780 241.700 ;
        RECT 2271.580 241.440 2271.840 241.700 ;
        RECT 115.560 45.600 115.820 45.860 ;
        RECT 2266.520 45.600 2266.780 45.860 ;
      LAYER met2 ;
        RECT 2271.530 260.000 2271.810 264.000 ;
        RECT 2271.640 241.730 2271.780 260.000 ;
        RECT 2266.520 241.410 2266.780 241.730 ;
        RECT 2271.580 241.410 2271.840 241.730 ;
        RECT 2266.580 45.890 2266.720 241.410 ;
        RECT 115.560 45.570 115.820 45.890 ;
        RECT 2266.520 45.570 2266.780 45.890 ;
        RECT 115.620 2.400 115.760 45.570 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 144.510 246.400 144.830 246.460 ;
        RECT 610.030 246.400 610.350 246.460 ;
        RECT 144.510 246.260 610.350 246.400 ;
        RECT 144.510 246.200 144.830 246.260 ;
        RECT 610.030 246.200 610.350 246.260 ;
        RECT 139.450 17.580 139.770 17.640 ;
        RECT 144.510 17.580 144.830 17.640 ;
        RECT 139.450 17.440 144.830 17.580 ;
        RECT 139.450 17.380 139.770 17.440 ;
        RECT 144.510 17.380 144.830 17.440 ;
      LAYER via ;
        RECT 144.540 246.200 144.800 246.460 ;
        RECT 610.060 246.200 610.320 246.460 ;
        RECT 139.480 17.380 139.740 17.640 ;
        RECT 144.540 17.380 144.800 17.640 ;
      LAYER met2 ;
        RECT 612.770 260.170 613.050 264.000 ;
        RECT 610.120 260.030 613.050 260.170 ;
        RECT 610.120 246.490 610.260 260.030 ;
        RECT 612.770 260.000 613.050 260.030 ;
        RECT 144.540 246.170 144.800 246.490 ;
        RECT 610.060 246.170 610.320 246.490 ;
        RECT 144.600 17.670 144.740 246.170 ;
        RECT 139.480 17.350 139.740 17.670 ;
        RECT 144.540 17.350 144.800 17.670 ;
        RECT 139.540 2.400 139.680 17.350 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 31.435 157.690 31.805 ;
        RECT 157.480 2.400 157.620 31.435 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 157.410 31.480 157.690 31.760 ;
      LAYER met3 ;
        RECT 2606.000 2051.370 2610.000 2051.760 ;
        RECT 2644.350 2051.370 2644.730 2051.380 ;
        RECT 2606.000 2051.160 2644.730 2051.370 ;
        RECT 2609.580 2051.070 2644.730 2051.160 ;
        RECT 2644.350 2051.060 2644.730 2051.070 ;
        RECT 157.385 31.770 157.715 31.785 ;
        RECT 2644.350 31.770 2644.730 31.780 ;
        RECT 157.385 31.470 2644.730 31.770 ;
        RECT 157.385 31.455 157.715 31.470 ;
        RECT 2644.350 31.460 2644.730 31.470 ;
      LAYER via3 ;
        RECT 2644.380 2051.060 2644.700 2051.380 ;
        RECT 2644.380 31.460 2644.700 31.780 ;
      LAYER met4 ;
        RECT 2644.375 2051.055 2644.705 2051.385 ;
        RECT 2644.390 31.785 2644.690 2051.055 ;
        RECT 2644.375 31.455 2644.705 31.785 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 555.290 245.380 555.610 245.440 ;
        RECT 1784.870 245.380 1785.190 245.440 ;
        RECT 555.290 245.240 1785.190 245.380 ;
        RECT 555.290 245.180 555.610 245.240 ;
        RECT 1784.870 245.180 1785.190 245.240 ;
        RECT 174.870 18.940 175.190 19.000 ;
        RECT 555.290 18.940 555.610 19.000 ;
        RECT 174.870 18.800 555.610 18.940 ;
        RECT 174.870 18.740 175.190 18.800 ;
        RECT 555.290 18.740 555.610 18.800 ;
      LAYER via ;
        RECT 555.320 245.180 555.580 245.440 ;
        RECT 1784.900 245.180 1785.160 245.440 ;
        RECT 174.900 18.740 175.160 19.000 ;
        RECT 555.320 18.740 555.580 19.000 ;
      LAYER met2 ;
        RECT 1784.850 260.000 1785.130 264.000 ;
        RECT 1784.960 245.470 1785.100 260.000 ;
        RECT 555.320 245.150 555.580 245.470 ;
        RECT 1784.900 245.150 1785.160 245.470 ;
        RECT 555.380 19.030 555.520 245.150 ;
        RECT 174.900 18.710 175.160 19.030 ;
        RECT 555.320 18.710 555.580 19.030 ;
        RECT 174.960 2.400 175.100 18.710 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 598.145 18.785 598.315 20.315 ;
      LAYER mcon ;
        RECT 598.145 20.145 598.315 20.315 ;
      LAYER met1 ;
        RECT 610.490 246.400 610.810 246.460 ;
        RECT 1342.350 246.400 1342.670 246.460 ;
        RECT 610.490 246.260 1342.670 246.400 ;
        RECT 610.490 246.200 610.810 246.260 ;
        RECT 1342.350 246.200 1342.670 246.260 ;
        RECT 192.350 20.300 192.670 20.360 ;
        RECT 598.085 20.300 598.375 20.345 ;
        RECT 192.350 20.160 598.375 20.300 ;
        RECT 192.350 20.100 192.670 20.160 ;
        RECT 598.085 20.115 598.375 20.160 ;
        RECT 607.270 20.300 607.590 20.360 ;
        RECT 610.490 20.300 610.810 20.360 ;
        RECT 607.270 20.160 610.810 20.300 ;
        RECT 607.270 20.100 607.590 20.160 ;
        RECT 610.490 20.100 610.810 20.160 ;
        RECT 598.085 18.940 598.375 18.985 ;
        RECT 607.270 18.940 607.590 19.000 ;
        RECT 598.085 18.800 607.590 18.940 ;
        RECT 598.085 18.755 598.375 18.800 ;
        RECT 607.270 18.740 607.590 18.800 ;
      LAYER via ;
        RECT 610.520 246.200 610.780 246.460 ;
        RECT 1342.380 246.200 1342.640 246.460 ;
        RECT 192.380 20.100 192.640 20.360 ;
        RECT 607.300 20.100 607.560 20.360 ;
        RECT 610.520 20.100 610.780 20.360 ;
        RECT 607.300 18.740 607.560 19.000 ;
      LAYER met2 ;
        RECT 1342.330 260.000 1342.610 264.000 ;
        RECT 1342.440 246.490 1342.580 260.000 ;
        RECT 610.520 246.170 610.780 246.490 ;
        RECT 1342.380 246.170 1342.640 246.490 ;
        RECT 610.580 20.390 610.720 246.170 ;
        RECT 192.380 20.070 192.640 20.390 ;
        RECT 607.300 20.070 607.560 20.390 ;
        RECT 610.520 20.070 610.780 20.390 ;
        RECT 192.440 10.610 192.580 20.070 ;
        RECT 607.360 19.030 607.500 20.070 ;
        RECT 607.300 18.710 607.560 19.030 ;
        RECT 192.440 10.470 193.040 10.610 ;
        RECT 192.900 2.400 193.040 10.470 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1642.345 247.605 1642.515 248.455 ;
      LAYER mcon ;
        RECT 1642.345 248.285 1642.515 248.455 ;
      LAYER met1 ;
        RECT 1617.890 248.440 1618.210 248.500 ;
        RECT 1642.285 248.440 1642.575 248.485 ;
        RECT 1617.890 248.300 1642.575 248.440 ;
        RECT 1617.890 248.240 1618.210 248.300 ;
        RECT 1642.285 248.255 1642.575 248.300 ;
        RECT 1796.830 248.100 1797.150 248.160 ;
        RECT 1704.460 247.960 1797.150 248.100 ;
        RECT 1642.285 247.760 1642.575 247.805 ;
        RECT 1704.460 247.760 1704.600 247.960 ;
        RECT 1796.830 247.900 1797.150 247.960 ;
        RECT 1642.285 247.620 1704.600 247.760 ;
        RECT 1642.285 247.575 1642.575 247.620 ;
        RECT 213.510 94.420 213.830 94.480 ;
        RECT 1617.890 94.420 1618.210 94.480 ;
        RECT 213.510 94.280 1618.210 94.420 ;
        RECT 213.510 94.220 213.830 94.280 ;
        RECT 1617.890 94.220 1618.210 94.280 ;
        RECT 210.750 17.580 211.070 17.640 ;
        RECT 213.510 17.580 213.830 17.640 ;
        RECT 210.750 17.440 213.830 17.580 ;
        RECT 210.750 17.380 211.070 17.440 ;
        RECT 213.510 17.380 213.830 17.440 ;
      LAYER via ;
        RECT 1617.920 248.240 1618.180 248.500 ;
        RECT 1796.860 247.900 1797.120 248.160 ;
        RECT 213.540 94.220 213.800 94.480 ;
        RECT 1617.920 94.220 1618.180 94.480 ;
        RECT 210.780 17.380 211.040 17.640 ;
        RECT 213.540 17.380 213.800 17.640 ;
      LAYER met2 ;
        RECT 1799.570 260.170 1799.850 264.000 ;
        RECT 1796.920 260.030 1799.850 260.170 ;
        RECT 1617.920 248.210 1618.180 248.530 ;
        RECT 1617.980 94.510 1618.120 248.210 ;
        RECT 1796.920 248.190 1797.060 260.030 ;
        RECT 1799.570 260.000 1799.850 260.030 ;
        RECT 1796.860 247.870 1797.120 248.190 ;
        RECT 213.540 94.190 213.800 94.510 ;
        RECT 1617.920 94.190 1618.180 94.510 ;
        RECT 213.600 17.670 213.740 94.190 ;
        RECT 210.780 17.350 211.040 17.670 ;
        RECT 213.540 17.350 213.800 17.670 ;
        RECT 210.840 2.400 210.980 17.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 230.990 2201.400 231.310 2201.460 ;
        RECT 296.770 2201.400 297.090 2201.460 ;
        RECT 230.990 2201.260 297.090 2201.400 ;
        RECT 230.990 2201.200 231.310 2201.260 ;
        RECT 296.770 2201.200 297.090 2201.260 ;
        RECT 228.690 17.580 229.010 17.640 ;
        RECT 230.990 17.580 231.310 17.640 ;
        RECT 228.690 17.440 231.310 17.580 ;
        RECT 228.690 17.380 229.010 17.440 ;
        RECT 230.990 17.380 231.310 17.440 ;
      LAYER via ;
        RECT 231.020 2201.200 231.280 2201.460 ;
        RECT 296.800 2201.200 297.060 2201.460 ;
        RECT 228.720 17.380 228.980 17.640 ;
        RECT 231.020 17.380 231.280 17.640 ;
      LAYER met2 ;
        RECT 296.790 2207.435 297.070 2207.805 ;
        RECT 296.860 2201.490 297.000 2207.435 ;
        RECT 231.020 2201.170 231.280 2201.490 ;
        RECT 296.800 2201.170 297.060 2201.490 ;
        RECT 231.080 17.670 231.220 2201.170 ;
        RECT 228.720 17.350 228.980 17.670 ;
        RECT 231.020 17.350 231.280 17.670 ;
        RECT 228.780 2.400 228.920 17.350 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 296.790 2207.480 297.070 2207.760 ;
      LAYER met3 ;
        RECT 296.765 2207.770 297.095 2207.785 ;
        RECT 310.000 2207.770 314.000 2208.160 ;
        RECT 296.765 2207.560 314.000 2207.770 ;
        RECT 296.765 2207.470 310.500 2207.560 ;
        RECT 296.765 2207.455 297.095 2207.470 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 44.780 50.530 44.840 ;
        RECT 2456.470 44.780 2456.790 44.840 ;
        RECT 50.210 44.640 2456.790 44.780 ;
        RECT 50.210 44.580 50.530 44.640 ;
        RECT 2456.470 44.580 2456.790 44.640 ;
      LAYER via ;
        RECT 50.240 44.580 50.500 44.840 ;
        RECT 2456.500 44.580 2456.760 44.840 ;
      LAYER met2 ;
        RECT 2457.370 260.170 2457.650 264.000 ;
        RECT 2456.560 260.030 2457.650 260.170 ;
        RECT 2456.560 44.870 2456.700 260.030 ;
        RECT 2457.370 260.000 2457.650 260.030 ;
        RECT 50.240 44.550 50.500 44.870 ;
        RECT 2456.500 44.550 2456.760 44.870 ;
        RECT 50.300 2.400 50.440 44.550 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.610 3275.035 1477.890 3275.405 ;
        RECT 1477.680 3260.000 1477.820 3275.035 ;
        RECT 1477.570 3256.000 1477.850 3260.000 ;
        RECT 252.630 17.155 252.910 17.525 ;
        RECT 252.700 2.400 252.840 17.155 ;
        RECT 252.490 -4.800 253.050 2.400 ;
      LAYER via2 ;
        RECT 1477.610 3275.080 1477.890 3275.360 ;
        RECT 252.630 17.200 252.910 17.480 ;
      LAYER met3 ;
        RECT 254.190 3275.370 254.570 3275.380 ;
        RECT 1477.585 3275.370 1477.915 3275.385 ;
        RECT 254.190 3275.070 1477.915 3275.370 ;
        RECT 254.190 3275.060 254.570 3275.070 ;
        RECT 1477.585 3275.055 1477.915 3275.070 ;
        RECT 252.605 17.490 252.935 17.505 ;
        RECT 254.190 17.490 254.570 17.500 ;
        RECT 252.605 17.190 254.570 17.490 ;
        RECT 252.605 17.175 252.935 17.190 ;
        RECT 254.190 17.180 254.570 17.190 ;
      LAYER via3 ;
        RECT 254.220 3275.060 254.540 3275.380 ;
        RECT 254.220 17.180 254.540 17.500 ;
      LAYER met4 ;
        RECT 254.215 3275.055 254.545 3275.385 ;
        RECT 254.230 17.505 254.530 3275.055 ;
        RECT 254.215 17.175 254.545 17.505 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 296.845 19.805 297.015 20.655 ;
      LAYER mcon ;
        RECT 296.845 20.485 297.015 20.655 ;
      LAYER met1 ;
        RECT 603.590 246.740 603.910 246.800 ;
        RECT 984.470 246.740 984.790 246.800 ;
        RECT 603.590 246.600 984.790 246.740 ;
        RECT 603.590 246.540 603.910 246.600 ;
        RECT 984.470 246.540 984.790 246.600 ;
        RECT 296.785 20.640 297.075 20.685 ;
        RECT 296.785 20.500 598.760 20.640 ;
        RECT 296.785 20.455 297.075 20.500 ;
        RECT 598.620 20.300 598.760 20.500 ;
        RECT 603.590 20.300 603.910 20.360 ;
        RECT 598.620 20.160 603.910 20.300 ;
        RECT 603.590 20.100 603.910 20.160 ;
        RECT 270.090 19.960 270.410 20.020 ;
        RECT 296.785 19.960 297.075 20.005 ;
        RECT 270.090 19.820 297.075 19.960 ;
        RECT 270.090 19.760 270.410 19.820 ;
        RECT 296.785 19.775 297.075 19.820 ;
      LAYER via ;
        RECT 603.620 246.540 603.880 246.800 ;
        RECT 984.500 246.540 984.760 246.800 ;
        RECT 603.620 20.100 603.880 20.360 ;
        RECT 270.120 19.760 270.380 20.020 ;
      LAYER met2 ;
        RECT 984.450 260.000 984.730 264.000 ;
        RECT 984.560 246.830 984.700 260.000 ;
        RECT 603.620 246.510 603.880 246.830 ;
        RECT 984.500 246.510 984.760 246.830 ;
        RECT 603.680 20.390 603.820 246.510 ;
        RECT 603.620 20.070 603.880 20.390 ;
        RECT 270.120 19.730 270.380 20.050 ;
        RECT 270.180 2.400 270.320 19.730 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 300.910 3273.080 301.230 3273.140 ;
        RECT 1034.150 3273.080 1034.470 3273.140 ;
        RECT 300.910 3272.940 1034.470 3273.080 ;
        RECT 300.910 3272.880 301.230 3272.940 ;
        RECT 1034.150 3272.880 1034.470 3272.940 ;
        RECT 285.270 982.840 285.590 982.900 ;
        RECT 300.910 982.840 301.230 982.900 ;
        RECT 285.270 982.700 301.230 982.840 ;
        RECT 285.270 982.640 285.590 982.700 ;
        RECT 300.910 982.640 301.230 982.700 ;
        RECT 285.270 20.640 285.590 20.700 ;
        RECT 288.030 20.640 288.350 20.700 ;
        RECT 285.270 20.500 288.350 20.640 ;
        RECT 285.270 20.440 285.590 20.500 ;
        RECT 288.030 20.440 288.350 20.500 ;
      LAYER via ;
        RECT 300.940 3272.880 301.200 3273.140 ;
        RECT 1034.180 3272.880 1034.440 3273.140 ;
        RECT 285.300 982.640 285.560 982.900 ;
        RECT 300.940 982.640 301.200 982.900 ;
        RECT 285.300 20.440 285.560 20.700 ;
        RECT 288.060 20.440 288.320 20.700 ;
      LAYER met2 ;
        RECT 300.940 3272.850 301.200 3273.170 ;
        RECT 1034.180 3272.850 1034.440 3273.170 ;
        RECT 301.000 982.930 301.140 3272.850 ;
        RECT 1034.240 3260.000 1034.380 3272.850 ;
        RECT 1034.130 3256.000 1034.410 3260.000 ;
        RECT 285.300 982.610 285.560 982.930 ;
        RECT 300.940 982.610 301.200 982.930 ;
        RECT 285.360 20.730 285.500 982.610 ;
        RECT 285.300 20.410 285.560 20.730 ;
        RECT 288.060 20.410 288.320 20.730 ;
        RECT 288.120 2.400 288.260 20.410 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 213.510 3269.000 213.830 3269.060 ;
        RECT 2192.430 3269.000 2192.750 3269.060 ;
        RECT 213.510 3268.860 2192.750 3269.000 ;
        RECT 213.510 3268.800 213.830 3268.860 ;
        RECT 2192.430 3268.800 2192.750 3268.860 ;
        RECT 213.510 252.180 213.830 252.240 ;
        RECT 303.670 252.180 303.990 252.240 ;
        RECT 213.510 252.040 303.990 252.180 ;
        RECT 213.510 251.980 213.830 252.040 ;
        RECT 303.670 251.980 303.990 252.040 ;
        RECT 303.670 16.220 303.990 16.280 ;
        RECT 305.970 16.220 306.290 16.280 ;
        RECT 303.670 16.080 306.290 16.220 ;
        RECT 303.670 16.020 303.990 16.080 ;
        RECT 305.970 16.020 306.290 16.080 ;
      LAYER via ;
        RECT 213.540 3268.800 213.800 3269.060 ;
        RECT 2192.460 3268.800 2192.720 3269.060 ;
        RECT 213.540 251.980 213.800 252.240 ;
        RECT 303.700 251.980 303.960 252.240 ;
        RECT 303.700 16.020 303.960 16.280 ;
        RECT 306.000 16.020 306.260 16.280 ;
      LAYER met2 ;
        RECT 213.540 3268.770 213.800 3269.090 ;
        RECT 2192.460 3268.770 2192.720 3269.090 ;
        RECT 213.600 252.270 213.740 3268.770 ;
        RECT 2192.520 3260.000 2192.660 3268.770 ;
        RECT 2192.410 3256.000 2192.690 3260.000 ;
        RECT 213.540 251.950 213.800 252.270 ;
        RECT 303.700 251.950 303.960 252.270 ;
        RECT 303.760 16.310 303.900 251.950 ;
        RECT 303.700 15.990 303.960 16.310 ;
        RECT 306.000 15.990 306.260 16.310 ;
        RECT 306.060 2.400 306.200 15.990 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.510 263.400 305.830 263.460 ;
        RECT 317.930 263.400 318.250 263.460 ;
        RECT 305.510 263.260 318.250 263.400 ;
        RECT 305.510 263.200 305.830 263.260 ;
        RECT 317.930 263.200 318.250 263.260 ;
        RECT 317.930 37.640 318.250 37.700 ;
        RECT 323.910 37.640 324.230 37.700 ;
        RECT 317.930 37.500 324.230 37.640 ;
        RECT 317.930 37.440 318.250 37.500 ;
        RECT 323.910 37.440 324.230 37.500 ;
      LAYER via ;
        RECT 305.540 263.200 305.800 263.460 ;
        RECT 317.960 263.200 318.220 263.460 ;
        RECT 317.960 37.440 318.220 37.700 ;
        RECT 323.940 37.440 324.200 37.700 ;
      LAYER met2 ;
        RECT 305.530 1932.715 305.810 1933.085 ;
        RECT 305.600 263.490 305.740 1932.715 ;
        RECT 305.540 263.170 305.800 263.490 ;
        RECT 317.960 263.170 318.220 263.490 ;
        RECT 318.020 37.730 318.160 263.170 ;
        RECT 317.960 37.410 318.220 37.730 ;
        RECT 323.940 37.410 324.200 37.730 ;
        RECT 324.000 2.400 324.140 37.410 ;
        RECT 323.790 -4.800 324.350 2.400 ;
      LAYER via2 ;
        RECT 305.530 1932.760 305.810 1933.040 ;
      LAYER met3 ;
        RECT 305.505 1933.050 305.835 1933.065 ;
        RECT 310.000 1933.050 314.000 1933.440 ;
        RECT 305.505 1932.840 314.000 1933.050 ;
        RECT 305.505 1932.750 310.500 1932.840 ;
        RECT 305.505 1932.735 305.835 1932.750 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 213.050 3271.720 213.370 3271.780 ;
        RECT 1162.950 3271.720 1163.270 3271.780 ;
        RECT 213.050 3271.580 1163.270 3271.720 ;
        RECT 213.050 3271.520 213.370 3271.580 ;
        RECT 1162.950 3271.520 1163.270 3271.580 ;
        RECT 213.050 261.020 213.370 261.080 ;
        RECT 338.170 261.020 338.490 261.080 ;
        RECT 213.050 260.880 338.490 261.020 ;
        RECT 213.050 260.820 213.370 260.880 ;
        RECT 338.170 260.820 338.490 260.880 ;
        RECT 338.170 18.600 338.490 18.660 ;
        RECT 341.390 18.600 341.710 18.660 ;
        RECT 338.170 18.460 341.710 18.600 ;
        RECT 338.170 18.400 338.490 18.460 ;
        RECT 341.390 18.400 341.710 18.460 ;
      LAYER via ;
        RECT 213.080 3271.520 213.340 3271.780 ;
        RECT 1162.980 3271.520 1163.240 3271.780 ;
        RECT 213.080 260.820 213.340 261.080 ;
        RECT 338.200 260.820 338.460 261.080 ;
        RECT 338.200 18.400 338.460 18.660 ;
        RECT 341.420 18.400 341.680 18.660 ;
      LAYER met2 ;
        RECT 213.080 3271.490 213.340 3271.810 ;
        RECT 1162.980 3271.490 1163.240 3271.810 ;
        RECT 213.140 261.110 213.280 3271.490 ;
        RECT 1163.040 3260.000 1163.180 3271.490 ;
        RECT 1162.930 3256.000 1163.210 3260.000 ;
        RECT 213.080 260.790 213.340 261.110 ;
        RECT 338.200 260.790 338.460 261.110 ;
        RECT 338.260 18.690 338.400 260.790 ;
        RECT 338.200 18.370 338.460 18.690 ;
        RECT 341.420 18.370 341.680 18.690 ;
        RECT 341.480 2.400 341.620 18.370 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 45.460 359.650 45.520 ;
        RECT 2525.470 45.460 2525.790 45.520 ;
        RECT 359.330 45.320 2525.790 45.460 ;
        RECT 359.330 45.260 359.650 45.320 ;
        RECT 2525.470 45.260 2525.790 45.320 ;
      LAYER via ;
        RECT 359.360 45.260 359.620 45.520 ;
        RECT 2525.500 45.260 2525.760 45.520 ;
      LAYER met2 ;
        RECT 2529.130 260.170 2529.410 264.000 ;
        RECT 2525.560 260.030 2529.410 260.170 ;
        RECT 2525.560 45.550 2525.700 260.030 ;
        RECT 2529.130 260.000 2529.410 260.030 ;
        RECT 359.360 45.230 359.620 45.550 ;
        RECT 2525.500 45.230 2525.760 45.550 ;
        RECT 359.420 2.400 359.560 45.230 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 301.830 393.280 302.150 393.340 ;
        RECT 313.790 393.280 314.110 393.340 ;
        RECT 301.830 393.140 314.110 393.280 ;
        RECT 301.830 393.080 302.150 393.140 ;
        RECT 313.790 393.080 314.110 393.140 ;
        RECT 313.790 15.880 314.110 15.940 ;
        RECT 377.270 15.880 377.590 15.940 ;
        RECT 313.790 15.740 377.590 15.880 ;
        RECT 313.790 15.680 314.110 15.740 ;
        RECT 377.270 15.680 377.590 15.740 ;
      LAYER via ;
        RECT 301.860 393.080 302.120 393.340 ;
        RECT 313.820 393.080 314.080 393.340 ;
        RECT 313.820 15.680 314.080 15.940 ;
        RECT 377.300 15.680 377.560 15.940 ;
      LAYER met2 ;
        RECT 301.850 1595.435 302.130 1595.805 ;
        RECT 301.920 393.370 302.060 1595.435 ;
        RECT 301.860 393.050 302.120 393.370 ;
        RECT 313.820 393.050 314.080 393.370 ;
        RECT 313.880 15.970 314.020 393.050 ;
        RECT 313.820 15.650 314.080 15.970 ;
        RECT 377.300 15.650 377.560 15.970 ;
        RECT 377.360 2.400 377.500 15.650 ;
        RECT 377.150 -4.800 377.710 2.400 ;
      LAYER via2 ;
        RECT 301.850 1595.480 302.130 1595.760 ;
      LAYER met3 ;
        RECT 301.825 1595.770 302.155 1595.785 ;
        RECT 310.000 1595.770 314.000 1596.160 ;
        RECT 301.825 1595.560 314.000 1595.770 ;
        RECT 301.825 1595.470 310.500 1595.560 ;
        RECT 301.825 1595.455 302.155 1595.470 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 59.060 395.530 59.120 ;
        RECT 2619.770 59.060 2620.090 59.120 ;
        RECT 395.210 58.920 2620.090 59.060 ;
        RECT 395.210 58.860 395.530 58.920 ;
        RECT 2619.770 58.860 2620.090 58.920 ;
      LAYER via ;
        RECT 395.240 58.860 395.500 59.120 ;
        RECT 2619.800 58.860 2620.060 59.120 ;
      LAYER met2 ;
        RECT 2619.790 443.515 2620.070 443.885 ;
        RECT 2619.860 59.150 2620.000 443.515 ;
        RECT 395.240 58.830 395.500 59.150 ;
        RECT 2619.800 58.830 2620.060 59.150 ;
        RECT 395.300 2.400 395.440 58.830 ;
        RECT 395.090 -4.800 395.650 2.400 ;
      LAYER via2 ;
        RECT 2619.790 443.560 2620.070 443.840 ;
      LAYER met3 ;
        RECT 2606.000 443.850 2610.000 444.240 ;
        RECT 2619.765 443.850 2620.095 443.865 ;
        RECT 2606.000 443.640 2620.095 443.850 ;
        RECT 2609.580 443.550 2620.095 443.640 ;
        RECT 2619.765 443.535 2620.095 443.550 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1238.390 247.760 1238.710 247.820 ;
        RECT 1570.510 247.760 1570.830 247.820 ;
        RECT 1238.390 247.620 1570.830 247.760 ;
        RECT 1238.390 247.560 1238.710 247.620 ;
        RECT 1570.510 247.560 1570.830 247.620 ;
        RECT 413.150 101.220 413.470 101.280 ;
        RECT 1238.390 101.220 1238.710 101.280 ;
        RECT 413.150 101.080 1238.710 101.220 ;
        RECT 413.150 101.020 413.470 101.080 ;
        RECT 1238.390 101.020 1238.710 101.080 ;
      LAYER via ;
        RECT 1238.420 247.560 1238.680 247.820 ;
        RECT 1570.540 247.560 1570.800 247.820 ;
        RECT 413.180 101.020 413.440 101.280 ;
        RECT 1238.420 101.020 1238.680 101.280 ;
      LAYER met2 ;
        RECT 1570.490 260.000 1570.770 264.000 ;
        RECT 1570.600 247.850 1570.740 260.000 ;
        RECT 1238.420 247.530 1238.680 247.850 ;
        RECT 1570.540 247.530 1570.800 247.850 ;
        RECT 1238.480 101.310 1238.620 247.530 ;
        RECT 413.180 100.990 413.440 101.310 ;
        RECT 1238.420 100.990 1238.680 101.310 ;
        RECT 413.240 2.400 413.380 100.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 1042.000 75.830 1042.060 ;
        RECT 296.770 1042.000 297.090 1042.060 ;
        RECT 75.510 1041.860 297.090 1042.000 ;
        RECT 75.510 1041.800 75.830 1041.860 ;
        RECT 296.770 1041.800 297.090 1041.860 ;
      LAYER via ;
        RECT 75.540 1041.800 75.800 1042.060 ;
        RECT 296.800 1041.800 297.060 1042.060 ;
      LAYER met2 ;
        RECT 296.790 1045.995 297.070 1046.365 ;
        RECT 296.860 1042.090 297.000 1045.995 ;
        RECT 75.540 1041.770 75.800 1042.090 ;
        RECT 296.800 1041.770 297.060 1042.090 ;
        RECT 75.600 17.410 75.740 1041.770 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 296.790 1046.040 297.070 1046.320 ;
      LAYER met3 ;
        RECT 296.765 1046.330 297.095 1046.345 ;
        RECT 310.000 1046.330 314.000 1046.720 ;
        RECT 296.765 1046.120 314.000 1046.330 ;
        RECT 296.765 1046.030 310.500 1046.120 ;
        RECT 296.765 1046.015 297.095 1046.030 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 307.810 244.700 308.130 244.760 ;
        RECT 427.870 244.700 428.190 244.760 ;
        RECT 307.810 244.560 428.190 244.700 ;
        RECT 307.810 244.500 308.130 244.560 ;
        RECT 427.870 244.500 428.190 244.560 ;
        RECT 427.870 2.960 428.190 3.020 ;
        RECT 430.630 2.960 430.950 3.020 ;
        RECT 427.870 2.820 430.950 2.960 ;
        RECT 427.870 2.760 428.190 2.820 ;
        RECT 430.630 2.760 430.950 2.820 ;
      LAYER via ;
        RECT 307.840 244.500 308.100 244.760 ;
        RECT 427.900 244.500 428.160 244.760 ;
        RECT 427.900 2.760 428.160 3.020 ;
        RECT 430.660 2.760 430.920 3.020 ;
      LAYER met2 ;
        RECT 307.830 3243.755 308.110 3244.125 ;
        RECT 307.900 244.790 308.040 3243.755 ;
        RECT 307.840 244.470 308.100 244.790 ;
        RECT 427.900 244.470 428.160 244.790 ;
        RECT 427.960 3.050 428.100 244.470 ;
        RECT 427.900 2.730 428.160 3.050 ;
        RECT 430.660 2.730 430.920 3.050 ;
        RECT 430.720 2.400 430.860 2.730 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 307.830 3243.800 308.110 3244.080 ;
      LAYER met3 ;
        RECT 307.805 3244.090 308.135 3244.105 ;
        RECT 310.000 3244.090 314.000 3244.480 ;
        RECT 307.805 3243.880 314.000 3244.090 ;
        RECT 307.805 3243.790 310.500 3243.880 ;
        RECT 307.805 3243.775 308.135 3243.790 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 455.010 210.700 455.330 210.760 ;
        RECT 2698.890 210.700 2699.210 210.760 ;
        RECT 455.010 210.560 2699.210 210.700 ;
        RECT 455.010 210.500 455.330 210.560 ;
        RECT 2698.890 210.500 2699.210 210.560 ;
        RECT 448.570 14.860 448.890 14.920 ;
        RECT 455.010 14.860 455.330 14.920 ;
        RECT 448.570 14.720 455.330 14.860 ;
        RECT 448.570 14.660 448.890 14.720 ;
        RECT 455.010 14.660 455.330 14.720 ;
      LAYER via ;
        RECT 455.040 210.500 455.300 210.760 ;
        RECT 2698.920 210.500 2699.180 210.760 ;
        RECT 448.600 14.660 448.860 14.920 ;
        RECT 455.040 14.660 455.300 14.920 ;
      LAYER met2 ;
        RECT 2535.610 3271.635 2535.890 3272.005 ;
        RECT 2698.910 3271.635 2699.190 3272.005 ;
        RECT 2535.680 3260.000 2535.820 3271.635 ;
        RECT 2535.570 3256.000 2535.850 3260.000 ;
        RECT 2698.980 210.790 2699.120 3271.635 ;
        RECT 455.040 210.470 455.300 210.790 ;
        RECT 2698.920 210.470 2699.180 210.790 ;
        RECT 455.100 14.950 455.240 210.470 ;
        RECT 448.600 14.630 448.860 14.950 ;
        RECT 455.040 14.630 455.300 14.950 ;
        RECT 448.660 2.400 448.800 14.630 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 2535.610 3271.680 2535.890 3271.960 ;
        RECT 2698.910 3271.680 2699.190 3271.960 ;
      LAYER met3 ;
        RECT 2535.585 3271.970 2535.915 3271.985 ;
        RECT 2698.885 3271.970 2699.215 3271.985 ;
        RECT 2535.585 3271.670 2699.215 3271.970 ;
        RECT 2535.585 3271.655 2535.915 3271.670 ;
        RECT 2698.885 3271.655 2699.215 3271.670 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 483.145 16.065 483.315 19.635 ;
      LAYER mcon ;
        RECT 483.145 19.465 483.315 19.635 ;
      LAYER met1 ;
        RECT 1707.590 241.640 1707.910 241.700 ;
        RECT 1714.030 241.640 1714.350 241.700 ;
        RECT 1707.590 241.500 1714.350 241.640 ;
        RECT 1707.590 241.440 1707.910 241.500 ;
        RECT 1714.030 241.440 1714.350 241.500 ;
        RECT 483.085 19.620 483.375 19.665 ;
        RECT 1707.590 19.620 1707.910 19.680 ;
        RECT 483.085 19.480 1707.910 19.620 ;
        RECT 483.085 19.435 483.375 19.480 ;
        RECT 1707.590 19.420 1707.910 19.480 ;
        RECT 466.510 16.220 466.830 16.280 ;
        RECT 483.085 16.220 483.375 16.265 ;
        RECT 466.510 16.080 483.375 16.220 ;
        RECT 466.510 16.020 466.830 16.080 ;
        RECT 483.085 16.035 483.375 16.080 ;
      LAYER via ;
        RECT 1707.620 241.440 1707.880 241.700 ;
        RECT 1714.060 241.440 1714.320 241.700 ;
        RECT 1707.620 19.420 1707.880 19.680 ;
        RECT 466.540 16.020 466.800 16.280 ;
      LAYER met2 ;
        RECT 1714.010 260.000 1714.290 264.000 ;
        RECT 1714.120 241.730 1714.260 260.000 ;
        RECT 1707.620 241.410 1707.880 241.730 ;
        RECT 1714.060 241.410 1714.320 241.730 ;
        RECT 1707.680 19.710 1707.820 241.410 ;
        RECT 1707.620 19.390 1707.880 19.710 ;
        RECT 466.540 15.990 466.800 16.310 ;
        RECT 466.600 2.400 466.740 15.990 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.510 244.700 489.830 244.760 ;
        RECT 567.710 244.700 568.030 244.760 ;
        RECT 489.510 244.560 568.030 244.700 ;
        RECT 489.510 244.500 489.830 244.560 ;
        RECT 567.710 244.500 568.030 244.560 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 489.510 15.200 489.830 15.260 ;
        RECT 484.450 15.060 489.830 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
        RECT 489.510 15.000 489.830 15.060 ;
      LAYER via ;
        RECT 489.540 244.500 489.800 244.760 ;
        RECT 567.740 244.500 568.000 244.760 ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 489.540 15.000 489.800 15.260 ;
      LAYER met2 ;
        RECT 569.530 260.170 569.810 264.000 ;
        RECT 567.800 260.030 569.810 260.170 ;
        RECT 567.800 244.790 567.940 260.030 ;
        RECT 569.530 260.000 569.810 260.030 ;
        RECT 489.540 244.470 489.800 244.790 ;
        RECT 567.740 244.470 568.000 244.790 ;
        RECT 489.600 15.290 489.740 244.470 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 489.540 14.970 489.800 15.290 ;
        RECT 484.540 2.400 484.680 14.970 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 497.330 16.560 497.650 16.620 ;
        RECT 502.390 16.560 502.710 16.620 ;
        RECT 497.330 16.420 502.710 16.560 ;
        RECT 497.330 16.360 497.650 16.420 ;
        RECT 502.390 16.360 502.710 16.420 ;
      LAYER via ;
        RECT 497.360 16.360 497.620 16.620 ;
        RECT 502.420 16.360 502.680 16.620 ;
      LAYER met2 ;
        RECT 2232.930 3256.930 2233.210 3257.045 ;
        RECT 2234.730 3256.930 2235.010 3260.000 ;
        RECT 2232.930 3256.790 2235.010 3256.930 ;
        RECT 2232.930 3256.675 2233.210 3256.790 ;
        RECT 2234.730 3256.000 2235.010 3256.790 ;
        RECT 497.350 259.235 497.630 259.605 ;
        RECT 497.420 16.650 497.560 259.235 ;
        RECT 497.360 16.330 497.620 16.650 ;
        RECT 502.420 16.330 502.680 16.650 ;
        RECT 502.480 2.400 502.620 16.330 ;
        RECT 502.270 -4.800 502.830 2.400 ;
      LAYER via2 ;
        RECT 2232.930 3256.720 2233.210 3257.000 ;
        RECT 497.350 259.280 497.630 259.560 ;
      LAYER met3 ;
        RECT 265.230 3257.010 265.610 3257.020 ;
        RECT 2232.905 3257.010 2233.235 3257.025 ;
        RECT 265.230 3256.710 2233.235 3257.010 ;
        RECT 265.230 3256.700 265.610 3256.710 ;
        RECT 2232.905 3256.695 2233.235 3256.710 ;
        RECT 265.230 259.570 265.610 259.580 ;
        RECT 497.325 259.570 497.655 259.585 ;
        RECT 265.230 259.270 497.655 259.570 ;
        RECT 265.230 259.260 265.610 259.270 ;
        RECT 497.325 259.255 497.655 259.270 ;
      LAYER via3 ;
        RECT 265.260 3256.700 265.580 3257.020 ;
        RECT 265.260 259.260 265.580 259.580 ;
      LAYER met4 ;
        RECT 265.255 3256.695 265.585 3257.025 ;
        RECT 265.270 259.585 265.570 3256.695 ;
        RECT 265.255 259.255 265.585 259.585 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 278.370 3258.120 278.690 3258.180 ;
        RECT 617.390 3258.120 617.710 3258.180 ;
        RECT 278.370 3257.980 617.710 3258.120 ;
        RECT 278.370 3257.920 278.690 3257.980 ;
        RECT 617.390 3257.920 617.710 3257.980 ;
        RECT 278.370 263.740 278.690 263.800 ;
        RECT 517.570 263.740 517.890 263.800 ;
        RECT 278.370 263.600 517.890 263.740 ;
        RECT 278.370 263.540 278.690 263.600 ;
        RECT 517.570 263.540 517.890 263.600 ;
        RECT 517.570 16.560 517.890 16.620 ;
        RECT 519.870 16.560 520.190 16.620 ;
        RECT 517.570 16.420 520.190 16.560 ;
        RECT 517.570 16.360 517.890 16.420 ;
        RECT 519.870 16.360 520.190 16.420 ;
      LAYER via ;
        RECT 278.400 3257.920 278.660 3258.180 ;
        RECT 617.420 3257.920 617.680 3258.180 ;
        RECT 278.400 263.540 278.660 263.800 ;
        RECT 517.600 263.540 517.860 263.800 ;
        RECT 517.600 16.360 517.860 16.620 ;
        RECT 519.900 16.360 520.160 16.620 ;
      LAYER met2 ;
        RECT 619.210 3258.290 619.490 3260.000 ;
        RECT 617.480 3258.210 619.490 3258.290 ;
        RECT 278.400 3257.890 278.660 3258.210 ;
        RECT 617.420 3258.150 619.490 3258.210 ;
        RECT 617.420 3257.890 617.680 3258.150 ;
        RECT 278.460 263.830 278.600 3257.890 ;
        RECT 619.210 3256.000 619.490 3258.150 ;
        RECT 278.400 263.510 278.660 263.830 ;
        RECT 517.600 263.510 517.860 263.830 ;
        RECT 517.660 16.650 517.800 263.510 ;
        RECT 517.600 16.330 517.860 16.650 ;
        RECT 519.900 16.330 520.160 16.650 ;
        RECT 519.960 2.400 520.100 16.330 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 253.990 3261.180 254.310 3261.240 ;
        RECT 948.590 3261.180 948.910 3261.240 ;
        RECT 253.990 3261.040 948.910 3261.180 ;
        RECT 253.990 3260.980 254.310 3261.040 ;
        RECT 948.590 3260.980 948.910 3261.040 ;
        RECT 253.990 245.380 254.310 245.440 ;
        RECT 531.830 245.380 532.150 245.440 ;
        RECT 253.990 245.240 532.150 245.380 ;
        RECT 253.990 245.180 254.310 245.240 ;
        RECT 531.830 245.180 532.150 245.240 ;
        RECT 531.830 16.560 532.150 16.620 ;
        RECT 537.810 16.560 538.130 16.620 ;
        RECT 531.830 16.420 538.130 16.560 ;
        RECT 531.830 16.360 532.150 16.420 ;
        RECT 537.810 16.360 538.130 16.420 ;
      LAYER via ;
        RECT 254.020 3260.980 254.280 3261.240 ;
        RECT 948.620 3260.980 948.880 3261.240 ;
        RECT 254.020 245.180 254.280 245.440 ;
        RECT 531.860 245.180 532.120 245.440 ;
        RECT 531.860 16.360 532.120 16.620 ;
        RECT 537.840 16.360 538.100 16.620 ;
      LAYER met2 ;
        RECT 254.020 3260.950 254.280 3261.270 ;
        RECT 948.620 3260.950 948.880 3261.270 ;
        RECT 254.080 245.470 254.220 3260.950 ;
        RECT 948.680 3260.000 948.820 3260.950 ;
        RECT 948.570 3256.000 948.850 3260.000 ;
        RECT 254.020 245.150 254.280 245.470 ;
        RECT 531.860 245.150 532.120 245.470 ;
        RECT 531.920 16.650 532.060 245.150 ;
        RECT 531.860 16.330 532.120 16.650 ;
        RECT 537.840 16.330 538.100 16.650 ;
        RECT 537.900 2.400 538.040 16.330 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 569.090 244.700 569.410 244.760 ;
        RECT 641.310 244.700 641.630 244.760 ;
        RECT 569.090 244.560 641.630 244.700 ;
        RECT 569.090 244.500 569.410 244.560 ;
        RECT 641.310 244.500 641.630 244.560 ;
        RECT 555.750 18.940 556.070 19.000 ;
        RECT 569.090 18.940 569.410 19.000 ;
        RECT 555.750 18.800 569.410 18.940 ;
        RECT 555.750 18.740 556.070 18.800 ;
        RECT 569.090 18.740 569.410 18.800 ;
      LAYER via ;
        RECT 569.120 244.500 569.380 244.760 ;
        RECT 641.340 244.500 641.600 244.760 ;
        RECT 555.780 18.740 556.040 19.000 ;
        RECT 569.120 18.740 569.380 19.000 ;
      LAYER met2 ;
        RECT 641.290 260.000 641.570 264.000 ;
        RECT 641.400 244.790 641.540 260.000 ;
        RECT 569.120 244.470 569.380 244.790 ;
        RECT 641.340 244.470 641.600 244.790 ;
        RECT 569.180 19.030 569.320 244.470 ;
        RECT 555.780 18.710 556.040 19.030 ;
        RECT 569.120 18.710 569.380 19.030 ;
        RECT 555.840 2.400 555.980 18.710 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.710 17.155 573.990 17.525 ;
        RECT 573.780 2.400 573.920 17.155 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 573.710 17.200 573.990 17.480 ;
      LAYER met3 ;
        RECT 2606.000 1881.370 2610.000 1881.760 ;
        RECT 2645.270 1881.370 2645.650 1881.380 ;
        RECT 2606.000 1881.160 2645.650 1881.370 ;
        RECT 2609.580 1881.070 2645.650 1881.160 ;
        RECT 2645.270 1881.060 2645.650 1881.070 ;
        RECT 573.685 17.490 574.015 17.505 ;
        RECT 2645.270 17.490 2645.650 17.500 ;
        RECT 573.685 17.190 2645.650 17.490 ;
        RECT 573.685 17.175 574.015 17.190 ;
        RECT 2645.270 17.180 2645.650 17.190 ;
      LAYER via3 ;
        RECT 2645.300 1881.060 2645.620 1881.380 ;
        RECT 2645.300 17.180 2645.620 17.500 ;
      LAYER met4 ;
        RECT 2645.295 1881.055 2645.625 1881.385 ;
        RECT 2645.310 17.505 2645.610 1881.055 ;
        RECT 2645.295 17.175 2645.625 17.505 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 734.765 244.545 734.935 247.095 ;
      LAYER mcon ;
        RECT 734.765 246.925 734.935 247.095 ;
      LAYER met1 ;
        RECT 734.705 247.080 734.995 247.125 ;
        RECT 999.190 247.080 999.510 247.140 ;
        RECT 734.705 246.940 999.510 247.080 ;
        RECT 734.705 246.895 734.995 246.940 ;
        RECT 999.190 246.880 999.510 246.940 ;
        RECT 686.390 244.700 686.710 244.760 ;
        RECT 734.705 244.700 734.995 244.745 ;
        RECT 686.390 244.560 734.995 244.700 ;
        RECT 686.390 244.500 686.710 244.560 ;
        RECT 734.705 244.515 734.995 244.560 ;
        RECT 685.930 16.560 686.250 16.620 ;
        RECT 629.440 16.420 686.250 16.560 ;
        RECT 591.170 16.220 591.490 16.280 ;
        RECT 629.440 16.220 629.580 16.420 ;
        RECT 685.930 16.360 686.250 16.420 ;
        RECT 591.170 16.080 629.580 16.220 ;
        RECT 591.170 16.020 591.490 16.080 ;
      LAYER via ;
        RECT 999.220 246.880 999.480 247.140 ;
        RECT 686.420 244.500 686.680 244.760 ;
        RECT 591.200 16.020 591.460 16.280 ;
        RECT 685.960 16.360 686.220 16.620 ;
      LAYER met2 ;
        RECT 999.170 260.000 999.450 264.000 ;
        RECT 999.280 247.170 999.420 260.000 ;
        RECT 999.220 246.850 999.480 247.170 ;
        RECT 686.420 244.470 686.680 244.790 ;
        RECT 686.480 26.250 686.620 244.470 ;
        RECT 686.020 26.110 686.620 26.250 ;
        RECT 686.020 16.650 686.160 26.110 ;
        RECT 685.960 16.330 686.220 16.650 ;
        RECT 591.200 15.990 591.460 16.310 ;
        RECT 591.260 2.400 591.400 15.990 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1555.790 247.420 1556.110 247.480 ;
        RECT 1956.910 247.420 1957.230 247.480 ;
        RECT 1555.790 247.280 1957.230 247.420 ;
        RECT 1555.790 247.220 1556.110 247.280 ;
        RECT 1956.910 247.220 1957.230 247.280 ;
        RECT 97.590 19.280 97.910 19.340 ;
        RECT 1555.790 19.280 1556.110 19.340 ;
        RECT 97.590 19.140 1556.110 19.280 ;
        RECT 97.590 19.080 97.910 19.140 ;
        RECT 1555.790 19.080 1556.110 19.140 ;
      LAYER via ;
        RECT 1555.820 247.220 1556.080 247.480 ;
        RECT 1956.940 247.220 1957.200 247.480 ;
        RECT 97.620 19.080 97.880 19.340 ;
        RECT 1555.820 19.080 1556.080 19.340 ;
      LAYER met2 ;
        RECT 1956.890 260.000 1957.170 264.000 ;
        RECT 1957.000 247.510 1957.140 260.000 ;
        RECT 1555.820 247.190 1556.080 247.510 ;
        RECT 1956.940 247.190 1957.200 247.510 ;
        RECT 1555.880 19.370 1556.020 247.190 ;
        RECT 97.620 19.050 97.880 19.370 ;
        RECT 1555.820 19.050 1556.080 19.370 ;
        RECT 97.680 2.400 97.820 19.050 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2155.245 17.765 2155.415 18.955 ;
      LAYER mcon ;
        RECT 2155.245 18.785 2155.415 18.955 ;
      LAYER met1 ;
        RECT 2176.790 243.680 2177.110 243.740 ;
        RECT 2185.990 243.680 2186.310 243.740 ;
        RECT 2176.790 243.540 2186.310 243.680 ;
        RECT 2176.790 243.480 2177.110 243.540 ;
        RECT 2185.990 243.480 2186.310 243.540 ;
        RECT 609.110 18.940 609.430 19.000 ;
        RECT 2155.185 18.940 2155.475 18.985 ;
        RECT 609.110 18.800 2155.475 18.940 ;
        RECT 609.110 18.740 609.430 18.800 ;
        RECT 2155.185 18.755 2155.475 18.800 ;
        RECT 2155.185 17.920 2155.475 17.965 ;
        RECT 2176.790 17.920 2177.110 17.980 ;
        RECT 2155.185 17.780 2177.110 17.920 ;
        RECT 2155.185 17.735 2155.475 17.780 ;
        RECT 2176.790 17.720 2177.110 17.780 ;
      LAYER via ;
        RECT 2176.820 243.480 2177.080 243.740 ;
        RECT 2186.020 243.480 2186.280 243.740 ;
        RECT 609.140 18.740 609.400 19.000 ;
        RECT 2176.820 17.720 2177.080 17.980 ;
      LAYER met2 ;
        RECT 2185.970 260.000 2186.250 264.000 ;
        RECT 2186.080 243.770 2186.220 260.000 ;
        RECT 2176.820 243.450 2177.080 243.770 ;
        RECT 2186.020 243.450 2186.280 243.770 ;
        RECT 609.140 18.710 609.400 19.030 ;
        RECT 609.200 2.400 609.340 18.710 ;
        RECT 2176.880 18.010 2177.020 243.450 ;
        RECT 2176.820 17.690 2177.080 18.010 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 302.290 262.720 302.610 262.780 ;
        RECT 320.690 262.720 321.010 262.780 ;
        RECT 302.290 262.580 321.010 262.720 ;
        RECT 302.290 262.520 302.610 262.580 ;
        RECT 320.690 262.520 321.010 262.580 ;
        RECT 320.690 16.900 321.010 16.960 ;
        RECT 627.050 16.900 627.370 16.960 ;
        RECT 320.690 16.760 627.370 16.900 ;
        RECT 320.690 16.700 321.010 16.760 ;
        RECT 627.050 16.700 627.370 16.760 ;
      LAYER via ;
        RECT 302.320 262.520 302.580 262.780 ;
        RECT 320.720 262.520 320.980 262.780 ;
        RECT 320.720 16.700 320.980 16.960 ;
        RECT 627.080 16.700 627.340 16.960 ;
      LAYER met2 ;
        RECT 302.310 2123.115 302.590 2123.485 ;
        RECT 302.380 262.810 302.520 2123.115 ;
        RECT 302.320 262.490 302.580 262.810 ;
        RECT 320.720 262.490 320.980 262.810 ;
        RECT 320.780 16.990 320.920 262.490 ;
        RECT 320.720 16.670 320.980 16.990 ;
        RECT 627.080 16.670 627.340 16.990 ;
        RECT 627.140 2.400 627.280 16.670 ;
        RECT 626.930 -4.800 627.490 2.400 ;
      LAYER via2 ;
        RECT 302.310 2123.160 302.590 2123.440 ;
      LAYER met3 ;
        RECT 302.285 2123.450 302.615 2123.465 ;
        RECT 310.000 2123.450 314.000 2123.840 ;
        RECT 302.285 2123.240 314.000 2123.450 ;
        RECT 302.285 2123.150 310.500 2123.240 ;
        RECT 302.285 2123.135 302.615 2123.150 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 123.810 3273.420 124.130 3273.480 ;
        RECT 805.070 3273.420 805.390 3273.480 ;
        RECT 123.810 3273.280 805.390 3273.420 ;
        RECT 123.810 3273.220 124.130 3273.280 ;
        RECT 805.070 3273.220 805.390 3273.280 ;
        RECT 121.510 16.900 121.830 16.960 ;
        RECT 123.810 16.900 124.130 16.960 ;
        RECT 121.510 16.760 124.130 16.900 ;
        RECT 121.510 16.700 121.830 16.760 ;
        RECT 123.810 16.700 124.130 16.760 ;
      LAYER via ;
        RECT 123.840 3273.220 124.100 3273.480 ;
        RECT 805.100 3273.220 805.360 3273.480 ;
        RECT 121.540 16.700 121.800 16.960 ;
        RECT 123.840 16.700 124.100 16.960 ;
      LAYER met2 ;
        RECT 123.840 3273.190 124.100 3273.510 ;
        RECT 805.100 3273.190 805.360 3273.510 ;
        RECT 123.900 16.990 124.040 3273.190 ;
        RECT 805.160 3260.000 805.300 3273.190 ;
        RECT 805.050 3256.000 805.330 3260.000 ;
        RECT 121.540 16.670 121.800 16.990 ;
        RECT 123.840 16.670 124.100 16.990 ;
        RECT 121.600 2.400 121.740 16.670 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 734.690 244.020 735.010 244.080 ;
        RECT 755.390 244.020 755.710 244.080 ;
        RECT 734.690 243.880 755.710 244.020 ;
        RECT 734.690 243.820 735.010 243.880 ;
        RECT 755.390 243.820 755.710 243.880 ;
        RECT 150.950 79.460 151.270 79.520 ;
        RECT 734.690 79.460 735.010 79.520 ;
        RECT 150.950 79.320 735.010 79.460 ;
        RECT 150.950 79.260 151.270 79.320 ;
        RECT 734.690 79.260 735.010 79.320 ;
        RECT 145.430 17.580 145.750 17.640 ;
        RECT 150.950 17.580 151.270 17.640 ;
        RECT 145.430 17.440 151.270 17.580 ;
        RECT 145.430 17.380 145.750 17.440 ;
        RECT 150.950 17.380 151.270 17.440 ;
      LAYER via ;
        RECT 734.720 243.820 734.980 244.080 ;
        RECT 755.420 243.820 755.680 244.080 ;
        RECT 150.980 79.260 151.240 79.520 ;
        RECT 734.720 79.260 734.980 79.520 ;
        RECT 145.460 17.380 145.720 17.640 ;
        RECT 150.980 17.380 151.240 17.640 ;
      LAYER met2 ;
        RECT 755.370 260.000 755.650 264.000 ;
        RECT 755.480 244.110 755.620 260.000 ;
        RECT 734.720 243.790 734.980 244.110 ;
        RECT 755.420 243.790 755.680 244.110 ;
        RECT 734.780 79.550 734.920 243.790 ;
        RECT 150.980 79.230 151.240 79.550 ;
        RECT 734.720 79.230 734.980 79.550 ;
        RECT 151.040 17.670 151.180 79.230 ;
        RECT 145.460 17.350 145.720 17.670 ;
        RECT 150.980 17.350 151.240 17.670 ;
        RECT 145.520 2.400 145.660 17.350 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 165.210 2180.660 165.530 2180.720 ;
        RECT 296.770 2180.660 297.090 2180.720 ;
        RECT 165.210 2180.520 297.090 2180.660 ;
        RECT 165.210 2180.460 165.530 2180.520 ;
        RECT 296.770 2180.460 297.090 2180.520 ;
      LAYER via ;
        RECT 165.240 2180.460 165.500 2180.720 ;
        RECT 296.800 2180.460 297.060 2180.720 ;
      LAYER met2 ;
        RECT 296.790 2187.035 297.070 2187.405 ;
        RECT 296.860 2180.750 297.000 2187.035 ;
        RECT 165.240 2180.430 165.500 2180.750 ;
        RECT 296.800 2180.430 297.060 2180.750 ;
        RECT 165.300 16.730 165.440 2180.430 ;
        RECT 163.460 16.590 165.440 16.730 ;
        RECT 163.460 2.400 163.600 16.590 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 296.790 2187.080 297.070 2187.360 ;
      LAYER met3 ;
        RECT 296.765 2187.370 297.095 2187.385 ;
        RECT 310.000 2187.370 314.000 2187.760 ;
        RECT 296.765 2187.160 314.000 2187.370 ;
        RECT 296.765 2187.070 310.500 2187.160 ;
        RECT 296.765 2187.055 297.095 2187.070 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 17.580 181.170 17.640 ;
        RECT 185.910 17.580 186.230 17.640 ;
        RECT 180.850 17.440 186.230 17.580 ;
        RECT 180.850 17.380 181.170 17.440 ;
        RECT 185.910 17.380 186.230 17.440 ;
      LAYER via ;
        RECT 180.880 17.380 181.140 17.640 ;
        RECT 185.940 17.380 186.200 17.640 ;
      LAYER met2 ;
        RECT 185.930 64.755 186.210 65.125 ;
        RECT 186.000 17.670 186.140 64.755 ;
        RECT 180.880 17.350 181.140 17.670 ;
        RECT 185.940 17.350 186.200 17.670 ;
        RECT 180.940 2.400 181.080 17.350 ;
        RECT 180.730 -4.800 181.290 2.400 ;
      LAYER via2 ;
        RECT 185.930 64.800 186.210 65.080 ;
      LAYER met3 ;
        RECT 2606.000 2853.770 2610.000 2854.160 ;
        RECT 2642.510 2853.770 2642.890 2853.780 ;
        RECT 2606.000 2853.560 2642.890 2853.770 ;
        RECT 2609.580 2853.470 2642.890 2853.560 ;
        RECT 2642.510 2853.460 2642.890 2853.470 ;
        RECT 185.905 65.090 186.235 65.105 ;
        RECT 2642.510 65.090 2642.890 65.100 ;
        RECT 185.905 64.790 2642.890 65.090 ;
        RECT 185.905 64.775 186.235 64.790 ;
        RECT 2642.510 64.780 2642.890 64.790 ;
      LAYER via3 ;
        RECT 2642.540 2853.460 2642.860 2853.780 ;
        RECT 2642.540 64.780 2642.860 65.100 ;
      LAYER met4 ;
        RECT 2642.535 2853.455 2642.865 2853.785 ;
        RECT 2642.550 65.105 2642.850 2853.455 ;
        RECT 2642.535 64.775 2642.865 65.105 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 3272.400 200.030 3272.460 ;
        RECT 1005.630 3272.400 1005.950 3272.460 ;
        RECT 199.710 3272.260 1005.950 3272.400 ;
        RECT 199.710 3272.200 200.030 3272.260 ;
        RECT 1005.630 3272.200 1005.950 3272.260 ;
      LAYER via ;
        RECT 199.740 3272.200 200.000 3272.460 ;
        RECT 1005.660 3272.200 1005.920 3272.460 ;
      LAYER met2 ;
        RECT 199.740 3272.170 200.000 3272.490 ;
        RECT 1005.660 3272.170 1005.920 3272.490 ;
        RECT 199.800 16.730 199.940 3272.170 ;
        RECT 1005.720 3260.000 1005.860 3272.170 ;
        RECT 1005.610 3256.000 1005.890 3260.000 ;
        RECT 198.880 16.590 199.940 16.730 ;
        RECT 198.880 2.400 199.020 16.590 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 219.490 246.060 219.810 246.120 ;
        RECT 369.910 246.060 370.230 246.120 ;
        RECT 219.490 245.920 370.230 246.060 ;
        RECT 219.490 245.860 219.810 245.920 ;
        RECT 369.910 245.860 370.230 245.920 ;
        RECT 216.730 17.580 217.050 17.640 ;
        RECT 219.490 17.580 219.810 17.640 ;
        RECT 216.730 17.440 219.810 17.580 ;
        RECT 216.730 17.380 217.050 17.440 ;
        RECT 219.490 17.380 219.810 17.440 ;
      LAYER via ;
        RECT 219.520 245.860 219.780 246.120 ;
        RECT 369.940 245.860 370.200 246.120 ;
        RECT 216.760 17.380 217.020 17.640 ;
        RECT 219.520 17.380 219.780 17.640 ;
      LAYER met2 ;
        RECT 369.890 260.000 370.170 264.000 ;
        RECT 370.000 246.150 370.140 260.000 ;
        RECT 219.520 245.830 219.780 246.150 ;
        RECT 369.940 245.830 370.200 246.150 ;
        RECT 219.580 17.670 219.720 245.830 ;
        RECT 216.760 17.350 217.020 17.670 ;
        RECT 219.520 17.350 219.780 17.670 ;
        RECT 216.820 2.400 216.960 17.350 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 257.670 828.140 257.990 828.200 ;
        RECT 296.770 828.140 297.090 828.200 ;
        RECT 257.670 828.000 297.090 828.140 ;
        RECT 257.670 827.940 257.990 828.000 ;
        RECT 296.770 827.940 297.090 828.000 ;
        RECT 234.670 20.980 234.990 21.040 ;
        RECT 257.670 20.980 257.990 21.040 ;
        RECT 234.670 20.840 257.990 20.980 ;
        RECT 234.670 20.780 234.990 20.840 ;
        RECT 257.670 20.780 257.990 20.840 ;
      LAYER via ;
        RECT 257.700 827.940 257.960 828.200 ;
        RECT 296.800 827.940 297.060 828.200 ;
        RECT 234.700 20.780 234.960 21.040 ;
        RECT 257.700 20.780 257.960 21.040 ;
      LAYER met2 ;
        RECT 296.790 833.835 297.070 834.205 ;
        RECT 296.860 828.230 297.000 833.835 ;
        RECT 257.700 827.910 257.960 828.230 ;
        RECT 296.800 827.910 297.060 828.230 ;
        RECT 257.760 21.070 257.900 827.910 ;
        RECT 234.700 20.750 234.960 21.070 ;
        RECT 257.700 20.750 257.960 21.070 ;
        RECT 234.760 2.400 234.900 20.750 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 296.790 833.880 297.070 834.160 ;
      LAYER met3 ;
        RECT 296.765 834.170 297.095 834.185 ;
        RECT 310.000 834.170 314.000 834.560 ;
        RECT 296.765 833.960 314.000 834.170 ;
        RECT 296.765 833.870 310.500 833.960 ;
        RECT 296.765 833.855 297.095 833.870 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 135.845 17.765 136.015 18.615 ;
      LAYER mcon ;
        RECT 135.845 18.445 136.015 18.615 ;
      LAYER met1 ;
        RECT 155.090 3133.000 155.410 3133.060 ;
        RECT 296.770 3133.000 297.090 3133.060 ;
        RECT 155.090 3132.860 297.090 3133.000 ;
        RECT 155.090 3132.800 155.410 3132.860 ;
        RECT 296.770 3132.800 297.090 3132.860 ;
        RECT 135.785 18.600 136.075 18.645 ;
        RECT 155.090 18.600 155.410 18.660 ;
        RECT 135.785 18.460 155.410 18.600 ;
        RECT 135.785 18.415 136.075 18.460 ;
        RECT 155.090 18.400 155.410 18.460 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 135.785 17.920 136.075 17.965 ;
        RECT 56.190 17.780 136.075 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 135.785 17.735 136.075 17.780 ;
      LAYER via ;
        RECT 155.120 3132.800 155.380 3133.060 ;
        RECT 296.800 3132.800 297.060 3133.060 ;
        RECT 155.120 18.400 155.380 18.660 ;
        RECT 56.220 17.720 56.480 17.980 ;
      LAYER met2 ;
        RECT 296.790 3137.675 297.070 3138.045 ;
        RECT 296.860 3133.090 297.000 3137.675 ;
        RECT 155.120 3132.770 155.380 3133.090 ;
        RECT 296.800 3132.770 297.060 3133.090 ;
        RECT 155.180 18.690 155.320 3132.770 ;
        RECT 155.120 18.370 155.380 18.690 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 296.790 3137.720 297.070 3138.000 ;
      LAYER met3 ;
        RECT 296.765 3138.010 297.095 3138.025 ;
        RECT 310.000 3138.010 314.000 3138.400 ;
        RECT 296.765 3137.800 314.000 3138.010 ;
        RECT 296.765 3137.710 310.500 3137.800 ;
        RECT 296.765 3137.695 297.095 3137.710 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 3272.740 82.730 3272.800 ;
        RECT 848.310 3272.740 848.630 3272.800 ;
        RECT 82.410 3272.600 848.630 3272.740 ;
        RECT 82.410 3272.540 82.730 3272.600 ;
        RECT 848.310 3272.540 848.630 3272.600 ;
        RECT 80.110 16.900 80.430 16.960 ;
        RECT 82.410 16.900 82.730 16.960 ;
        RECT 80.110 16.760 82.730 16.900 ;
        RECT 80.110 16.700 80.430 16.760 ;
        RECT 82.410 16.700 82.730 16.760 ;
      LAYER via ;
        RECT 82.440 3272.540 82.700 3272.800 ;
        RECT 848.340 3272.540 848.600 3272.800 ;
        RECT 80.140 16.700 80.400 16.960 ;
        RECT 82.440 16.700 82.700 16.960 ;
      LAYER met2 ;
        RECT 82.440 3272.510 82.700 3272.830 ;
        RECT 848.340 3272.510 848.600 3272.830 ;
        RECT 82.500 16.990 82.640 3272.510 ;
        RECT 848.400 3260.000 848.540 3272.510 ;
        RECT 848.290 3256.000 848.570 3260.000 ;
        RECT 80.140 16.670 80.400 16.990 ;
        RECT 82.440 16.670 82.700 16.990 ;
        RECT 80.200 2.400 80.340 16.670 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 489.970 3274.780 490.290 3274.840 ;
        RECT 2020.390 3274.780 2020.710 3274.840 ;
        RECT 489.970 3274.640 2020.710 3274.780 ;
        RECT 489.970 3274.580 490.290 3274.640 ;
        RECT 2020.390 3274.580 2020.710 3274.640 ;
        RECT 103.570 15.540 103.890 15.600 ;
        RECT 110.010 15.540 110.330 15.600 ;
        RECT 103.570 15.400 110.330 15.540 ;
        RECT 103.570 15.340 103.890 15.400 ;
        RECT 110.010 15.340 110.330 15.400 ;
      LAYER via ;
        RECT 490.000 3274.580 490.260 3274.840 ;
        RECT 2020.420 3274.580 2020.680 3274.840 ;
        RECT 103.600 15.340 103.860 15.600 ;
        RECT 110.040 15.340 110.300 15.600 ;
      LAYER met2 ;
        RECT 490.000 3274.550 490.260 3274.870 ;
        RECT 2020.420 3274.550 2020.680 3274.870 ;
        RECT 490.060 3271.325 490.200 3274.550 ;
        RECT 110.030 3270.955 110.310 3271.325 ;
        RECT 489.990 3270.955 490.270 3271.325 ;
        RECT 110.100 15.630 110.240 3270.955 ;
        RECT 2020.480 3260.000 2020.620 3274.550 ;
        RECT 2020.370 3256.000 2020.650 3260.000 ;
        RECT 103.600 15.310 103.860 15.630 ;
        RECT 110.040 15.310 110.300 15.630 ;
        RECT 103.660 2.400 103.800 15.310 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 110.030 3271.000 110.310 3271.280 ;
        RECT 489.990 3271.000 490.270 3271.280 ;
      LAYER met3 ;
        RECT 110.005 3271.290 110.335 3271.305 ;
        RECT 489.965 3271.290 490.295 3271.305 ;
        RECT 110.005 3270.990 490.295 3271.290 ;
        RECT 110.005 3270.975 110.335 3270.990 ;
        RECT 489.965 3270.975 490.295 3270.990 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 16.560 127.810 16.620 ;
        RECT 130.710 16.560 131.030 16.620 ;
        RECT 127.490 16.420 131.030 16.560 ;
        RECT 127.490 16.360 127.810 16.420 ;
        RECT 130.710 16.360 131.030 16.420 ;
      LAYER via ;
        RECT 127.520 16.360 127.780 16.620 ;
        RECT 130.740 16.360 131.000 16.620 ;
      LAYER met2 ;
        RECT 130.730 3272.315 131.010 3272.685 ;
        RECT 1677.250 3272.315 1677.530 3272.685 ;
        RECT 130.800 16.650 130.940 3272.315 ;
        RECT 1677.320 3260.000 1677.460 3272.315 ;
        RECT 1677.210 3256.000 1677.490 3260.000 ;
        RECT 127.520 16.330 127.780 16.650 ;
        RECT 130.740 16.330 131.000 16.650 ;
        RECT 127.580 2.400 127.720 16.330 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 130.730 3272.360 131.010 3272.640 ;
        RECT 1677.250 3272.360 1677.530 3272.640 ;
      LAYER met3 ;
        RECT 130.705 3272.650 131.035 3272.665 ;
        RECT 1677.225 3272.650 1677.555 3272.665 ;
        RECT 130.705 3272.350 1677.555 3272.650 ;
        RECT 130.705 3272.335 131.035 3272.350 ;
        RECT 1677.225 3272.335 1677.555 3272.350 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 217.190 3271.380 217.510 3271.440 ;
        RECT 518.950 3271.380 519.270 3271.440 ;
        RECT 217.190 3271.240 519.270 3271.380 ;
        RECT 217.190 3271.180 217.510 3271.240 ;
        RECT 518.950 3271.180 519.270 3271.240 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 217.190 17.240 217.510 17.300 ;
        RECT 26.290 17.100 217.510 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 217.190 17.040 217.510 17.100 ;
      LAYER via ;
        RECT 217.220 3271.180 217.480 3271.440 ;
        RECT 518.980 3271.180 519.240 3271.440 ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 217.220 17.040 217.480 17.300 ;
      LAYER met2 ;
        RECT 217.220 3271.150 217.480 3271.470 ;
        RECT 518.980 3271.150 519.240 3271.470 ;
        RECT 217.280 17.330 217.420 3271.150 ;
        RECT 519.040 3260.000 519.180 3271.150 ;
        RECT 518.930 3256.000 519.210 3260.000 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 217.220 17.010 217.480 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1755.890 246.400 1756.210 246.460 ;
        RECT 1814.310 246.400 1814.630 246.460 ;
        RECT 1755.890 246.260 1814.630 246.400 ;
        RECT 1755.890 246.200 1756.210 246.260 ;
        RECT 1814.310 246.200 1814.630 246.260 ;
        RECT 32.270 18.260 32.590 18.320 ;
        RECT 1755.890 18.260 1756.210 18.320 ;
        RECT 32.270 18.120 1756.210 18.260 ;
        RECT 32.270 18.060 32.590 18.120 ;
        RECT 1755.890 18.060 1756.210 18.120 ;
      LAYER via ;
        RECT 1755.920 246.200 1756.180 246.460 ;
        RECT 1814.340 246.200 1814.600 246.460 ;
        RECT 32.300 18.060 32.560 18.320 ;
        RECT 1755.920 18.060 1756.180 18.320 ;
      LAYER met2 ;
        RECT 1814.290 260.000 1814.570 264.000 ;
        RECT 1814.400 246.490 1814.540 260.000 ;
        RECT 1755.920 246.170 1756.180 246.490 ;
        RECT 1814.340 246.170 1814.600 246.490 ;
        RECT 1755.980 18.350 1756.120 246.170 ;
        RECT 32.300 18.030 32.560 18.350 ;
        RECT 1755.920 18.030 1756.180 18.350 ;
        RECT 32.360 2.400 32.500 18.030 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 3260.000 457.020 3528.900 ;
        RECT 634.020 3260.000 637.020 3528.900 ;
        RECT 814.020 3260.000 817.020 3528.900 ;
        RECT 994.020 3260.000 997.020 3528.900 ;
        RECT 1174.020 3260.000 1177.020 3528.900 ;
        RECT 1354.020 3260.000 1357.020 3528.900 ;
        RECT 1534.020 3260.000 1537.020 3528.900 ;
        RECT 1714.020 3260.000 1717.020 3528.900 ;
        RECT 1894.020 3260.000 1897.020 3528.900 ;
        RECT 2074.020 3260.000 2077.020 3528.900 ;
        RECT 2254.020 3260.000 2257.020 3528.900 ;
        RECT 2434.020 3260.000 2437.020 3528.900 ;
        RECT 454.020 -9.220 457.020 260.000 ;
        RECT 634.020 -9.220 637.020 260.000 ;
        RECT 814.020 -9.220 817.020 260.000 ;
        RECT 994.020 -9.220 997.020 260.000 ;
        RECT 1174.020 -9.220 1177.020 260.000 ;
        RECT 1354.020 -9.220 1357.020 260.000 ;
        RECT 1534.020 -9.220 1537.020 260.000 ;
        RECT 1714.020 -9.220 1717.020 260.000 ;
        RECT 1894.020 -9.220 1897.020 260.000 ;
        RECT 2074.020 -9.220 2077.020 260.000 ;
        RECT 2254.020 -9.220 2257.020 260.000 ;
        RECT 2434.020 -9.220 2437.020 260.000 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 3260.000 385.020 3538.100 ;
        RECT 562.020 3260.000 565.020 3538.100 ;
        RECT 742.020 3260.000 745.020 3538.100 ;
        RECT 922.020 3260.000 925.020 3538.100 ;
        RECT 1102.020 3260.000 1105.020 3538.100 ;
        RECT 1282.020 3260.000 1285.020 3538.100 ;
        RECT 1462.020 3260.000 1465.020 3538.100 ;
        RECT 1642.020 3260.000 1645.020 3538.100 ;
        RECT 1822.020 3260.000 1825.020 3538.100 ;
        RECT 2002.020 3260.000 2005.020 3538.100 ;
        RECT 2182.020 3260.000 2185.020 3538.100 ;
        RECT 2362.020 3260.000 2365.020 3538.100 ;
        RECT 2542.020 3260.000 2545.020 3538.100 ;
        RECT 382.020 -18.420 385.020 260.000 ;
        RECT 562.020 -18.420 565.020 260.000 ;
        RECT 742.020 -18.420 745.020 260.000 ;
        RECT 922.020 -18.420 925.020 260.000 ;
        RECT 1102.020 -18.420 1105.020 260.000 ;
        RECT 1282.020 -18.420 1285.020 260.000 ;
        RECT 1462.020 -18.420 1465.020 260.000 ;
        RECT 1642.020 -18.420 1645.020 260.000 ;
        RECT 1822.020 -18.420 1825.020 260.000 ;
        RECT 2002.020 -18.420 2005.020 260.000 ;
        RECT 2182.020 -18.420 2185.020 260.000 ;
        RECT 2362.020 -18.420 2365.020 260.000 ;
        RECT 2542.020 -18.420 2545.020 260.000 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 3260.000 475.020 3538.100 ;
        RECT 652.020 3260.000 655.020 3538.100 ;
        RECT 832.020 3260.000 835.020 3538.100 ;
        RECT 1012.020 3260.000 1015.020 3538.100 ;
        RECT 1192.020 3260.000 1195.020 3538.100 ;
        RECT 1372.020 3260.000 1375.020 3538.100 ;
        RECT 1552.020 3260.000 1555.020 3538.100 ;
        RECT 1732.020 3260.000 1735.020 3538.100 ;
        RECT 1912.020 3260.000 1915.020 3538.100 ;
        RECT 2092.020 3260.000 2095.020 3538.100 ;
        RECT 2272.020 3260.000 2275.020 3538.100 ;
        RECT 2452.020 3260.000 2455.020 3538.100 ;
        RECT 472.020 -18.420 475.020 260.000 ;
        RECT 652.020 -18.420 655.020 260.000 ;
        RECT 832.020 -18.420 835.020 260.000 ;
        RECT 1012.020 -18.420 1015.020 260.000 ;
        RECT 1192.020 -18.420 1195.020 260.000 ;
        RECT 1372.020 -18.420 1375.020 260.000 ;
        RECT 1552.020 -18.420 1555.020 260.000 ;
        RECT 1732.020 -18.420 1735.020 260.000 ;
        RECT 1912.020 -18.420 1915.020 260.000 ;
        RECT 2092.020 -18.420 2095.020 260.000 ;
        RECT 2272.020 -18.420 2275.020 260.000 ;
        RECT 2452.020 -18.420 2455.020 260.000 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 3260.000 403.020 3547.300 ;
        RECT 580.020 3260.000 583.020 3547.300 ;
        RECT 760.020 3260.000 763.020 3547.300 ;
        RECT 940.020 3260.000 943.020 3547.300 ;
        RECT 1120.020 3260.000 1123.020 3547.300 ;
        RECT 1300.020 3260.000 1303.020 3547.300 ;
        RECT 1480.020 3260.000 1483.020 3547.300 ;
        RECT 1660.020 3260.000 1663.020 3547.300 ;
        RECT 1840.020 3260.000 1843.020 3547.300 ;
        RECT 2020.020 3260.000 2023.020 3547.300 ;
        RECT 2200.020 3260.000 2203.020 3547.300 ;
        RECT 2380.020 3260.000 2383.020 3547.300 ;
        RECT 2560.020 3260.000 2563.020 3547.300 ;
        RECT 400.020 -27.620 403.020 260.000 ;
        RECT 580.020 -27.620 583.020 260.000 ;
        RECT 760.020 -27.620 763.020 260.000 ;
        RECT 940.020 -27.620 943.020 260.000 ;
        RECT 1120.020 -27.620 1123.020 260.000 ;
        RECT 1300.020 -27.620 1303.020 260.000 ;
        RECT 1480.020 -27.620 1483.020 260.000 ;
        RECT 1660.020 -27.620 1663.020 260.000 ;
        RECT 1840.020 -27.620 1843.020 260.000 ;
        RECT 2020.020 -27.620 2023.020 260.000 ;
        RECT 2200.020 -27.620 2203.020 260.000 ;
        RECT 2380.020 -27.620 2383.020 260.000 ;
        RECT 2560.020 -27.620 2563.020 260.000 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 3260.000 313.020 3547.300 ;
        RECT 490.020 3260.000 493.020 3547.300 ;
        RECT 670.020 3260.000 673.020 3547.300 ;
        RECT 850.020 3260.000 853.020 3547.300 ;
        RECT 1030.020 3260.000 1033.020 3547.300 ;
        RECT 1210.020 3260.000 1213.020 3547.300 ;
        RECT 1390.020 3260.000 1393.020 3547.300 ;
        RECT 1570.020 3260.000 1573.020 3547.300 ;
        RECT 1750.020 3260.000 1753.020 3547.300 ;
        RECT 1930.020 3260.000 1933.020 3547.300 ;
        RECT 2110.020 3260.000 2113.020 3547.300 ;
        RECT 2290.020 3260.000 2293.020 3547.300 ;
        RECT 2470.020 3260.000 2473.020 3547.300 ;
        RECT 310.020 -27.620 313.020 260.000 ;
        RECT 490.020 -27.620 493.020 260.000 ;
        RECT 670.020 -27.620 673.020 260.000 ;
        RECT 850.020 -27.620 853.020 260.000 ;
        RECT 1030.020 -27.620 1033.020 260.000 ;
        RECT 1210.020 -27.620 1213.020 260.000 ;
        RECT 1390.020 -27.620 1393.020 260.000 ;
        RECT 1570.020 -27.620 1573.020 260.000 ;
        RECT 1750.020 -27.620 1753.020 260.000 ;
        RECT 1930.020 -27.620 1933.020 260.000 ;
        RECT 2110.020 -27.620 2113.020 260.000 ;
        RECT 2290.020 -27.620 2293.020 260.000 ;
        RECT 2470.020 -27.620 2473.020 260.000 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 3260.000 421.020 3556.500 ;
        RECT 598.020 3260.000 601.020 3556.500 ;
        RECT 778.020 3260.000 781.020 3556.500 ;
        RECT 958.020 3260.000 961.020 3556.500 ;
        RECT 1138.020 3260.000 1141.020 3556.500 ;
        RECT 1318.020 3260.000 1321.020 3556.500 ;
        RECT 1498.020 3260.000 1501.020 3556.500 ;
        RECT 1678.020 3260.000 1681.020 3556.500 ;
        RECT 1858.020 3260.000 1861.020 3556.500 ;
        RECT 2038.020 3260.000 2041.020 3556.500 ;
        RECT 2218.020 3260.000 2221.020 3556.500 ;
        RECT 2398.020 3260.000 2401.020 3556.500 ;
        RECT 2578.020 3260.000 2581.020 3556.500 ;
        RECT 418.020 -36.820 421.020 260.000 ;
        RECT 598.020 -36.820 601.020 260.000 ;
        RECT 778.020 -36.820 781.020 260.000 ;
        RECT 958.020 -36.820 961.020 260.000 ;
        RECT 1138.020 -36.820 1141.020 260.000 ;
        RECT 1318.020 -36.820 1321.020 260.000 ;
        RECT 1498.020 -36.820 1501.020 260.000 ;
        RECT 1678.020 -36.820 1681.020 260.000 ;
        RECT 1858.020 -36.820 1861.020 260.000 ;
        RECT 2038.020 -36.820 2041.020 260.000 ;
        RECT 2218.020 -36.820 2221.020 260.000 ;
        RECT 2398.020 -36.820 2401.020 260.000 ;
        RECT 2578.020 -36.820 2581.020 260.000 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 3260.000 331.020 3556.500 ;
        RECT 508.020 3260.000 511.020 3556.500 ;
        RECT 688.020 3260.000 691.020 3556.500 ;
        RECT 868.020 3260.000 871.020 3556.500 ;
        RECT 1048.020 3260.000 1051.020 3556.500 ;
        RECT 1228.020 3260.000 1231.020 3556.500 ;
        RECT 1408.020 3260.000 1411.020 3556.500 ;
        RECT 1588.020 3260.000 1591.020 3556.500 ;
        RECT 1768.020 3260.000 1771.020 3556.500 ;
        RECT 1948.020 3260.000 1951.020 3556.500 ;
        RECT 2128.020 3260.000 2131.020 3556.500 ;
        RECT 2308.020 3260.000 2311.020 3556.500 ;
        RECT 2488.020 3260.000 2491.020 3556.500 ;
        RECT 328.020 -36.820 331.020 260.000 ;
        RECT 508.020 -36.820 511.020 260.000 ;
        RECT 688.020 -36.820 691.020 260.000 ;
        RECT 868.020 -36.820 871.020 260.000 ;
        RECT 1048.020 -36.820 1051.020 260.000 ;
        RECT 1228.020 -36.820 1231.020 260.000 ;
        RECT 1408.020 -36.820 1411.020 260.000 ;
        RECT 1588.020 -36.820 1591.020 260.000 ;
        RECT 1768.020 -36.820 1771.020 260.000 ;
        RECT 1948.020 -36.820 1951.020 260.000 ;
        RECT 2128.020 -36.820 2131.020 260.000 ;
        RECT 2308.020 -36.820 2311.020 260.000 ;
        RECT 2488.020 -36.820 2491.020 260.000 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 315.520 270.795 2604.480 3246.645 ;
      LAYER met1 ;
        RECT 315.520 264.460 2604.480 3252.300 ;
      LAYER met2 ;
        RECT 316.080 3255.720 319.010 3256.000 ;
        RECT 319.850 3255.720 332.810 3256.000 ;
        RECT 333.650 3255.720 347.530 3256.000 ;
        RECT 348.370 3255.720 361.330 3256.000 ;
        RECT 362.170 3255.720 376.050 3256.000 ;
        RECT 376.890 3255.720 389.850 3256.000 ;
        RECT 390.690 3255.720 404.570 3256.000 ;
        RECT 405.410 3255.720 418.370 3256.000 ;
        RECT 419.210 3255.720 433.090 3256.000 ;
        RECT 433.930 3255.720 446.890 3256.000 ;
        RECT 447.730 3255.720 461.610 3256.000 ;
        RECT 462.450 3255.720 476.330 3256.000 ;
        RECT 477.170 3255.720 490.130 3256.000 ;
        RECT 490.970 3255.720 504.850 3256.000 ;
        RECT 505.690 3255.720 518.650 3256.000 ;
        RECT 519.490 3255.720 533.370 3256.000 ;
        RECT 534.210 3255.720 547.170 3256.000 ;
        RECT 548.010 3255.720 561.890 3256.000 ;
        RECT 562.730 3255.720 575.690 3256.000 ;
        RECT 576.530 3255.720 590.410 3256.000 ;
        RECT 591.250 3255.720 604.210 3256.000 ;
        RECT 605.050 3255.720 618.930 3256.000 ;
        RECT 619.770 3255.720 633.650 3256.000 ;
        RECT 634.490 3255.720 647.450 3256.000 ;
        RECT 648.290 3255.720 662.170 3256.000 ;
        RECT 663.010 3255.720 675.970 3256.000 ;
        RECT 676.810 3255.720 690.690 3256.000 ;
        RECT 691.530 3255.720 704.490 3256.000 ;
        RECT 705.330 3255.720 719.210 3256.000 ;
        RECT 720.050 3255.720 733.010 3256.000 ;
        RECT 733.850 3255.720 747.730 3256.000 ;
        RECT 748.570 3255.720 761.530 3256.000 ;
        RECT 762.370 3255.720 776.250 3256.000 ;
        RECT 777.090 3255.720 790.970 3256.000 ;
        RECT 791.810 3255.720 804.770 3256.000 ;
        RECT 805.610 3255.720 819.490 3256.000 ;
        RECT 820.330 3255.720 833.290 3256.000 ;
        RECT 834.130 3255.720 848.010 3256.000 ;
        RECT 848.850 3255.720 861.810 3256.000 ;
        RECT 862.650 3255.720 876.530 3256.000 ;
        RECT 877.370 3255.720 890.330 3256.000 ;
        RECT 891.170 3255.720 905.050 3256.000 ;
        RECT 905.890 3255.720 918.850 3256.000 ;
        RECT 919.690 3255.720 933.570 3256.000 ;
        RECT 934.410 3255.720 948.290 3256.000 ;
        RECT 949.130 3255.720 962.090 3256.000 ;
        RECT 962.930 3255.720 976.810 3256.000 ;
        RECT 977.650 3255.720 990.610 3256.000 ;
        RECT 991.450 3255.720 1005.330 3256.000 ;
        RECT 1006.170 3255.720 1019.130 3256.000 ;
        RECT 1019.970 3255.720 1033.850 3256.000 ;
        RECT 1034.690 3255.720 1047.650 3256.000 ;
        RECT 1048.490 3255.720 1062.370 3256.000 ;
        RECT 1063.210 3255.720 1076.170 3256.000 ;
        RECT 1077.010 3255.720 1090.890 3256.000 ;
        RECT 1091.730 3255.720 1104.690 3256.000 ;
        RECT 1105.530 3255.720 1119.410 3256.000 ;
        RECT 1120.250 3255.720 1134.130 3256.000 ;
        RECT 1134.970 3255.720 1147.930 3256.000 ;
        RECT 1148.770 3255.720 1162.650 3256.000 ;
        RECT 1163.490 3255.720 1176.450 3256.000 ;
        RECT 1177.290 3255.720 1191.170 3256.000 ;
        RECT 1192.010 3255.720 1204.970 3256.000 ;
        RECT 1205.810 3255.720 1219.690 3256.000 ;
        RECT 1220.530 3255.720 1233.490 3256.000 ;
        RECT 1234.330 3255.720 1248.210 3256.000 ;
        RECT 1249.050 3255.720 1262.010 3256.000 ;
        RECT 1262.850 3255.720 1276.730 3256.000 ;
        RECT 1277.570 3255.720 1291.450 3256.000 ;
        RECT 1292.290 3255.720 1305.250 3256.000 ;
        RECT 1306.090 3255.720 1319.970 3256.000 ;
        RECT 1320.810 3255.720 1333.770 3256.000 ;
        RECT 1334.610 3255.720 1348.490 3256.000 ;
        RECT 1349.330 3255.720 1362.290 3256.000 ;
        RECT 1363.130 3255.720 1377.010 3256.000 ;
        RECT 1377.850 3255.720 1390.810 3256.000 ;
        RECT 1391.650 3255.720 1405.530 3256.000 ;
        RECT 1406.370 3255.720 1419.330 3256.000 ;
        RECT 1420.170 3255.720 1434.050 3256.000 ;
        RECT 1434.890 3255.720 1448.770 3256.000 ;
        RECT 1449.610 3255.720 1462.570 3256.000 ;
        RECT 1463.410 3255.720 1477.290 3256.000 ;
        RECT 1478.130 3255.720 1491.090 3256.000 ;
        RECT 1491.930 3255.720 1505.810 3256.000 ;
        RECT 1506.650 3255.720 1519.610 3256.000 ;
        RECT 1520.450 3255.720 1534.330 3256.000 ;
        RECT 1535.170 3255.720 1548.130 3256.000 ;
        RECT 1548.970 3255.720 1562.850 3256.000 ;
        RECT 1563.690 3255.720 1576.650 3256.000 ;
        RECT 1577.490 3255.720 1591.370 3256.000 ;
        RECT 1592.210 3255.720 1605.170 3256.000 ;
        RECT 1606.010 3255.720 1619.890 3256.000 ;
        RECT 1620.730 3255.720 1634.610 3256.000 ;
        RECT 1635.450 3255.720 1648.410 3256.000 ;
        RECT 1649.250 3255.720 1663.130 3256.000 ;
        RECT 1663.970 3255.720 1676.930 3256.000 ;
        RECT 1677.770 3255.720 1691.650 3256.000 ;
        RECT 1692.490 3255.720 1705.450 3256.000 ;
        RECT 1706.290 3255.720 1720.170 3256.000 ;
        RECT 1721.010 3255.720 1733.970 3256.000 ;
        RECT 1734.810 3255.720 1748.690 3256.000 ;
        RECT 1749.530 3255.720 1762.490 3256.000 ;
        RECT 1763.330 3255.720 1777.210 3256.000 ;
        RECT 1778.050 3255.720 1791.930 3256.000 ;
        RECT 1792.770 3255.720 1805.730 3256.000 ;
        RECT 1806.570 3255.720 1820.450 3256.000 ;
        RECT 1821.290 3255.720 1834.250 3256.000 ;
        RECT 1835.090 3255.720 1848.970 3256.000 ;
        RECT 1849.810 3255.720 1862.770 3256.000 ;
        RECT 1863.610 3255.720 1877.490 3256.000 ;
        RECT 1878.330 3255.720 1891.290 3256.000 ;
        RECT 1892.130 3255.720 1906.010 3256.000 ;
        RECT 1906.850 3255.720 1919.810 3256.000 ;
        RECT 1920.650 3255.720 1934.530 3256.000 ;
        RECT 1935.370 3255.720 1949.250 3256.000 ;
        RECT 1950.090 3255.720 1963.050 3256.000 ;
        RECT 1963.890 3255.720 1977.770 3256.000 ;
        RECT 1978.610 3255.720 1991.570 3256.000 ;
        RECT 1992.410 3255.720 2006.290 3256.000 ;
        RECT 2007.130 3255.720 2020.090 3256.000 ;
        RECT 2020.930 3255.720 2034.810 3256.000 ;
        RECT 2035.650 3255.720 2048.610 3256.000 ;
        RECT 2049.450 3255.720 2063.330 3256.000 ;
        RECT 2064.170 3255.720 2077.130 3256.000 ;
        RECT 2077.970 3255.720 2091.850 3256.000 ;
        RECT 2092.690 3255.720 2105.650 3256.000 ;
        RECT 2106.490 3255.720 2120.370 3256.000 ;
        RECT 2121.210 3255.720 2135.090 3256.000 ;
        RECT 2135.930 3255.720 2148.890 3256.000 ;
        RECT 2149.730 3255.720 2163.610 3256.000 ;
        RECT 2164.450 3255.720 2177.410 3256.000 ;
        RECT 2178.250 3255.720 2192.130 3256.000 ;
        RECT 2192.970 3255.720 2205.930 3256.000 ;
        RECT 2206.770 3255.720 2220.650 3256.000 ;
        RECT 2221.490 3255.720 2234.450 3256.000 ;
        RECT 2235.290 3255.720 2249.170 3256.000 ;
        RECT 2250.010 3255.720 2262.970 3256.000 ;
        RECT 2263.810 3255.720 2277.690 3256.000 ;
        RECT 2278.530 3255.720 2292.410 3256.000 ;
        RECT 2293.250 3255.720 2306.210 3256.000 ;
        RECT 2307.050 3255.720 2320.930 3256.000 ;
        RECT 2321.770 3255.720 2334.730 3256.000 ;
        RECT 2335.570 3255.720 2349.450 3256.000 ;
        RECT 2350.290 3255.720 2363.250 3256.000 ;
        RECT 2364.090 3255.720 2377.970 3256.000 ;
        RECT 2378.810 3255.720 2391.770 3256.000 ;
        RECT 2392.610 3255.720 2406.490 3256.000 ;
        RECT 2407.330 3255.720 2420.290 3256.000 ;
        RECT 2421.130 3255.720 2435.010 3256.000 ;
        RECT 2435.850 3255.720 2449.730 3256.000 ;
        RECT 2450.570 3255.720 2463.530 3256.000 ;
        RECT 2464.370 3255.720 2478.250 3256.000 ;
        RECT 2479.090 3255.720 2492.050 3256.000 ;
        RECT 2492.890 3255.720 2506.770 3256.000 ;
        RECT 2507.610 3255.720 2520.570 3256.000 ;
        RECT 2521.410 3255.720 2535.290 3256.000 ;
        RECT 2536.130 3255.720 2549.090 3256.000 ;
        RECT 2549.930 3255.720 2563.810 3256.000 ;
        RECT 2564.650 3255.720 2577.610 3256.000 ;
        RECT 2578.450 3255.720 2592.330 3256.000 ;
        RECT 2593.170 3255.720 2606.130 3256.000 ;
        RECT 316.080 264.280 2606.620 3255.720 ;
        RECT 316.080 264.000 326.370 264.280 ;
        RECT 327.210 264.000 341.090 264.280 ;
        RECT 341.930 264.000 354.890 264.280 ;
        RECT 355.730 264.000 369.610 264.280 ;
        RECT 370.450 264.000 383.410 264.280 ;
        RECT 384.250 264.000 398.130 264.280 ;
        RECT 398.970 264.000 411.930 264.280 ;
        RECT 412.770 264.000 426.650 264.280 ;
        RECT 427.490 264.000 440.450 264.280 ;
        RECT 441.290 264.000 455.170 264.280 ;
        RECT 456.010 264.000 468.970 264.280 ;
        RECT 469.810 264.000 483.690 264.280 ;
        RECT 484.530 264.000 498.410 264.280 ;
        RECT 499.250 264.000 512.210 264.280 ;
        RECT 513.050 264.000 526.930 264.280 ;
        RECT 527.770 264.000 540.730 264.280 ;
        RECT 541.570 264.000 555.450 264.280 ;
        RECT 556.290 264.000 569.250 264.280 ;
        RECT 570.090 264.000 583.970 264.280 ;
        RECT 584.810 264.000 597.770 264.280 ;
        RECT 598.610 264.000 612.490 264.280 ;
        RECT 613.330 264.000 626.290 264.280 ;
        RECT 627.130 264.000 641.010 264.280 ;
        RECT 641.850 264.000 655.730 264.280 ;
        RECT 656.570 264.000 669.530 264.280 ;
        RECT 670.370 264.000 684.250 264.280 ;
        RECT 685.090 264.000 698.050 264.280 ;
        RECT 698.890 264.000 712.770 264.280 ;
        RECT 713.610 264.000 726.570 264.280 ;
        RECT 727.410 264.000 741.290 264.280 ;
        RECT 742.130 264.000 755.090 264.280 ;
        RECT 755.930 264.000 769.810 264.280 ;
        RECT 770.650 264.000 783.610 264.280 ;
        RECT 784.450 264.000 798.330 264.280 ;
        RECT 799.170 264.000 813.050 264.280 ;
        RECT 813.890 264.000 826.850 264.280 ;
        RECT 827.690 264.000 841.570 264.280 ;
        RECT 842.410 264.000 855.370 264.280 ;
        RECT 856.210 264.000 870.090 264.280 ;
        RECT 870.930 264.000 883.890 264.280 ;
        RECT 884.730 264.000 898.610 264.280 ;
        RECT 899.450 264.000 912.410 264.280 ;
        RECT 913.250 264.000 927.130 264.280 ;
        RECT 927.970 264.000 940.930 264.280 ;
        RECT 941.770 264.000 955.650 264.280 ;
        RECT 956.490 264.000 969.450 264.280 ;
        RECT 970.290 264.000 984.170 264.280 ;
        RECT 985.010 264.000 998.890 264.280 ;
        RECT 999.730 264.000 1012.690 264.280 ;
        RECT 1013.530 264.000 1027.410 264.280 ;
        RECT 1028.250 264.000 1041.210 264.280 ;
        RECT 1042.050 264.000 1055.930 264.280 ;
        RECT 1056.770 264.000 1069.730 264.280 ;
        RECT 1070.570 264.000 1084.450 264.280 ;
        RECT 1085.290 264.000 1098.250 264.280 ;
        RECT 1099.090 264.000 1112.970 264.280 ;
        RECT 1113.810 264.000 1126.770 264.280 ;
        RECT 1127.610 264.000 1141.490 264.280 ;
        RECT 1142.330 264.000 1156.210 264.280 ;
        RECT 1157.050 264.000 1170.010 264.280 ;
        RECT 1170.850 264.000 1184.730 264.280 ;
        RECT 1185.570 264.000 1198.530 264.280 ;
        RECT 1199.370 264.000 1213.250 264.280 ;
        RECT 1214.090 264.000 1227.050 264.280 ;
        RECT 1227.890 264.000 1241.770 264.280 ;
        RECT 1242.610 264.000 1255.570 264.280 ;
        RECT 1256.410 264.000 1270.290 264.280 ;
        RECT 1271.130 264.000 1284.090 264.280 ;
        RECT 1284.930 264.000 1298.810 264.280 ;
        RECT 1299.650 264.000 1313.530 264.280 ;
        RECT 1314.370 264.000 1327.330 264.280 ;
        RECT 1328.170 264.000 1342.050 264.280 ;
        RECT 1342.890 264.000 1355.850 264.280 ;
        RECT 1356.690 264.000 1370.570 264.280 ;
        RECT 1371.410 264.000 1384.370 264.280 ;
        RECT 1385.210 264.000 1399.090 264.280 ;
        RECT 1399.930 264.000 1412.890 264.280 ;
        RECT 1413.730 264.000 1427.610 264.280 ;
        RECT 1428.450 264.000 1441.410 264.280 ;
        RECT 1442.250 264.000 1456.130 264.280 ;
        RECT 1456.970 264.000 1469.930 264.280 ;
        RECT 1470.770 264.000 1484.650 264.280 ;
        RECT 1485.490 264.000 1499.370 264.280 ;
        RECT 1500.210 264.000 1513.170 264.280 ;
        RECT 1514.010 264.000 1527.890 264.280 ;
        RECT 1528.730 264.000 1541.690 264.280 ;
        RECT 1542.530 264.000 1556.410 264.280 ;
        RECT 1557.250 264.000 1570.210 264.280 ;
        RECT 1571.050 264.000 1584.930 264.280 ;
        RECT 1585.770 264.000 1598.730 264.280 ;
        RECT 1599.570 264.000 1613.450 264.280 ;
        RECT 1614.290 264.000 1627.250 264.280 ;
        RECT 1628.090 264.000 1641.970 264.280 ;
        RECT 1642.810 264.000 1656.690 264.280 ;
        RECT 1657.530 264.000 1670.490 264.280 ;
        RECT 1671.330 264.000 1685.210 264.280 ;
        RECT 1686.050 264.000 1699.010 264.280 ;
        RECT 1699.850 264.000 1713.730 264.280 ;
        RECT 1714.570 264.000 1727.530 264.280 ;
        RECT 1728.370 264.000 1742.250 264.280 ;
        RECT 1743.090 264.000 1756.050 264.280 ;
        RECT 1756.890 264.000 1770.770 264.280 ;
        RECT 1771.610 264.000 1784.570 264.280 ;
        RECT 1785.410 264.000 1799.290 264.280 ;
        RECT 1800.130 264.000 1814.010 264.280 ;
        RECT 1814.850 264.000 1827.810 264.280 ;
        RECT 1828.650 264.000 1842.530 264.280 ;
        RECT 1843.370 264.000 1856.330 264.280 ;
        RECT 1857.170 264.000 1871.050 264.280 ;
        RECT 1871.890 264.000 1884.850 264.280 ;
        RECT 1885.690 264.000 1899.570 264.280 ;
        RECT 1900.410 264.000 1913.370 264.280 ;
        RECT 1914.210 264.000 1928.090 264.280 ;
        RECT 1928.930 264.000 1941.890 264.280 ;
        RECT 1942.730 264.000 1956.610 264.280 ;
        RECT 1957.450 264.000 1970.410 264.280 ;
        RECT 1971.250 264.000 1985.130 264.280 ;
        RECT 1985.970 264.000 1999.850 264.280 ;
        RECT 2000.690 264.000 2013.650 264.280 ;
        RECT 2014.490 264.000 2028.370 264.280 ;
        RECT 2029.210 264.000 2042.170 264.280 ;
        RECT 2043.010 264.000 2056.890 264.280 ;
        RECT 2057.730 264.000 2070.690 264.280 ;
        RECT 2071.530 264.000 2085.410 264.280 ;
        RECT 2086.250 264.000 2099.210 264.280 ;
        RECT 2100.050 264.000 2113.930 264.280 ;
        RECT 2114.770 264.000 2127.730 264.280 ;
        RECT 2128.570 264.000 2142.450 264.280 ;
        RECT 2143.290 264.000 2157.170 264.280 ;
        RECT 2158.010 264.000 2170.970 264.280 ;
        RECT 2171.810 264.000 2185.690 264.280 ;
        RECT 2186.530 264.000 2199.490 264.280 ;
        RECT 2200.330 264.000 2214.210 264.280 ;
        RECT 2215.050 264.000 2228.010 264.280 ;
        RECT 2228.850 264.000 2242.730 264.280 ;
        RECT 2243.570 264.000 2256.530 264.280 ;
        RECT 2257.370 264.000 2271.250 264.280 ;
        RECT 2272.090 264.000 2285.050 264.280 ;
        RECT 2285.890 264.000 2299.770 264.280 ;
        RECT 2300.610 264.000 2314.490 264.280 ;
        RECT 2315.330 264.000 2328.290 264.280 ;
        RECT 2329.130 264.000 2343.010 264.280 ;
        RECT 2343.850 264.000 2356.810 264.280 ;
        RECT 2357.650 264.000 2371.530 264.280 ;
        RECT 2372.370 264.000 2385.330 264.280 ;
        RECT 2386.170 264.000 2400.050 264.280 ;
        RECT 2400.890 264.000 2413.850 264.280 ;
        RECT 2414.690 264.000 2428.570 264.280 ;
        RECT 2429.410 264.000 2442.370 264.280 ;
        RECT 2443.210 264.000 2457.090 264.280 ;
        RECT 2457.930 264.000 2471.810 264.280 ;
        RECT 2472.650 264.000 2485.610 264.280 ;
        RECT 2486.450 264.000 2500.330 264.280 ;
        RECT 2501.170 264.000 2514.130 264.280 ;
        RECT 2514.970 264.000 2528.850 264.280 ;
        RECT 2529.690 264.000 2542.650 264.280 ;
        RECT 2543.490 264.000 2557.370 264.280 ;
        RECT 2558.210 264.000 2571.170 264.280 ;
        RECT 2572.010 264.000 2585.890 264.280 ;
        RECT 2586.730 264.000 2599.690 264.280 ;
        RECT 2600.530 264.000 2606.620 264.280 ;
      LAYER met3 ;
        RECT 314.000 3244.880 2606.000 3247.745 ;
        RECT 314.400 3243.480 2606.000 3244.880 ;
        RECT 314.000 3235.360 2606.000 3243.480 ;
        RECT 314.000 3233.960 2605.600 3235.360 ;
        RECT 314.000 3224.480 2606.000 3233.960 ;
        RECT 314.400 3223.080 2606.000 3224.480 ;
        RECT 314.000 3213.600 2606.000 3223.080 ;
        RECT 314.000 3212.200 2605.600 3213.600 ;
        RECT 314.000 3202.720 2606.000 3212.200 ;
        RECT 314.400 3201.320 2606.000 3202.720 ;
        RECT 314.000 3193.200 2606.000 3201.320 ;
        RECT 314.000 3191.800 2605.600 3193.200 ;
        RECT 314.000 3180.960 2606.000 3191.800 ;
        RECT 314.400 3179.560 2606.000 3180.960 ;
        RECT 314.000 3171.440 2606.000 3179.560 ;
        RECT 314.000 3170.040 2605.600 3171.440 ;
        RECT 314.000 3160.560 2606.000 3170.040 ;
        RECT 314.400 3159.160 2606.000 3160.560 ;
        RECT 314.000 3151.040 2606.000 3159.160 ;
        RECT 314.000 3149.640 2605.600 3151.040 ;
        RECT 314.000 3138.800 2606.000 3149.640 ;
        RECT 314.400 3137.400 2606.000 3138.800 ;
        RECT 314.000 3129.280 2606.000 3137.400 ;
        RECT 314.000 3127.880 2605.600 3129.280 ;
        RECT 314.000 3118.400 2606.000 3127.880 ;
        RECT 314.400 3117.000 2606.000 3118.400 ;
        RECT 314.000 3108.880 2606.000 3117.000 ;
        RECT 314.000 3107.480 2605.600 3108.880 ;
        RECT 314.000 3096.640 2606.000 3107.480 ;
        RECT 314.400 3095.240 2606.000 3096.640 ;
        RECT 314.000 3087.120 2606.000 3095.240 ;
        RECT 314.000 3085.720 2605.600 3087.120 ;
        RECT 314.000 3076.240 2606.000 3085.720 ;
        RECT 314.400 3074.840 2606.000 3076.240 ;
        RECT 314.000 3066.720 2606.000 3074.840 ;
        RECT 314.000 3065.320 2605.600 3066.720 ;
        RECT 314.000 3054.480 2606.000 3065.320 ;
        RECT 314.400 3053.080 2606.000 3054.480 ;
        RECT 314.000 3044.960 2606.000 3053.080 ;
        RECT 314.000 3043.560 2605.600 3044.960 ;
        RECT 314.000 3034.080 2606.000 3043.560 ;
        RECT 314.400 3032.680 2606.000 3034.080 ;
        RECT 314.000 3024.560 2606.000 3032.680 ;
        RECT 314.000 3023.160 2605.600 3024.560 ;
        RECT 314.000 3012.320 2606.000 3023.160 ;
        RECT 314.400 3010.920 2606.000 3012.320 ;
        RECT 314.000 3002.800 2606.000 3010.920 ;
        RECT 314.000 3001.400 2605.600 3002.800 ;
        RECT 314.000 2991.920 2606.000 3001.400 ;
        RECT 314.400 2990.520 2606.000 2991.920 ;
        RECT 314.000 2981.040 2606.000 2990.520 ;
        RECT 314.000 2979.640 2605.600 2981.040 ;
        RECT 314.000 2970.160 2606.000 2979.640 ;
        RECT 314.400 2968.760 2606.000 2970.160 ;
        RECT 314.000 2960.640 2606.000 2968.760 ;
        RECT 314.000 2959.240 2605.600 2960.640 ;
        RECT 314.000 2948.400 2606.000 2959.240 ;
        RECT 314.400 2947.000 2606.000 2948.400 ;
        RECT 314.000 2938.880 2606.000 2947.000 ;
        RECT 314.000 2937.480 2605.600 2938.880 ;
        RECT 314.000 2928.000 2606.000 2937.480 ;
        RECT 314.400 2926.600 2606.000 2928.000 ;
        RECT 314.000 2918.480 2606.000 2926.600 ;
        RECT 314.000 2917.080 2605.600 2918.480 ;
        RECT 314.000 2906.240 2606.000 2917.080 ;
        RECT 314.400 2904.840 2606.000 2906.240 ;
        RECT 314.000 2896.720 2606.000 2904.840 ;
        RECT 314.000 2895.320 2605.600 2896.720 ;
        RECT 314.000 2885.840 2606.000 2895.320 ;
        RECT 314.400 2884.440 2606.000 2885.840 ;
        RECT 314.000 2876.320 2606.000 2884.440 ;
        RECT 314.000 2874.920 2605.600 2876.320 ;
        RECT 314.000 2864.080 2606.000 2874.920 ;
        RECT 314.400 2862.680 2606.000 2864.080 ;
        RECT 314.000 2854.560 2606.000 2862.680 ;
        RECT 314.000 2853.160 2605.600 2854.560 ;
        RECT 314.000 2843.680 2606.000 2853.160 ;
        RECT 314.400 2842.280 2606.000 2843.680 ;
        RECT 314.000 2834.160 2606.000 2842.280 ;
        RECT 314.000 2832.760 2605.600 2834.160 ;
        RECT 314.000 2821.920 2606.000 2832.760 ;
        RECT 314.400 2820.520 2606.000 2821.920 ;
        RECT 314.000 2812.400 2606.000 2820.520 ;
        RECT 314.000 2811.000 2605.600 2812.400 ;
        RECT 314.000 2801.520 2606.000 2811.000 ;
        RECT 314.400 2800.120 2606.000 2801.520 ;
        RECT 314.000 2792.000 2606.000 2800.120 ;
        RECT 314.000 2790.600 2605.600 2792.000 ;
        RECT 314.000 2779.760 2606.000 2790.600 ;
        RECT 314.400 2778.360 2606.000 2779.760 ;
        RECT 314.000 2770.240 2606.000 2778.360 ;
        RECT 314.000 2768.840 2605.600 2770.240 ;
        RECT 314.000 2759.360 2606.000 2768.840 ;
        RECT 314.400 2757.960 2606.000 2759.360 ;
        RECT 314.000 2748.480 2606.000 2757.960 ;
        RECT 314.000 2747.080 2605.600 2748.480 ;
        RECT 314.000 2737.600 2606.000 2747.080 ;
        RECT 314.400 2736.200 2606.000 2737.600 ;
        RECT 314.000 2728.080 2606.000 2736.200 ;
        RECT 314.000 2726.680 2605.600 2728.080 ;
        RECT 314.000 2715.840 2606.000 2726.680 ;
        RECT 314.400 2714.440 2606.000 2715.840 ;
        RECT 314.000 2706.320 2606.000 2714.440 ;
        RECT 314.000 2704.920 2605.600 2706.320 ;
        RECT 314.000 2695.440 2606.000 2704.920 ;
        RECT 314.400 2694.040 2606.000 2695.440 ;
        RECT 314.000 2685.920 2606.000 2694.040 ;
        RECT 314.000 2684.520 2605.600 2685.920 ;
        RECT 314.000 2673.680 2606.000 2684.520 ;
        RECT 314.400 2672.280 2606.000 2673.680 ;
        RECT 314.000 2664.160 2606.000 2672.280 ;
        RECT 314.000 2662.760 2605.600 2664.160 ;
        RECT 314.000 2653.280 2606.000 2662.760 ;
        RECT 314.400 2651.880 2606.000 2653.280 ;
        RECT 314.000 2643.760 2606.000 2651.880 ;
        RECT 314.000 2642.360 2605.600 2643.760 ;
        RECT 314.000 2631.520 2606.000 2642.360 ;
        RECT 314.400 2630.120 2606.000 2631.520 ;
        RECT 314.000 2622.000 2606.000 2630.120 ;
        RECT 314.000 2620.600 2605.600 2622.000 ;
        RECT 314.000 2611.120 2606.000 2620.600 ;
        RECT 314.400 2609.720 2606.000 2611.120 ;
        RECT 314.000 2601.600 2606.000 2609.720 ;
        RECT 314.000 2600.200 2605.600 2601.600 ;
        RECT 314.000 2589.360 2606.000 2600.200 ;
        RECT 314.400 2587.960 2606.000 2589.360 ;
        RECT 314.000 2579.840 2606.000 2587.960 ;
        RECT 314.000 2578.440 2605.600 2579.840 ;
        RECT 314.000 2568.960 2606.000 2578.440 ;
        RECT 314.400 2567.560 2606.000 2568.960 ;
        RECT 314.000 2559.440 2606.000 2567.560 ;
        RECT 314.000 2558.040 2605.600 2559.440 ;
        RECT 314.000 2547.200 2606.000 2558.040 ;
        RECT 314.400 2545.800 2606.000 2547.200 ;
        RECT 314.000 2537.680 2606.000 2545.800 ;
        RECT 314.000 2536.280 2605.600 2537.680 ;
        RECT 314.000 2526.800 2606.000 2536.280 ;
        RECT 314.400 2525.400 2606.000 2526.800 ;
        RECT 314.000 2515.920 2606.000 2525.400 ;
        RECT 314.000 2514.520 2605.600 2515.920 ;
        RECT 314.000 2505.040 2606.000 2514.520 ;
        RECT 314.400 2503.640 2606.000 2505.040 ;
        RECT 314.000 2495.520 2606.000 2503.640 ;
        RECT 314.000 2494.120 2605.600 2495.520 ;
        RECT 314.000 2484.640 2606.000 2494.120 ;
        RECT 314.400 2483.240 2606.000 2484.640 ;
        RECT 314.000 2473.760 2606.000 2483.240 ;
        RECT 314.000 2472.360 2605.600 2473.760 ;
        RECT 314.000 2462.880 2606.000 2472.360 ;
        RECT 314.400 2461.480 2606.000 2462.880 ;
        RECT 314.000 2453.360 2606.000 2461.480 ;
        RECT 314.000 2451.960 2605.600 2453.360 ;
        RECT 314.000 2441.120 2606.000 2451.960 ;
        RECT 314.400 2439.720 2606.000 2441.120 ;
        RECT 314.000 2431.600 2606.000 2439.720 ;
        RECT 314.000 2430.200 2605.600 2431.600 ;
        RECT 314.000 2420.720 2606.000 2430.200 ;
        RECT 314.400 2419.320 2606.000 2420.720 ;
        RECT 314.000 2411.200 2606.000 2419.320 ;
        RECT 314.000 2409.800 2605.600 2411.200 ;
        RECT 314.000 2398.960 2606.000 2409.800 ;
        RECT 314.400 2397.560 2606.000 2398.960 ;
        RECT 314.000 2389.440 2606.000 2397.560 ;
        RECT 314.000 2388.040 2605.600 2389.440 ;
        RECT 314.000 2378.560 2606.000 2388.040 ;
        RECT 314.400 2377.160 2606.000 2378.560 ;
        RECT 314.000 2369.040 2606.000 2377.160 ;
        RECT 314.000 2367.640 2605.600 2369.040 ;
        RECT 314.000 2356.800 2606.000 2367.640 ;
        RECT 314.400 2355.400 2606.000 2356.800 ;
        RECT 314.000 2347.280 2606.000 2355.400 ;
        RECT 314.000 2345.880 2605.600 2347.280 ;
        RECT 314.000 2336.400 2606.000 2345.880 ;
        RECT 314.400 2335.000 2606.000 2336.400 ;
        RECT 314.000 2326.880 2606.000 2335.000 ;
        RECT 314.000 2325.480 2605.600 2326.880 ;
        RECT 314.000 2314.640 2606.000 2325.480 ;
        RECT 314.400 2313.240 2606.000 2314.640 ;
        RECT 314.000 2305.120 2606.000 2313.240 ;
        RECT 314.000 2303.720 2605.600 2305.120 ;
        RECT 314.000 2294.240 2606.000 2303.720 ;
        RECT 314.400 2292.840 2606.000 2294.240 ;
        RECT 314.000 2284.720 2606.000 2292.840 ;
        RECT 314.000 2283.320 2605.600 2284.720 ;
        RECT 314.000 2272.480 2606.000 2283.320 ;
        RECT 314.400 2271.080 2606.000 2272.480 ;
        RECT 314.000 2262.960 2606.000 2271.080 ;
        RECT 314.000 2261.560 2605.600 2262.960 ;
        RECT 314.000 2252.080 2606.000 2261.560 ;
        RECT 314.400 2250.680 2606.000 2252.080 ;
        RECT 314.000 2241.200 2606.000 2250.680 ;
        RECT 314.000 2239.800 2605.600 2241.200 ;
        RECT 314.000 2230.320 2606.000 2239.800 ;
        RECT 314.400 2228.920 2606.000 2230.320 ;
        RECT 314.000 2220.800 2606.000 2228.920 ;
        RECT 314.000 2219.400 2605.600 2220.800 ;
        RECT 314.000 2208.560 2606.000 2219.400 ;
        RECT 314.400 2207.160 2606.000 2208.560 ;
        RECT 314.000 2199.040 2606.000 2207.160 ;
        RECT 314.000 2197.640 2605.600 2199.040 ;
        RECT 314.000 2188.160 2606.000 2197.640 ;
        RECT 314.400 2186.760 2606.000 2188.160 ;
        RECT 314.000 2178.640 2606.000 2186.760 ;
        RECT 314.000 2177.240 2605.600 2178.640 ;
        RECT 314.000 2166.400 2606.000 2177.240 ;
        RECT 314.400 2165.000 2606.000 2166.400 ;
        RECT 314.000 2156.880 2606.000 2165.000 ;
        RECT 314.000 2155.480 2605.600 2156.880 ;
        RECT 314.000 2146.000 2606.000 2155.480 ;
        RECT 314.400 2144.600 2606.000 2146.000 ;
        RECT 314.000 2136.480 2606.000 2144.600 ;
        RECT 314.000 2135.080 2605.600 2136.480 ;
        RECT 314.000 2124.240 2606.000 2135.080 ;
        RECT 314.400 2122.840 2606.000 2124.240 ;
        RECT 314.000 2114.720 2606.000 2122.840 ;
        RECT 314.000 2113.320 2605.600 2114.720 ;
        RECT 314.000 2103.840 2606.000 2113.320 ;
        RECT 314.400 2102.440 2606.000 2103.840 ;
        RECT 314.000 2094.320 2606.000 2102.440 ;
        RECT 314.000 2092.920 2605.600 2094.320 ;
        RECT 314.000 2082.080 2606.000 2092.920 ;
        RECT 314.400 2080.680 2606.000 2082.080 ;
        RECT 314.000 2072.560 2606.000 2080.680 ;
        RECT 314.000 2071.160 2605.600 2072.560 ;
        RECT 314.000 2061.680 2606.000 2071.160 ;
        RECT 314.400 2060.280 2606.000 2061.680 ;
        RECT 314.000 2052.160 2606.000 2060.280 ;
        RECT 314.000 2050.760 2605.600 2052.160 ;
        RECT 314.000 2039.920 2606.000 2050.760 ;
        RECT 314.400 2038.520 2606.000 2039.920 ;
        RECT 314.000 2030.400 2606.000 2038.520 ;
        RECT 314.000 2029.000 2605.600 2030.400 ;
        RECT 314.000 2019.520 2606.000 2029.000 ;
        RECT 314.400 2018.120 2606.000 2019.520 ;
        RECT 314.000 2008.640 2606.000 2018.120 ;
        RECT 314.000 2007.240 2605.600 2008.640 ;
        RECT 314.000 1997.760 2606.000 2007.240 ;
        RECT 314.400 1996.360 2606.000 1997.760 ;
        RECT 314.000 1988.240 2606.000 1996.360 ;
        RECT 314.000 1986.840 2605.600 1988.240 ;
        RECT 314.000 1976.000 2606.000 1986.840 ;
        RECT 314.400 1974.600 2606.000 1976.000 ;
        RECT 314.000 1966.480 2606.000 1974.600 ;
        RECT 314.000 1965.080 2605.600 1966.480 ;
        RECT 314.000 1955.600 2606.000 1965.080 ;
        RECT 314.400 1954.200 2606.000 1955.600 ;
        RECT 314.000 1946.080 2606.000 1954.200 ;
        RECT 314.000 1944.680 2605.600 1946.080 ;
        RECT 314.000 1933.840 2606.000 1944.680 ;
        RECT 314.400 1932.440 2606.000 1933.840 ;
        RECT 314.000 1924.320 2606.000 1932.440 ;
        RECT 314.000 1922.920 2605.600 1924.320 ;
        RECT 314.000 1913.440 2606.000 1922.920 ;
        RECT 314.400 1912.040 2606.000 1913.440 ;
        RECT 314.000 1903.920 2606.000 1912.040 ;
        RECT 314.000 1902.520 2605.600 1903.920 ;
        RECT 314.000 1891.680 2606.000 1902.520 ;
        RECT 314.400 1890.280 2606.000 1891.680 ;
        RECT 314.000 1882.160 2606.000 1890.280 ;
        RECT 314.000 1880.760 2605.600 1882.160 ;
        RECT 314.000 1871.280 2606.000 1880.760 ;
        RECT 314.400 1869.880 2606.000 1871.280 ;
        RECT 314.000 1861.760 2606.000 1869.880 ;
        RECT 314.000 1860.360 2605.600 1861.760 ;
        RECT 314.000 1849.520 2606.000 1860.360 ;
        RECT 314.400 1848.120 2606.000 1849.520 ;
        RECT 314.000 1840.000 2606.000 1848.120 ;
        RECT 314.000 1838.600 2605.600 1840.000 ;
        RECT 314.000 1829.120 2606.000 1838.600 ;
        RECT 314.400 1827.720 2606.000 1829.120 ;
        RECT 314.000 1819.600 2606.000 1827.720 ;
        RECT 314.000 1818.200 2605.600 1819.600 ;
        RECT 314.000 1807.360 2606.000 1818.200 ;
        RECT 314.400 1805.960 2606.000 1807.360 ;
        RECT 314.000 1797.840 2606.000 1805.960 ;
        RECT 314.000 1796.440 2605.600 1797.840 ;
        RECT 314.000 1786.960 2606.000 1796.440 ;
        RECT 314.400 1785.560 2606.000 1786.960 ;
        RECT 314.000 1776.080 2606.000 1785.560 ;
        RECT 314.000 1774.680 2605.600 1776.080 ;
        RECT 314.000 1765.200 2606.000 1774.680 ;
        RECT 314.400 1763.800 2606.000 1765.200 ;
        RECT 314.000 1755.680 2606.000 1763.800 ;
        RECT 314.000 1754.280 2605.600 1755.680 ;
        RECT 314.000 1744.800 2606.000 1754.280 ;
        RECT 314.400 1743.400 2606.000 1744.800 ;
        RECT 314.000 1733.920 2606.000 1743.400 ;
        RECT 314.000 1732.520 2605.600 1733.920 ;
        RECT 314.000 1723.040 2606.000 1732.520 ;
        RECT 314.400 1721.640 2606.000 1723.040 ;
        RECT 314.000 1713.520 2606.000 1721.640 ;
        RECT 314.000 1712.120 2605.600 1713.520 ;
        RECT 314.000 1701.280 2606.000 1712.120 ;
        RECT 314.400 1699.880 2606.000 1701.280 ;
        RECT 314.000 1691.760 2606.000 1699.880 ;
        RECT 314.000 1690.360 2605.600 1691.760 ;
        RECT 314.000 1680.880 2606.000 1690.360 ;
        RECT 314.400 1679.480 2606.000 1680.880 ;
        RECT 314.000 1671.360 2606.000 1679.480 ;
        RECT 314.000 1669.960 2605.600 1671.360 ;
        RECT 314.000 1659.120 2606.000 1669.960 ;
        RECT 314.400 1657.720 2606.000 1659.120 ;
        RECT 314.000 1649.600 2606.000 1657.720 ;
        RECT 314.000 1648.200 2605.600 1649.600 ;
        RECT 314.000 1638.720 2606.000 1648.200 ;
        RECT 314.400 1637.320 2606.000 1638.720 ;
        RECT 314.000 1629.200 2606.000 1637.320 ;
        RECT 314.000 1627.800 2605.600 1629.200 ;
        RECT 314.000 1616.960 2606.000 1627.800 ;
        RECT 314.400 1615.560 2606.000 1616.960 ;
        RECT 314.000 1607.440 2606.000 1615.560 ;
        RECT 314.000 1606.040 2605.600 1607.440 ;
        RECT 314.000 1596.560 2606.000 1606.040 ;
        RECT 314.400 1595.160 2606.000 1596.560 ;
        RECT 314.000 1587.040 2606.000 1595.160 ;
        RECT 314.000 1585.640 2605.600 1587.040 ;
        RECT 314.000 1574.800 2606.000 1585.640 ;
        RECT 314.400 1573.400 2606.000 1574.800 ;
        RECT 314.000 1565.280 2606.000 1573.400 ;
        RECT 314.000 1563.880 2605.600 1565.280 ;
        RECT 314.000 1554.400 2606.000 1563.880 ;
        RECT 314.400 1553.000 2606.000 1554.400 ;
        RECT 314.000 1544.880 2606.000 1553.000 ;
        RECT 314.000 1543.480 2605.600 1544.880 ;
        RECT 314.000 1532.640 2606.000 1543.480 ;
        RECT 314.400 1531.240 2606.000 1532.640 ;
        RECT 314.000 1523.120 2606.000 1531.240 ;
        RECT 314.000 1521.720 2605.600 1523.120 ;
        RECT 314.000 1512.240 2606.000 1521.720 ;
        RECT 314.400 1510.840 2606.000 1512.240 ;
        RECT 314.000 1501.360 2606.000 1510.840 ;
        RECT 314.000 1499.960 2605.600 1501.360 ;
        RECT 314.000 1490.480 2606.000 1499.960 ;
        RECT 314.400 1489.080 2606.000 1490.480 ;
        RECT 314.000 1480.960 2606.000 1489.080 ;
        RECT 314.000 1479.560 2605.600 1480.960 ;
        RECT 314.000 1468.720 2606.000 1479.560 ;
        RECT 314.400 1467.320 2606.000 1468.720 ;
        RECT 314.000 1459.200 2606.000 1467.320 ;
        RECT 314.000 1457.800 2605.600 1459.200 ;
        RECT 314.000 1448.320 2606.000 1457.800 ;
        RECT 314.400 1446.920 2606.000 1448.320 ;
        RECT 314.000 1438.800 2606.000 1446.920 ;
        RECT 314.000 1437.400 2605.600 1438.800 ;
        RECT 314.000 1426.560 2606.000 1437.400 ;
        RECT 314.400 1425.160 2606.000 1426.560 ;
        RECT 314.000 1417.040 2606.000 1425.160 ;
        RECT 314.000 1415.640 2605.600 1417.040 ;
        RECT 314.000 1406.160 2606.000 1415.640 ;
        RECT 314.400 1404.760 2606.000 1406.160 ;
        RECT 314.000 1396.640 2606.000 1404.760 ;
        RECT 314.000 1395.240 2605.600 1396.640 ;
        RECT 314.000 1384.400 2606.000 1395.240 ;
        RECT 314.400 1383.000 2606.000 1384.400 ;
        RECT 314.000 1374.880 2606.000 1383.000 ;
        RECT 314.000 1373.480 2605.600 1374.880 ;
        RECT 314.000 1364.000 2606.000 1373.480 ;
        RECT 314.400 1362.600 2606.000 1364.000 ;
        RECT 314.000 1354.480 2606.000 1362.600 ;
        RECT 314.000 1353.080 2605.600 1354.480 ;
        RECT 314.000 1342.240 2606.000 1353.080 ;
        RECT 314.400 1340.840 2606.000 1342.240 ;
        RECT 314.000 1332.720 2606.000 1340.840 ;
        RECT 314.000 1331.320 2605.600 1332.720 ;
        RECT 314.000 1321.840 2606.000 1331.320 ;
        RECT 314.400 1320.440 2606.000 1321.840 ;
        RECT 314.000 1312.320 2606.000 1320.440 ;
        RECT 314.000 1310.920 2605.600 1312.320 ;
        RECT 314.000 1300.080 2606.000 1310.920 ;
        RECT 314.400 1298.680 2606.000 1300.080 ;
        RECT 314.000 1290.560 2606.000 1298.680 ;
        RECT 314.000 1289.160 2605.600 1290.560 ;
        RECT 314.000 1279.680 2606.000 1289.160 ;
        RECT 314.400 1278.280 2606.000 1279.680 ;
        RECT 314.000 1268.800 2606.000 1278.280 ;
        RECT 314.000 1267.400 2605.600 1268.800 ;
        RECT 314.000 1257.920 2606.000 1267.400 ;
        RECT 314.400 1256.520 2606.000 1257.920 ;
        RECT 314.000 1248.400 2606.000 1256.520 ;
        RECT 314.000 1247.000 2605.600 1248.400 ;
        RECT 314.000 1236.160 2606.000 1247.000 ;
        RECT 314.400 1234.760 2606.000 1236.160 ;
        RECT 314.000 1226.640 2606.000 1234.760 ;
        RECT 314.000 1225.240 2605.600 1226.640 ;
        RECT 314.000 1215.760 2606.000 1225.240 ;
        RECT 314.400 1214.360 2606.000 1215.760 ;
        RECT 314.000 1206.240 2606.000 1214.360 ;
        RECT 314.000 1204.840 2605.600 1206.240 ;
        RECT 314.000 1194.000 2606.000 1204.840 ;
        RECT 314.400 1192.600 2606.000 1194.000 ;
        RECT 314.000 1184.480 2606.000 1192.600 ;
        RECT 314.000 1183.080 2605.600 1184.480 ;
        RECT 314.000 1173.600 2606.000 1183.080 ;
        RECT 314.400 1172.200 2606.000 1173.600 ;
        RECT 314.000 1164.080 2606.000 1172.200 ;
        RECT 314.000 1162.680 2605.600 1164.080 ;
        RECT 314.000 1151.840 2606.000 1162.680 ;
        RECT 314.400 1150.440 2606.000 1151.840 ;
        RECT 314.000 1142.320 2606.000 1150.440 ;
        RECT 314.000 1140.920 2605.600 1142.320 ;
        RECT 314.000 1131.440 2606.000 1140.920 ;
        RECT 314.400 1130.040 2606.000 1131.440 ;
        RECT 314.000 1121.920 2606.000 1130.040 ;
        RECT 314.000 1120.520 2605.600 1121.920 ;
        RECT 314.000 1109.680 2606.000 1120.520 ;
        RECT 314.400 1108.280 2606.000 1109.680 ;
        RECT 314.000 1100.160 2606.000 1108.280 ;
        RECT 314.000 1098.760 2605.600 1100.160 ;
        RECT 314.000 1089.280 2606.000 1098.760 ;
        RECT 314.400 1087.880 2606.000 1089.280 ;
        RECT 314.000 1079.760 2606.000 1087.880 ;
        RECT 314.000 1078.360 2605.600 1079.760 ;
        RECT 314.000 1067.520 2606.000 1078.360 ;
        RECT 314.400 1066.120 2606.000 1067.520 ;
        RECT 314.000 1058.000 2606.000 1066.120 ;
        RECT 314.000 1056.600 2605.600 1058.000 ;
        RECT 314.000 1047.120 2606.000 1056.600 ;
        RECT 314.400 1045.720 2606.000 1047.120 ;
        RECT 314.000 1036.240 2606.000 1045.720 ;
        RECT 314.000 1034.840 2605.600 1036.240 ;
        RECT 314.000 1025.360 2606.000 1034.840 ;
        RECT 314.400 1023.960 2606.000 1025.360 ;
        RECT 314.000 1015.840 2606.000 1023.960 ;
        RECT 314.000 1014.440 2605.600 1015.840 ;
        RECT 314.000 1004.960 2606.000 1014.440 ;
        RECT 314.400 1003.560 2606.000 1004.960 ;
        RECT 314.000 994.080 2606.000 1003.560 ;
        RECT 314.000 992.680 2605.600 994.080 ;
        RECT 314.000 983.200 2606.000 992.680 ;
        RECT 314.400 981.800 2606.000 983.200 ;
        RECT 314.000 973.680 2606.000 981.800 ;
        RECT 314.000 972.280 2605.600 973.680 ;
        RECT 314.000 961.440 2606.000 972.280 ;
        RECT 314.400 960.040 2606.000 961.440 ;
        RECT 314.000 951.920 2606.000 960.040 ;
        RECT 314.000 950.520 2605.600 951.920 ;
        RECT 314.000 941.040 2606.000 950.520 ;
        RECT 314.400 939.640 2606.000 941.040 ;
        RECT 314.000 931.520 2606.000 939.640 ;
        RECT 314.000 930.120 2605.600 931.520 ;
        RECT 314.000 919.280 2606.000 930.120 ;
        RECT 314.400 917.880 2606.000 919.280 ;
        RECT 314.000 909.760 2606.000 917.880 ;
        RECT 314.000 908.360 2605.600 909.760 ;
        RECT 314.000 898.880 2606.000 908.360 ;
        RECT 314.400 897.480 2606.000 898.880 ;
        RECT 314.000 889.360 2606.000 897.480 ;
        RECT 314.000 887.960 2605.600 889.360 ;
        RECT 314.000 877.120 2606.000 887.960 ;
        RECT 314.400 875.720 2606.000 877.120 ;
        RECT 314.000 867.600 2606.000 875.720 ;
        RECT 314.000 866.200 2605.600 867.600 ;
        RECT 314.000 856.720 2606.000 866.200 ;
        RECT 314.400 855.320 2606.000 856.720 ;
        RECT 314.000 847.200 2606.000 855.320 ;
        RECT 314.000 845.800 2605.600 847.200 ;
        RECT 314.000 834.960 2606.000 845.800 ;
        RECT 314.400 833.560 2606.000 834.960 ;
        RECT 314.000 825.440 2606.000 833.560 ;
        RECT 314.000 824.040 2605.600 825.440 ;
        RECT 314.000 814.560 2606.000 824.040 ;
        RECT 314.400 813.160 2606.000 814.560 ;
        RECT 314.000 805.040 2606.000 813.160 ;
        RECT 314.000 803.640 2605.600 805.040 ;
        RECT 314.000 792.800 2606.000 803.640 ;
        RECT 314.400 791.400 2606.000 792.800 ;
        RECT 314.000 783.280 2606.000 791.400 ;
        RECT 314.000 781.880 2605.600 783.280 ;
        RECT 314.000 772.400 2606.000 781.880 ;
        RECT 314.400 771.000 2606.000 772.400 ;
        RECT 314.000 761.520 2606.000 771.000 ;
        RECT 314.000 760.120 2605.600 761.520 ;
        RECT 314.000 750.640 2606.000 760.120 ;
        RECT 314.400 749.240 2606.000 750.640 ;
        RECT 314.000 741.120 2606.000 749.240 ;
        RECT 314.000 739.720 2605.600 741.120 ;
        RECT 314.000 728.880 2606.000 739.720 ;
        RECT 314.400 727.480 2606.000 728.880 ;
        RECT 314.000 719.360 2606.000 727.480 ;
        RECT 314.000 717.960 2605.600 719.360 ;
        RECT 314.000 708.480 2606.000 717.960 ;
        RECT 314.400 707.080 2606.000 708.480 ;
        RECT 314.000 698.960 2606.000 707.080 ;
        RECT 314.000 697.560 2605.600 698.960 ;
        RECT 314.000 686.720 2606.000 697.560 ;
        RECT 314.400 685.320 2606.000 686.720 ;
        RECT 314.000 677.200 2606.000 685.320 ;
        RECT 314.000 675.800 2605.600 677.200 ;
        RECT 314.000 666.320 2606.000 675.800 ;
        RECT 314.400 664.920 2606.000 666.320 ;
        RECT 314.000 656.800 2606.000 664.920 ;
        RECT 314.000 655.400 2605.600 656.800 ;
        RECT 314.000 644.560 2606.000 655.400 ;
        RECT 314.400 643.160 2606.000 644.560 ;
        RECT 314.000 635.040 2606.000 643.160 ;
        RECT 314.000 633.640 2605.600 635.040 ;
        RECT 314.000 624.160 2606.000 633.640 ;
        RECT 314.400 622.760 2606.000 624.160 ;
        RECT 314.000 614.640 2606.000 622.760 ;
        RECT 314.000 613.240 2605.600 614.640 ;
        RECT 314.000 602.400 2606.000 613.240 ;
        RECT 314.400 601.000 2606.000 602.400 ;
        RECT 314.000 592.880 2606.000 601.000 ;
        RECT 314.000 591.480 2605.600 592.880 ;
        RECT 314.000 582.000 2606.000 591.480 ;
        RECT 314.400 580.600 2606.000 582.000 ;
        RECT 314.000 572.480 2606.000 580.600 ;
        RECT 314.000 571.080 2605.600 572.480 ;
        RECT 314.000 560.240 2606.000 571.080 ;
        RECT 314.400 558.840 2606.000 560.240 ;
        RECT 314.000 550.720 2606.000 558.840 ;
        RECT 314.000 549.320 2605.600 550.720 ;
        RECT 314.000 539.840 2606.000 549.320 ;
        RECT 314.400 538.440 2606.000 539.840 ;
        RECT 314.000 528.960 2606.000 538.440 ;
        RECT 314.000 527.560 2605.600 528.960 ;
        RECT 314.000 518.080 2606.000 527.560 ;
        RECT 314.400 516.680 2606.000 518.080 ;
        RECT 314.000 508.560 2606.000 516.680 ;
        RECT 314.000 507.160 2605.600 508.560 ;
        RECT 314.000 496.320 2606.000 507.160 ;
        RECT 314.400 494.920 2606.000 496.320 ;
        RECT 314.000 486.800 2606.000 494.920 ;
        RECT 314.000 485.400 2605.600 486.800 ;
        RECT 314.000 475.920 2606.000 485.400 ;
        RECT 314.400 474.520 2606.000 475.920 ;
        RECT 314.000 466.400 2606.000 474.520 ;
        RECT 314.000 465.000 2605.600 466.400 ;
        RECT 314.000 454.160 2606.000 465.000 ;
        RECT 314.400 452.760 2606.000 454.160 ;
        RECT 314.000 444.640 2606.000 452.760 ;
        RECT 314.000 443.240 2605.600 444.640 ;
        RECT 314.000 433.760 2606.000 443.240 ;
        RECT 314.400 432.360 2606.000 433.760 ;
        RECT 314.000 424.240 2606.000 432.360 ;
        RECT 314.000 422.840 2605.600 424.240 ;
        RECT 314.000 412.000 2606.000 422.840 ;
        RECT 314.400 410.600 2606.000 412.000 ;
        RECT 314.000 402.480 2606.000 410.600 ;
        RECT 314.000 401.080 2605.600 402.480 ;
        RECT 314.000 391.600 2606.000 401.080 ;
        RECT 314.400 390.200 2606.000 391.600 ;
        RECT 314.000 382.080 2606.000 390.200 ;
        RECT 314.000 380.680 2605.600 382.080 ;
        RECT 314.000 369.840 2606.000 380.680 ;
        RECT 314.400 368.440 2606.000 369.840 ;
        RECT 314.000 360.320 2606.000 368.440 ;
        RECT 314.000 358.920 2605.600 360.320 ;
        RECT 314.000 349.440 2606.000 358.920 ;
        RECT 314.400 348.040 2606.000 349.440 ;
        RECT 314.000 339.920 2606.000 348.040 ;
        RECT 314.000 338.520 2605.600 339.920 ;
        RECT 314.000 327.680 2606.000 338.520 ;
        RECT 314.400 326.280 2606.000 327.680 ;
        RECT 314.000 318.160 2606.000 326.280 ;
        RECT 314.000 316.760 2605.600 318.160 ;
        RECT 314.000 307.280 2606.000 316.760 ;
        RECT 314.400 305.880 2606.000 307.280 ;
        RECT 314.000 296.400 2606.000 305.880 ;
        RECT 314.000 295.000 2605.600 296.400 ;
        RECT 314.000 285.520 2606.000 295.000 ;
        RECT 314.400 284.120 2606.000 285.520 ;
        RECT 314.000 276.000 2606.000 284.120 ;
        RECT 314.000 274.600 2605.600 276.000 ;
        RECT 314.000 264.255 2606.000 274.600 ;
      LAYER met4 ;
        RECT 317.655 270.640 330.640 3246.800 ;
      LAYER met4 ;
        RECT 331.040 270.640 332.640 3246.800 ;
      LAYER met4 ;
        RECT 333.040 2970.490 407.440 3246.800 ;
        RECT 333.040 2969.310 407.430 2970.490 ;
        RECT 333.040 2797.090 407.440 2969.310 ;
        RECT 333.040 2795.910 407.430 2797.090 ;
        RECT 333.040 2599.890 407.440 2795.910 ;
        RECT 333.040 2598.710 407.430 2599.890 ;
        RECT 333.040 2236.090 407.440 2598.710 ;
        RECT 333.040 2234.910 407.430 2236.090 ;
        RECT 333.040 2168.090 407.440 2234.910 ;
        RECT 333.040 2166.910 407.430 2168.090 ;
        RECT 333.040 2072.890 407.440 2166.910 ;
        RECT 333.040 2071.710 407.430 2072.890 ;
        RECT 333.040 2059.290 407.440 2071.710 ;
        RECT 333.040 2058.110 407.430 2059.290 ;
        RECT 333.040 1797.490 407.440 2058.110 ;
        RECT 333.040 1796.310 407.430 1797.490 ;
        RECT 333.040 1787.290 407.440 1796.310 ;
        RECT 333.040 1786.110 407.430 1787.290 ;
        RECT 333.040 1250.090 407.440 1786.110 ;
        RECT 333.040 1248.910 407.430 1250.090 ;
        RECT 333.040 971.290 407.440 1248.910 ;
        RECT 333.040 970.110 407.430 971.290 ;
        RECT 333.040 631.290 407.440 970.110 ;
        RECT 333.040 630.110 407.430 631.290 ;
        RECT 333.040 621.090 407.440 630.110 ;
        RECT 333.040 619.910 407.430 621.090 ;
        RECT 333.040 529.290 407.440 619.910 ;
        RECT 333.040 528.110 407.430 529.290 ;
        RECT 333.040 270.640 407.440 528.110 ;
        RECT 409.840 270.640 2590.385 3246.800 ;
  END
END user_project_wrapper
END LIBRARY

