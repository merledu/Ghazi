VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 89.660 2619.170 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2618.850 89.520 2899.310 89.660 ;
        RECT 2618.850 89.460 2619.170 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2618.880 89.460 2619.140 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2618.870 249.715 2619.150 250.085 ;
        RECT 2618.940 89.750 2619.080 249.715 ;
        RECT 2618.880 89.430 2619.140 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2618.870 249.760 2619.150 250.040 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2618.845 250.050 2619.175 250.065 ;
        RECT 2609.580 249.960 2619.175 250.050 ;
        RECT 2606.000 249.750 2619.175 249.960 ;
        RECT 2606.000 249.360 2610.000 249.750 ;
        RECT 2618.845 249.735 2619.175 249.750 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2429.200 2619.170 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2618.850 2429.060 2901.150 2429.200 ;
        RECT 2618.850 2429.000 2619.170 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
      LAYER via ;
        RECT 2618.880 2429.000 2619.140 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2618.880 2428.970 2619.140 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2618.940 2249.965 2619.080 2428.970 ;
        RECT 2618.870 2249.595 2619.150 2249.965 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2618.870 2249.640 2619.150 2249.920 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2618.845 2249.930 2619.175 2249.945 ;
        RECT 2609.580 2249.840 2619.175 2249.930 ;
        RECT 2606.000 2249.630 2619.175 2249.840 ;
        RECT 2606.000 2249.240 2610.000 2249.630 ;
        RECT 2618.845 2249.615 2619.175 2249.630 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 2456.400 2621.930 2456.460 ;
        RECT 2901.750 2456.400 2902.070 2456.460 ;
        RECT 2621.610 2456.260 2902.070 2456.400 ;
        RECT 2621.610 2456.200 2621.930 2456.260 ;
        RECT 2901.750 2456.200 2902.070 2456.260 ;
      LAYER via ;
        RECT 2621.640 2456.200 2621.900 2456.460 ;
        RECT 2901.780 2456.200 2902.040 2456.460 ;
      LAYER met2 ;
        RECT 2901.770 2669.155 2902.050 2669.525 ;
        RECT 2901.840 2456.490 2901.980 2669.155 ;
        RECT 2621.640 2456.170 2621.900 2456.490 ;
        RECT 2901.780 2456.170 2902.040 2456.490 ;
        RECT 2621.700 2449.885 2621.840 2456.170 ;
        RECT 2621.630 2449.515 2621.910 2449.885 ;
      LAYER via2 ;
        RECT 2901.770 2669.200 2902.050 2669.480 ;
        RECT 2621.630 2449.560 2621.910 2449.840 ;
      LAYER met3 ;
        RECT 2901.745 2669.490 2902.075 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2901.745 2669.190 2924.800 2669.490 ;
        RECT 2901.745 2669.175 2902.075 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2621.605 2449.850 2621.935 2449.865 ;
        RECT 2609.580 2449.760 2621.935 2449.850 ;
        RECT 2606.000 2449.550 2621.935 2449.760 ;
        RECT 2606.000 2449.160 2610.000 2449.550 ;
        RECT 2621.605 2449.535 2621.935 2449.550 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2616.090 2656.320 2616.410 2656.380 ;
        RECT 2901.290 2656.320 2901.610 2656.380 ;
        RECT 2616.090 2656.180 2901.610 2656.320 ;
        RECT 2616.090 2656.120 2616.410 2656.180 ;
        RECT 2901.290 2656.120 2901.610 2656.180 ;
      LAYER via ;
        RECT 2616.120 2656.120 2616.380 2656.380 ;
        RECT 2901.320 2656.120 2901.580 2656.380 ;
      LAYER met2 ;
        RECT 2901.310 2903.755 2901.590 2904.125 ;
        RECT 2901.380 2656.410 2901.520 2903.755 ;
        RECT 2616.120 2656.090 2616.380 2656.410 ;
        RECT 2901.320 2656.090 2901.580 2656.410 ;
        RECT 2616.180 2649.805 2616.320 2656.090 ;
        RECT 2616.110 2649.435 2616.390 2649.805 ;
      LAYER via2 ;
        RECT 2901.310 2903.800 2901.590 2904.080 ;
        RECT 2616.110 2649.480 2616.390 2649.760 ;
      LAYER met3 ;
        RECT 2901.285 2904.090 2901.615 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2901.285 2903.790 2924.800 2904.090 ;
        RECT 2901.285 2903.775 2901.615 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2616.085 2649.770 2616.415 2649.785 ;
        RECT 2609.580 2649.680 2616.415 2649.770 ;
        RECT 2606.000 2649.470 2616.415 2649.680 ;
        RECT 2606.000 2649.080 2610.000 2649.470 ;
        RECT 2616.085 2649.455 2616.415 2649.470 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 2849.440 2621.930 2849.500 ;
        RECT 2901.750 2849.440 2902.070 2849.500 ;
        RECT 2621.610 2849.300 2902.070 2849.440 ;
        RECT 2621.610 2849.240 2621.930 2849.300 ;
        RECT 2901.750 2849.240 2902.070 2849.300 ;
      LAYER via ;
        RECT 2621.640 2849.240 2621.900 2849.500 ;
        RECT 2901.780 2849.240 2902.040 2849.500 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 2621.630 2849.355 2621.910 2849.725 ;
        RECT 2901.840 2849.530 2901.980 3138.355 ;
        RECT 2621.640 2849.210 2621.900 2849.355 ;
        RECT 2901.780 2849.210 2902.040 2849.530 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
        RECT 2621.630 2849.400 2621.910 2849.680 ;
      LAYER met3 ;
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2621.605 2849.690 2621.935 2849.705 ;
        RECT 2609.580 2849.600 2621.935 2849.690 ;
        RECT 2606.000 2849.390 2621.935 2849.600 ;
        RECT 2606.000 2849.000 2610.000 2849.390 ;
        RECT 2621.605 2849.375 2621.935 2849.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 3049.700 2621.930 3049.760 ;
        RECT 2901.290 3049.700 2901.610 3049.760 ;
        RECT 2621.610 3049.560 2901.610 3049.700 ;
        RECT 2621.610 3049.500 2621.930 3049.560 ;
        RECT 2901.290 3049.500 2901.610 3049.560 ;
      LAYER via ;
        RECT 2621.640 3049.500 2621.900 3049.760 ;
        RECT 2901.320 3049.500 2901.580 3049.760 ;
      LAYER met2 ;
        RECT 2901.310 3372.955 2901.590 3373.325 ;
        RECT 2901.380 3049.790 2901.520 3372.955 ;
        RECT 2621.640 3049.645 2621.900 3049.790 ;
        RECT 2621.630 3049.275 2621.910 3049.645 ;
        RECT 2901.320 3049.470 2901.580 3049.790 ;
      LAYER via2 ;
        RECT 2901.310 3373.000 2901.590 3373.280 ;
        RECT 2621.630 3049.320 2621.910 3049.600 ;
      LAYER met3 ;
        RECT 2901.285 3373.290 2901.615 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2901.285 3372.990 2924.800 3373.290 ;
        RECT 2901.285 3372.975 2901.615 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2621.605 3049.610 2621.935 3049.625 ;
        RECT 2609.580 3049.520 2621.935 3049.610 ;
        RECT 2606.000 3049.310 2621.935 3049.520 ;
        RECT 2606.000 3048.920 2610.000 3049.310 ;
        RECT 2621.605 3049.295 2621.935 3049.310 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 3502.240 2573.630 3502.300 ;
        RECT 2798.250 3502.240 2798.570 3502.300 ;
        RECT 2573.310 3502.100 2798.570 3502.240 ;
        RECT 2573.310 3502.040 2573.630 3502.100 ;
        RECT 2798.250 3502.040 2798.570 3502.100 ;
        RECT 2566.870 3228.200 2567.190 3228.260 ;
        RECT 2573.310 3228.200 2573.630 3228.260 ;
        RECT 2566.870 3228.060 2573.630 3228.200 ;
        RECT 2566.870 3228.000 2567.190 3228.060 ;
        RECT 2573.310 3228.000 2573.630 3228.060 ;
      LAYER via ;
        RECT 2573.340 3502.040 2573.600 3502.300 ;
        RECT 2798.280 3502.040 2798.540 3502.300 ;
        RECT 2566.900 3228.000 2567.160 3228.260 ;
        RECT 2573.340 3228.000 2573.600 3228.260 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3502.330 2798.480 3517.600 ;
        RECT 2573.340 3502.010 2573.600 3502.330 ;
        RECT 2798.280 3502.010 2798.540 3502.330 ;
        RECT 2573.400 3228.290 2573.540 3502.010 ;
        RECT 2566.900 3227.970 2567.160 3228.290 ;
        RECT 2573.340 3227.970 2573.600 3228.290 ;
        RECT 2566.960 3216.000 2567.100 3227.970 ;
        RECT 2566.850 3212.000 2567.130 3216.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2318.010 3502.240 2318.330 3502.300 ;
        RECT 2473.950 3502.240 2474.270 3502.300 ;
        RECT 2318.010 3502.100 2474.270 3502.240 ;
        RECT 2318.010 3502.040 2318.330 3502.100 ;
        RECT 2473.950 3502.040 2474.270 3502.100 ;
        RECT 2311.570 3229.220 2311.890 3229.280 ;
        RECT 2318.010 3229.220 2318.330 3229.280 ;
        RECT 2311.570 3229.080 2318.330 3229.220 ;
        RECT 2311.570 3229.020 2311.890 3229.080 ;
        RECT 2318.010 3229.020 2318.330 3229.080 ;
      LAYER via ;
        RECT 2318.040 3502.040 2318.300 3502.300 ;
        RECT 2473.980 3502.040 2474.240 3502.300 ;
        RECT 2311.600 3229.020 2311.860 3229.280 ;
        RECT 2318.040 3229.020 2318.300 3229.280 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3502.330 2474.180 3517.600 ;
        RECT 2318.040 3502.010 2318.300 3502.330 ;
        RECT 2473.980 3502.010 2474.240 3502.330 ;
        RECT 2318.100 3229.310 2318.240 3502.010 ;
        RECT 2311.600 3228.990 2311.860 3229.310 ;
        RECT 2318.040 3228.990 2318.300 3229.310 ;
        RECT 2311.660 3216.000 2311.800 3228.990 ;
        RECT 2311.550 3212.000 2311.830 3216.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 3501.900 2056.130 3501.960 ;
        RECT 2149.190 3501.900 2149.510 3501.960 ;
        RECT 2055.810 3501.760 2149.510 3501.900 ;
        RECT 2055.810 3501.700 2056.130 3501.760 ;
        RECT 2149.190 3501.700 2149.510 3501.760 ;
      LAYER via ;
        RECT 2055.840 3501.700 2056.100 3501.960 ;
        RECT 2149.220 3501.700 2149.480 3501.960 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3501.990 2149.420 3517.600 ;
        RECT 2055.840 3501.670 2056.100 3501.990 ;
        RECT 2149.220 3501.670 2149.480 3501.990 ;
        RECT 2055.900 3216.000 2056.040 3501.670 ;
        RECT 2055.790 3212.000 2056.070 3216.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.510 3498.500 1800.830 3498.560 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1800.510 3498.360 1825.210 3498.500 ;
        RECT 1800.510 3498.300 1800.830 3498.360 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
      LAYER via ;
        RECT 1800.540 3498.300 1800.800 3498.560 ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1800.540 3498.270 1800.800 3498.590 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1800.600 3216.000 1800.740 3498.270 ;
        RECT 1800.490 3212.000 1800.770 3216.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 3224.460 1504.130 3224.520 ;
        RECT 1544.750 3224.460 1545.070 3224.520 ;
        RECT 1503.810 3224.320 1545.070 3224.460 ;
        RECT 1503.810 3224.260 1504.130 3224.320 ;
        RECT 1544.750 3224.260 1545.070 3224.320 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 3224.260 1504.100 3224.520 ;
        RECT 1544.780 3224.260 1545.040 3224.520 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3224.550 1504.040 3498.270 ;
        RECT 1503.840 3224.230 1504.100 3224.550 ;
        RECT 1544.780 3224.230 1545.040 3224.550 ;
        RECT 1544.840 3216.000 1544.980 3224.230 ;
        RECT 1544.730 3212.000 1545.010 3216.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 324.260 2619.630 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2619.310 324.120 2899.310 324.260 ;
        RECT 2619.310 324.060 2619.630 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2619.340 324.060 2619.600 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2619.330 449.635 2619.610 450.005 ;
        RECT 2619.400 324.350 2619.540 449.635 ;
        RECT 2619.340 324.030 2619.600 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2619.330 449.680 2619.610 449.960 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2619.305 449.970 2619.635 449.985 ;
        RECT 2609.580 449.880 2619.635 449.970 ;
        RECT 2606.000 449.670 2619.635 449.880 ;
        RECT 2606.000 449.280 2610.000 449.670 ;
        RECT 2619.305 449.655 2619.635 449.670 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3225.820 1179.830 3225.880 ;
        RECT 1289.450 3225.820 1289.770 3225.880 ;
        RECT 1179.510 3225.680 1289.770 3225.820 ;
        RECT 1179.510 3225.620 1179.830 3225.680 ;
        RECT 1289.450 3225.620 1289.770 3225.680 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3225.620 1179.800 3225.880 ;
        RECT 1289.480 3225.620 1289.740 3225.880 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3225.910 1179.740 3498.270 ;
        RECT 1179.540 3225.590 1179.800 3225.910 ;
        RECT 1289.480 3225.590 1289.740 3225.910 ;
        RECT 1289.540 3216.000 1289.680 3225.590 ;
        RECT 1289.430 3212.000 1289.710 3216.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 855.210 3501.220 855.530 3501.280 ;
        RECT 851.530 3501.080 855.530 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 855.210 3501.020 855.530 3501.080 ;
        RECT 855.210 3226.160 855.530 3226.220 ;
        RECT 1033.690 3226.160 1034.010 3226.220 ;
        RECT 855.210 3226.020 1034.010 3226.160 ;
        RECT 855.210 3225.960 855.530 3226.020 ;
        RECT 1033.690 3225.960 1034.010 3226.020 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 855.240 3501.020 855.500 3501.280 ;
        RECT 855.240 3225.960 855.500 3226.220 ;
        RECT 1033.720 3225.960 1033.980 3226.220 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 855.240 3500.990 855.500 3501.310 ;
        RECT 855.300 3226.250 855.440 3500.990 ;
        RECT 855.240 3225.930 855.500 3226.250 ;
        RECT 1033.720 3225.930 1033.980 3226.250 ;
        RECT 1033.780 3216.000 1033.920 3225.930 ;
        RECT 1033.670 3212.000 1033.950 3216.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 3226.160 531.230 3226.220 ;
        RECT 777.930 3226.160 778.250 3226.220 ;
        RECT 530.910 3226.020 778.250 3226.160 ;
        RECT 530.910 3225.960 531.230 3226.020 ;
        RECT 777.930 3225.960 778.250 3226.020 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 3225.960 531.200 3226.220 ;
        RECT 777.960 3225.960 778.220 3226.220 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 3226.250 531.140 3498.270 ;
        RECT 530.940 3225.930 531.200 3226.250 ;
        RECT 777.960 3225.930 778.220 3226.250 ;
        RECT 778.020 3216.000 778.160 3225.930 ;
        RECT 777.910 3212.000 778.190 3216.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 3226.500 206.930 3226.560 ;
        RECT 522.630 3226.500 522.950 3226.560 ;
        RECT 206.610 3226.360 522.950 3226.500 ;
        RECT 206.610 3226.300 206.930 3226.360 ;
        RECT 522.630 3226.300 522.950 3226.360 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 3226.300 206.900 3226.560 ;
        RECT 522.660 3226.300 522.920 3226.560 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 3226.590 206.840 3501.670 ;
        RECT 206.640 3226.270 206.900 3226.590 ;
        RECT 522.660 3226.270 522.920 3226.590 ;
        RECT 522.720 3216.000 522.860 3226.270 ;
        RECT 522.610 3212.000 522.890 3216.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3180.940 17.410 3181.000 ;
        RECT 296.770 3180.940 297.090 3181.000 ;
        RECT 17.090 3180.800 297.090 3180.940 ;
        RECT 17.090 3180.740 17.410 3180.800 ;
        RECT 296.770 3180.740 297.090 3180.800 ;
      LAYER via ;
        RECT 17.120 3180.740 17.380 3181.000 ;
        RECT 296.800 3180.740 297.060 3181.000 ;
      LAYER met2 ;
        RECT 17.110 3411.035 17.390 3411.405 ;
        RECT 17.180 3181.030 17.320 3411.035 ;
        RECT 17.120 3180.710 17.380 3181.030 ;
        RECT 296.800 3180.710 297.060 3181.030 ;
        RECT 296.860 3180.205 297.000 3180.710 ;
        RECT 296.790 3179.835 297.070 3180.205 ;
      LAYER via2 ;
        RECT 17.110 3411.080 17.390 3411.360 ;
        RECT 296.790 3179.880 297.070 3180.160 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.085 3411.370 17.415 3411.385 ;
        RECT -4.800 3411.070 17.415 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.085 3411.055 17.415 3411.070 ;
        RECT 296.765 3180.170 297.095 3180.185 ;
        RECT 296.765 3180.080 310.500 3180.170 ;
        RECT 296.765 3179.870 314.000 3180.080 ;
        RECT 296.765 3179.855 297.095 3179.870 ;
        RECT 310.000 3179.480 314.000 3179.870 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2966.740 17.410 2966.800 ;
        RECT 296.770 2966.740 297.090 2966.800 ;
        RECT 17.090 2966.600 297.090 2966.740 ;
        RECT 17.090 2966.540 17.410 2966.600 ;
        RECT 296.770 2966.540 297.090 2966.600 ;
      LAYER via ;
        RECT 17.120 2966.540 17.380 2966.800 ;
        RECT 296.800 2966.540 297.060 2966.800 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 2966.830 17.320 3124.075 ;
        RECT 17.120 2966.510 17.380 2966.830 ;
        RECT 296.800 2966.510 297.060 2966.830 ;
        RECT 296.860 2966.005 297.000 2966.510 ;
        RECT 296.790 2965.635 297.070 2966.005 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
        RECT 296.790 2965.680 297.070 2965.960 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
        RECT 296.765 2965.970 297.095 2965.985 ;
        RECT 296.765 2965.880 310.500 2965.970 ;
        RECT 296.765 2965.670 314.000 2965.880 ;
        RECT 296.765 2965.655 297.095 2965.670 ;
        RECT 310.000 2965.280 314.000 2965.670 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2752.880 17.410 2752.940 ;
        RECT 296.770 2752.880 297.090 2752.940 ;
        RECT 17.090 2752.740 297.090 2752.880 ;
        RECT 17.090 2752.680 17.410 2752.740 ;
        RECT 296.770 2752.680 297.090 2752.740 ;
      LAYER via ;
        RECT 17.120 2752.680 17.380 2752.940 ;
        RECT 296.800 2752.680 297.060 2752.940 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2752.970 17.320 2836.435 ;
        RECT 17.120 2752.650 17.380 2752.970 ;
        RECT 296.800 2752.650 297.060 2752.970 ;
        RECT 296.860 2751.805 297.000 2752.650 ;
        RECT 296.790 2751.435 297.070 2751.805 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
        RECT 296.790 2751.480 297.070 2751.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
        RECT 296.765 2751.770 297.095 2751.785 ;
        RECT 296.765 2751.680 310.500 2751.770 ;
        RECT 296.765 2751.470 314.000 2751.680 ;
        RECT 296.765 2751.455 297.095 2751.470 ;
        RECT 310.000 2751.080 314.000 2751.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2539.020 16.950 2539.080 ;
        RECT 296.770 2539.020 297.090 2539.080 ;
        RECT 16.630 2538.880 297.090 2539.020 ;
        RECT 16.630 2538.820 16.950 2538.880 ;
        RECT 296.770 2538.820 297.090 2538.880 ;
      LAYER via ;
        RECT 16.660 2538.820 16.920 2539.080 ;
        RECT 296.800 2538.820 297.060 2539.080 ;
      LAYER met2 ;
        RECT 16.650 2549.475 16.930 2549.845 ;
        RECT 16.720 2539.110 16.860 2549.475 ;
        RECT 16.660 2538.790 16.920 2539.110 ;
        RECT 296.800 2538.790 297.060 2539.110 ;
        RECT 296.860 2537.605 297.000 2538.790 ;
        RECT 296.790 2537.235 297.070 2537.605 ;
      LAYER via2 ;
        RECT 16.650 2549.520 16.930 2549.800 ;
        RECT 296.790 2537.280 297.070 2537.560 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.625 2549.810 16.955 2549.825 ;
        RECT -4.800 2549.510 16.955 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.625 2549.495 16.955 2549.510 ;
        RECT 296.765 2537.570 297.095 2537.585 ;
        RECT 296.765 2537.480 310.500 2537.570 ;
        RECT 296.765 2537.270 314.000 2537.480 ;
        RECT 296.765 2537.255 297.095 2537.270 ;
        RECT 310.000 2536.880 314.000 2537.270 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2262.940 17.410 2263.000 ;
        RECT 299.990 2262.940 300.310 2263.000 ;
        RECT 17.090 2262.800 300.310 2262.940 ;
        RECT 17.090 2262.740 17.410 2262.800 ;
        RECT 299.990 2262.740 300.310 2262.800 ;
      LAYER via ;
        RECT 17.120 2262.740 17.380 2263.000 ;
        RECT 300.020 2262.740 300.280 2263.000 ;
      LAYER met2 ;
        RECT 300.010 2323.035 300.290 2323.405 ;
        RECT 300.080 2263.030 300.220 2323.035 ;
        RECT 17.120 2262.710 17.380 2263.030 ;
        RECT 300.020 2262.710 300.280 2263.030 ;
        RECT 17.180 2262.205 17.320 2262.710 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
      LAYER via2 ;
        RECT 300.010 2323.080 300.290 2323.360 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
        RECT 299.985 2323.370 300.315 2323.385 ;
        RECT 299.985 2323.280 310.500 2323.370 ;
        RECT 299.985 2323.070 314.000 2323.280 ;
        RECT 299.985 2323.055 300.315 2323.070 ;
        RECT 310.000 2322.680 314.000 2323.070 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 300.450 1980.060 300.770 1980.120 ;
        RECT 15.710 1979.920 300.770 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 300.450 1979.860 300.770 1979.920 ;
      LAYER via ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 300.480 1979.860 300.740 1980.120 ;
      LAYER met2 ;
        RECT 300.470 2108.835 300.750 2109.205 ;
        RECT 300.540 1980.150 300.680 2108.835 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 300.480 1979.830 300.740 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 300.470 2108.880 300.750 2109.160 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT 300.445 2109.170 300.775 2109.185 ;
        RECT 300.445 2109.080 310.500 2109.170 ;
        RECT 300.445 2108.870 314.000 2109.080 ;
        RECT 300.445 2108.855 300.775 2108.870 ;
        RECT 310.000 2108.480 314.000 2108.870 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 558.860 2619.630 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2619.310 558.720 2899.310 558.860 ;
        RECT 2619.310 558.660 2619.630 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2619.340 558.660 2619.600 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2619.330 649.555 2619.610 649.925 ;
        RECT 2619.400 558.950 2619.540 649.555 ;
        RECT 2619.340 558.630 2619.600 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2619.330 649.600 2619.610 649.880 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2619.305 649.890 2619.635 649.905 ;
        RECT 2609.580 649.800 2619.635 649.890 ;
        RECT 2606.000 649.590 2619.635 649.800 ;
        RECT 2606.000 649.200 2610.000 649.590 ;
        RECT 2619.305 649.575 2619.635 649.590 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 299.990 1690.380 300.310 1690.440 ;
        RECT 17.090 1690.240 300.310 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 299.990 1690.180 300.310 1690.240 ;
      LAYER via ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 300.020 1690.180 300.280 1690.440 ;
      LAYER met2 ;
        RECT 300.010 1894.635 300.290 1895.005 ;
        RECT 300.080 1690.470 300.220 1894.635 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 300.020 1690.150 300.280 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 300.010 1894.680 300.290 1894.960 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT 299.985 1894.970 300.315 1894.985 ;
        RECT 299.985 1894.880 310.500 1894.970 ;
        RECT 299.985 1894.670 314.000 1894.880 ;
        RECT 299.985 1894.655 300.315 1894.670 ;
        RECT 310.000 1894.280 314.000 1894.670 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1476.520 17.410 1476.580 ;
        RECT 301.370 1476.520 301.690 1476.580 ;
        RECT 17.090 1476.380 301.690 1476.520 ;
        RECT 17.090 1476.320 17.410 1476.380 ;
        RECT 301.370 1476.320 301.690 1476.380 ;
      LAYER via ;
        RECT 17.120 1476.320 17.380 1476.580 ;
        RECT 301.400 1476.320 301.660 1476.580 ;
      LAYER met2 ;
        RECT 301.390 1679.755 301.670 1680.125 ;
        RECT 301.460 1476.610 301.600 1679.755 ;
        RECT 17.120 1476.290 17.380 1476.610 ;
        RECT 301.400 1476.290 301.660 1476.610 ;
        RECT 17.180 1472.045 17.320 1476.290 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 301.390 1679.800 301.670 1680.080 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT 301.365 1680.090 301.695 1680.105 ;
        RECT 301.365 1680.000 310.500 1680.090 ;
        RECT 301.365 1679.790 314.000 1680.000 ;
        RECT 301.365 1679.775 301.695 1679.790 ;
        RECT 310.000 1679.400 314.000 1679.790 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1262.660 17.410 1262.720 ;
        RECT 301.370 1262.660 301.690 1262.720 ;
        RECT 17.090 1262.520 301.690 1262.660 ;
        RECT 17.090 1262.460 17.410 1262.520 ;
        RECT 301.370 1262.460 301.690 1262.520 ;
      LAYER via ;
        RECT 17.120 1262.460 17.380 1262.720 ;
        RECT 301.400 1262.460 301.660 1262.720 ;
      LAYER met2 ;
        RECT 301.390 1465.555 301.670 1465.925 ;
        RECT 301.460 1262.750 301.600 1465.555 ;
        RECT 17.120 1262.430 17.380 1262.750 ;
        RECT 301.400 1262.430 301.660 1262.750 ;
        RECT 17.180 1256.485 17.320 1262.430 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
      LAYER via2 ;
        RECT 301.390 1465.600 301.670 1465.880 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
      LAYER met3 ;
        RECT 301.365 1465.890 301.695 1465.905 ;
        RECT 301.365 1465.800 310.500 1465.890 ;
        RECT 301.365 1465.590 314.000 1465.800 ;
        RECT 301.365 1465.575 301.695 1465.590 ;
        RECT 310.000 1465.200 314.000 1465.590 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 299.990 1041.660 300.310 1041.720 ;
        RECT 17.090 1041.520 300.310 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 299.990 1041.460 300.310 1041.520 ;
      LAYER via ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 300.020 1041.460 300.280 1041.720 ;
      LAYER met2 ;
        RECT 300.010 1251.355 300.290 1251.725 ;
        RECT 300.080 1041.750 300.220 1251.355 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 300.020 1041.430 300.280 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 300.010 1251.400 300.290 1251.680 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT 299.985 1251.690 300.315 1251.705 ;
        RECT 299.985 1251.600 310.500 1251.690 ;
        RECT 299.985 1251.390 314.000 1251.600 ;
        RECT 299.985 1251.375 300.315 1251.390 ;
        RECT 310.000 1251.000 314.000 1251.390 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 300.450 827.800 300.770 827.860 ;
        RECT 17.550 827.660 300.770 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 300.450 827.600 300.770 827.660 ;
      LAYER via ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 300.480 827.600 300.740 827.860 ;
      LAYER met2 ;
        RECT 300.470 1037.155 300.750 1037.525 ;
        RECT 300.540 827.890 300.680 1037.155 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 300.480 827.570 300.740 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 300.470 1037.200 300.750 1037.480 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT 300.445 1037.490 300.775 1037.505 ;
        RECT 300.445 1037.400 310.500 1037.490 ;
        RECT 300.445 1037.190 314.000 1037.400 ;
        RECT 300.445 1037.175 300.775 1037.190 ;
        RECT 310.000 1036.800 314.000 1037.190 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 613.940 17.410 614.000 ;
        RECT 299.990 613.940 300.310 614.000 ;
        RECT 17.090 613.800 300.310 613.940 ;
        RECT 17.090 613.740 17.410 613.800 ;
        RECT 299.990 613.740 300.310 613.800 ;
      LAYER via ;
        RECT 17.120 613.740 17.380 614.000 ;
        RECT 300.020 613.740 300.280 614.000 ;
      LAYER met2 ;
        RECT 300.010 822.955 300.290 823.325 ;
        RECT 300.080 614.030 300.220 822.955 ;
        RECT 17.120 613.710 17.380 614.030 ;
        RECT 300.020 613.710 300.280 614.030 ;
        RECT 17.180 610.485 17.320 613.710 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 300.010 823.000 300.290 823.280 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT 299.985 823.290 300.315 823.305 ;
        RECT 299.985 823.200 310.500 823.290 ;
        RECT 299.985 822.990 314.000 823.200 ;
        RECT 299.985 822.975 300.315 822.990 ;
        RECT 310.000 822.600 314.000 822.990 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 400.080 17.410 400.140 ;
        RECT 300.450 400.080 300.770 400.140 ;
        RECT 17.090 399.940 300.770 400.080 ;
        RECT 17.090 399.880 17.410 399.940 ;
        RECT 300.450 399.880 300.770 399.940 ;
      LAYER via ;
        RECT 17.120 399.880 17.380 400.140 ;
        RECT 300.480 399.880 300.740 400.140 ;
      LAYER met2 ;
        RECT 300.470 608.755 300.750 609.125 ;
        RECT 300.540 400.170 300.680 608.755 ;
        RECT 17.120 399.850 17.380 400.170 ;
        RECT 300.480 399.850 300.740 400.170 ;
        RECT 17.180 394.925 17.320 399.850 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 300.470 608.800 300.750 609.080 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT 300.445 609.090 300.775 609.105 ;
        RECT 300.445 609.000 310.500 609.090 ;
        RECT 300.445 608.790 314.000 609.000 ;
        RECT 300.445 608.775 300.775 608.790 ;
        RECT 310.000 608.400 314.000 608.790 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 299.990 179.420 300.310 179.480 ;
        RECT 17.090 179.280 300.310 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 299.990 179.220 300.310 179.280 ;
      LAYER via ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 300.020 179.220 300.280 179.480 ;
      LAYER met2 ;
        RECT 300.010 394.555 300.290 394.925 ;
        RECT 300.080 179.510 300.220 394.555 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 300.020 179.190 300.280 179.510 ;
      LAYER via2 ;
        RECT 300.010 394.600 300.290 394.880 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 299.985 394.890 300.315 394.905 ;
        RECT 299.985 394.800 310.500 394.890 ;
        RECT 299.985 394.590 314.000 394.800 ;
        RECT 299.985 394.575 300.315 394.590 ;
        RECT 310.000 394.200 314.000 394.590 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 793.460 2618.710 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2618.390 793.320 2899.310 793.460 ;
        RECT 2618.390 793.260 2618.710 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2618.420 793.260 2618.680 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2618.410 849.475 2618.690 849.845 ;
        RECT 2618.480 793.550 2618.620 849.475 ;
        RECT 2618.420 793.230 2618.680 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2618.410 849.520 2618.690 849.800 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2618.385 849.810 2618.715 849.825 ;
        RECT 2609.580 849.720 2618.715 849.810 ;
        RECT 2606.000 849.510 2618.715 849.720 ;
        RECT 2606.000 849.120 2610.000 849.510 ;
        RECT 2618.385 849.495 2618.715 849.510 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2617.010 1028.060 2617.330 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2617.010 1027.920 2899.310 1028.060 ;
        RECT 2617.010 1027.860 2617.330 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2617.040 1027.860 2617.300 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2617.030 1049.395 2617.310 1049.765 ;
        RECT 2617.100 1028.150 2617.240 1049.395 ;
        RECT 2617.040 1027.830 2617.300 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2617.030 1049.440 2617.310 1049.720 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2617.005 1049.730 2617.335 1049.745 ;
        RECT 2609.580 1049.640 2617.335 1049.730 ;
        RECT 2606.000 1049.430 2617.335 1049.640 ;
        RECT 2606.000 1049.040 2610.000 1049.430 ;
        RECT 2617.005 1049.415 2617.335 1049.430 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.770 1256.200 2620.090 1256.260 ;
        RECT 2900.830 1256.200 2901.150 1256.260 ;
        RECT 2619.770 1256.060 2901.150 1256.200 ;
        RECT 2619.770 1256.000 2620.090 1256.060 ;
        RECT 2900.830 1256.000 2901.150 1256.060 ;
      LAYER via ;
        RECT 2619.800 1256.000 2620.060 1256.260 ;
        RECT 2900.860 1256.000 2901.120 1256.260 ;
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 1256.290 2901.060 1260.875 ;
        RECT 2619.800 1255.970 2620.060 1256.290 ;
        RECT 2900.860 1255.970 2901.120 1256.290 ;
        RECT 2619.860 1249.685 2620.000 1255.970 ;
        RECT 2619.790 1249.315 2620.070 1249.685 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 2619.790 1249.360 2620.070 1249.640 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2619.765 1249.650 2620.095 1249.665 ;
        RECT 2609.580 1249.560 2620.095 1249.650 ;
        RECT 2606.000 1249.350 2620.095 1249.560 ;
        RECT 2606.000 1248.960 2610.000 1249.350 ;
        RECT 2619.765 1249.335 2620.095 1249.350 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2616.090 1490.800 2616.410 1490.860 ;
        RECT 2900.830 1490.800 2901.150 1490.860 ;
        RECT 2616.090 1490.660 2901.150 1490.800 ;
        RECT 2616.090 1490.600 2616.410 1490.660 ;
        RECT 2900.830 1490.600 2901.150 1490.660 ;
      LAYER via ;
        RECT 2616.120 1490.600 2616.380 1490.860 ;
        RECT 2900.860 1490.600 2901.120 1490.860 ;
      LAYER met2 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
        RECT 2900.920 1490.890 2901.060 1495.475 ;
        RECT 2616.120 1490.570 2616.380 1490.890 ;
        RECT 2900.860 1490.570 2901.120 1490.890 ;
        RECT 2616.180 1449.605 2616.320 1490.570 ;
        RECT 2616.110 1449.235 2616.390 1449.605 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
        RECT 2616.110 1449.280 2616.390 1449.560 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2616.085 1449.570 2616.415 1449.585 ;
        RECT 2609.580 1449.480 2616.415 1449.570 ;
        RECT 2606.000 1449.270 2616.415 1449.480 ;
        RECT 2606.000 1448.880 2610.000 1449.270 ;
        RECT 2616.085 1449.255 2616.415 1449.270 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1725.400 2618.710 1725.460 ;
        RECT 2900.830 1725.400 2901.150 1725.460 ;
        RECT 2618.390 1725.260 2901.150 1725.400 ;
        RECT 2618.390 1725.200 2618.710 1725.260 ;
        RECT 2900.830 1725.200 2901.150 1725.260 ;
      LAYER via ;
        RECT 2618.420 1725.200 2618.680 1725.460 ;
        RECT 2900.860 1725.200 2901.120 1725.460 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 2900.920 1725.490 2901.060 1730.075 ;
        RECT 2618.420 1725.170 2618.680 1725.490 ;
        RECT 2900.860 1725.170 2901.120 1725.490 ;
        RECT 2618.480 1649.525 2618.620 1725.170 ;
        RECT 2618.410 1649.155 2618.690 1649.525 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
        RECT 2618.410 1649.200 2618.690 1649.480 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2618.385 1649.490 2618.715 1649.505 ;
        RECT 2609.580 1649.400 2618.715 1649.490 ;
        RECT 2606.000 1649.190 2618.715 1649.400 ;
        RECT 2606.000 1648.800 2610.000 1649.190 ;
        RECT 2618.385 1649.175 2618.715 1649.190 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1960.000 2619.170 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 2618.850 1959.860 2901.150 1960.000 ;
        RECT 2618.850 1959.800 2619.170 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
      LAYER via ;
        RECT 2618.880 1959.800 2619.140 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 2618.880 1959.770 2619.140 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 2618.940 1850.125 2619.080 1959.770 ;
        RECT 2618.870 1849.755 2619.150 1850.125 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
        RECT 2618.870 1849.800 2619.150 1850.080 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2618.845 1850.090 2619.175 1850.105 ;
        RECT 2609.580 1850.000 2619.175 1850.090 ;
        RECT 2606.000 1849.790 2619.175 1850.000 ;
        RECT 2606.000 1849.400 2610.000 1849.790 ;
        RECT 2618.845 1849.775 2619.175 1849.790 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2194.600 2618.710 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2618.390 2194.460 2901.150 2194.600 ;
        RECT 2618.390 2194.400 2618.710 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
      LAYER via ;
        RECT 2618.420 2194.400 2618.680 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2618.420 2194.370 2618.680 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2618.480 2050.045 2618.620 2194.370 ;
        RECT 2618.410 2049.675 2618.690 2050.045 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2618.410 2049.720 2618.690 2050.000 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2618.385 2050.010 2618.715 2050.025 ;
        RECT 2609.580 2049.920 2618.715 2050.010 ;
        RECT 2606.000 2049.710 2618.715 2049.920 ;
        RECT 2606.000 2049.320 2610.000 2049.710 ;
        RECT 2618.385 2049.695 2618.715 2049.710 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 206.960 2618.710 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2618.390 206.820 2901.150 206.960 ;
        RECT 2618.390 206.760 2618.710 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2618.420 206.760 2618.680 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2618.410 382.995 2618.690 383.365 ;
        RECT 2618.480 207.050 2618.620 382.995 ;
        RECT 2618.420 206.730 2618.680 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2618.410 383.040 2618.690 383.320 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2618.385 383.330 2618.715 383.345 ;
        RECT 2609.580 383.240 2618.715 383.330 ;
        RECT 2606.000 383.030 2618.715 383.240 ;
        RECT 2606.000 382.640 2610.000 383.030 ;
        RECT 2618.385 383.015 2618.715 383.030 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.310 2546.500 2619.630 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2619.310 2546.360 2901.150 2546.500 ;
        RECT 2619.310 2546.300 2619.630 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
      LAYER via ;
        RECT 2619.340 2546.300 2619.600 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2619.340 2546.270 2619.600 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2619.400 2383.245 2619.540 2546.270 ;
        RECT 2619.330 2382.875 2619.610 2383.245 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2619.330 2382.920 2619.610 2383.200 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2619.305 2383.210 2619.635 2383.225 ;
        RECT 2609.580 2383.120 2619.635 2383.210 ;
        RECT 2606.000 2382.910 2619.635 2383.120 ;
        RECT 2606.000 2382.520 2610.000 2382.910 ;
        RECT 2619.305 2382.895 2619.635 2382.910 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.310 2781.100 2619.630 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2619.310 2780.960 2901.150 2781.100 ;
        RECT 2619.310 2780.900 2619.630 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 2619.340 2780.900 2619.600 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2619.340 2780.870 2619.600 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2619.400 2583.165 2619.540 2780.870 ;
        RECT 2619.330 2582.795 2619.610 2583.165 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2619.330 2582.840 2619.610 2583.120 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2619.305 2583.130 2619.635 2583.145 ;
        RECT 2609.580 2583.040 2619.635 2583.130 ;
        RECT 2606.000 2582.830 2619.635 2583.040 ;
        RECT 2606.000 2582.440 2610.000 2582.830 ;
        RECT 2619.305 2582.815 2619.635 2582.830 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3015.700 2619.170 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2618.850 3015.560 2901.150 3015.700 ;
        RECT 2618.850 3015.500 2619.170 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 2618.880 3015.500 2619.140 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2618.880 3015.470 2619.140 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 2618.940 2783.085 2619.080 3015.470 ;
        RECT 2618.870 2782.715 2619.150 2783.085 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 2618.870 2782.760 2619.150 2783.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2618.845 2783.050 2619.175 2783.065 ;
        RECT 2609.580 2782.960 2619.175 2783.050 ;
        RECT 2606.000 2782.750 2619.175 2782.960 ;
        RECT 2606.000 2782.360 2610.000 2782.750 ;
        RECT 2618.845 2782.735 2619.175 2782.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2987.480 2618.710 2987.540 ;
        RECT 2902.210 2987.480 2902.530 2987.540 ;
        RECT 2618.390 2987.340 2902.530 2987.480 ;
        RECT 2618.390 2987.280 2618.710 2987.340 ;
        RECT 2902.210 2987.280 2902.530 2987.340 ;
      LAYER via ;
        RECT 2618.420 2987.280 2618.680 2987.540 ;
        RECT 2902.240 2987.280 2902.500 2987.540 ;
      LAYER met2 ;
        RECT 2902.230 3255.315 2902.510 3255.685 ;
        RECT 2902.300 2987.570 2902.440 3255.315 ;
        RECT 2618.420 2987.250 2618.680 2987.570 ;
        RECT 2902.240 2987.250 2902.500 2987.570 ;
        RECT 2618.480 2983.005 2618.620 2987.250 ;
        RECT 2618.410 2982.635 2618.690 2983.005 ;
      LAYER via2 ;
        RECT 2902.230 3255.360 2902.510 3255.640 ;
        RECT 2618.410 2982.680 2618.690 2982.960 ;
      LAYER met3 ;
        RECT 2902.205 3255.650 2902.535 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2902.205 3255.350 2924.800 3255.650 ;
        RECT 2902.205 3255.335 2902.535 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2618.385 2982.970 2618.715 2982.985 ;
        RECT 2609.580 2982.880 2618.715 2982.970 ;
        RECT 2606.000 2982.670 2618.715 2982.880 ;
        RECT 2606.000 2982.280 2610.000 2982.670 ;
        RECT 2618.385 2982.655 2618.715 2982.670 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3484.900 2619.170 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2618.850 3484.760 2901.150 3484.900 ;
        RECT 2618.850 3484.700 2619.170 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 2618.880 3484.700 2619.140 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2618.880 3484.670 2619.140 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2618.940 3182.925 2619.080 3484.670 ;
        RECT 2618.870 3182.555 2619.150 3182.925 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2618.870 3182.600 2619.150 3182.880 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2618.845 3182.890 2619.175 3182.905 ;
        RECT 2609.580 3182.800 2619.175 3182.890 ;
        RECT 2606.000 3182.590 2619.175 3182.800 ;
        RECT 2606.000 3182.200 2610.000 3182.590 ;
        RECT 2618.845 3182.575 2619.175 3182.590 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2400.810 3501.560 2401.130 3501.620 ;
        RECT 2635.870 3501.560 2636.190 3501.620 ;
        RECT 2400.810 3501.420 2636.190 3501.560 ;
        RECT 2400.810 3501.360 2401.130 3501.420 ;
        RECT 2635.870 3501.360 2636.190 3501.420 ;
        RECT 2396.670 3229.220 2396.990 3229.280 ;
        RECT 2400.810 3229.220 2401.130 3229.280 ;
        RECT 2396.670 3229.080 2401.130 3229.220 ;
        RECT 2396.670 3229.020 2396.990 3229.080 ;
        RECT 2400.810 3229.020 2401.130 3229.080 ;
      LAYER via ;
        RECT 2400.840 3501.360 2401.100 3501.620 ;
        RECT 2635.900 3501.360 2636.160 3501.620 ;
        RECT 2396.700 3229.020 2396.960 3229.280 ;
        RECT 2400.840 3229.020 2401.100 3229.280 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.650 2636.100 3517.600 ;
        RECT 2400.840 3501.330 2401.100 3501.650 ;
        RECT 2635.900 3501.330 2636.160 3501.650 ;
        RECT 2400.900 3229.310 2401.040 3501.330 ;
        RECT 2396.700 3228.990 2396.960 3229.310 ;
        RECT 2400.840 3228.990 2401.100 3229.310 ;
        RECT 2396.760 3216.000 2396.900 3228.990 ;
        RECT 2396.650 3212.000 2396.930 3216.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2145.510 3501.560 2145.830 3501.620 ;
        RECT 2311.570 3501.560 2311.890 3501.620 ;
        RECT 2145.510 3501.420 2311.890 3501.560 ;
        RECT 2145.510 3501.360 2145.830 3501.420 ;
        RECT 2311.570 3501.360 2311.890 3501.420 ;
        RECT 2140.910 3229.220 2141.230 3229.280 ;
        RECT 2145.510 3229.220 2145.830 3229.280 ;
        RECT 2140.910 3229.080 2145.830 3229.220 ;
        RECT 2140.910 3229.020 2141.230 3229.080 ;
        RECT 2145.510 3229.020 2145.830 3229.080 ;
      LAYER via ;
        RECT 2145.540 3501.360 2145.800 3501.620 ;
        RECT 2311.600 3501.360 2311.860 3501.620 ;
        RECT 2140.940 3229.020 2141.200 3229.280 ;
        RECT 2145.540 3229.020 2145.800 3229.280 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.650 2311.800 3517.600 ;
        RECT 2145.540 3501.330 2145.800 3501.650 ;
        RECT 2311.600 3501.330 2311.860 3501.650 ;
        RECT 2145.600 3229.310 2145.740 3501.330 ;
        RECT 2140.940 3228.990 2141.200 3229.310 ;
        RECT 2145.540 3228.990 2145.800 3229.310 ;
        RECT 2141.000 3216.000 2141.140 3228.990 ;
        RECT 2140.890 3212.000 2141.170 3216.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1890.210 3501.560 1890.530 3501.620 ;
        RECT 1987.270 3501.560 1987.590 3501.620 ;
        RECT 1890.210 3501.420 1987.590 3501.560 ;
        RECT 1890.210 3501.360 1890.530 3501.420 ;
        RECT 1987.270 3501.360 1987.590 3501.420 ;
        RECT 1885.610 3229.220 1885.930 3229.280 ;
        RECT 1890.210 3229.220 1890.530 3229.280 ;
        RECT 1885.610 3229.080 1890.530 3229.220 ;
        RECT 1885.610 3229.020 1885.930 3229.080 ;
        RECT 1890.210 3229.020 1890.530 3229.080 ;
      LAYER via ;
        RECT 1890.240 3501.360 1890.500 3501.620 ;
        RECT 1987.300 3501.360 1987.560 3501.620 ;
        RECT 1885.640 3229.020 1885.900 3229.280 ;
        RECT 1890.240 3229.020 1890.500 3229.280 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3501.650 1987.500 3517.600 ;
        RECT 1890.240 3501.330 1890.500 3501.650 ;
        RECT 1987.300 3501.330 1987.560 3501.650 ;
        RECT 1890.300 3229.310 1890.440 3501.330 ;
        RECT 1885.640 3228.990 1885.900 3229.310 ;
        RECT 1890.240 3228.990 1890.500 3229.310 ;
        RECT 1885.700 3216.000 1885.840 3228.990 ;
        RECT 1885.590 3212.000 1885.870 3216.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1634.910 3498.500 1635.230 3498.560 ;
        RECT 1662.510 3498.500 1662.830 3498.560 ;
        RECT 1634.910 3498.360 1662.830 3498.500 ;
        RECT 1634.910 3498.300 1635.230 3498.360 ;
        RECT 1662.510 3498.300 1662.830 3498.360 ;
        RECT 1629.850 3227.520 1630.170 3227.580 ;
        RECT 1634.910 3227.520 1635.230 3227.580 ;
        RECT 1629.850 3227.380 1635.230 3227.520 ;
        RECT 1629.850 3227.320 1630.170 3227.380 ;
        RECT 1634.910 3227.320 1635.230 3227.380 ;
      LAYER via ;
        RECT 1634.940 3498.300 1635.200 3498.560 ;
        RECT 1662.540 3498.300 1662.800 3498.560 ;
        RECT 1629.880 3227.320 1630.140 3227.580 ;
        RECT 1634.940 3227.320 1635.200 3227.580 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3498.590 1662.740 3517.600 ;
        RECT 1634.940 3498.270 1635.200 3498.590 ;
        RECT 1662.540 3498.270 1662.800 3498.590 ;
        RECT 1635.000 3227.610 1635.140 3498.270 ;
        RECT 1629.880 3227.290 1630.140 3227.610 ;
        RECT 1634.940 3227.290 1635.200 3227.610 ;
        RECT 1629.940 3216.000 1630.080 3227.290 ;
        RECT 1629.830 3212.000 1630.110 3216.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3225.820 1338.530 3225.880 ;
        RECT 1374.550 3225.820 1374.870 3225.880 ;
        RECT 1338.210 3225.680 1374.870 3225.820 ;
        RECT 1338.210 3225.620 1338.530 3225.680 ;
        RECT 1374.550 3225.620 1374.870 3225.680 ;
      LAYER via ;
        RECT 1338.240 3225.620 1338.500 3225.880 ;
        RECT 1374.580 3225.620 1374.840 3225.880 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3225.910 1338.440 3517.600 ;
        RECT 1338.240 3225.590 1338.500 3225.910 ;
        RECT 1374.580 3225.590 1374.840 3225.910 ;
        RECT 1374.640 3216.000 1374.780 3225.590 ;
        RECT 1374.530 3212.000 1374.810 3216.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 441.560 2618.710 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2618.390 441.420 2901.150 441.560 ;
        RECT 2618.390 441.360 2618.710 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2618.420 441.360 2618.680 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2618.410 582.915 2618.690 583.285 ;
        RECT 2618.480 441.650 2618.620 582.915 ;
        RECT 2618.420 441.330 2618.680 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2618.410 582.960 2618.690 583.240 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2618.385 583.250 2618.715 583.265 ;
        RECT 2609.580 583.160 2618.715 583.250 ;
        RECT 2606.000 582.950 2618.715 583.160 ;
        RECT 2606.000 582.560 2610.000 582.950 ;
        RECT 2618.385 582.935 2618.715 582.950 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3225.820 1014.230 3225.880 ;
        RECT 1118.790 3225.820 1119.110 3225.880 ;
        RECT 1013.910 3225.680 1119.110 3225.820 ;
        RECT 1013.910 3225.620 1014.230 3225.680 ;
        RECT 1118.790 3225.620 1119.110 3225.680 ;
      LAYER via ;
        RECT 1013.940 3225.620 1014.200 3225.880 ;
        RECT 1118.820 3225.620 1119.080 3225.880 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3225.910 1014.140 3517.600 ;
        RECT 1013.940 3225.590 1014.200 3225.910 ;
        RECT 1118.820 3225.590 1119.080 3225.910 ;
        RECT 1118.880 3216.000 1119.020 3225.590 ;
        RECT 1118.770 3212.000 1119.050 3216.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 689.225 3429.325 689.395 3477.435 ;
      LAYER mcon ;
        RECT 689.225 3477.265 689.395 3477.435 ;
      LAYER met1 ;
        RECT 688.690 3491.360 689.010 3491.420 ;
        RECT 689.610 3491.360 689.930 3491.420 ;
        RECT 688.690 3491.220 689.930 3491.360 ;
        RECT 688.690 3491.160 689.010 3491.220 ;
        RECT 689.610 3491.160 689.930 3491.220 ;
        RECT 689.165 3477.420 689.455 3477.465 ;
        RECT 689.610 3477.420 689.930 3477.480 ;
        RECT 689.165 3477.280 689.930 3477.420 ;
        RECT 689.165 3477.235 689.455 3477.280 ;
        RECT 689.610 3477.220 689.930 3477.280 ;
        RECT 689.150 3429.480 689.470 3429.540 ;
        RECT 688.955 3429.340 689.470 3429.480 ;
        RECT 689.150 3429.280 689.470 3429.340 ;
        RECT 689.150 3395.140 689.470 3395.200 ;
        RECT 688.780 3395.000 689.470 3395.140 ;
        RECT 688.780 3394.860 688.920 3395.000 ;
        RECT 689.150 3394.940 689.470 3395.000 ;
        RECT 688.690 3394.600 689.010 3394.860 ;
        RECT 688.690 3367.600 689.010 3367.660 ;
        RECT 689.610 3367.600 689.930 3367.660 ;
        RECT 688.690 3367.460 689.930 3367.600 ;
        RECT 688.690 3367.400 689.010 3367.460 ;
        RECT 689.610 3367.400 689.930 3367.460 ;
        RECT 688.690 3270.700 689.010 3270.760 ;
        RECT 689.610 3270.700 689.930 3270.760 ;
        RECT 688.690 3270.560 689.930 3270.700 ;
        RECT 688.690 3270.500 689.010 3270.560 ;
        RECT 689.610 3270.500 689.930 3270.560 ;
        RECT 689.610 3226.500 689.930 3226.560 ;
        RECT 863.490 3226.500 863.810 3226.560 ;
        RECT 689.610 3226.360 863.810 3226.500 ;
        RECT 689.610 3226.300 689.930 3226.360 ;
        RECT 863.490 3226.300 863.810 3226.360 ;
      LAYER via ;
        RECT 688.720 3491.160 688.980 3491.420 ;
        RECT 689.640 3491.160 689.900 3491.420 ;
        RECT 689.640 3477.220 689.900 3477.480 ;
        RECT 689.180 3429.280 689.440 3429.540 ;
        RECT 689.180 3394.940 689.440 3395.200 ;
        RECT 688.720 3394.600 688.980 3394.860 ;
        RECT 688.720 3367.400 688.980 3367.660 ;
        RECT 689.640 3367.400 689.900 3367.660 ;
        RECT 688.720 3270.500 688.980 3270.760 ;
        RECT 689.640 3270.500 689.900 3270.760 ;
        RECT 689.640 3226.300 689.900 3226.560 ;
        RECT 863.520 3226.300 863.780 3226.560 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.780 3517.230 689.380 3517.370 ;
        RECT 688.780 3491.450 688.920 3517.230 ;
        RECT 688.720 3491.130 688.980 3491.450 ;
        RECT 689.640 3491.130 689.900 3491.450 ;
        RECT 689.700 3477.510 689.840 3491.130 ;
        RECT 689.640 3477.190 689.900 3477.510 ;
        RECT 689.180 3429.250 689.440 3429.570 ;
        RECT 689.240 3395.230 689.380 3429.250 ;
        RECT 689.180 3394.910 689.440 3395.230 ;
        RECT 688.720 3394.570 688.980 3394.890 ;
        RECT 688.780 3367.690 688.920 3394.570 ;
        RECT 688.720 3367.370 688.980 3367.690 ;
        RECT 689.640 3367.370 689.900 3367.690 ;
        RECT 689.700 3318.810 689.840 3367.370 ;
        RECT 688.780 3318.670 689.840 3318.810 ;
        RECT 688.780 3270.790 688.920 3318.670 ;
        RECT 688.720 3270.470 688.980 3270.790 ;
        RECT 689.640 3270.470 689.900 3270.790 ;
        RECT 689.700 3226.590 689.840 3270.470 ;
        RECT 689.640 3226.270 689.900 3226.590 ;
        RECT 863.520 3226.270 863.780 3226.590 ;
        RECT 863.580 3216.000 863.720 3226.270 ;
        RECT 863.470 3212.000 863.750 3216.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 362.625 3422.865 362.795 3470.635 ;
        RECT 364.005 3380.365 364.175 3422.355 ;
      LAYER mcon ;
        RECT 362.625 3470.465 362.795 3470.635 ;
        RECT 364.005 3422.185 364.175 3422.355 ;
      LAYER met1 ;
        RECT 362.565 3470.620 362.855 3470.665 ;
        RECT 363.470 3470.620 363.790 3470.680 ;
        RECT 362.565 3470.480 363.790 3470.620 ;
        RECT 362.565 3470.435 362.855 3470.480 ;
        RECT 363.470 3470.420 363.790 3470.480 ;
        RECT 362.550 3423.020 362.870 3423.080 ;
        RECT 362.355 3422.880 362.870 3423.020 ;
        RECT 362.550 3422.820 362.870 3422.880 ;
        RECT 362.550 3422.340 362.870 3422.400 ;
        RECT 363.945 3422.340 364.235 3422.385 ;
        RECT 362.550 3422.200 364.235 3422.340 ;
        RECT 362.550 3422.140 362.870 3422.200 ;
        RECT 363.945 3422.155 364.235 3422.200 ;
        RECT 363.930 3380.520 364.250 3380.580 ;
        RECT 363.735 3380.380 364.250 3380.520 ;
        RECT 363.930 3380.320 364.250 3380.380 ;
        RECT 363.930 3346.660 364.250 3346.920 ;
        RECT 364.020 3346.240 364.160 3346.660 ;
        RECT 363.930 3345.980 364.250 3346.240 ;
        RECT 365.310 3226.840 365.630 3226.900 ;
        RECT 607.730 3226.840 608.050 3226.900 ;
        RECT 365.310 3226.700 608.050 3226.840 ;
        RECT 365.310 3226.640 365.630 3226.700 ;
        RECT 607.730 3226.640 608.050 3226.700 ;
      LAYER via ;
        RECT 363.500 3470.420 363.760 3470.680 ;
        RECT 362.580 3422.820 362.840 3423.080 ;
        RECT 362.580 3422.140 362.840 3422.400 ;
        RECT 363.960 3380.320 364.220 3380.580 ;
        RECT 363.960 3346.660 364.220 3346.920 ;
        RECT 363.960 3345.980 364.220 3346.240 ;
        RECT 365.340 3226.640 365.600 3226.900 ;
        RECT 607.760 3226.640 608.020 3226.900 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3470.710 363.700 3491.390 ;
        RECT 363.500 3470.390 363.760 3470.710 ;
        RECT 362.580 3422.790 362.840 3423.110 ;
        RECT 362.640 3422.430 362.780 3422.790 ;
        RECT 362.580 3422.110 362.840 3422.430 ;
        RECT 363.960 3380.290 364.220 3380.610 ;
        RECT 364.020 3346.950 364.160 3380.290 ;
        RECT 363.960 3346.630 364.220 3346.950 ;
        RECT 363.960 3345.950 364.220 3346.270 ;
        RECT 364.020 3298.410 364.160 3345.950 ;
        RECT 364.020 3298.270 365.080 3298.410 ;
        RECT 364.940 3250.130 365.080 3298.270 ;
        RECT 364.940 3249.990 365.540 3250.130 ;
        RECT 365.400 3226.930 365.540 3249.990 ;
        RECT 365.340 3226.610 365.600 3226.930 ;
        RECT 607.760 3226.610 608.020 3226.930 ;
        RECT 607.820 3216.000 607.960 3226.610 ;
        RECT 607.710 3212.000 607.990 3216.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 41.010 3226.160 41.330 3226.220 ;
        RECT 352.430 3226.160 352.750 3226.220 ;
        RECT 41.010 3226.020 352.750 3226.160 ;
        RECT 41.010 3225.960 41.330 3226.020 ;
        RECT 352.430 3225.960 352.750 3226.020 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 41.040 3225.960 41.300 3226.220 ;
        RECT 352.460 3225.960 352.720 3226.220 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3226.250 41.240 3270.470 ;
        RECT 41.040 3225.930 41.300 3226.250 ;
        RECT 352.460 3225.930 352.720 3226.250 ;
        RECT 352.520 3216.000 352.660 3225.930 ;
        RECT 352.410 3212.000 352.690 3216.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 3042.900 18.330 3042.960 ;
        RECT 296.770 3042.900 297.090 3042.960 ;
        RECT 18.010 3042.760 297.090 3042.900 ;
        RECT 18.010 3042.700 18.330 3042.760 ;
        RECT 296.770 3042.700 297.090 3042.760 ;
      LAYER via ;
        RECT 18.040 3042.700 18.300 3042.960 ;
        RECT 296.800 3042.700 297.060 3042.960 ;
      LAYER met2 ;
        RECT 18.030 3267.555 18.310 3267.925 ;
        RECT 18.100 3042.990 18.240 3267.555 ;
        RECT 18.040 3042.670 18.300 3042.990 ;
        RECT 296.800 3042.670 297.060 3042.990 ;
        RECT 296.860 3037.405 297.000 3042.670 ;
        RECT 296.790 3037.035 297.070 3037.405 ;
      LAYER via2 ;
        RECT 18.030 3267.600 18.310 3267.880 ;
        RECT 296.790 3037.080 297.070 3037.360 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 18.005 3267.890 18.335 3267.905 ;
        RECT -4.800 3267.590 18.335 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 18.005 3267.575 18.335 3267.590 ;
        RECT 296.765 3037.370 297.095 3037.385 ;
        RECT 296.765 3037.280 310.500 3037.370 ;
        RECT 296.765 3037.070 314.000 3037.280 ;
        RECT 296.765 3037.055 297.095 3037.070 ;
        RECT 310.000 3036.680 314.000 3037.070 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 2829.040 18.330 2829.100 ;
        RECT 296.770 2829.040 297.090 2829.100 ;
        RECT 18.010 2828.900 297.090 2829.040 ;
        RECT 18.010 2828.840 18.330 2828.900 ;
        RECT 296.770 2828.840 297.090 2828.900 ;
      LAYER via ;
        RECT 18.040 2828.840 18.300 2829.100 ;
        RECT 296.800 2828.840 297.060 2829.100 ;
      LAYER met2 ;
        RECT 18.030 2979.915 18.310 2980.285 ;
        RECT 18.100 2829.130 18.240 2979.915 ;
        RECT 18.040 2828.810 18.300 2829.130 ;
        RECT 296.800 2828.810 297.060 2829.130 ;
        RECT 296.860 2823.205 297.000 2828.810 ;
        RECT 296.790 2822.835 297.070 2823.205 ;
      LAYER via2 ;
        RECT 18.030 2979.960 18.310 2980.240 ;
        RECT 296.790 2822.880 297.070 2823.160 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 18.005 2980.250 18.335 2980.265 ;
        RECT -4.800 2979.950 18.335 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 18.005 2979.935 18.335 2979.950 ;
        RECT 296.765 2823.170 297.095 2823.185 ;
        RECT 296.765 2823.080 310.500 2823.170 ;
        RECT 296.765 2822.870 314.000 2823.080 ;
        RECT 296.765 2822.855 297.095 2822.870 ;
        RECT 310.000 2822.480 314.000 2822.870 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2614.840 17.410 2614.900 ;
        RECT 296.770 2614.840 297.090 2614.900 ;
        RECT 17.090 2614.700 297.090 2614.840 ;
        RECT 17.090 2614.640 17.410 2614.700 ;
        RECT 296.770 2614.640 297.090 2614.700 ;
      LAYER via ;
        RECT 17.120 2614.640 17.380 2614.900 ;
        RECT 296.800 2614.640 297.060 2614.900 ;
      LAYER met2 ;
        RECT 17.110 2692.955 17.390 2693.325 ;
        RECT 17.180 2614.930 17.320 2692.955 ;
        RECT 17.120 2614.610 17.380 2614.930 ;
        RECT 296.800 2614.610 297.060 2614.930 ;
        RECT 296.860 2609.005 297.000 2614.610 ;
        RECT 296.790 2608.635 297.070 2609.005 ;
      LAYER via2 ;
        RECT 17.110 2693.000 17.390 2693.280 ;
        RECT 296.790 2608.680 297.070 2608.960 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.085 2693.290 17.415 2693.305 ;
        RECT -4.800 2692.990 17.415 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.085 2692.975 17.415 2692.990 ;
        RECT 296.765 2608.970 297.095 2608.985 ;
        RECT 296.765 2608.880 310.500 2608.970 ;
        RECT 296.765 2608.670 314.000 2608.880 ;
        RECT 296.765 2608.655 297.095 2608.670 ;
        RECT 310.000 2608.280 314.000 2608.670 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 2400.980 18.330 2401.040 ;
        RECT 296.770 2400.980 297.090 2401.040 ;
        RECT 18.010 2400.840 297.090 2400.980 ;
        RECT 18.010 2400.780 18.330 2400.840 ;
        RECT 296.770 2400.780 297.090 2400.840 ;
      LAYER via ;
        RECT 18.040 2400.780 18.300 2401.040 ;
        RECT 296.800 2400.780 297.060 2401.040 ;
      LAYER met2 ;
        RECT 18.030 2405.315 18.310 2405.685 ;
        RECT 18.100 2401.070 18.240 2405.315 ;
        RECT 18.040 2400.750 18.300 2401.070 ;
        RECT 296.800 2400.750 297.060 2401.070 ;
        RECT 296.860 2394.805 297.000 2400.750 ;
        RECT 296.790 2394.435 297.070 2394.805 ;
      LAYER via2 ;
        RECT 18.030 2405.360 18.310 2405.640 ;
        RECT 296.790 2394.480 297.070 2394.760 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 18.005 2405.650 18.335 2405.665 ;
        RECT -4.800 2405.350 18.335 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 18.005 2405.335 18.335 2405.350 ;
        RECT 296.765 2394.770 297.095 2394.785 ;
        RECT 296.765 2394.680 310.500 2394.770 ;
        RECT 296.765 2394.470 314.000 2394.680 ;
        RECT 296.765 2394.455 297.095 2394.470 ;
        RECT 310.000 2394.080 314.000 2394.470 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2125.240 16.490 2125.300 ;
        RECT 299.990 2125.240 300.310 2125.300 ;
        RECT 16.170 2125.100 300.310 2125.240 ;
        RECT 16.170 2125.040 16.490 2125.100 ;
        RECT 299.990 2125.040 300.310 2125.100 ;
      LAYER via ;
        RECT 16.200 2125.040 16.460 2125.300 ;
        RECT 300.020 2125.040 300.280 2125.300 ;
      LAYER met2 ;
        RECT 300.010 2180.235 300.290 2180.605 ;
        RECT 300.080 2125.330 300.220 2180.235 ;
        RECT 16.200 2125.010 16.460 2125.330 ;
        RECT 300.020 2125.010 300.280 2125.330 ;
        RECT 16.260 2118.725 16.400 2125.010 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
      LAYER via2 ;
        RECT 300.010 2180.280 300.290 2180.560 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
      LAYER met3 ;
        RECT 299.985 2180.570 300.315 2180.585 ;
        RECT 299.985 2180.480 310.500 2180.570 ;
        RECT 299.985 2180.270 314.000 2180.480 ;
        RECT 299.985 2180.255 300.315 2180.270 ;
        RECT 310.000 2179.880 314.000 2180.270 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 300.450 1835.220 300.770 1835.280 ;
        RECT 15.710 1835.080 300.770 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 300.450 1835.020 300.770 1835.080 ;
      LAYER via ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 300.480 1835.020 300.740 1835.280 ;
      LAYER met2 ;
        RECT 300.470 1966.035 300.750 1966.405 ;
        RECT 300.540 1835.310 300.680 1966.035 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 300.480 1834.990 300.740 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 300.470 1966.080 300.750 1966.360 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT 300.445 1966.370 300.775 1966.385 ;
        RECT 300.445 1966.280 310.500 1966.370 ;
        RECT 300.445 1966.070 314.000 1966.280 ;
        RECT 300.445 1966.055 300.775 1966.070 ;
        RECT 310.000 1965.680 314.000 1966.070 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 676.160 2618.710 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2618.390 676.020 2901.150 676.160 ;
        RECT 2618.390 675.960 2618.710 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2618.420 675.960 2618.680 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2618.410 782.835 2618.690 783.205 ;
        RECT 2618.480 676.250 2618.620 782.835 ;
        RECT 2618.420 675.930 2618.680 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2618.410 782.880 2618.690 783.160 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2618.385 783.170 2618.715 783.185 ;
        RECT 2609.580 783.080 2618.715 783.170 ;
        RECT 2606.000 782.870 2618.715 783.080 ;
        RECT 2606.000 782.480 2610.000 782.870 ;
        RECT 2618.385 782.855 2618.715 782.870 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 300.450 1545.540 300.770 1545.600 ;
        RECT 16.630 1545.400 300.770 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 300.450 1545.340 300.770 1545.400 ;
      LAYER via ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 300.480 1545.340 300.740 1545.600 ;
      LAYER met2 ;
        RECT 300.470 1751.835 300.750 1752.205 ;
        RECT 300.540 1545.630 300.680 1751.835 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 300.480 1545.310 300.740 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 300.470 1751.880 300.750 1752.160 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 300.445 1752.170 300.775 1752.185 ;
        RECT 300.445 1752.080 310.500 1752.170 ;
        RECT 300.445 1751.870 314.000 1752.080 ;
        RECT 300.445 1751.855 300.775 1751.870 ;
        RECT 310.000 1751.480 314.000 1751.870 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1331.680 16.030 1331.740 ;
        RECT 300.910 1331.680 301.230 1331.740 ;
        RECT 15.710 1331.540 301.230 1331.680 ;
        RECT 15.710 1331.480 16.030 1331.540 ;
        RECT 300.910 1331.480 301.230 1331.540 ;
      LAYER via ;
        RECT 15.740 1331.480 16.000 1331.740 ;
        RECT 300.940 1331.480 301.200 1331.740 ;
      LAYER met2 ;
        RECT 300.930 1536.955 301.210 1537.325 ;
        RECT 301.000 1331.770 301.140 1536.955 ;
        RECT 15.740 1331.450 16.000 1331.770 ;
        RECT 300.940 1331.450 301.200 1331.770 ;
        RECT 15.800 1328.565 15.940 1331.450 ;
        RECT 15.730 1328.195 16.010 1328.565 ;
      LAYER via2 ;
        RECT 300.930 1537.000 301.210 1537.280 ;
        RECT 15.730 1328.240 16.010 1328.520 ;
      LAYER met3 ;
        RECT 300.905 1537.290 301.235 1537.305 ;
        RECT 300.905 1537.200 310.500 1537.290 ;
        RECT 300.905 1536.990 314.000 1537.200 ;
        RECT 300.905 1536.975 301.235 1536.990 ;
        RECT 310.000 1536.600 314.000 1536.990 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 15.705 1328.530 16.035 1328.545 ;
        RECT -4.800 1328.230 16.035 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 15.705 1328.215 16.035 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 301.830 1117.820 302.150 1117.880 ;
        RECT 15.710 1117.680 302.150 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 301.830 1117.620 302.150 1117.680 ;
      LAYER via ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 301.860 1117.620 302.120 1117.880 ;
      LAYER met2 ;
        RECT 301.850 1322.755 302.130 1323.125 ;
        RECT 301.920 1117.910 302.060 1322.755 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 301.860 1117.590 302.120 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 301.850 1322.800 302.130 1323.080 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 301.825 1323.090 302.155 1323.105 ;
        RECT 301.825 1323.000 310.500 1323.090 ;
        RECT 301.825 1322.790 314.000 1323.000 ;
        RECT 301.825 1322.775 302.155 1322.790 ;
        RECT 310.000 1322.400 314.000 1322.790 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 301.370 903.960 301.690 904.020 ;
        RECT 16.170 903.820 301.690 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 301.370 903.760 301.690 903.820 ;
      LAYER via ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 301.400 903.760 301.660 904.020 ;
      LAYER met2 ;
        RECT 301.390 1108.555 301.670 1108.925 ;
        RECT 301.460 904.050 301.600 1108.555 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 301.400 903.730 301.660 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 301.390 1108.600 301.670 1108.880 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 301.365 1108.890 301.695 1108.905 ;
        RECT 301.365 1108.800 310.500 1108.890 ;
        RECT 301.365 1108.590 314.000 1108.800 ;
        RECT 301.365 1108.575 301.695 1108.590 ;
        RECT 310.000 1108.200 314.000 1108.590 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 301.370 682.960 301.690 683.020 ;
        RECT 16.170 682.820 301.690 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 301.370 682.760 301.690 682.820 ;
      LAYER via ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 301.400 682.760 301.660 683.020 ;
      LAYER met2 ;
        RECT 301.390 894.355 301.670 894.725 ;
        RECT 301.460 683.050 301.600 894.355 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 301.400 682.730 301.660 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 301.390 894.400 301.670 894.680 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 301.365 894.690 301.695 894.705 ;
        RECT 301.365 894.600 310.500 894.690 ;
        RECT 301.365 894.390 314.000 894.600 ;
        RECT 301.365 894.375 301.695 894.390 ;
        RECT 310.000 894.000 314.000 894.390 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 300.910 469.100 301.230 469.160 ;
        RECT 17.090 468.960 301.230 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 300.910 468.900 301.230 468.960 ;
      LAYER via ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 300.940 468.900 301.200 469.160 ;
      LAYER met2 ;
        RECT 300.930 680.155 301.210 680.525 ;
        RECT 301.000 469.190 301.140 680.155 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 300.940 468.870 301.200 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 300.930 680.200 301.210 680.480 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 300.905 680.490 301.235 680.505 ;
        RECT 300.905 680.400 310.500 680.490 ;
        RECT 300.905 680.190 314.000 680.400 ;
        RECT 300.905 680.175 301.235 680.190 ;
        RECT 310.000 679.800 314.000 680.190 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 301.370 255.240 301.690 255.300 ;
        RECT 17.090 255.100 301.690 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 301.370 255.040 301.690 255.100 ;
      LAYER via ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 301.400 255.040 301.660 255.300 ;
      LAYER met2 ;
        RECT 301.390 465.955 301.670 466.325 ;
        RECT 301.460 255.330 301.600 465.955 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 301.400 255.010 301.660 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 301.390 466.000 301.670 466.280 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 301.365 466.290 301.695 466.305 ;
        RECT 301.365 466.200 310.500 466.290 ;
        RECT 301.365 465.990 314.000 466.200 ;
        RECT 301.365 465.975 301.695 465.990 ;
        RECT 310.000 465.600 314.000 465.990 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 300.450 41.380 300.770 41.440 ;
        RECT 17.090 41.240 300.770 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 300.450 41.180 300.770 41.240 ;
      LAYER via ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 300.480 41.180 300.740 41.440 ;
      LAYER met2 ;
        RECT 300.470 251.755 300.750 252.125 ;
        RECT 300.540 41.470 300.680 251.755 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 300.480 41.150 300.740 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 300.470 251.800 300.750 252.080 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 300.445 252.090 300.775 252.105 ;
        RECT 300.445 252.000 310.500 252.090 ;
        RECT 300.445 251.790 314.000 252.000 ;
        RECT 300.445 251.775 300.775 251.790 ;
        RECT 310.000 251.400 314.000 251.790 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 910.760 2618.710 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2618.390 910.620 2901.150 910.760 ;
        RECT 2618.390 910.560 2618.710 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2618.420 910.560 2618.680 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2618.410 982.755 2618.690 983.125 ;
        RECT 2618.480 910.850 2618.620 982.755 ;
        RECT 2618.420 910.530 2618.680 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2618.410 982.800 2618.690 983.080 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2618.385 983.090 2618.715 983.105 ;
        RECT 2609.580 983.000 2618.715 983.090 ;
        RECT 2606.000 982.790 2618.715 983.000 ;
        RECT 2606.000 982.400 2610.000 982.790 ;
        RECT 2618.385 982.775 2618.715 982.790 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1145.360 2618.710 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2618.390 1145.220 2901.150 1145.360 ;
        RECT 2618.390 1145.160 2618.710 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2618.420 1145.160 2618.680 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2618.410 1182.675 2618.690 1183.045 ;
        RECT 2618.480 1145.450 2618.620 1182.675 ;
        RECT 2618.420 1145.130 2618.680 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2618.410 1182.720 2618.690 1183.000 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2618.385 1183.010 2618.715 1183.025 ;
        RECT 2609.580 1182.920 2618.715 1183.010 ;
        RECT 2606.000 1182.710 2618.715 1182.920 ;
        RECT 2606.000 1182.320 2610.000 1182.710 ;
        RECT 2618.385 1182.695 2618.715 1182.710 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1379.960 2621.930 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2621.610 1379.820 2901.150 1379.960 ;
        RECT 2621.610 1379.760 2621.930 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 2621.640 1379.760 2621.900 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 2621.630 1382.595 2621.910 1382.965 ;
        RECT 2621.700 1380.050 2621.840 1382.595 ;
        RECT 2621.640 1379.730 2621.900 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2621.630 1382.640 2621.910 1382.920 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2621.605 1382.930 2621.935 1382.945 ;
        RECT 2609.580 1382.840 2621.935 1382.930 ;
        RECT 2606.000 1382.630 2621.935 1382.840 ;
        RECT 2606.000 1382.240 2610.000 1382.630 ;
        RECT 2621.605 1382.615 2621.935 1382.630 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2617.470 1608.100 2617.790 1608.160 ;
        RECT 2900.830 1608.100 2901.150 1608.160 ;
        RECT 2617.470 1607.960 2901.150 1608.100 ;
        RECT 2617.470 1607.900 2617.790 1607.960 ;
        RECT 2900.830 1607.900 2901.150 1607.960 ;
      LAYER via ;
        RECT 2617.500 1607.900 2617.760 1608.160 ;
        RECT 2900.860 1607.900 2901.120 1608.160 ;
      LAYER met2 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
        RECT 2900.920 1608.190 2901.060 1613.115 ;
        RECT 2617.500 1607.870 2617.760 1608.190 ;
        RECT 2900.860 1607.870 2901.120 1608.190 ;
        RECT 2617.560 1582.885 2617.700 1607.870 ;
        RECT 2617.490 1582.515 2617.770 1582.885 ;
      LAYER via2 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
        RECT 2617.490 1582.560 2617.770 1582.840 ;
      LAYER met3 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 2617.465 1582.850 2617.795 1582.865 ;
        RECT 2609.580 1582.760 2617.795 1582.850 ;
        RECT 2606.000 1582.550 2617.795 1582.760 ;
        RECT 2606.000 1582.160 2610.000 1582.550 ;
        RECT 2617.465 1582.535 2617.795 1582.550 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1842.700 2618.710 1842.760 ;
        RECT 2900.830 1842.700 2901.150 1842.760 ;
        RECT 2618.390 1842.560 2901.150 1842.700 ;
        RECT 2618.390 1842.500 2618.710 1842.560 ;
        RECT 2900.830 1842.500 2901.150 1842.560 ;
      LAYER via ;
        RECT 2618.420 1842.500 2618.680 1842.760 ;
        RECT 2900.860 1842.500 2901.120 1842.760 ;
      LAYER met2 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
        RECT 2900.920 1842.790 2901.060 1847.715 ;
        RECT 2618.420 1842.470 2618.680 1842.790 ;
        RECT 2900.860 1842.470 2901.120 1842.790 ;
        RECT 2618.480 1783.485 2618.620 1842.470 ;
        RECT 2618.410 1783.115 2618.690 1783.485 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
        RECT 2618.410 1783.160 2618.690 1783.440 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2618.385 1783.450 2618.715 1783.465 ;
        RECT 2609.580 1783.360 2618.715 1783.450 ;
        RECT 2606.000 1783.150 2618.715 1783.360 ;
        RECT 2606.000 1782.760 2610.000 1783.150 ;
        RECT 2618.385 1783.135 2618.715 1783.150 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2077.300 2619.170 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 2618.850 2077.160 2901.150 2077.300 ;
        RECT 2618.850 2077.100 2619.170 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
      LAYER via ;
        RECT 2618.880 2077.100 2619.140 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 2618.880 2077.070 2619.140 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 2618.940 1983.405 2619.080 2077.070 ;
        RECT 2618.870 1983.035 2619.150 1983.405 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
        RECT 2618.870 1983.080 2619.150 1983.360 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2618.845 1983.370 2619.175 1983.385 ;
        RECT 2609.580 1983.280 2619.175 1983.370 ;
        RECT 2606.000 1983.070 2619.175 1983.280 ;
        RECT 2606.000 1982.680 2610.000 1983.070 ;
        RECT 2618.845 1983.055 2619.175 1983.070 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.770 2311.900 2620.090 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2619.770 2311.760 2901.150 2311.900 ;
        RECT 2619.770 2311.700 2620.090 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
      LAYER via ;
        RECT 2619.800 2311.700 2620.060 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2619.800 2311.670 2620.060 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2619.860 2183.325 2620.000 2311.670 ;
        RECT 2619.790 2182.955 2620.070 2183.325 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2619.790 2183.000 2620.070 2183.280 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2619.765 2183.290 2620.095 2183.305 ;
        RECT 2609.580 2183.200 2620.095 2183.290 ;
        RECT 2606.000 2182.990 2620.095 2183.200 ;
        RECT 2606.000 2182.600 2610.000 2182.990 ;
        RECT 2619.765 2182.975 2620.095 2182.990 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.310 151.540 2619.630 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2619.310 151.400 2901.150 151.540 ;
        RECT 2619.310 151.340 2619.630 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2619.340 151.340 2619.600 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2619.330 316.355 2619.610 316.725 ;
        RECT 2619.400 151.630 2619.540 316.355 ;
        RECT 2619.340 151.310 2619.600 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2619.330 316.400 2619.610 316.680 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2619.305 316.690 2619.635 316.705 ;
        RECT 2609.580 316.600 2619.635 316.690 ;
        RECT 2606.000 316.390 2619.635 316.600 ;
        RECT 2606.000 316.000 2610.000 316.390 ;
        RECT 2619.305 316.375 2619.635 316.390 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2491.080 2618.710 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 2618.390 2490.940 2901.150 2491.080 ;
        RECT 2618.390 2490.880 2618.710 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
      LAYER via ;
        RECT 2618.420 2490.880 2618.680 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 2618.420 2490.850 2618.680 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 2618.480 2316.605 2618.620 2490.850 ;
        RECT 2618.410 2316.235 2618.690 2316.605 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 2618.410 2316.280 2618.690 2316.560 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2618.385 2316.570 2618.715 2316.585 ;
        RECT 2609.580 2316.480 2618.715 2316.570 ;
        RECT 2606.000 2316.270 2618.715 2316.480 ;
        RECT 2606.000 2315.880 2610.000 2316.270 ;
        RECT 2618.385 2316.255 2618.715 2316.270 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2725.680 2619.170 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2618.850 2725.540 2901.150 2725.680 ;
        RECT 2618.850 2725.480 2619.170 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 2618.880 2725.480 2619.140 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2618.880 2725.450 2619.140 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 2618.940 2516.525 2619.080 2725.450 ;
        RECT 2618.870 2516.155 2619.150 2516.525 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 2618.870 2516.200 2619.150 2516.480 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2618.845 2516.490 2619.175 2516.505 ;
        RECT 2609.580 2516.400 2619.175 2516.490 ;
        RECT 2606.000 2516.190 2619.175 2516.400 ;
        RECT 2606.000 2515.800 2610.000 2516.190 ;
        RECT 2618.845 2516.175 2619.175 2516.190 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2960.280 2618.710 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 2618.390 2960.140 2901.150 2960.280 ;
        RECT 2618.390 2960.080 2618.710 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 2618.420 2960.080 2618.680 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 2618.420 2960.050 2618.680 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 2618.480 2716.445 2618.620 2960.050 ;
        RECT 2618.410 2716.075 2618.690 2716.445 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 2618.410 2716.120 2618.690 2716.400 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2618.385 2716.410 2618.715 2716.425 ;
        RECT 2609.580 2716.320 2618.715 2716.410 ;
        RECT 2606.000 2716.110 2618.715 2716.320 ;
        RECT 2606.000 2715.720 2610.000 2716.110 ;
        RECT 2618.385 2716.095 2618.715 2716.110 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.310 3194.880 2619.630 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2619.310 3194.740 2901.150 3194.880 ;
        RECT 2619.310 3194.680 2619.630 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 2619.340 3194.680 2619.600 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2619.340 3194.650 2619.600 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 2619.400 2916.365 2619.540 3194.650 ;
        RECT 2619.330 2915.995 2619.610 2916.365 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 2619.330 2916.040 2619.610 2916.320 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2619.305 2916.330 2619.635 2916.345 ;
        RECT 2609.580 2916.240 2619.635 2916.330 ;
        RECT 2606.000 2916.030 2619.635 2916.240 ;
        RECT 2606.000 2915.640 2610.000 2916.030 ;
        RECT 2619.305 2916.015 2619.635 2916.030 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 3429.480 2618.710 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2618.390 3429.340 2901.150 3429.480 ;
        RECT 2618.390 3429.280 2618.710 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 2618.420 3429.280 2618.680 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 2618.420 3429.250 2618.680 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 2618.480 3116.285 2618.620 3429.250 ;
        RECT 2618.410 3115.915 2618.690 3116.285 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 2618.410 3115.960 2618.690 3116.240 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2618.385 3116.250 2618.715 3116.265 ;
        RECT 2609.580 3116.160 2618.715 3116.250 ;
        RECT 2606.000 3115.950 2618.715 3116.160 ;
        RECT 2606.000 3115.560 2610.000 3115.950 ;
        RECT 2618.385 3115.935 2618.715 3115.950 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2483.610 3501.900 2483.930 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 2483.610 3501.760 2717.610 3501.900 ;
        RECT 2483.610 3501.700 2483.930 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 2483.640 3501.700 2483.900 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 2483.640 3501.670 2483.900 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 2481.750 3215.450 2482.030 3216.000 ;
        RECT 2483.700 3215.450 2483.840 3501.670 ;
        RECT 2481.750 3215.310 2483.840 3215.450 ;
        RECT 2481.750 3212.000 2482.030 3215.310 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2228.310 3501.900 2228.630 3501.960 ;
        RECT 2392.530 3501.900 2392.850 3501.960 ;
        RECT 2228.310 3501.760 2392.850 3501.900 ;
        RECT 2228.310 3501.700 2228.630 3501.760 ;
        RECT 2392.530 3501.700 2392.850 3501.760 ;
      LAYER via ;
        RECT 2228.340 3501.700 2228.600 3501.960 ;
        RECT 2392.560 3501.700 2392.820 3501.960 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.990 2392.760 3517.600 ;
        RECT 2228.340 3501.670 2228.600 3501.990 ;
        RECT 2392.560 3501.670 2392.820 3501.990 ;
        RECT 2226.450 3215.450 2226.730 3216.000 ;
        RECT 2228.400 3215.450 2228.540 3501.670 ;
        RECT 2226.450 3215.310 2228.540 3215.450 ;
        RECT 2226.450 3212.000 2226.730 3215.310 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 3502.240 1973.330 3502.300 ;
        RECT 2068.230 3502.240 2068.550 3502.300 ;
        RECT 1973.010 3502.100 2068.550 3502.240 ;
        RECT 1973.010 3502.040 1973.330 3502.100 ;
        RECT 2068.230 3502.040 2068.550 3502.100 ;
      LAYER via ;
        RECT 1973.040 3502.040 1973.300 3502.300 ;
        RECT 2068.260 3502.040 2068.520 3502.300 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3502.330 2068.460 3517.600 ;
        RECT 1973.040 3502.010 1973.300 3502.330 ;
        RECT 2068.260 3502.010 2068.520 3502.330 ;
        RECT 1970.690 3214.770 1970.970 3216.000 ;
        RECT 1973.100 3214.770 1973.240 3502.010 ;
        RECT 1970.690 3214.630 1973.240 3214.770 ;
        RECT 1970.690 3212.000 1970.970 3214.630 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1721.390 3501.560 1721.710 3501.620 ;
        RECT 1743.930 3501.560 1744.250 3501.620 ;
        RECT 1721.390 3501.420 1744.250 3501.560 ;
        RECT 1721.390 3501.360 1721.710 3501.420 ;
        RECT 1743.930 3501.360 1744.250 3501.420 ;
        RECT 1714.950 3229.220 1715.270 3229.280 ;
        RECT 1721.390 3229.220 1721.710 3229.280 ;
        RECT 1714.950 3229.080 1721.710 3229.220 ;
        RECT 1714.950 3229.020 1715.270 3229.080 ;
        RECT 1721.390 3229.020 1721.710 3229.080 ;
      LAYER via ;
        RECT 1721.420 3501.360 1721.680 3501.620 ;
        RECT 1743.960 3501.360 1744.220 3501.620 ;
        RECT 1714.980 3229.020 1715.240 3229.280 ;
        RECT 1721.420 3229.020 1721.680 3229.280 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3501.650 1744.160 3517.600 ;
        RECT 1721.420 3501.330 1721.680 3501.650 ;
        RECT 1743.960 3501.330 1744.220 3501.650 ;
        RECT 1721.480 3229.310 1721.620 3501.330 ;
        RECT 1714.980 3228.990 1715.240 3229.310 ;
        RECT 1721.420 3228.990 1721.680 3229.310 ;
        RECT 1715.040 3216.000 1715.180 3228.990 ;
        RECT 1714.930 3212.000 1715.210 3216.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1420.165 3381.045 1420.335 3429.155 ;
      LAYER mcon ;
        RECT 1420.165 3428.985 1420.335 3429.155 ;
      LAYER met1 ;
        RECT 1419.170 3477.760 1419.490 3477.820 ;
        RECT 1419.630 3477.760 1419.950 3477.820 ;
        RECT 1419.170 3477.620 1419.950 3477.760 ;
        RECT 1419.170 3477.560 1419.490 3477.620 ;
        RECT 1419.630 3477.560 1419.950 3477.620 ;
        RECT 1419.630 3443.080 1419.950 3443.140 ;
        RECT 1420.550 3443.080 1420.870 3443.140 ;
        RECT 1419.630 3442.940 1420.870 3443.080 ;
        RECT 1419.630 3442.880 1419.950 3442.940 ;
        RECT 1420.550 3442.880 1420.870 3442.940 ;
        RECT 1420.105 3429.140 1420.395 3429.185 ;
        RECT 1420.550 3429.140 1420.870 3429.200 ;
        RECT 1420.105 3429.000 1420.870 3429.140 ;
        RECT 1420.105 3428.955 1420.395 3429.000 ;
        RECT 1420.550 3428.940 1420.870 3429.000 ;
        RECT 1420.090 3381.200 1420.410 3381.260 ;
        RECT 1419.895 3381.060 1420.410 3381.200 ;
        RECT 1420.090 3381.000 1420.410 3381.060 ;
        RECT 1420.090 3367.600 1420.410 3367.660 ;
        RECT 1421.010 3367.600 1421.330 3367.660 ;
        RECT 1420.090 3367.460 1421.330 3367.600 ;
        RECT 1420.090 3367.400 1420.410 3367.460 ;
        RECT 1421.010 3367.400 1421.330 3367.460 ;
        RECT 1420.090 3270.700 1420.410 3270.760 ;
        RECT 1421.010 3270.700 1421.330 3270.760 ;
        RECT 1420.090 3270.560 1421.330 3270.700 ;
        RECT 1420.090 3270.500 1420.410 3270.560 ;
        RECT 1421.010 3270.500 1421.330 3270.560 ;
        RECT 1421.010 3225.820 1421.330 3225.880 ;
        RECT 1459.650 3225.820 1459.970 3225.880 ;
        RECT 1421.010 3225.680 1459.970 3225.820 ;
        RECT 1421.010 3225.620 1421.330 3225.680 ;
        RECT 1459.650 3225.620 1459.970 3225.680 ;
      LAYER via ;
        RECT 1419.200 3477.560 1419.460 3477.820 ;
        RECT 1419.660 3477.560 1419.920 3477.820 ;
        RECT 1419.660 3442.880 1419.920 3443.140 ;
        RECT 1420.580 3442.880 1420.840 3443.140 ;
        RECT 1420.580 3428.940 1420.840 3429.200 ;
        RECT 1420.120 3381.000 1420.380 3381.260 ;
        RECT 1420.120 3367.400 1420.380 3367.660 ;
        RECT 1421.040 3367.400 1421.300 3367.660 ;
        RECT 1420.120 3270.500 1420.380 3270.760 ;
        RECT 1421.040 3270.500 1421.300 3270.760 ;
        RECT 1421.040 3225.620 1421.300 3225.880 ;
        RECT 1459.680 3225.620 1459.940 3225.880 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3477.850 1419.400 3517.600 ;
        RECT 1419.200 3477.530 1419.460 3477.850 ;
        RECT 1419.660 3477.530 1419.920 3477.850 ;
        RECT 1419.720 3443.170 1419.860 3477.530 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3270.790 1420.320 3318.670 ;
        RECT 1420.120 3270.470 1420.380 3270.790 ;
        RECT 1421.040 3270.470 1421.300 3270.790 ;
        RECT 1421.100 3225.910 1421.240 3270.470 ;
        RECT 1421.040 3225.590 1421.300 3225.910 ;
        RECT 1459.680 3225.590 1459.940 3225.910 ;
        RECT 1459.740 3216.000 1459.880 3225.590 ;
        RECT 1459.630 3212.000 1459.910 3216.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 386.140 2619.170 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2618.850 386.000 2901.150 386.140 ;
        RECT 2618.850 385.940 2619.170 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2618.880 385.940 2619.140 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2618.870 516.275 2619.150 516.645 ;
        RECT 2618.940 386.230 2619.080 516.275 ;
        RECT 2618.880 385.910 2619.140 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2618.870 516.320 2619.150 516.600 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 2618.845 516.610 2619.175 516.625 ;
        RECT 2609.580 516.520 2619.175 516.610 ;
        RECT 2606.000 516.310 2619.175 516.520 ;
        RECT 2606.000 515.920 2610.000 516.310 ;
        RECT 2618.845 516.295 2619.175 516.310 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1094.945 3332.765 1095.115 3380.875 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1094.945 3380.705 1095.115 3380.875 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1094.870 3380.860 1095.190 3380.920 ;
        RECT 1094.675 3380.720 1095.190 3380.860 ;
        RECT 1094.870 3380.660 1095.190 3380.720 ;
        RECT 1094.885 3332.920 1095.175 3332.965 ;
        RECT 1095.330 3332.920 1095.650 3332.980 ;
        RECT 1094.885 3332.780 1095.650 3332.920 ;
        RECT 1094.885 3332.735 1095.175 3332.780 ;
        RECT 1095.330 3332.720 1095.650 3332.780 ;
        RECT 1096.710 3226.160 1097.030 3226.220 ;
        RECT 1203.890 3226.160 1204.210 3226.220 ;
        RECT 1096.710 3226.020 1204.210 3226.160 ;
        RECT 1096.710 3225.960 1097.030 3226.020 ;
        RECT 1203.890 3225.960 1204.210 3226.020 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1094.900 3380.660 1095.160 3380.920 ;
        RECT 1095.360 3332.720 1095.620 3332.980 ;
        RECT 1096.740 3225.960 1097.000 3226.220 ;
        RECT 1203.920 3225.960 1204.180 3226.220 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3394.970 1095.560 3429.250 ;
        RECT 1094.960 3394.830 1095.560 3394.970 ;
        RECT 1094.960 3380.950 1095.100 3394.830 ;
        RECT 1094.900 3380.630 1095.160 3380.950 ;
        RECT 1095.360 3332.690 1095.620 3333.010 ;
        RECT 1095.420 3298.410 1095.560 3332.690 ;
        RECT 1095.420 3298.270 1096.480 3298.410 ;
        RECT 1096.340 3250.130 1096.480 3298.270 ;
        RECT 1096.340 3249.990 1096.940 3250.130 ;
        RECT 1096.800 3226.250 1096.940 3249.990 ;
        RECT 1096.740 3225.930 1097.000 3226.250 ;
        RECT 1203.920 3225.930 1204.180 3226.250 ;
        RECT 1203.980 3216.000 1204.120 3225.930 ;
        RECT 1203.870 3212.000 1204.150 3216.000 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 772.410 3225.820 772.730 3225.880 ;
        RECT 948.590 3225.820 948.910 3225.880 ;
        RECT 772.410 3225.680 948.910 3225.820 ;
        RECT 772.410 3225.620 772.730 3225.680 ;
        RECT 948.590 3225.620 948.910 3225.680 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 772.440 3225.620 772.700 3225.880 ;
        RECT 948.620 3225.620 948.880 3225.880 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3225.910 772.640 3270.470 ;
        RECT 772.440 3225.590 772.700 3225.910 ;
        RECT 948.620 3225.590 948.880 3225.910 ;
        RECT 948.680 3216.000 948.820 3225.590 ;
        RECT 948.570 3212.000 948.850 3216.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 3225.820 448.430 3225.880 ;
        RECT 692.830 3225.820 693.150 3225.880 ;
        RECT 448.110 3225.680 693.150 3225.820 ;
        RECT 448.110 3225.620 448.430 3225.680 ;
        RECT 692.830 3225.620 693.150 3225.680 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 3225.620 448.400 3225.880 ;
        RECT 692.860 3225.620 693.120 3225.880 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 3225.910 448.340 3498.270 ;
        RECT 448.140 3225.590 448.400 3225.910 ;
        RECT 692.860 3225.590 693.120 3225.910 ;
        RECT 692.920 3216.000 693.060 3225.590 ;
        RECT 692.810 3212.000 693.090 3216.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 3225.820 124.130 3225.880 ;
        RECT 437.530 3225.820 437.850 3225.880 ;
        RECT 123.810 3225.680 437.850 3225.820 ;
        RECT 123.810 3225.620 124.130 3225.680 ;
        RECT 437.530 3225.620 437.850 3225.680 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 3225.620 124.100 3225.880 ;
        RECT 437.560 3225.620 437.820 3225.880 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 3225.910 124.040 3498.270 ;
        RECT 123.840 3225.590 124.100 3225.910 ;
        RECT 437.560 3225.590 437.820 3225.910 ;
        RECT 437.620 3216.000 437.760 3225.590 ;
        RECT 437.510 3212.000 437.790 3216.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 3111.920 17.870 3111.980 ;
        RECT 296.770 3111.920 297.090 3111.980 ;
        RECT 17.550 3111.780 297.090 3111.920 ;
        RECT 17.550 3111.720 17.870 3111.780 ;
        RECT 296.770 3111.720 297.090 3111.780 ;
      LAYER via ;
        RECT 17.580 3111.720 17.840 3111.980 ;
        RECT 296.800 3111.720 297.060 3111.980 ;
      LAYER met2 ;
        RECT 17.570 3339.635 17.850 3340.005 ;
        RECT 17.640 3112.010 17.780 3339.635 ;
        RECT 17.580 3111.690 17.840 3112.010 ;
        RECT 296.800 3111.690 297.060 3112.010 ;
        RECT 296.860 3108.805 297.000 3111.690 ;
        RECT 296.790 3108.435 297.070 3108.805 ;
      LAYER via2 ;
        RECT 17.570 3339.680 17.850 3339.960 ;
        RECT 296.790 3108.480 297.070 3108.760 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.545 3339.970 17.875 3339.985 ;
        RECT -4.800 3339.670 17.875 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.545 3339.655 17.875 3339.670 ;
        RECT 296.765 3108.770 297.095 3108.785 ;
        RECT 296.765 3108.680 310.500 3108.770 ;
        RECT 296.765 3108.470 314.000 3108.680 ;
        RECT 296.765 3108.455 297.095 3108.470 ;
        RECT 310.000 3108.080 314.000 3108.470 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2898.060 17.870 2898.120 ;
        RECT 296.770 2898.060 297.090 2898.120 ;
        RECT 17.550 2897.920 297.090 2898.060 ;
        RECT 17.550 2897.860 17.870 2897.920 ;
        RECT 296.770 2897.860 297.090 2897.920 ;
      LAYER via ;
        RECT 17.580 2897.860 17.840 2898.120 ;
        RECT 296.800 2897.860 297.060 2898.120 ;
      LAYER met2 ;
        RECT 17.570 3051.995 17.850 3052.365 ;
        RECT 17.640 2898.150 17.780 3051.995 ;
        RECT 17.580 2897.830 17.840 2898.150 ;
        RECT 296.800 2897.830 297.060 2898.150 ;
        RECT 296.860 2894.605 297.000 2897.830 ;
        RECT 296.790 2894.235 297.070 2894.605 ;
      LAYER via2 ;
        RECT 17.570 3052.040 17.850 3052.320 ;
        RECT 296.790 2894.280 297.070 2894.560 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.545 3052.330 17.875 3052.345 ;
        RECT -4.800 3052.030 17.875 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.545 3052.015 17.875 3052.030 ;
        RECT 296.765 2894.570 297.095 2894.585 ;
        RECT 296.765 2894.480 310.500 2894.570 ;
        RECT 296.765 2894.270 314.000 2894.480 ;
        RECT 296.765 2894.255 297.095 2894.270 ;
        RECT 310.000 2893.880 314.000 2894.270 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2683.860 17.870 2683.920 ;
        RECT 296.770 2683.860 297.090 2683.920 ;
        RECT 17.550 2683.720 297.090 2683.860 ;
        RECT 17.550 2683.660 17.870 2683.720 ;
        RECT 296.770 2683.660 297.090 2683.720 ;
      LAYER via ;
        RECT 17.580 2683.660 17.840 2683.920 ;
        RECT 296.800 2683.660 297.060 2683.920 ;
      LAYER met2 ;
        RECT 17.570 2765.035 17.850 2765.405 ;
        RECT 17.640 2683.950 17.780 2765.035 ;
        RECT 17.580 2683.630 17.840 2683.950 ;
        RECT 296.800 2683.630 297.060 2683.950 ;
        RECT 296.860 2680.405 297.000 2683.630 ;
        RECT 296.790 2680.035 297.070 2680.405 ;
      LAYER via2 ;
        RECT 17.570 2765.080 17.850 2765.360 ;
        RECT 296.790 2680.080 297.070 2680.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 17.545 2765.370 17.875 2765.385 ;
        RECT -4.800 2765.070 17.875 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 17.545 2765.055 17.875 2765.070 ;
        RECT 296.765 2680.370 297.095 2680.385 ;
        RECT 296.765 2680.280 310.500 2680.370 ;
        RECT 296.765 2680.070 314.000 2680.280 ;
        RECT 296.765 2680.055 297.095 2680.070 ;
        RECT 310.000 2679.680 314.000 2680.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2470.000 16.950 2470.060 ;
        RECT 296.770 2470.000 297.090 2470.060 ;
        RECT 16.630 2469.860 297.090 2470.000 ;
        RECT 16.630 2469.800 16.950 2469.860 ;
        RECT 296.770 2469.800 297.090 2469.860 ;
      LAYER via ;
        RECT 16.660 2469.800 16.920 2470.060 ;
        RECT 296.800 2469.800 297.060 2470.060 ;
      LAYER met2 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 16.720 2470.090 16.860 2477.395 ;
        RECT 16.660 2469.770 16.920 2470.090 ;
        RECT 296.800 2469.770 297.060 2470.090 ;
        RECT 296.860 2466.205 297.000 2469.770 ;
        RECT 296.790 2465.835 297.070 2466.205 ;
      LAYER via2 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
        RECT 296.790 2465.880 297.070 2466.160 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
        RECT 296.765 2466.170 297.095 2466.185 ;
        RECT 296.765 2466.080 310.500 2466.170 ;
        RECT 296.765 2465.870 314.000 2466.080 ;
        RECT 296.765 2465.855 297.095 2465.870 ;
        RECT 310.000 2465.480 314.000 2465.870 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2194.260 16.030 2194.320 ;
        RECT 299.990 2194.260 300.310 2194.320 ;
        RECT 15.710 2194.120 300.310 2194.260 ;
        RECT 15.710 2194.060 16.030 2194.120 ;
        RECT 299.990 2194.060 300.310 2194.120 ;
      LAYER via ;
        RECT 15.740 2194.060 16.000 2194.320 ;
        RECT 300.020 2194.060 300.280 2194.320 ;
      LAYER met2 ;
        RECT 300.010 2251.635 300.290 2252.005 ;
        RECT 300.080 2194.350 300.220 2251.635 ;
        RECT 15.740 2194.030 16.000 2194.350 ;
        RECT 300.020 2194.030 300.280 2194.350 ;
        RECT 15.800 2190.125 15.940 2194.030 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
      LAYER via2 ;
        RECT 300.010 2251.680 300.290 2251.960 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
      LAYER met3 ;
        RECT 299.985 2251.970 300.315 2251.985 ;
        RECT 299.985 2251.880 310.500 2251.970 ;
        RECT 299.985 2251.670 314.000 2251.880 ;
        RECT 299.985 2251.655 300.315 2251.670 ;
        RECT 310.000 2251.280 314.000 2251.670 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.800 2189.790 16.035 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1904.240 16.490 1904.300 ;
        RECT 299.990 1904.240 300.310 1904.300 ;
        RECT 16.170 1904.100 300.310 1904.240 ;
        RECT 16.170 1904.040 16.490 1904.100 ;
        RECT 299.990 1904.040 300.310 1904.100 ;
      LAYER via ;
        RECT 16.200 1904.040 16.460 1904.300 ;
        RECT 300.020 1904.040 300.280 1904.300 ;
      LAYER met2 ;
        RECT 300.010 2037.435 300.290 2037.805 ;
        RECT 300.080 1904.330 300.220 2037.435 ;
        RECT 16.200 1904.010 16.460 1904.330 ;
        RECT 300.020 1904.010 300.280 1904.330 ;
        RECT 16.260 1903.165 16.400 1904.010 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
      LAYER via2 ;
        RECT 300.010 2037.480 300.290 2037.760 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT 299.985 2037.770 300.315 2037.785 ;
        RECT 299.985 2037.680 310.500 2037.770 ;
        RECT 299.985 2037.470 314.000 2037.680 ;
        RECT 299.985 2037.455 300.315 2037.470 ;
        RECT 310.000 2037.080 314.000 2037.470 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 620.740 2619.170 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2618.850 620.600 2901.150 620.740 ;
        RECT 2618.850 620.540 2619.170 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2618.880 620.540 2619.140 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2618.870 716.195 2619.150 716.565 ;
        RECT 2618.940 620.830 2619.080 716.195 ;
        RECT 2618.880 620.510 2619.140 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2618.870 716.240 2619.150 716.520 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2618.845 716.530 2619.175 716.545 ;
        RECT 2609.580 716.440 2619.175 716.530 ;
        RECT 2606.000 716.230 2619.175 716.440 ;
        RECT 2606.000 715.840 2610.000 716.230 ;
        RECT 2618.845 716.215 2619.175 716.230 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 300.910 1621.360 301.230 1621.420 ;
        RECT 16.170 1621.220 301.230 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 300.910 1621.160 301.230 1621.220 ;
      LAYER via ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 300.940 1621.160 301.200 1621.420 ;
      LAYER met2 ;
        RECT 300.930 1823.235 301.210 1823.605 ;
        RECT 301.000 1621.450 301.140 1823.235 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 300.940 1621.130 301.200 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 300.930 1823.280 301.210 1823.560 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT 300.905 1823.570 301.235 1823.585 ;
        RECT 300.905 1823.480 310.500 1823.570 ;
        RECT 300.905 1823.270 314.000 1823.480 ;
        RECT 300.905 1823.255 301.235 1823.270 ;
        RECT 310.000 1822.880 314.000 1823.270 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 299.990 1400.700 300.310 1400.760 ;
        RECT 17.090 1400.560 300.310 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 299.990 1400.500 300.310 1400.560 ;
      LAYER via ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 300.020 1400.500 300.280 1400.760 ;
      LAYER met2 ;
        RECT 300.010 1608.355 300.290 1608.725 ;
        RECT 300.080 1400.790 300.220 1608.355 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 300.020 1400.470 300.280 1400.790 ;
      LAYER via2 ;
        RECT 300.010 1608.400 300.290 1608.680 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 299.985 1608.690 300.315 1608.705 ;
        RECT 299.985 1608.600 310.500 1608.690 ;
        RECT 299.985 1608.390 314.000 1608.600 ;
        RECT 299.985 1608.375 300.315 1608.390 ;
        RECT 310.000 1608.000 314.000 1608.390 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 300.450 1186.840 300.770 1186.900 ;
        RECT 17.090 1186.700 300.770 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 300.450 1186.640 300.770 1186.700 ;
      LAYER via ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 300.480 1186.640 300.740 1186.900 ;
      LAYER met2 ;
        RECT 300.470 1394.155 300.750 1394.525 ;
        RECT 300.540 1186.930 300.680 1394.155 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 300.480 1186.610 300.740 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 300.470 1394.200 300.750 1394.480 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT 300.445 1394.490 300.775 1394.505 ;
        RECT 300.445 1394.400 310.500 1394.490 ;
        RECT 300.445 1394.190 314.000 1394.400 ;
        RECT 300.445 1394.175 300.775 1394.190 ;
        RECT 310.000 1393.800 314.000 1394.190 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 300.910 972.640 301.230 972.700 ;
        RECT 15.710 972.500 301.230 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 300.910 972.440 301.230 972.500 ;
      LAYER via ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 300.940 972.440 301.200 972.700 ;
      LAYER met2 ;
        RECT 300.930 1179.955 301.210 1180.325 ;
        RECT 301.000 972.730 301.140 1179.955 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 300.940 972.410 301.200 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 300.930 1180.000 301.210 1180.280 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT 300.905 1180.290 301.235 1180.305 ;
        RECT 300.905 1180.200 310.500 1180.290 ;
        RECT 300.905 1179.990 314.000 1180.200 ;
        RECT 300.905 1179.975 301.235 1179.990 ;
        RECT 310.000 1179.600 314.000 1179.990 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 300.910 758.780 301.230 758.840 ;
        RECT 15.710 758.640 301.230 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 300.910 758.580 301.230 758.640 ;
      LAYER via ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 300.940 758.580 301.200 758.840 ;
      LAYER met2 ;
        RECT 300.930 965.755 301.210 966.125 ;
        RECT 301.000 758.870 301.140 965.755 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 300.940 758.550 301.200 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 300.930 965.800 301.210 966.080 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 300.905 966.090 301.235 966.105 ;
        RECT 300.905 966.000 310.500 966.090 ;
        RECT 300.905 965.790 314.000 966.000 ;
        RECT 300.905 965.775 301.235 965.790 ;
        RECT 310.000 965.400 314.000 965.790 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 301.830 544.920 302.150 544.980 ;
        RECT 16.170 544.780 302.150 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 301.830 544.720 302.150 544.780 ;
      LAYER via ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 301.860 544.720 302.120 544.980 ;
      LAYER met2 ;
        RECT 301.850 751.555 302.130 751.925 ;
        RECT 301.920 545.010 302.060 751.555 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 301.860 544.690 302.120 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 301.850 751.600 302.130 751.880 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 301.825 751.890 302.155 751.905 ;
        RECT 301.825 751.800 310.500 751.890 ;
        RECT 301.825 751.590 314.000 751.800 ;
        RECT 301.825 751.575 302.155 751.590 ;
        RECT 310.000 751.200 314.000 751.590 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 301.830 324.260 302.150 324.320 ;
        RECT 16.630 324.120 302.150 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 301.830 324.060 302.150 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 301.860 324.060 302.120 324.320 ;
      LAYER met2 ;
        RECT 301.850 537.355 302.130 537.725 ;
        RECT 301.920 324.350 302.060 537.355 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 301.860 324.030 302.120 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 301.850 537.400 302.130 537.680 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 301.825 537.690 302.155 537.705 ;
        RECT 301.825 537.600 310.500 537.690 ;
        RECT 301.825 537.390 314.000 537.600 ;
        RECT 301.825 537.375 302.155 537.390 ;
        RECT 310.000 537.000 314.000 537.390 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 300.910 110.400 301.230 110.460 ;
        RECT 15.710 110.260 301.230 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 300.910 110.200 301.230 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 300.940 110.200 301.200 110.460 ;
      LAYER met2 ;
        RECT 300.930 323.155 301.210 323.525 ;
        RECT 301.000 110.490 301.140 323.155 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 300.940 110.170 301.200 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 300.930 323.200 301.210 323.480 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 300.905 323.490 301.235 323.505 ;
        RECT 300.905 323.400 310.500 323.490 ;
        RECT 300.905 323.190 314.000 323.400 ;
        RECT 300.905 323.175 301.235 323.190 ;
        RECT 310.000 322.800 314.000 323.190 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 855.340 2619.170 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2618.850 855.200 2901.150 855.340 ;
        RECT 2618.850 855.140 2619.170 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2618.880 855.140 2619.140 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2618.870 916.115 2619.150 916.485 ;
        RECT 2618.940 855.430 2619.080 916.115 ;
        RECT 2618.880 855.110 2619.140 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2618.870 916.160 2619.150 916.440 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2618.845 916.450 2619.175 916.465 ;
        RECT 2609.580 916.360 2619.175 916.450 ;
        RECT 2606.000 916.150 2619.175 916.360 ;
        RECT 2606.000 915.760 2610.000 916.150 ;
        RECT 2618.845 916.135 2619.175 916.150 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1089.940 2618.710 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2618.390 1089.800 2901.150 1089.940 ;
        RECT 2618.390 1089.740 2618.710 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2618.420 1089.740 2618.680 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2618.410 1116.035 2618.690 1116.405 ;
        RECT 2618.480 1090.030 2618.620 1116.035 ;
        RECT 2618.420 1089.710 2618.680 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2618.410 1116.080 2618.690 1116.360 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2618.385 1116.370 2618.715 1116.385 ;
        RECT 2609.580 1116.280 2618.715 1116.370 ;
        RECT 2606.000 1116.070 2618.715 1116.280 ;
        RECT 2606.000 1115.680 2610.000 1116.070 ;
        RECT 2618.385 1116.055 2618.715 1116.070 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1318.080 2621.930 1318.140 ;
        RECT 2898.990 1318.080 2899.310 1318.140 ;
        RECT 2621.610 1317.940 2899.310 1318.080 ;
        RECT 2621.610 1317.880 2621.930 1317.940 ;
        RECT 2898.990 1317.880 2899.310 1317.940 ;
      LAYER via ;
        RECT 2621.640 1317.880 2621.900 1318.140 ;
        RECT 2899.020 1317.880 2899.280 1318.140 ;
      LAYER met2 ;
        RECT 2899.010 1319.355 2899.290 1319.725 ;
        RECT 2899.080 1318.170 2899.220 1319.355 ;
        RECT 2621.640 1317.850 2621.900 1318.170 ;
        RECT 2899.020 1317.850 2899.280 1318.170 ;
        RECT 2621.700 1316.325 2621.840 1317.850 ;
        RECT 2621.630 1315.955 2621.910 1316.325 ;
      LAYER via2 ;
        RECT 2899.010 1319.400 2899.290 1319.680 ;
        RECT 2621.630 1316.000 2621.910 1316.280 ;
      LAYER met3 ;
        RECT 2898.985 1319.690 2899.315 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2898.985 1319.390 2924.800 1319.690 ;
        RECT 2898.985 1319.375 2899.315 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 2621.605 1316.290 2621.935 1316.305 ;
        RECT 2609.580 1316.200 2621.935 1316.290 ;
        RECT 2606.000 1315.990 2621.935 1316.200 ;
        RECT 2606.000 1315.600 2610.000 1315.990 ;
        RECT 2621.605 1315.975 2621.935 1315.990 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1552.680 2618.710 1552.740 ;
        RECT 2898.990 1552.680 2899.310 1552.740 ;
        RECT 2618.390 1552.540 2899.310 1552.680 ;
        RECT 2618.390 1552.480 2618.710 1552.540 ;
        RECT 2898.990 1552.480 2899.310 1552.540 ;
      LAYER via ;
        RECT 2618.420 1552.480 2618.680 1552.740 ;
        RECT 2899.020 1552.480 2899.280 1552.740 ;
      LAYER met2 ;
        RECT 2899.010 1553.955 2899.290 1554.325 ;
        RECT 2899.080 1552.770 2899.220 1553.955 ;
        RECT 2618.420 1552.450 2618.680 1552.770 ;
        RECT 2899.020 1552.450 2899.280 1552.770 ;
        RECT 2618.480 1516.245 2618.620 1552.450 ;
        RECT 2618.410 1515.875 2618.690 1516.245 ;
      LAYER via2 ;
        RECT 2899.010 1554.000 2899.290 1554.280 ;
        RECT 2618.410 1515.920 2618.690 1516.200 ;
      LAYER met3 ;
        RECT 2898.985 1554.290 2899.315 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2898.985 1553.990 2924.800 1554.290 ;
        RECT 2898.985 1553.975 2899.315 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 2618.385 1516.210 2618.715 1516.225 ;
        RECT 2609.580 1516.120 2618.715 1516.210 ;
        RECT 2606.000 1515.910 2618.715 1516.120 ;
        RECT 2606.000 1515.520 2610.000 1515.910 ;
        RECT 2618.385 1515.895 2618.715 1515.910 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1787.280 2619.170 1787.340 ;
        RECT 2900.830 1787.280 2901.150 1787.340 ;
        RECT 2618.850 1787.140 2901.150 1787.280 ;
        RECT 2618.850 1787.080 2619.170 1787.140 ;
        RECT 2900.830 1787.080 2901.150 1787.140 ;
      LAYER via ;
        RECT 2618.880 1787.080 2619.140 1787.340 ;
        RECT 2900.860 1787.080 2901.120 1787.340 ;
      LAYER met2 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
        RECT 2900.920 1787.370 2901.060 1789.235 ;
        RECT 2618.880 1787.050 2619.140 1787.370 ;
        RECT 2900.860 1787.050 2901.120 1787.370 ;
        RECT 2618.940 1716.165 2619.080 1787.050 ;
        RECT 2618.870 1715.795 2619.150 1716.165 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
        RECT 2618.870 1715.840 2619.150 1716.120 ;
      LAYER met3 ;
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2618.845 1716.130 2619.175 1716.145 ;
        RECT 2609.580 1716.040 2619.175 1716.130 ;
        RECT 2606.000 1715.830 2619.175 1716.040 ;
        RECT 2606.000 1715.440 2610.000 1715.830 ;
        RECT 2618.845 1715.815 2619.175 1715.830 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2021.880 2618.710 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 2618.390 2021.740 2901.150 2021.880 ;
        RECT 2618.390 2021.680 2618.710 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 2618.420 2021.680 2618.680 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 2618.420 2021.650 2618.680 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 2618.480 1916.765 2618.620 2021.650 ;
        RECT 2618.410 1916.395 2618.690 1916.765 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
        RECT 2618.410 1916.440 2618.690 1916.720 ;
      LAYER met3 ;
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2618.385 1916.730 2618.715 1916.745 ;
        RECT 2609.580 1916.640 2618.715 1916.730 ;
        RECT 2606.000 1916.430 2618.715 1916.640 ;
        RECT 2606.000 1916.040 2610.000 1916.430 ;
        RECT 2618.385 1916.415 2618.715 1916.430 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.310 2256.480 2619.630 2256.540 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 2619.310 2256.340 2901.150 2256.480 ;
        RECT 2619.310 2256.280 2619.630 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
      LAYER via ;
        RECT 2619.340 2256.280 2619.600 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 2619.340 2256.250 2619.600 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 2619.400 2116.685 2619.540 2256.250 ;
        RECT 2619.330 2116.315 2619.610 2116.685 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
        RECT 2619.330 2116.360 2619.610 2116.640 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2619.305 2116.650 2619.635 2116.665 ;
        RECT 2609.580 2116.560 2619.635 2116.650 ;
        RECT 2606.000 2116.350 2619.635 2116.560 ;
        RECT 2606.000 2115.960 2610.000 2116.350 ;
        RECT 2619.305 2116.335 2619.635 2116.350 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 324.370 200.840 324.690 200.900 ;
        RECT 330.810 200.840 331.130 200.900 ;
        RECT 324.370 200.700 331.130 200.840 ;
        RECT 324.370 200.640 324.690 200.700 ;
        RECT 330.810 200.640 331.130 200.700 ;
        RECT 330.810 24.380 331.130 24.440 ;
        RECT 633.030 24.380 633.350 24.440 ;
        RECT 330.810 24.240 633.350 24.380 ;
        RECT 330.810 24.180 331.130 24.240 ;
        RECT 633.030 24.180 633.350 24.240 ;
      LAYER via ;
        RECT 324.400 200.640 324.660 200.900 ;
        RECT 330.840 200.640 331.100 200.900 ;
        RECT 330.840 24.180 331.100 24.440 ;
        RECT 633.060 24.180 633.320 24.440 ;
      LAYER met2 ;
        RECT 324.350 216.000 324.630 220.000 ;
        RECT 324.460 200.930 324.600 216.000 ;
        RECT 324.400 200.610 324.660 200.930 ;
        RECT 330.840 200.610 331.100 200.930 ;
        RECT 330.900 24.470 331.040 200.610 ;
        RECT 330.840 24.150 331.100 24.470 ;
        RECT 633.060 24.150 633.320 24.470 ;
        RECT 633.120 2.400 633.260 24.150 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2111.930 200.500 2112.250 200.560 ;
        RECT 2117.910 200.500 2118.230 200.560 ;
        RECT 2111.930 200.360 2118.230 200.500 ;
        RECT 2111.930 200.300 2112.250 200.360 ;
        RECT 2117.910 200.300 2118.230 200.360 ;
        RECT 2117.910 31.180 2118.230 31.240 ;
        RECT 2417.370 31.180 2417.690 31.240 ;
        RECT 2117.910 31.040 2417.690 31.180 ;
        RECT 2117.910 30.980 2118.230 31.040 ;
        RECT 2417.370 30.980 2417.690 31.040 ;
      LAYER via ;
        RECT 2111.960 200.300 2112.220 200.560 ;
        RECT 2117.940 200.300 2118.200 200.560 ;
        RECT 2117.940 30.980 2118.200 31.240 ;
        RECT 2417.400 30.980 2417.660 31.240 ;
      LAYER met2 ;
        RECT 2111.910 216.000 2112.190 220.000 ;
        RECT 2112.020 200.590 2112.160 216.000 ;
        RECT 2111.960 200.270 2112.220 200.590 ;
        RECT 2117.940 200.270 2118.200 200.590 ;
        RECT 2118.000 31.270 2118.140 200.270 ;
        RECT 2117.940 30.950 2118.200 31.270 ;
        RECT 2417.400 30.950 2417.660 31.270 ;
        RECT 2417.460 2.400 2417.600 30.950 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 37.980 2132.030 38.040 ;
        RECT 2434.850 37.980 2435.170 38.040 ;
        RECT 2131.710 37.840 2435.170 37.980 ;
        RECT 2131.710 37.780 2132.030 37.840 ;
        RECT 2434.850 37.780 2435.170 37.840 ;
      LAYER via ;
        RECT 2131.740 37.780 2132.000 38.040 ;
        RECT 2434.880 37.780 2435.140 38.040 ;
      LAYER met2 ;
        RECT 2129.850 216.650 2130.130 220.000 ;
        RECT 2129.850 216.510 2131.940 216.650 ;
        RECT 2129.850 216.000 2130.130 216.510 ;
        RECT 2131.800 38.070 2131.940 216.510 ;
        RECT 2131.740 37.750 2132.000 38.070 ;
        RECT 2434.880 37.750 2435.140 38.070 ;
        RECT 2434.940 2.400 2435.080 37.750 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2147.810 200.500 2148.130 200.560 ;
        RECT 2152.410 200.500 2152.730 200.560 ;
        RECT 2147.810 200.360 2152.730 200.500 ;
        RECT 2147.810 200.300 2148.130 200.360 ;
        RECT 2152.410 200.300 2152.730 200.360 ;
        RECT 2152.410 44.780 2152.730 44.840 ;
        RECT 2452.790 44.780 2453.110 44.840 ;
        RECT 2152.410 44.640 2453.110 44.780 ;
        RECT 2152.410 44.580 2152.730 44.640 ;
        RECT 2452.790 44.580 2453.110 44.640 ;
      LAYER via ;
        RECT 2147.840 200.300 2148.100 200.560 ;
        RECT 2152.440 200.300 2152.700 200.560 ;
        RECT 2152.440 44.580 2152.700 44.840 ;
        RECT 2452.820 44.580 2453.080 44.840 ;
      LAYER met2 ;
        RECT 2147.790 216.000 2148.070 220.000 ;
        RECT 2147.900 200.590 2148.040 216.000 ;
        RECT 2147.840 200.270 2148.100 200.590 ;
        RECT 2152.440 200.270 2152.700 200.590 ;
        RECT 2152.500 44.870 2152.640 200.270 ;
        RECT 2152.440 44.550 2152.700 44.870 ;
        RECT 2452.820 44.550 2453.080 44.870 ;
        RECT 2452.880 2.400 2453.020 44.550 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.210 196.760 2166.530 196.820 ;
        RECT 2470.270 196.760 2470.590 196.820 ;
        RECT 2166.210 196.620 2470.590 196.760 ;
        RECT 2166.210 196.560 2166.530 196.620 ;
        RECT 2470.270 196.560 2470.590 196.620 ;
      LAYER via ;
        RECT 2166.240 196.560 2166.500 196.820 ;
        RECT 2470.300 196.560 2470.560 196.820 ;
      LAYER met2 ;
        RECT 2165.730 216.650 2166.010 220.000 ;
        RECT 2165.730 216.510 2166.440 216.650 ;
        RECT 2165.730 216.000 2166.010 216.510 ;
        RECT 2166.300 196.850 2166.440 216.510 ;
        RECT 2166.240 196.530 2166.500 196.850 ;
        RECT 2470.300 196.530 2470.560 196.850 ;
        RECT 2470.360 17.410 2470.500 196.530 ;
        RECT 2470.360 17.270 2470.960 17.410 ;
        RECT 2470.820 2.400 2470.960 17.270 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 51.580 2187.230 51.640 ;
        RECT 2484.070 51.580 2484.390 51.640 ;
        RECT 2186.910 51.440 2484.390 51.580 ;
        RECT 2186.910 51.380 2187.230 51.440 ;
        RECT 2484.070 51.380 2484.390 51.440 ;
      LAYER via ;
        RECT 2186.940 51.380 2187.200 51.640 ;
        RECT 2484.100 51.380 2484.360 51.640 ;
      LAYER met2 ;
        RECT 2183.670 216.650 2183.950 220.000 ;
        RECT 2183.670 216.510 2187.140 216.650 ;
        RECT 2183.670 216.000 2183.950 216.510 ;
        RECT 2187.000 51.670 2187.140 216.510 ;
        RECT 2186.940 51.350 2187.200 51.670 ;
        RECT 2484.100 51.350 2484.360 51.670 ;
        RECT 2484.160 17.410 2484.300 51.350 ;
        RECT 2484.160 17.270 2488.900 17.410 ;
        RECT 2488.760 2.400 2488.900 17.270 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2201.630 200.500 2201.950 200.560 ;
        RECT 2207.610 200.500 2207.930 200.560 ;
        RECT 2201.630 200.360 2207.930 200.500 ;
        RECT 2201.630 200.300 2201.950 200.360 ;
        RECT 2207.610 200.300 2207.930 200.360 ;
        RECT 2207.610 59.060 2207.930 59.120 ;
        RECT 2504.770 59.060 2505.090 59.120 ;
        RECT 2207.610 58.920 2505.090 59.060 ;
        RECT 2207.610 58.860 2207.930 58.920 ;
        RECT 2504.770 58.860 2505.090 58.920 ;
      LAYER via ;
        RECT 2201.660 200.300 2201.920 200.560 ;
        RECT 2207.640 200.300 2207.900 200.560 ;
        RECT 2207.640 58.860 2207.900 59.120 ;
        RECT 2504.800 58.860 2505.060 59.120 ;
      LAYER met2 ;
        RECT 2201.610 216.000 2201.890 220.000 ;
        RECT 2201.720 200.590 2201.860 216.000 ;
        RECT 2201.660 200.270 2201.920 200.590 ;
        RECT 2207.640 200.270 2207.900 200.590 ;
        RECT 2207.700 59.150 2207.840 200.270 ;
        RECT 2207.640 58.830 2207.900 59.150 ;
        RECT 2504.800 58.830 2505.060 59.150 ;
        RECT 2504.860 16.730 2505.000 58.830 ;
        RECT 2504.860 16.590 2506.380 16.730 ;
        RECT 2506.240 2.400 2506.380 16.590 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2221.410 65.860 2221.730 65.920 ;
        RECT 2518.570 65.860 2518.890 65.920 ;
        RECT 2221.410 65.720 2518.890 65.860 ;
        RECT 2221.410 65.660 2221.730 65.720 ;
        RECT 2518.570 65.660 2518.890 65.720 ;
      LAYER via ;
        RECT 2221.440 65.660 2221.700 65.920 ;
        RECT 2518.600 65.660 2518.860 65.920 ;
      LAYER met2 ;
        RECT 2219.550 216.650 2219.830 220.000 ;
        RECT 2219.550 216.510 2221.640 216.650 ;
        RECT 2219.550 216.000 2219.830 216.510 ;
        RECT 2221.500 65.950 2221.640 216.510 ;
        RECT 2221.440 65.630 2221.700 65.950 ;
        RECT 2518.600 65.630 2518.860 65.950 ;
        RECT 2518.660 16.730 2518.800 65.630 ;
        RECT 2518.660 16.590 2524.320 16.730 ;
        RECT 2524.180 2.400 2524.320 16.590 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2237.050 200.500 2237.370 200.560 ;
        RECT 2242.110 200.500 2242.430 200.560 ;
        RECT 2237.050 200.360 2242.430 200.500 ;
        RECT 2237.050 200.300 2237.370 200.360 ;
        RECT 2242.110 200.300 2242.430 200.360 ;
        RECT 2242.110 72.320 2242.430 72.380 ;
        RECT 2539.270 72.320 2539.590 72.380 ;
        RECT 2242.110 72.180 2539.590 72.320 ;
        RECT 2242.110 72.120 2242.430 72.180 ;
        RECT 2539.270 72.120 2539.590 72.180 ;
      LAYER via ;
        RECT 2237.080 200.300 2237.340 200.560 ;
        RECT 2242.140 200.300 2242.400 200.560 ;
        RECT 2242.140 72.120 2242.400 72.380 ;
        RECT 2539.300 72.120 2539.560 72.380 ;
      LAYER met2 ;
        RECT 2237.030 216.000 2237.310 220.000 ;
        RECT 2237.140 200.590 2237.280 216.000 ;
        RECT 2237.080 200.270 2237.340 200.590 ;
        RECT 2242.140 200.270 2242.400 200.590 ;
        RECT 2242.200 72.410 2242.340 200.270 ;
        RECT 2242.140 72.090 2242.400 72.410 ;
        RECT 2539.300 72.090 2539.560 72.410 ;
        RECT 2539.360 16.730 2539.500 72.090 ;
        RECT 2539.360 16.590 2542.260 16.730 ;
        RECT 2542.120 2.400 2542.260 16.590 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2254.990 189.960 2255.310 190.020 ;
        RECT 2559.970 189.960 2560.290 190.020 ;
        RECT 2254.990 189.820 2560.290 189.960 ;
        RECT 2254.990 189.760 2255.310 189.820 ;
        RECT 2559.970 189.760 2560.290 189.820 ;
      LAYER via ;
        RECT 2255.020 189.760 2255.280 190.020 ;
        RECT 2560.000 189.760 2560.260 190.020 ;
      LAYER met2 ;
        RECT 2254.970 216.000 2255.250 220.000 ;
        RECT 2255.080 190.050 2255.220 216.000 ;
        RECT 2255.020 189.730 2255.280 190.050 ;
        RECT 2560.000 189.730 2560.260 190.050 ;
        RECT 2560.060 2.400 2560.200 189.730 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2276.610 25.740 2276.930 25.800 ;
        RECT 2577.910 25.740 2578.230 25.800 ;
        RECT 2276.610 25.600 2578.230 25.740 ;
        RECT 2276.610 25.540 2276.930 25.600 ;
        RECT 2577.910 25.540 2578.230 25.600 ;
      LAYER via ;
        RECT 2276.640 25.540 2276.900 25.800 ;
        RECT 2577.940 25.540 2578.200 25.800 ;
      LAYER met2 ;
        RECT 2272.910 216.650 2273.190 220.000 ;
        RECT 2272.910 216.510 2276.840 216.650 ;
        RECT 2272.910 216.000 2273.190 216.510 ;
        RECT 2276.700 25.830 2276.840 216.510 ;
        RECT 2276.640 25.510 2276.900 25.830 ;
        RECT 2577.940 25.510 2578.200 25.830 ;
        RECT 2578.000 2.400 2578.140 25.510 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 502.850 30.840 503.170 30.900 ;
        RECT 811.510 30.840 811.830 30.900 ;
        RECT 502.850 30.700 811.830 30.840 ;
        RECT 502.850 30.640 503.170 30.700 ;
        RECT 811.510 30.640 811.830 30.700 ;
      LAYER via ;
        RECT 502.880 30.640 503.140 30.900 ;
        RECT 811.540 30.640 811.800 30.900 ;
      LAYER met2 ;
        RECT 503.290 216.650 503.570 220.000 ;
        RECT 502.940 216.510 503.570 216.650 ;
        RECT 502.940 30.930 503.080 216.510 ;
        RECT 503.290 216.000 503.570 216.510 ;
        RECT 502.880 30.610 503.140 30.930 ;
        RECT 811.540 30.610 811.800 30.930 ;
        RECT 811.600 2.400 811.740 30.610 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2290.870 200.500 2291.190 200.560 ;
        RECT 2297.310 200.500 2297.630 200.560 ;
        RECT 2290.870 200.360 2297.630 200.500 ;
        RECT 2290.870 200.300 2291.190 200.360 ;
        RECT 2297.310 200.300 2297.630 200.360 ;
        RECT 2297.310 24.380 2297.630 24.440 ;
        RECT 2595.390 24.380 2595.710 24.440 ;
        RECT 2297.310 24.240 2595.710 24.380 ;
        RECT 2297.310 24.180 2297.630 24.240 ;
        RECT 2595.390 24.180 2595.710 24.240 ;
      LAYER via ;
        RECT 2290.900 200.300 2291.160 200.560 ;
        RECT 2297.340 200.300 2297.600 200.560 ;
        RECT 2297.340 24.180 2297.600 24.440 ;
        RECT 2595.420 24.180 2595.680 24.440 ;
      LAYER met2 ;
        RECT 2290.850 216.000 2291.130 220.000 ;
        RECT 2290.960 200.590 2291.100 216.000 ;
        RECT 2290.900 200.270 2291.160 200.590 ;
        RECT 2297.340 200.270 2297.600 200.590 ;
        RECT 2297.400 24.470 2297.540 200.270 ;
        RECT 2297.340 24.150 2297.600 24.470 ;
        RECT 2595.420 24.150 2595.680 24.470 ;
        RECT 2595.480 2.400 2595.620 24.150 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2311.110 24.720 2311.430 24.780 ;
        RECT 2613.330 24.720 2613.650 24.780 ;
        RECT 2311.110 24.580 2613.650 24.720 ;
        RECT 2311.110 24.520 2311.430 24.580 ;
        RECT 2613.330 24.520 2613.650 24.580 ;
      LAYER via ;
        RECT 2311.140 24.520 2311.400 24.780 ;
        RECT 2613.360 24.520 2613.620 24.780 ;
      LAYER met2 ;
        RECT 2308.790 216.650 2309.070 220.000 ;
        RECT 2308.790 216.510 2311.340 216.650 ;
        RECT 2308.790 216.000 2309.070 216.510 ;
        RECT 2311.200 24.810 2311.340 216.510 ;
        RECT 2311.140 24.490 2311.400 24.810 ;
        RECT 2613.360 24.490 2613.620 24.810 ;
        RECT 2613.420 2.400 2613.560 24.490 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2326.750 200.500 2327.070 200.560 ;
        RECT 2331.810 200.500 2332.130 200.560 ;
        RECT 2326.750 200.360 2332.130 200.500 ;
        RECT 2326.750 200.300 2327.070 200.360 ;
        RECT 2331.810 200.300 2332.130 200.360 ;
        RECT 2331.810 26.080 2332.130 26.140 ;
        RECT 2631.270 26.080 2631.590 26.140 ;
        RECT 2331.810 25.940 2631.590 26.080 ;
        RECT 2331.810 25.880 2332.130 25.940 ;
        RECT 2631.270 25.880 2631.590 25.940 ;
      LAYER via ;
        RECT 2326.780 200.300 2327.040 200.560 ;
        RECT 2331.840 200.300 2332.100 200.560 ;
        RECT 2331.840 25.880 2332.100 26.140 ;
        RECT 2631.300 25.880 2631.560 26.140 ;
      LAYER met2 ;
        RECT 2326.730 216.000 2327.010 220.000 ;
        RECT 2326.840 200.590 2326.980 216.000 ;
        RECT 2326.780 200.270 2327.040 200.590 ;
        RECT 2331.840 200.270 2332.100 200.590 ;
        RECT 2331.900 26.170 2332.040 200.270 ;
        RECT 2331.840 25.850 2332.100 26.170 ;
        RECT 2631.300 25.850 2631.560 26.170 ;
        RECT 2631.360 2.400 2631.500 25.850 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 79.460 2345.930 79.520 ;
        RECT 2643.230 79.460 2643.550 79.520 ;
        RECT 2345.610 79.320 2643.550 79.460 ;
        RECT 2345.610 79.260 2345.930 79.320 ;
        RECT 2643.230 79.260 2643.550 79.320 ;
        RECT 2643.230 18.260 2643.550 18.320 ;
        RECT 2649.210 18.260 2649.530 18.320 ;
        RECT 2643.230 18.120 2649.530 18.260 ;
        RECT 2643.230 18.060 2643.550 18.120 ;
        RECT 2649.210 18.060 2649.530 18.120 ;
      LAYER via ;
        RECT 2345.640 79.260 2345.900 79.520 ;
        RECT 2643.260 79.260 2643.520 79.520 ;
        RECT 2643.260 18.060 2643.520 18.320 ;
        RECT 2649.240 18.060 2649.500 18.320 ;
      LAYER met2 ;
        RECT 2344.670 216.650 2344.950 220.000 ;
        RECT 2344.670 216.510 2345.840 216.650 ;
        RECT 2344.670 216.000 2344.950 216.510 ;
        RECT 2345.700 79.550 2345.840 216.510 ;
        RECT 2345.640 79.230 2345.900 79.550 ;
        RECT 2643.260 79.230 2643.520 79.550 ;
        RECT 2643.320 18.350 2643.460 79.230 ;
        RECT 2643.260 18.030 2643.520 18.350 ;
        RECT 2649.240 18.030 2649.500 18.350 ;
        RECT 2649.300 2.400 2649.440 18.030 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2362.170 200.500 2362.490 200.560 ;
        RECT 2366.310 200.500 2366.630 200.560 ;
        RECT 2362.170 200.360 2366.630 200.500 ;
        RECT 2362.170 200.300 2362.490 200.360 ;
        RECT 2366.310 200.300 2366.630 200.360 ;
        RECT 2366.310 26.420 2366.630 26.480 ;
        RECT 2667.150 26.420 2667.470 26.480 ;
        RECT 2366.310 26.280 2667.470 26.420 ;
        RECT 2366.310 26.220 2366.630 26.280 ;
        RECT 2667.150 26.220 2667.470 26.280 ;
      LAYER via ;
        RECT 2362.200 200.300 2362.460 200.560 ;
        RECT 2366.340 200.300 2366.600 200.560 ;
        RECT 2366.340 26.220 2366.600 26.480 ;
        RECT 2667.180 26.220 2667.440 26.480 ;
      LAYER met2 ;
        RECT 2362.150 216.000 2362.430 220.000 ;
        RECT 2362.260 200.590 2362.400 216.000 ;
        RECT 2362.200 200.270 2362.460 200.590 ;
        RECT 2366.340 200.270 2366.600 200.590 ;
        RECT 2366.400 26.510 2366.540 200.270 ;
        RECT 2366.340 26.190 2366.600 26.510 ;
        RECT 2667.180 26.190 2667.440 26.510 ;
        RECT 2667.240 2.400 2667.380 26.190 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2380.110 24.040 2380.430 24.100 ;
        RECT 2684.630 24.040 2684.950 24.100 ;
        RECT 2380.110 23.900 2684.950 24.040 ;
        RECT 2380.110 23.840 2380.430 23.900 ;
        RECT 2684.630 23.840 2684.950 23.900 ;
      LAYER via ;
        RECT 2380.140 23.840 2380.400 24.100 ;
        RECT 2684.660 23.840 2684.920 24.100 ;
      LAYER met2 ;
        RECT 2380.090 216.000 2380.370 220.000 ;
        RECT 2380.200 24.130 2380.340 216.000 ;
        RECT 2380.140 23.810 2380.400 24.130 ;
        RECT 2684.660 23.810 2684.920 24.130 ;
        RECT 2684.720 2.400 2684.860 23.810 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.810 25.060 2401.130 25.120 ;
        RECT 2702.570 25.060 2702.890 25.120 ;
        RECT 2400.810 24.920 2702.890 25.060 ;
        RECT 2400.810 24.860 2401.130 24.920 ;
        RECT 2702.570 24.860 2702.890 24.920 ;
      LAYER via ;
        RECT 2400.840 24.860 2401.100 25.120 ;
        RECT 2702.600 24.860 2702.860 25.120 ;
      LAYER met2 ;
        RECT 2398.030 216.650 2398.310 220.000 ;
        RECT 2398.030 216.510 2401.040 216.650 ;
        RECT 2398.030 216.000 2398.310 216.510 ;
        RECT 2400.900 25.150 2401.040 216.510 ;
        RECT 2400.840 24.830 2401.100 25.150 ;
        RECT 2702.600 24.830 2702.860 25.150 ;
        RECT 2702.660 2.400 2702.800 24.830 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2415.990 200.500 2416.310 200.560 ;
        RECT 2421.510 200.500 2421.830 200.560 ;
        RECT 2415.990 200.360 2421.830 200.500 ;
        RECT 2415.990 200.300 2416.310 200.360 ;
        RECT 2421.510 200.300 2421.830 200.360 ;
        RECT 2421.510 27.100 2421.830 27.160 ;
        RECT 2720.510 27.100 2720.830 27.160 ;
        RECT 2421.510 26.960 2720.830 27.100 ;
        RECT 2421.510 26.900 2421.830 26.960 ;
        RECT 2720.510 26.900 2720.830 26.960 ;
      LAYER via ;
        RECT 2416.020 200.300 2416.280 200.560 ;
        RECT 2421.540 200.300 2421.800 200.560 ;
        RECT 2421.540 26.900 2421.800 27.160 ;
        RECT 2720.540 26.900 2720.800 27.160 ;
      LAYER met2 ;
        RECT 2415.970 216.000 2416.250 220.000 ;
        RECT 2416.080 200.590 2416.220 216.000 ;
        RECT 2416.020 200.270 2416.280 200.590 ;
        RECT 2421.540 200.270 2421.800 200.590 ;
        RECT 2421.600 27.190 2421.740 200.270 ;
        RECT 2421.540 26.870 2421.800 27.190 ;
        RECT 2720.540 26.870 2720.800 27.190 ;
        RECT 2720.600 2.400 2720.740 26.870 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2435.310 26.760 2435.630 26.820 ;
        RECT 2738.450 26.760 2738.770 26.820 ;
        RECT 2435.310 26.620 2738.770 26.760 ;
        RECT 2435.310 26.560 2435.630 26.620 ;
        RECT 2738.450 26.560 2738.770 26.620 ;
      LAYER via ;
        RECT 2435.340 26.560 2435.600 26.820 ;
        RECT 2738.480 26.560 2738.740 26.820 ;
      LAYER met2 ;
        RECT 2433.910 216.650 2434.190 220.000 ;
        RECT 2433.910 216.510 2435.540 216.650 ;
        RECT 2433.910 216.000 2434.190 216.510 ;
        RECT 2435.400 26.850 2435.540 216.510 ;
        RECT 2435.340 26.530 2435.600 26.850 ;
        RECT 2738.480 26.530 2738.740 26.850 ;
        RECT 2738.540 2.400 2738.680 26.530 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2451.870 200.500 2452.190 200.560 ;
        RECT 2456.010 200.500 2456.330 200.560 ;
        RECT 2451.870 200.360 2456.330 200.500 ;
        RECT 2451.870 200.300 2452.190 200.360 ;
        RECT 2456.010 200.300 2456.330 200.360 ;
        RECT 2456.010 44.780 2456.330 44.840 ;
        RECT 2755.930 44.780 2756.250 44.840 ;
        RECT 2456.010 44.640 2756.250 44.780 ;
        RECT 2456.010 44.580 2456.330 44.640 ;
        RECT 2755.930 44.580 2756.250 44.640 ;
      LAYER via ;
        RECT 2451.900 200.300 2452.160 200.560 ;
        RECT 2456.040 200.300 2456.300 200.560 ;
        RECT 2456.040 44.580 2456.300 44.840 ;
        RECT 2755.960 44.580 2756.220 44.840 ;
      LAYER met2 ;
        RECT 2451.850 216.000 2452.130 220.000 ;
        RECT 2451.960 200.590 2452.100 216.000 ;
        RECT 2451.900 200.270 2452.160 200.590 ;
        RECT 2456.040 200.270 2456.300 200.590 ;
        RECT 2456.100 44.870 2456.240 200.270 ;
        RECT 2456.040 44.550 2456.300 44.870 ;
        RECT 2755.960 44.550 2756.220 44.870 ;
        RECT 2756.020 2.400 2756.160 44.550 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 524.010 38.320 524.330 38.380 ;
        RECT 829.450 38.320 829.770 38.380 ;
        RECT 524.010 38.180 829.770 38.320 ;
        RECT 524.010 38.120 524.330 38.180 ;
        RECT 829.450 38.120 829.770 38.180 ;
      LAYER via ;
        RECT 524.040 38.120 524.300 38.380 ;
        RECT 829.480 38.120 829.740 38.380 ;
      LAYER met2 ;
        RECT 521.230 216.650 521.510 220.000 ;
        RECT 521.230 216.510 524.240 216.650 ;
        RECT 521.230 216.000 521.510 216.510 ;
        RECT 524.100 38.410 524.240 216.510 ;
        RECT 524.040 38.090 524.300 38.410 ;
        RECT 829.480 38.090 829.740 38.410 ;
        RECT 829.540 2.400 829.680 38.090 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2469.350 182.820 2469.670 182.880 ;
        RECT 2773.870 182.820 2774.190 182.880 ;
        RECT 2469.350 182.680 2774.190 182.820 ;
        RECT 2469.350 182.620 2469.670 182.680 ;
        RECT 2773.870 182.620 2774.190 182.680 ;
      LAYER via ;
        RECT 2469.380 182.620 2469.640 182.880 ;
        RECT 2773.900 182.620 2774.160 182.880 ;
      LAYER met2 ;
        RECT 2469.790 216.650 2470.070 220.000 ;
        RECT 2469.440 216.510 2470.070 216.650 ;
        RECT 2469.440 182.910 2469.580 216.510 ;
        RECT 2469.790 216.000 2470.070 216.510 ;
        RECT 2469.380 182.590 2469.640 182.910 ;
        RECT 2773.900 182.590 2774.160 182.910 ;
        RECT 2773.960 2.400 2774.100 182.590 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2490.510 51.580 2490.830 51.640 ;
        RECT 2787.670 51.580 2787.990 51.640 ;
        RECT 2490.510 51.440 2787.990 51.580 ;
        RECT 2490.510 51.380 2490.830 51.440 ;
        RECT 2787.670 51.380 2787.990 51.440 ;
      LAYER via ;
        RECT 2490.540 51.380 2490.800 51.640 ;
        RECT 2787.700 51.380 2787.960 51.640 ;
      LAYER met2 ;
        RECT 2487.270 216.650 2487.550 220.000 ;
        RECT 2487.270 216.510 2490.740 216.650 ;
        RECT 2487.270 216.000 2487.550 216.510 ;
        RECT 2490.600 51.670 2490.740 216.510 ;
        RECT 2490.540 51.350 2490.800 51.670 ;
        RECT 2787.700 51.350 2787.960 51.670 ;
        RECT 2787.760 17.410 2787.900 51.350 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2505.230 196.760 2505.550 196.820 ;
        RECT 2808.370 196.760 2808.690 196.820 ;
        RECT 2505.230 196.620 2808.690 196.760 ;
        RECT 2505.230 196.560 2505.550 196.620 ;
        RECT 2808.370 196.560 2808.690 196.620 ;
      LAYER via ;
        RECT 2505.260 196.560 2505.520 196.820 ;
        RECT 2808.400 196.560 2808.660 196.820 ;
      LAYER met2 ;
        RECT 2505.210 216.000 2505.490 220.000 ;
        RECT 2505.320 196.850 2505.460 216.000 ;
        RECT 2505.260 196.530 2505.520 196.850 ;
        RECT 2808.400 196.530 2808.660 196.850 ;
        RECT 2808.460 17.410 2808.600 196.530 ;
        RECT 2808.460 17.270 2809.980 17.410 ;
        RECT 2809.840 2.400 2809.980 17.270 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2525.010 65.520 2525.330 65.580 ;
        RECT 2822.170 65.520 2822.490 65.580 ;
        RECT 2525.010 65.380 2822.490 65.520 ;
        RECT 2525.010 65.320 2525.330 65.380 ;
        RECT 2822.170 65.320 2822.490 65.380 ;
      LAYER via ;
        RECT 2525.040 65.320 2525.300 65.580 ;
        RECT 2822.200 65.320 2822.460 65.580 ;
      LAYER met2 ;
        RECT 2523.150 216.650 2523.430 220.000 ;
        RECT 2523.150 216.510 2525.240 216.650 ;
        RECT 2523.150 216.000 2523.430 216.510 ;
        RECT 2525.100 65.610 2525.240 216.510 ;
        RECT 2525.040 65.290 2525.300 65.610 ;
        RECT 2822.200 65.290 2822.460 65.610 ;
        RECT 2822.260 17.410 2822.400 65.290 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2541.110 200.500 2541.430 200.560 ;
        RECT 2545.710 200.500 2546.030 200.560 ;
        RECT 2541.110 200.360 2546.030 200.500 ;
        RECT 2541.110 200.300 2541.430 200.360 ;
        RECT 2545.710 200.300 2546.030 200.360 ;
        RECT 2545.710 72.320 2546.030 72.380 ;
        RECT 2842.870 72.320 2843.190 72.380 ;
        RECT 2545.710 72.180 2843.190 72.320 ;
        RECT 2545.710 72.120 2546.030 72.180 ;
        RECT 2842.870 72.120 2843.190 72.180 ;
      LAYER via ;
        RECT 2541.140 200.300 2541.400 200.560 ;
        RECT 2545.740 200.300 2546.000 200.560 ;
        RECT 2545.740 72.120 2546.000 72.380 ;
        RECT 2842.900 72.120 2843.160 72.380 ;
      LAYER met2 ;
        RECT 2541.090 216.000 2541.370 220.000 ;
        RECT 2541.200 200.590 2541.340 216.000 ;
        RECT 2541.140 200.270 2541.400 200.590 ;
        RECT 2545.740 200.270 2546.000 200.590 ;
        RECT 2545.800 72.410 2545.940 200.270 ;
        RECT 2545.740 72.090 2546.000 72.410 ;
        RECT 2842.900 72.090 2843.160 72.410 ;
        RECT 2842.960 17.410 2843.100 72.090 ;
        RECT 2842.960 17.270 2845.400 17.410 ;
        RECT 2845.260 2.400 2845.400 17.270 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2559.050 176.020 2559.370 176.080 ;
        RECT 2857.130 176.020 2857.450 176.080 ;
        RECT 2559.050 175.880 2857.450 176.020 ;
        RECT 2559.050 175.820 2559.370 175.880 ;
        RECT 2857.130 175.820 2857.450 175.880 ;
        RECT 2857.130 17.580 2857.450 17.640 ;
        RECT 2863.110 17.580 2863.430 17.640 ;
        RECT 2857.130 17.440 2863.430 17.580 ;
        RECT 2857.130 17.380 2857.450 17.440 ;
        RECT 2863.110 17.380 2863.430 17.440 ;
      LAYER via ;
        RECT 2559.080 175.820 2559.340 176.080 ;
        RECT 2857.160 175.820 2857.420 176.080 ;
        RECT 2857.160 17.380 2857.420 17.640 ;
        RECT 2863.140 17.380 2863.400 17.640 ;
      LAYER met2 ;
        RECT 2559.030 216.000 2559.310 220.000 ;
        RECT 2559.140 176.110 2559.280 216.000 ;
        RECT 2559.080 175.790 2559.340 176.110 ;
        RECT 2857.160 175.790 2857.420 176.110 ;
        RECT 2857.220 17.670 2857.360 175.790 ;
        RECT 2857.160 17.350 2857.420 17.670 ;
        RECT 2863.140 17.350 2863.400 17.670 ;
        RECT 2863.200 2.400 2863.340 17.350 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2580.210 30.840 2580.530 30.900 ;
        RECT 2881.050 30.840 2881.370 30.900 ;
        RECT 2580.210 30.700 2881.370 30.840 ;
        RECT 2580.210 30.640 2580.530 30.700 ;
        RECT 2881.050 30.640 2881.370 30.700 ;
      LAYER via ;
        RECT 2580.240 30.640 2580.500 30.900 ;
        RECT 2881.080 30.640 2881.340 30.900 ;
      LAYER met2 ;
        RECT 2576.970 216.650 2577.250 220.000 ;
        RECT 2576.970 216.510 2580.440 216.650 ;
        RECT 2576.970 216.000 2577.250 216.510 ;
        RECT 2580.300 30.930 2580.440 216.510 ;
        RECT 2580.240 30.610 2580.500 30.930 ;
        RECT 2881.080 30.610 2881.340 30.930 ;
        RECT 2881.140 2.400 2881.280 30.610 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2594.930 200.500 2595.250 200.560 ;
        RECT 2600.450 200.500 2600.770 200.560 ;
        RECT 2594.930 200.360 2600.770 200.500 ;
        RECT 2594.930 200.300 2595.250 200.360 ;
        RECT 2600.450 200.300 2600.770 200.360 ;
        RECT 2600.450 37.980 2600.770 38.040 ;
        RECT 2898.990 37.980 2899.310 38.040 ;
        RECT 2600.450 37.840 2899.310 37.980 ;
        RECT 2600.450 37.780 2600.770 37.840 ;
        RECT 2898.990 37.780 2899.310 37.840 ;
      LAYER via ;
        RECT 2594.960 200.300 2595.220 200.560 ;
        RECT 2600.480 200.300 2600.740 200.560 ;
        RECT 2600.480 37.780 2600.740 38.040 ;
        RECT 2899.020 37.780 2899.280 38.040 ;
      LAYER met2 ;
        RECT 2594.910 216.000 2595.190 220.000 ;
        RECT 2595.020 200.590 2595.160 216.000 ;
        RECT 2594.960 200.270 2595.220 200.590 ;
        RECT 2600.480 200.270 2600.740 200.590 ;
        RECT 2600.540 38.070 2600.680 200.270 ;
        RECT 2600.480 37.750 2600.740 38.070 ;
        RECT 2899.020 37.750 2899.280 38.070 ;
        RECT 2899.080 2.400 2899.220 37.750 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 539.190 200.500 539.510 200.560 ;
        RECT 544.710 200.500 545.030 200.560 ;
        RECT 539.190 200.360 545.030 200.500 ;
        RECT 539.190 200.300 539.510 200.360 ;
        RECT 544.710 200.300 545.030 200.360 ;
        RECT 544.710 44.780 545.030 44.840 ;
        RECT 846.930 44.780 847.250 44.840 ;
        RECT 544.710 44.640 847.250 44.780 ;
        RECT 544.710 44.580 545.030 44.640 ;
        RECT 846.930 44.580 847.250 44.640 ;
      LAYER via ;
        RECT 539.220 200.300 539.480 200.560 ;
        RECT 544.740 200.300 545.000 200.560 ;
        RECT 544.740 44.580 545.000 44.840 ;
        RECT 846.960 44.580 847.220 44.840 ;
      LAYER met2 ;
        RECT 539.170 216.000 539.450 220.000 ;
        RECT 539.280 200.590 539.420 216.000 ;
        RECT 539.220 200.270 539.480 200.590 ;
        RECT 544.740 200.270 545.000 200.590 ;
        RECT 544.800 44.870 544.940 200.270 ;
        RECT 544.740 44.550 545.000 44.870 ;
        RECT 846.960 44.550 847.220 44.870 ;
        RECT 847.020 2.400 847.160 44.550 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.510 51.580 558.830 51.640 ;
        RECT 862.570 51.580 862.890 51.640 ;
        RECT 558.510 51.440 862.890 51.580 ;
        RECT 558.510 51.380 558.830 51.440 ;
        RECT 862.570 51.380 862.890 51.440 ;
      LAYER via ;
        RECT 558.540 51.380 558.800 51.640 ;
        RECT 862.600 51.380 862.860 51.640 ;
      LAYER met2 ;
        RECT 557.110 216.650 557.390 220.000 ;
        RECT 557.110 216.510 558.740 216.650 ;
        RECT 557.110 216.000 557.390 216.510 ;
        RECT 558.600 51.670 558.740 216.510 ;
        RECT 558.540 51.350 558.800 51.670 ;
        RECT 862.600 51.350 862.860 51.670 ;
        RECT 862.660 16.730 862.800 51.350 ;
        RECT 862.660 16.590 865.100 16.730 ;
        RECT 864.960 2.400 865.100 16.590 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 574.610 200.500 574.930 200.560 ;
        RECT 579.210 200.500 579.530 200.560 ;
        RECT 574.610 200.360 579.530 200.500 ;
        RECT 574.610 200.300 574.930 200.360 ;
        RECT 579.210 200.300 579.530 200.360 ;
        RECT 579.210 58.720 579.530 58.780 ;
        RECT 876.830 58.720 877.150 58.780 ;
        RECT 579.210 58.580 877.150 58.720 ;
        RECT 579.210 58.520 579.530 58.580 ;
        RECT 876.830 58.520 877.150 58.580 ;
        RECT 876.830 16.560 877.150 16.620 ;
        RECT 882.810 16.560 883.130 16.620 ;
        RECT 876.830 16.420 883.130 16.560 ;
        RECT 876.830 16.360 877.150 16.420 ;
        RECT 882.810 16.360 883.130 16.420 ;
      LAYER via ;
        RECT 574.640 200.300 574.900 200.560 ;
        RECT 579.240 200.300 579.500 200.560 ;
        RECT 579.240 58.520 579.500 58.780 ;
        RECT 876.860 58.520 877.120 58.780 ;
        RECT 876.860 16.360 877.120 16.620 ;
        RECT 882.840 16.360 883.100 16.620 ;
      LAYER met2 ;
        RECT 574.590 216.000 574.870 220.000 ;
        RECT 574.700 200.590 574.840 216.000 ;
        RECT 574.640 200.270 574.900 200.590 ;
        RECT 579.240 200.270 579.500 200.590 ;
        RECT 579.300 58.810 579.440 200.270 ;
        RECT 579.240 58.490 579.500 58.810 ;
        RECT 876.860 58.490 877.120 58.810 ;
        RECT 876.920 16.650 877.060 58.490 ;
        RECT 876.860 16.330 877.120 16.650 ;
        RECT 882.840 16.330 883.100 16.650 ;
        RECT 882.900 2.400 883.040 16.330 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 592.550 65.520 592.870 65.580 ;
        RECT 897.070 65.520 897.390 65.580 ;
        RECT 592.550 65.380 897.390 65.520 ;
        RECT 592.550 65.320 592.870 65.380 ;
        RECT 897.070 65.320 897.390 65.380 ;
      LAYER via ;
        RECT 592.580 65.320 592.840 65.580 ;
        RECT 897.100 65.320 897.360 65.580 ;
      LAYER met2 ;
        RECT 592.530 216.000 592.810 220.000 ;
        RECT 592.640 65.610 592.780 216.000 ;
        RECT 592.580 65.290 592.840 65.610 ;
        RECT 897.100 65.290 897.360 65.610 ;
        RECT 897.160 16.730 897.300 65.290 ;
        RECT 897.160 16.590 900.980 16.730 ;
        RECT 900.840 2.400 900.980 16.590 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 613.710 72.320 614.030 72.380 ;
        RECT 918.230 72.320 918.550 72.380 ;
        RECT 613.710 72.180 918.550 72.320 ;
        RECT 613.710 72.120 614.030 72.180 ;
        RECT 918.230 72.120 918.550 72.180 ;
      LAYER via ;
        RECT 613.740 72.120 614.000 72.380 ;
        RECT 918.260 72.120 918.520 72.380 ;
      LAYER met2 ;
        RECT 610.470 216.650 610.750 220.000 ;
        RECT 610.470 216.510 613.940 216.650 ;
        RECT 610.470 216.000 610.750 216.510 ;
        RECT 613.800 72.410 613.940 216.510 ;
        RECT 613.740 72.090 614.000 72.410 ;
        RECT 918.260 72.090 918.520 72.410 ;
        RECT 918.320 17.410 918.460 72.090 ;
        RECT 918.320 17.270 918.920 17.410 ;
        RECT 918.780 2.400 918.920 17.270 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 628.430 201.860 628.750 201.920 ;
        RECT 633.950 201.860 634.270 201.920 ;
        RECT 628.430 201.720 634.270 201.860 ;
        RECT 628.430 201.660 628.750 201.720 ;
        RECT 633.950 201.660 634.270 201.720 ;
        RECT 633.950 79.800 634.270 79.860 ;
        RECT 931.570 79.800 931.890 79.860 ;
        RECT 633.950 79.660 931.890 79.800 ;
        RECT 633.950 79.600 634.270 79.660 ;
        RECT 931.570 79.600 931.890 79.660 ;
      LAYER via ;
        RECT 628.460 201.660 628.720 201.920 ;
        RECT 633.980 201.660 634.240 201.920 ;
        RECT 633.980 79.600 634.240 79.860 ;
        RECT 931.600 79.600 931.860 79.860 ;
      LAYER met2 ;
        RECT 628.410 216.000 628.690 220.000 ;
        RECT 628.520 201.950 628.660 216.000 ;
        RECT 628.460 201.630 628.720 201.950 ;
        RECT 633.980 201.630 634.240 201.950 ;
        RECT 634.040 79.890 634.180 201.630 ;
        RECT 633.980 79.570 634.240 79.890 ;
        RECT 931.600 79.570 931.860 79.890 ;
        RECT 931.660 16.730 931.800 79.570 ;
        RECT 931.660 16.590 936.400 16.730 ;
        RECT 936.260 2.400 936.400 16.590 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 86.260 648.530 86.320 ;
        RECT 952.270 86.260 952.590 86.320 ;
        RECT 648.210 86.120 952.590 86.260 ;
        RECT 648.210 86.060 648.530 86.120 ;
        RECT 952.270 86.060 952.590 86.120 ;
      LAYER via ;
        RECT 648.240 86.060 648.500 86.320 ;
        RECT 952.300 86.060 952.560 86.320 ;
      LAYER met2 ;
        RECT 646.350 216.650 646.630 220.000 ;
        RECT 646.350 216.510 648.440 216.650 ;
        RECT 646.350 216.000 646.630 216.510 ;
        RECT 648.300 86.350 648.440 216.510 ;
        RECT 648.240 86.030 648.500 86.350 ;
        RECT 952.300 86.030 952.560 86.350 ;
        RECT 952.360 16.730 952.500 86.030 ;
        RECT 952.360 16.590 954.340 16.730 ;
        RECT 954.200 2.400 954.340 16.590 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 664.310 200.500 664.630 200.560 ;
        RECT 668.910 200.500 669.230 200.560 ;
        RECT 664.310 200.360 669.230 200.500 ;
        RECT 664.310 200.300 664.630 200.360 ;
        RECT 668.910 200.300 669.230 200.360 ;
        RECT 668.910 24.720 669.230 24.780 ;
        RECT 972.050 24.720 972.370 24.780 ;
        RECT 668.910 24.580 972.370 24.720 ;
        RECT 668.910 24.520 669.230 24.580 ;
        RECT 972.050 24.520 972.370 24.580 ;
      LAYER via ;
        RECT 664.340 200.300 664.600 200.560 ;
        RECT 668.940 200.300 669.200 200.560 ;
        RECT 668.940 24.520 669.200 24.780 ;
        RECT 972.080 24.520 972.340 24.780 ;
      LAYER met2 ;
        RECT 664.290 216.000 664.570 220.000 ;
        RECT 664.400 200.590 664.540 216.000 ;
        RECT 664.340 200.270 664.600 200.590 ;
        RECT 668.940 200.270 669.200 200.590 ;
        RECT 669.000 24.810 669.140 200.270 ;
        RECT 668.940 24.490 669.200 24.810 ;
        RECT 972.080 24.490 972.340 24.810 ;
        RECT 972.140 2.400 972.280 24.490 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 344.610 24.040 344.930 24.100 ;
        RECT 650.970 24.040 651.290 24.100 ;
        RECT 344.610 23.900 651.290 24.040 ;
        RECT 344.610 23.840 344.930 23.900 ;
        RECT 650.970 23.840 651.290 23.900 ;
      LAYER via ;
        RECT 344.640 23.840 344.900 24.100 ;
        RECT 651.000 23.840 651.260 24.100 ;
      LAYER met2 ;
        RECT 342.290 216.650 342.570 220.000 ;
        RECT 342.290 216.510 344.840 216.650 ;
        RECT 342.290 216.000 342.570 216.510 ;
        RECT 344.700 24.130 344.840 216.510 ;
        RECT 344.640 23.810 344.900 24.130 ;
        RECT 651.000 23.810 651.260 24.130 ;
        RECT 651.060 2.400 651.200 23.810 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.250 93.060 682.570 93.120 ;
        RECT 986.770 93.060 987.090 93.120 ;
        RECT 682.250 92.920 987.090 93.060 ;
        RECT 682.250 92.860 682.570 92.920 ;
        RECT 986.770 92.860 987.090 92.920 ;
      LAYER via ;
        RECT 682.280 92.860 682.540 93.120 ;
        RECT 986.800 92.860 987.060 93.120 ;
      LAYER met2 ;
        RECT 682.230 216.000 682.510 220.000 ;
        RECT 682.340 93.150 682.480 216.000 ;
        RECT 682.280 92.830 682.540 93.150 ;
        RECT 986.800 92.830 987.060 93.150 ;
        RECT 986.860 16.730 987.000 92.830 ;
        RECT 986.860 16.590 990.220 16.730 ;
        RECT 990.080 2.400 990.220 16.590 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 99.860 703.730 99.920 ;
        RECT 1007.930 99.860 1008.250 99.920 ;
        RECT 703.410 99.720 1008.250 99.860 ;
        RECT 703.410 99.660 703.730 99.720 ;
        RECT 1007.930 99.660 1008.250 99.720 ;
      LAYER via ;
        RECT 703.440 99.660 703.700 99.920 ;
        RECT 1007.960 99.660 1008.220 99.920 ;
      LAYER met2 ;
        RECT 699.710 216.650 699.990 220.000 ;
        RECT 699.710 216.510 703.640 216.650 ;
        RECT 699.710 216.000 699.990 216.510 ;
        RECT 703.500 99.950 703.640 216.510 ;
        RECT 703.440 99.630 703.700 99.950 ;
        RECT 1007.960 99.630 1008.220 99.950 ;
        RECT 1008.020 17.410 1008.160 99.630 ;
        RECT 1007.560 17.270 1008.160 17.410 ;
        RECT 1007.560 2.400 1007.700 17.270 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.670 201.180 717.990 201.240 ;
        RECT 724.110 201.180 724.430 201.240 ;
        RECT 717.670 201.040 724.430 201.180 ;
        RECT 717.670 200.980 717.990 201.040 ;
        RECT 724.110 200.980 724.430 201.040 ;
        RECT 724.110 107.000 724.430 107.060 ;
        RECT 1021.270 107.000 1021.590 107.060 ;
        RECT 724.110 106.860 1021.590 107.000 ;
        RECT 724.110 106.800 724.430 106.860 ;
        RECT 1021.270 106.800 1021.590 106.860 ;
      LAYER via ;
        RECT 717.700 200.980 717.960 201.240 ;
        RECT 724.140 200.980 724.400 201.240 ;
        RECT 724.140 106.800 724.400 107.060 ;
        RECT 1021.300 106.800 1021.560 107.060 ;
      LAYER met2 ;
        RECT 717.650 216.000 717.930 220.000 ;
        RECT 717.760 201.270 717.900 216.000 ;
        RECT 717.700 200.950 717.960 201.270 ;
        RECT 724.140 200.950 724.400 201.270 ;
        RECT 724.200 107.090 724.340 200.950 ;
        RECT 724.140 106.770 724.400 107.090 ;
        RECT 1021.300 106.770 1021.560 107.090 ;
        RECT 1021.360 16.730 1021.500 106.770 ;
        RECT 1021.360 16.590 1025.640 16.730 ;
        RECT 1025.500 2.400 1025.640 16.590 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 113.800 738.230 113.860 ;
        RECT 1041.970 113.800 1042.290 113.860 ;
        RECT 737.910 113.660 1042.290 113.800 ;
        RECT 737.910 113.600 738.230 113.660 ;
        RECT 1041.970 113.600 1042.290 113.660 ;
      LAYER via ;
        RECT 737.940 113.600 738.200 113.860 ;
        RECT 1042.000 113.600 1042.260 113.860 ;
      LAYER met2 ;
        RECT 735.590 216.650 735.870 220.000 ;
        RECT 735.590 216.510 738.140 216.650 ;
        RECT 735.590 216.000 735.870 216.510 ;
        RECT 738.000 113.890 738.140 216.510 ;
        RECT 737.940 113.570 738.200 113.890 ;
        RECT 1042.000 113.570 1042.260 113.890 ;
        RECT 1042.060 16.730 1042.200 113.570 ;
        RECT 1042.060 16.590 1043.580 16.730 ;
        RECT 1043.440 2.400 1043.580 16.590 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 753.550 200.500 753.870 200.560 ;
        RECT 758.610 200.500 758.930 200.560 ;
        RECT 753.550 200.360 758.930 200.500 ;
        RECT 753.550 200.300 753.870 200.360 ;
        RECT 758.610 200.300 758.930 200.360 ;
        RECT 758.610 120.600 758.930 120.660 ;
        RECT 1055.770 120.600 1056.090 120.660 ;
        RECT 758.610 120.460 1056.090 120.600 ;
        RECT 758.610 120.400 758.930 120.460 ;
        RECT 1055.770 120.400 1056.090 120.460 ;
      LAYER via ;
        RECT 753.580 200.300 753.840 200.560 ;
        RECT 758.640 200.300 758.900 200.560 ;
        RECT 758.640 120.400 758.900 120.660 ;
        RECT 1055.800 120.400 1056.060 120.660 ;
      LAYER met2 ;
        RECT 753.530 216.000 753.810 220.000 ;
        RECT 753.640 200.590 753.780 216.000 ;
        RECT 753.580 200.270 753.840 200.590 ;
        RECT 758.640 200.270 758.900 200.590 ;
        RECT 758.700 120.690 758.840 200.270 ;
        RECT 758.640 120.370 758.900 120.690 ;
        RECT 1055.800 120.370 1056.060 120.690 ;
        RECT 1055.860 16.730 1056.000 120.370 ;
        RECT 1055.860 16.590 1061.520 16.730 ;
        RECT 1061.380 2.400 1061.520 16.590 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 772.410 127.740 772.730 127.800 ;
        RECT 1076.470 127.740 1076.790 127.800 ;
        RECT 772.410 127.600 1076.790 127.740 ;
        RECT 772.410 127.540 772.730 127.600 ;
        RECT 1076.470 127.540 1076.790 127.600 ;
      LAYER via ;
        RECT 772.440 127.540 772.700 127.800 ;
        RECT 1076.500 127.540 1076.760 127.800 ;
      LAYER met2 ;
        RECT 771.470 216.650 771.750 220.000 ;
        RECT 771.470 216.510 772.640 216.650 ;
        RECT 771.470 216.000 771.750 216.510 ;
        RECT 772.500 127.830 772.640 216.510 ;
        RECT 772.440 127.510 772.700 127.830 ;
        RECT 1076.500 127.510 1076.760 127.830 ;
        RECT 1076.560 16.730 1076.700 127.510 ;
        RECT 1076.560 16.590 1079.460 16.730 ;
        RECT 1079.320 2.400 1079.460 16.590 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 789.430 200.500 789.750 200.560 ;
        RECT 793.110 200.500 793.430 200.560 ;
        RECT 789.430 200.360 793.430 200.500 ;
        RECT 789.430 200.300 789.750 200.360 ;
        RECT 793.110 200.300 793.430 200.360 ;
        RECT 793.110 134.540 793.430 134.600 ;
        RECT 1090.730 134.540 1091.050 134.600 ;
        RECT 793.110 134.400 1091.050 134.540 ;
        RECT 793.110 134.340 793.430 134.400 ;
        RECT 1090.730 134.340 1091.050 134.400 ;
        RECT 1090.730 17.580 1091.050 17.640 ;
        RECT 1096.710 17.580 1097.030 17.640 ;
        RECT 1090.730 17.440 1097.030 17.580 ;
        RECT 1090.730 17.380 1091.050 17.440 ;
        RECT 1096.710 17.380 1097.030 17.440 ;
      LAYER via ;
        RECT 789.460 200.300 789.720 200.560 ;
        RECT 793.140 200.300 793.400 200.560 ;
        RECT 793.140 134.340 793.400 134.600 ;
        RECT 1090.760 134.340 1091.020 134.600 ;
        RECT 1090.760 17.380 1091.020 17.640 ;
        RECT 1096.740 17.380 1097.000 17.640 ;
      LAYER met2 ;
        RECT 789.410 216.000 789.690 220.000 ;
        RECT 789.520 200.590 789.660 216.000 ;
        RECT 789.460 200.270 789.720 200.590 ;
        RECT 793.140 200.270 793.400 200.590 ;
        RECT 793.200 134.630 793.340 200.270 ;
        RECT 793.140 134.310 793.400 134.630 ;
        RECT 1090.760 134.310 1091.020 134.630 ;
        RECT 1090.820 17.670 1090.960 134.310 ;
        RECT 1090.760 17.350 1091.020 17.670 ;
        RECT 1096.740 17.350 1097.000 17.670 ;
        RECT 1096.800 2.400 1096.940 17.350 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 807.370 200.500 807.690 200.560 ;
        RECT 813.810 200.500 814.130 200.560 ;
        RECT 807.370 200.360 814.130 200.500 ;
        RECT 807.370 200.300 807.690 200.360 ;
        RECT 813.810 200.300 814.130 200.360 ;
        RECT 813.810 31.520 814.130 31.580 ;
        RECT 1114.650 31.520 1114.970 31.580 ;
        RECT 813.810 31.380 1114.970 31.520 ;
        RECT 813.810 31.320 814.130 31.380 ;
        RECT 1114.650 31.320 1114.970 31.380 ;
      LAYER via ;
        RECT 807.400 200.300 807.660 200.560 ;
        RECT 813.840 200.300 814.100 200.560 ;
        RECT 813.840 31.320 814.100 31.580 ;
        RECT 1114.680 31.320 1114.940 31.580 ;
      LAYER met2 ;
        RECT 807.350 216.000 807.630 220.000 ;
        RECT 807.460 200.590 807.600 216.000 ;
        RECT 807.400 200.270 807.660 200.590 ;
        RECT 813.840 200.270 814.100 200.590 ;
        RECT 813.900 31.610 814.040 200.270 ;
        RECT 813.840 31.290 814.100 31.610 ;
        RECT 1114.680 31.290 1114.940 31.610 ;
        RECT 1114.740 2.400 1114.880 31.290 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 141.340 827.930 141.400 ;
        RECT 1131.670 141.340 1131.990 141.400 ;
        RECT 827.610 141.200 1131.990 141.340 ;
        RECT 827.610 141.140 827.930 141.200 ;
        RECT 1131.670 141.140 1131.990 141.200 ;
      LAYER via ;
        RECT 827.640 141.140 827.900 141.400 ;
        RECT 1131.700 141.140 1131.960 141.400 ;
      LAYER met2 ;
        RECT 824.830 216.650 825.110 220.000 ;
        RECT 824.830 216.510 827.840 216.650 ;
        RECT 824.830 216.000 825.110 216.510 ;
        RECT 827.700 141.430 827.840 216.510 ;
        RECT 827.640 141.110 827.900 141.430 ;
        RECT 1131.700 141.110 1131.960 141.430 ;
        RECT 1131.760 16.730 1131.900 141.110 ;
        RECT 1131.760 16.590 1132.820 16.730 ;
        RECT 1132.680 2.400 1132.820 16.590 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 842.790 200.500 843.110 200.560 ;
        RECT 848.310 200.500 848.630 200.560 ;
        RECT 842.790 200.360 848.630 200.500 ;
        RECT 842.790 200.300 843.110 200.360 ;
        RECT 848.310 200.300 848.630 200.360 ;
        RECT 848.310 38.320 848.630 38.380 ;
        RECT 1150.530 38.320 1150.850 38.380 ;
        RECT 848.310 38.180 1150.850 38.320 ;
        RECT 848.310 38.120 848.630 38.180 ;
        RECT 1150.530 38.120 1150.850 38.180 ;
      LAYER via ;
        RECT 842.820 200.300 843.080 200.560 ;
        RECT 848.340 200.300 848.600 200.560 ;
        RECT 848.340 38.120 848.600 38.380 ;
        RECT 1150.560 38.120 1150.820 38.380 ;
      LAYER met2 ;
        RECT 842.770 216.000 843.050 220.000 ;
        RECT 842.880 200.590 843.020 216.000 ;
        RECT 842.820 200.270 843.080 200.590 ;
        RECT 848.340 200.270 848.600 200.590 ;
        RECT 848.400 38.410 848.540 200.270 ;
        RECT 848.340 38.090 848.600 38.410 ;
        RECT 1150.560 38.090 1150.820 38.410 ;
        RECT 1150.620 2.400 1150.760 38.090 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 360.250 200.500 360.570 200.560 ;
        RECT 365.310 200.500 365.630 200.560 ;
        RECT 360.250 200.360 365.630 200.500 ;
        RECT 360.250 200.300 360.570 200.360 ;
        RECT 365.310 200.300 365.630 200.360 ;
        RECT 365.310 93.060 365.630 93.120 ;
        RECT 662.930 93.060 663.250 93.120 ;
        RECT 365.310 92.920 663.250 93.060 ;
        RECT 365.310 92.860 365.630 92.920 ;
        RECT 662.930 92.860 663.250 92.920 ;
        RECT 662.930 20.300 663.250 20.360 ;
        RECT 668.910 20.300 669.230 20.360 ;
        RECT 662.930 20.160 669.230 20.300 ;
        RECT 662.930 20.100 663.250 20.160 ;
        RECT 668.910 20.100 669.230 20.160 ;
      LAYER via ;
        RECT 360.280 200.300 360.540 200.560 ;
        RECT 365.340 200.300 365.600 200.560 ;
        RECT 365.340 92.860 365.600 93.120 ;
        RECT 662.960 92.860 663.220 93.120 ;
        RECT 662.960 20.100 663.220 20.360 ;
        RECT 668.940 20.100 669.200 20.360 ;
      LAYER met2 ;
        RECT 360.230 216.000 360.510 220.000 ;
        RECT 360.340 200.590 360.480 216.000 ;
        RECT 360.280 200.270 360.540 200.590 ;
        RECT 365.340 200.270 365.600 200.590 ;
        RECT 365.400 93.150 365.540 200.270 ;
        RECT 365.340 92.830 365.600 93.150 ;
        RECT 662.960 92.830 663.220 93.150 ;
        RECT 663.020 20.390 663.160 92.830 ;
        RECT 662.960 20.070 663.220 20.390 ;
        RECT 668.940 20.070 669.200 20.390 ;
        RECT 669.000 2.400 669.140 20.070 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 44.780 862.430 44.840 ;
        RECT 1168.470 44.780 1168.790 44.840 ;
        RECT 862.110 44.640 1168.790 44.780 ;
        RECT 862.110 44.580 862.430 44.640 ;
        RECT 1168.470 44.580 1168.790 44.640 ;
      LAYER via ;
        RECT 862.140 44.580 862.400 44.840 ;
        RECT 1168.500 44.580 1168.760 44.840 ;
      LAYER met2 ;
        RECT 860.710 216.650 860.990 220.000 ;
        RECT 860.710 216.510 862.340 216.650 ;
        RECT 860.710 216.000 860.990 216.510 ;
        RECT 862.200 44.870 862.340 216.510 ;
        RECT 862.140 44.550 862.400 44.870 ;
        RECT 1168.500 44.550 1168.760 44.870 ;
        RECT 1168.560 2.400 1168.700 44.550 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 878.670 200.500 878.990 200.560 ;
        RECT 882.810 200.500 883.130 200.560 ;
        RECT 878.670 200.360 883.130 200.500 ;
        RECT 878.670 200.300 878.990 200.360 ;
        RECT 882.810 200.300 883.130 200.360 ;
        RECT 882.810 51.920 883.130 51.980 ;
        RECT 1180.430 51.920 1180.750 51.980 ;
        RECT 882.810 51.780 1180.750 51.920 ;
        RECT 882.810 51.720 883.130 51.780 ;
        RECT 1180.430 51.720 1180.750 51.780 ;
        RECT 1180.430 17.920 1180.750 17.980 ;
        RECT 1185.950 17.920 1186.270 17.980 ;
        RECT 1180.430 17.780 1186.270 17.920 ;
        RECT 1180.430 17.720 1180.750 17.780 ;
        RECT 1185.950 17.720 1186.270 17.780 ;
      LAYER via ;
        RECT 878.700 200.300 878.960 200.560 ;
        RECT 882.840 200.300 883.100 200.560 ;
        RECT 882.840 51.720 883.100 51.980 ;
        RECT 1180.460 51.720 1180.720 51.980 ;
        RECT 1180.460 17.720 1180.720 17.980 ;
        RECT 1185.980 17.720 1186.240 17.980 ;
      LAYER met2 ;
        RECT 878.650 216.000 878.930 220.000 ;
        RECT 878.760 200.590 878.900 216.000 ;
        RECT 878.700 200.270 878.960 200.590 ;
        RECT 882.840 200.270 883.100 200.590 ;
        RECT 882.900 52.010 883.040 200.270 ;
        RECT 882.840 51.690 883.100 52.010 ;
        RECT 1180.460 51.690 1180.720 52.010 ;
        RECT 1180.520 18.010 1180.660 51.690 ;
        RECT 1180.460 17.690 1180.720 18.010 ;
        RECT 1185.980 17.690 1186.240 18.010 ;
        RECT 1186.040 2.400 1186.180 17.690 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.150 58.720 896.470 58.780 ;
        RECT 1200.670 58.720 1200.990 58.780 ;
        RECT 896.150 58.580 1200.990 58.720 ;
        RECT 896.150 58.520 896.470 58.580 ;
        RECT 1200.670 58.520 1200.990 58.580 ;
      LAYER via ;
        RECT 896.180 58.520 896.440 58.780 ;
        RECT 1200.700 58.520 1200.960 58.780 ;
      LAYER met2 ;
        RECT 896.590 216.650 896.870 220.000 ;
        RECT 896.240 216.510 896.870 216.650 ;
        RECT 896.240 58.810 896.380 216.510 ;
        RECT 896.590 216.000 896.870 216.510 ;
        RECT 896.180 58.490 896.440 58.810 ;
        RECT 1200.700 58.490 1200.960 58.810 ;
        RECT 1200.760 16.730 1200.900 58.490 ;
        RECT 1200.760 16.590 1204.120 16.730 ;
        RECT 1203.980 2.400 1204.120 16.590 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 65.520 917.630 65.580 ;
        RECT 1221.830 65.520 1222.150 65.580 ;
        RECT 917.310 65.380 1222.150 65.520 ;
        RECT 917.310 65.320 917.630 65.380 ;
        RECT 1221.830 65.320 1222.150 65.380 ;
      LAYER via ;
        RECT 917.340 65.320 917.600 65.580 ;
        RECT 1221.860 65.320 1222.120 65.580 ;
      LAYER met2 ;
        RECT 914.530 216.650 914.810 220.000 ;
        RECT 914.530 216.510 917.540 216.650 ;
        RECT 914.530 216.000 914.810 216.510 ;
        RECT 917.400 65.610 917.540 216.510 ;
        RECT 917.340 65.290 917.600 65.610 ;
        RECT 1221.860 65.290 1222.120 65.610 ;
        RECT 1221.920 2.400 1222.060 65.290 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 932.490 200.500 932.810 200.560 ;
        RECT 938.010 200.500 938.330 200.560 ;
        RECT 932.490 200.360 938.330 200.500 ;
        RECT 932.490 200.300 932.810 200.360 ;
        RECT 938.010 200.300 938.330 200.360 ;
        RECT 938.010 72.320 938.330 72.380 ;
        RECT 1235.170 72.320 1235.490 72.380 ;
        RECT 938.010 72.180 1235.490 72.320 ;
        RECT 938.010 72.120 938.330 72.180 ;
        RECT 1235.170 72.120 1235.490 72.180 ;
      LAYER via ;
        RECT 932.520 200.300 932.780 200.560 ;
        RECT 938.040 200.300 938.300 200.560 ;
        RECT 938.040 72.120 938.300 72.380 ;
        RECT 1235.200 72.120 1235.460 72.380 ;
      LAYER met2 ;
        RECT 932.470 216.000 932.750 220.000 ;
        RECT 932.580 200.590 932.720 216.000 ;
        RECT 932.520 200.270 932.780 200.590 ;
        RECT 938.040 200.270 938.300 200.590 ;
        RECT 938.100 72.410 938.240 200.270 ;
        RECT 938.040 72.090 938.300 72.410 ;
        RECT 1235.200 72.090 1235.460 72.410 ;
        RECT 1235.260 16.730 1235.400 72.090 ;
        RECT 1235.260 16.590 1240.000 16.730 ;
        RECT 1239.860 2.400 1240.000 16.590 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 24.380 952.130 24.440 ;
        RECT 1257.250 24.380 1257.570 24.440 ;
        RECT 951.810 24.240 1257.570 24.380 ;
        RECT 951.810 24.180 952.130 24.240 ;
        RECT 1257.250 24.180 1257.570 24.240 ;
      LAYER via ;
        RECT 951.840 24.180 952.100 24.440 ;
        RECT 1257.280 24.180 1257.540 24.440 ;
      LAYER met2 ;
        RECT 950.410 216.650 950.690 220.000 ;
        RECT 950.410 216.510 952.040 216.650 ;
        RECT 950.410 216.000 950.690 216.510 ;
        RECT 951.900 24.470 952.040 216.510 ;
        RECT 951.840 24.150 952.100 24.470 ;
        RECT 1257.280 24.150 1257.540 24.470 ;
        RECT 1257.340 2.400 1257.480 24.150 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 967.910 200.500 968.230 200.560 ;
        RECT 972.510 200.500 972.830 200.560 ;
        RECT 967.910 200.360 972.830 200.500 ;
        RECT 967.910 200.300 968.230 200.360 ;
        RECT 972.510 200.300 972.830 200.360 ;
        RECT 972.510 79.460 972.830 79.520 ;
        RECT 1269.670 79.460 1269.990 79.520 ;
        RECT 972.510 79.320 1269.990 79.460 ;
        RECT 972.510 79.260 972.830 79.320 ;
        RECT 1269.670 79.260 1269.990 79.320 ;
      LAYER via ;
        RECT 967.940 200.300 968.200 200.560 ;
        RECT 972.540 200.300 972.800 200.560 ;
        RECT 972.540 79.260 972.800 79.520 ;
        RECT 1269.700 79.260 1269.960 79.520 ;
      LAYER met2 ;
        RECT 967.890 216.000 968.170 220.000 ;
        RECT 968.000 200.590 968.140 216.000 ;
        RECT 967.940 200.270 968.200 200.590 ;
        RECT 972.540 200.270 972.800 200.590 ;
        RECT 972.600 79.550 972.740 200.270 ;
        RECT 972.540 79.230 972.800 79.550 ;
        RECT 1269.700 79.230 1269.960 79.550 ;
        RECT 1269.760 16.730 1269.900 79.230 ;
        RECT 1269.760 16.590 1275.420 16.730 ;
        RECT 1275.280 2.400 1275.420 16.590 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 985.850 86.260 986.170 86.320 ;
        RECT 1290.370 86.260 1290.690 86.320 ;
        RECT 985.850 86.120 1290.690 86.260 ;
        RECT 985.850 86.060 986.170 86.120 ;
        RECT 1290.370 86.060 1290.690 86.120 ;
      LAYER via ;
        RECT 985.880 86.060 986.140 86.320 ;
        RECT 1290.400 86.060 1290.660 86.320 ;
      LAYER met2 ;
        RECT 985.830 216.000 986.110 220.000 ;
        RECT 985.940 86.350 986.080 216.000 ;
        RECT 985.880 86.030 986.140 86.350 ;
        RECT 1290.400 86.030 1290.660 86.350 ;
        RECT 1290.460 17.410 1290.600 86.030 ;
        RECT 1290.460 17.270 1293.360 17.410 ;
        RECT 1293.220 2.400 1293.360 17.270 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 93.060 1007.330 93.120 ;
        RECT 1311.530 93.060 1311.850 93.120 ;
        RECT 1007.010 92.920 1311.850 93.060 ;
        RECT 1007.010 92.860 1007.330 92.920 ;
        RECT 1311.530 92.860 1311.850 92.920 ;
      LAYER via ;
        RECT 1007.040 92.860 1007.300 93.120 ;
        RECT 1311.560 92.860 1311.820 93.120 ;
      LAYER met2 ;
        RECT 1003.770 216.650 1004.050 220.000 ;
        RECT 1003.770 216.510 1007.240 216.650 ;
        RECT 1003.770 216.000 1004.050 216.510 ;
        RECT 1007.100 93.150 1007.240 216.510 ;
        RECT 1007.040 92.830 1007.300 93.150 ;
        RECT 1311.560 92.830 1311.820 93.150 ;
        RECT 1311.620 17.410 1311.760 92.830 ;
        RECT 1311.160 17.270 1311.760 17.410 ;
        RECT 1311.160 2.400 1311.300 17.270 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.730 200.500 1022.050 200.560 ;
        RECT 1027.710 200.500 1028.030 200.560 ;
        RECT 1021.730 200.360 1028.030 200.500 ;
        RECT 1021.730 200.300 1022.050 200.360 ;
        RECT 1027.710 200.300 1028.030 200.360 ;
        RECT 1027.710 107.000 1028.030 107.060 ;
        RECT 1324.870 107.000 1325.190 107.060 ;
        RECT 1027.710 106.860 1325.190 107.000 ;
        RECT 1027.710 106.800 1028.030 106.860 ;
        RECT 1324.870 106.800 1325.190 106.860 ;
      LAYER via ;
        RECT 1021.760 200.300 1022.020 200.560 ;
        RECT 1027.740 200.300 1028.000 200.560 ;
        RECT 1027.740 106.800 1028.000 107.060 ;
        RECT 1324.900 106.800 1325.160 107.060 ;
      LAYER met2 ;
        RECT 1021.710 216.000 1021.990 220.000 ;
        RECT 1021.820 200.590 1021.960 216.000 ;
        RECT 1021.760 200.270 1022.020 200.590 ;
        RECT 1027.740 200.270 1028.000 200.590 ;
        RECT 1027.800 107.090 1027.940 200.270 ;
        RECT 1027.740 106.770 1028.000 107.090 ;
        RECT 1324.900 106.770 1325.160 107.090 ;
        RECT 1324.960 17.410 1325.100 106.770 ;
        RECT 1324.960 17.270 1329.240 17.410 ;
        RECT 1329.100 2.400 1329.240 17.270 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 379.110 99.860 379.430 99.920 ;
        RECT 683.170 99.860 683.490 99.920 ;
        RECT 379.110 99.720 683.490 99.860 ;
        RECT 379.110 99.660 379.430 99.720 ;
        RECT 683.170 99.660 683.490 99.720 ;
      LAYER via ;
        RECT 379.140 99.660 379.400 99.920 ;
        RECT 683.200 99.660 683.460 99.920 ;
      LAYER met2 ;
        RECT 378.170 216.650 378.450 220.000 ;
        RECT 378.170 216.510 379.340 216.650 ;
        RECT 378.170 216.000 378.450 216.510 ;
        RECT 379.200 99.950 379.340 216.510 ;
        RECT 379.140 99.630 379.400 99.950 ;
        RECT 683.200 99.630 683.460 99.950 ;
        RECT 683.260 16.730 683.400 99.630 ;
        RECT 683.260 16.590 686.620 16.730 ;
        RECT 686.480 2.400 686.620 16.590 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 99.860 1041.830 99.920 ;
        RECT 1345.570 99.860 1345.890 99.920 ;
        RECT 1041.510 99.720 1345.890 99.860 ;
        RECT 1041.510 99.660 1041.830 99.720 ;
        RECT 1345.570 99.660 1345.890 99.720 ;
      LAYER via ;
        RECT 1041.540 99.660 1041.800 99.920 ;
        RECT 1345.600 99.660 1345.860 99.920 ;
      LAYER met2 ;
        RECT 1039.650 216.650 1039.930 220.000 ;
        RECT 1039.650 216.510 1041.740 216.650 ;
        RECT 1039.650 216.000 1039.930 216.510 ;
        RECT 1041.600 99.950 1041.740 216.510 ;
        RECT 1041.540 99.630 1041.800 99.950 ;
        RECT 1345.600 99.630 1345.860 99.950 ;
        RECT 1345.660 17.410 1345.800 99.630 ;
        RECT 1345.660 17.270 1346.720 17.410 ;
        RECT 1346.580 2.400 1346.720 17.270 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1057.610 200.500 1057.930 200.560 ;
        RECT 1062.210 200.500 1062.530 200.560 ;
        RECT 1057.610 200.360 1062.530 200.500 ;
        RECT 1057.610 200.300 1057.930 200.360 ;
        RECT 1062.210 200.300 1062.530 200.360 ;
        RECT 1062.210 120.600 1062.530 120.660 ;
        RECT 1359.370 120.600 1359.690 120.660 ;
        RECT 1062.210 120.460 1359.690 120.600 ;
        RECT 1062.210 120.400 1062.530 120.460 ;
        RECT 1359.370 120.400 1359.690 120.460 ;
      LAYER via ;
        RECT 1057.640 200.300 1057.900 200.560 ;
        RECT 1062.240 200.300 1062.500 200.560 ;
        RECT 1062.240 120.400 1062.500 120.660 ;
        RECT 1359.400 120.400 1359.660 120.660 ;
      LAYER met2 ;
        RECT 1057.590 216.000 1057.870 220.000 ;
        RECT 1057.700 200.590 1057.840 216.000 ;
        RECT 1057.640 200.270 1057.900 200.590 ;
        RECT 1062.240 200.270 1062.500 200.590 ;
        RECT 1062.300 120.690 1062.440 200.270 ;
        RECT 1062.240 120.370 1062.500 120.690 ;
        RECT 1359.400 120.370 1359.660 120.690 ;
        RECT 1359.460 17.410 1359.600 120.370 ;
        RECT 1359.460 17.270 1364.660 17.410 ;
        RECT 1364.520 2.400 1364.660 17.270 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1075.550 113.800 1075.870 113.860 ;
        RECT 1380.070 113.800 1380.390 113.860 ;
        RECT 1075.550 113.660 1380.390 113.800 ;
        RECT 1075.550 113.600 1075.870 113.660 ;
        RECT 1380.070 113.600 1380.390 113.660 ;
      LAYER via ;
        RECT 1075.580 113.600 1075.840 113.860 ;
        RECT 1380.100 113.600 1380.360 113.860 ;
      LAYER met2 ;
        RECT 1075.530 216.000 1075.810 220.000 ;
        RECT 1075.640 113.890 1075.780 216.000 ;
        RECT 1075.580 113.570 1075.840 113.890 ;
        RECT 1380.100 113.570 1380.360 113.890 ;
        RECT 1380.160 17.410 1380.300 113.570 ;
        RECT 1380.160 17.270 1382.600 17.410 ;
        RECT 1382.460 2.400 1382.600 17.270 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1093.030 200.500 1093.350 200.560 ;
        RECT 1096.710 200.500 1097.030 200.560 ;
        RECT 1093.030 200.360 1097.030 200.500 ;
        RECT 1093.030 200.300 1093.350 200.360 ;
        RECT 1096.710 200.300 1097.030 200.360 ;
        RECT 1096.710 31.180 1097.030 31.240 ;
        RECT 1399.850 31.180 1400.170 31.240 ;
        RECT 1096.710 31.040 1400.170 31.180 ;
        RECT 1096.710 30.980 1097.030 31.040 ;
        RECT 1399.850 30.980 1400.170 31.040 ;
      LAYER via ;
        RECT 1093.060 200.300 1093.320 200.560 ;
        RECT 1096.740 200.300 1097.000 200.560 ;
        RECT 1096.740 30.980 1097.000 31.240 ;
        RECT 1399.880 30.980 1400.140 31.240 ;
      LAYER met2 ;
        RECT 1093.010 216.000 1093.290 220.000 ;
        RECT 1093.120 200.590 1093.260 216.000 ;
        RECT 1093.060 200.270 1093.320 200.590 ;
        RECT 1096.740 200.270 1097.000 200.590 ;
        RECT 1096.800 31.270 1096.940 200.270 ;
        RECT 1096.740 30.950 1097.000 31.270 ;
        RECT 1399.880 30.950 1400.140 31.270 ;
        RECT 1399.940 30.330 1400.080 30.950 ;
        RECT 1399.940 30.190 1400.540 30.330 ;
        RECT 1400.400 2.400 1400.540 30.190 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.970 200.500 1111.290 200.560 ;
        RECT 1117.410 200.500 1117.730 200.560 ;
        RECT 1110.970 200.360 1117.730 200.500 ;
        RECT 1110.970 200.300 1111.290 200.360 ;
        RECT 1117.410 200.300 1117.730 200.360 ;
        RECT 1117.410 37.980 1117.730 38.040 ;
        RECT 1418.250 37.980 1418.570 38.040 ;
        RECT 1117.410 37.840 1418.570 37.980 ;
        RECT 1117.410 37.780 1117.730 37.840 ;
        RECT 1418.250 37.780 1418.570 37.840 ;
      LAYER via ;
        RECT 1111.000 200.300 1111.260 200.560 ;
        RECT 1117.440 200.300 1117.700 200.560 ;
        RECT 1117.440 37.780 1117.700 38.040 ;
        RECT 1418.280 37.780 1418.540 38.040 ;
      LAYER met2 ;
        RECT 1110.950 216.000 1111.230 220.000 ;
        RECT 1111.060 200.590 1111.200 216.000 ;
        RECT 1111.000 200.270 1111.260 200.590 ;
        RECT 1117.440 200.270 1117.700 200.590 ;
        RECT 1117.500 38.070 1117.640 200.270 ;
        RECT 1117.440 37.750 1117.700 38.070 ;
        RECT 1418.280 37.750 1418.540 38.070 ;
        RECT 1418.340 2.400 1418.480 37.750 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 127.740 1131.530 127.800 ;
        RECT 1435.730 127.740 1436.050 127.800 ;
        RECT 1131.210 127.600 1436.050 127.740 ;
        RECT 1131.210 127.540 1131.530 127.600 ;
        RECT 1435.730 127.540 1436.050 127.600 ;
      LAYER via ;
        RECT 1131.240 127.540 1131.500 127.800 ;
        RECT 1435.760 127.540 1436.020 127.800 ;
      LAYER met2 ;
        RECT 1128.890 216.650 1129.170 220.000 ;
        RECT 1128.890 216.510 1131.440 216.650 ;
        RECT 1128.890 216.000 1129.170 216.510 ;
        RECT 1131.300 127.830 1131.440 216.510 ;
        RECT 1131.240 127.510 1131.500 127.830 ;
        RECT 1435.760 127.510 1436.020 127.830 ;
        RECT 1435.820 2.400 1435.960 127.510 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1146.850 200.500 1147.170 200.560 ;
        RECT 1151.910 200.500 1152.230 200.560 ;
        RECT 1146.850 200.360 1152.230 200.500 ;
        RECT 1146.850 200.300 1147.170 200.360 ;
        RECT 1151.910 200.300 1152.230 200.360 ;
        RECT 1151.910 45.120 1152.230 45.180 ;
        RECT 1453.670 45.120 1453.990 45.180 ;
        RECT 1151.910 44.980 1453.990 45.120 ;
        RECT 1151.910 44.920 1152.230 44.980 ;
        RECT 1453.670 44.920 1453.990 44.980 ;
      LAYER via ;
        RECT 1146.880 200.300 1147.140 200.560 ;
        RECT 1151.940 200.300 1152.200 200.560 ;
        RECT 1151.940 44.920 1152.200 45.180 ;
        RECT 1453.700 44.920 1453.960 45.180 ;
      LAYER met2 ;
        RECT 1146.830 216.000 1147.110 220.000 ;
        RECT 1146.940 200.590 1147.080 216.000 ;
        RECT 1146.880 200.270 1147.140 200.590 ;
        RECT 1151.940 200.270 1152.200 200.590 ;
        RECT 1152.000 45.210 1152.140 200.270 ;
        RECT 1151.940 44.890 1152.200 45.210 ;
        RECT 1453.700 44.890 1453.960 45.210 ;
        RECT 1453.760 2.400 1453.900 44.890 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 51.580 1166.030 51.640 ;
        RECT 1469.770 51.580 1470.090 51.640 ;
        RECT 1165.710 51.440 1470.090 51.580 ;
        RECT 1165.710 51.380 1166.030 51.440 ;
        RECT 1469.770 51.380 1470.090 51.440 ;
      LAYER via ;
        RECT 1165.740 51.380 1166.000 51.640 ;
        RECT 1469.800 51.380 1470.060 51.640 ;
      LAYER met2 ;
        RECT 1164.770 216.650 1165.050 220.000 ;
        RECT 1164.770 216.510 1165.940 216.650 ;
        RECT 1164.770 216.000 1165.050 216.510 ;
        RECT 1165.800 51.670 1165.940 216.510 ;
        RECT 1165.740 51.350 1166.000 51.670 ;
        RECT 1469.800 51.350 1470.060 51.670 ;
        RECT 1469.860 17.410 1470.000 51.350 ;
        RECT 1469.860 17.270 1471.840 17.410 ;
        RECT 1471.700 2.400 1471.840 17.270 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 134.540 1186.730 134.600 ;
        RECT 1484.030 134.540 1484.350 134.600 ;
        RECT 1186.410 134.400 1484.350 134.540 ;
        RECT 1186.410 134.340 1186.730 134.400 ;
        RECT 1484.030 134.340 1484.350 134.400 ;
      LAYER via ;
        RECT 1186.440 134.340 1186.700 134.600 ;
        RECT 1484.060 134.340 1484.320 134.600 ;
      LAYER met2 ;
        RECT 1182.710 216.650 1182.990 220.000 ;
        RECT 1182.710 216.510 1186.640 216.650 ;
        RECT 1182.710 216.000 1182.990 216.510 ;
        RECT 1186.500 134.630 1186.640 216.510 ;
        RECT 1186.440 134.310 1186.700 134.630 ;
        RECT 1484.060 134.310 1484.320 134.630 ;
        RECT 1484.120 16.730 1484.260 134.310 ;
        RECT 1484.120 16.590 1489.780 16.730 ;
        RECT 1489.640 2.400 1489.780 16.590 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.670 200.500 1200.990 200.560 ;
        RECT 1207.110 200.500 1207.430 200.560 ;
        RECT 1200.670 200.360 1207.430 200.500 ;
        RECT 1200.670 200.300 1200.990 200.360 ;
        RECT 1207.110 200.300 1207.430 200.360 ;
        RECT 1207.110 58.720 1207.430 58.780 ;
        RECT 1504.270 58.720 1504.590 58.780 ;
        RECT 1207.110 58.580 1504.590 58.720 ;
        RECT 1207.110 58.520 1207.430 58.580 ;
        RECT 1504.270 58.520 1504.590 58.580 ;
      LAYER via ;
        RECT 1200.700 200.300 1200.960 200.560 ;
        RECT 1207.140 200.300 1207.400 200.560 ;
        RECT 1207.140 58.520 1207.400 58.780 ;
        RECT 1504.300 58.520 1504.560 58.780 ;
      LAYER met2 ;
        RECT 1200.650 216.000 1200.930 220.000 ;
        RECT 1200.760 200.590 1200.900 216.000 ;
        RECT 1200.700 200.270 1200.960 200.590 ;
        RECT 1207.140 200.270 1207.400 200.590 ;
        RECT 1207.200 58.810 1207.340 200.270 ;
        RECT 1207.140 58.490 1207.400 58.810 ;
        RECT 1504.300 58.490 1504.560 58.810 ;
        RECT 1504.360 16.730 1504.500 58.490 ;
        RECT 1504.360 16.590 1507.260 16.730 ;
        RECT 1507.120 2.400 1507.260 16.590 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 399.810 107.000 400.130 107.060 ;
        RECT 703.870 107.000 704.190 107.060 ;
        RECT 399.810 106.860 704.190 107.000 ;
        RECT 399.810 106.800 400.130 106.860 ;
        RECT 703.870 106.800 704.190 106.860 ;
      LAYER via ;
        RECT 399.840 106.800 400.100 107.060 ;
        RECT 703.900 106.800 704.160 107.060 ;
      LAYER met2 ;
        RECT 396.110 216.650 396.390 220.000 ;
        RECT 396.110 216.510 400.040 216.650 ;
        RECT 396.110 216.000 396.390 216.510 ;
        RECT 399.900 107.090 400.040 216.510 ;
        RECT 399.840 106.770 400.100 107.090 ;
        RECT 703.900 106.770 704.160 107.090 ;
        RECT 703.960 17.410 704.100 106.770 ;
        RECT 703.960 17.270 704.560 17.410 ;
        RECT 704.420 2.400 704.560 17.270 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 141.340 1221.230 141.400 ;
        RECT 1525.430 141.340 1525.750 141.400 ;
        RECT 1220.910 141.200 1525.750 141.340 ;
        RECT 1220.910 141.140 1221.230 141.200 ;
        RECT 1525.430 141.140 1525.750 141.200 ;
      LAYER via ;
        RECT 1220.940 141.140 1221.200 141.400 ;
        RECT 1525.460 141.140 1525.720 141.400 ;
      LAYER met2 ;
        RECT 1218.130 216.650 1218.410 220.000 ;
        RECT 1218.130 216.510 1221.140 216.650 ;
        RECT 1218.130 216.000 1218.410 216.510 ;
        RECT 1221.000 141.430 1221.140 216.510 ;
        RECT 1220.940 141.110 1221.200 141.430 ;
        RECT 1525.460 141.110 1525.720 141.430 ;
        RECT 1525.520 7.890 1525.660 141.110 ;
        RECT 1525.060 7.750 1525.660 7.890 ;
        RECT 1525.060 2.400 1525.200 7.750 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1236.090 202.880 1236.410 202.940 ;
        RECT 1241.610 202.880 1241.930 202.940 ;
        RECT 1236.090 202.740 1241.930 202.880 ;
        RECT 1236.090 202.680 1236.410 202.740 ;
        RECT 1241.610 202.680 1241.930 202.740 ;
        RECT 1241.610 65.860 1241.930 65.920 ;
        RECT 1538.770 65.860 1539.090 65.920 ;
        RECT 1241.610 65.720 1539.090 65.860 ;
        RECT 1241.610 65.660 1241.930 65.720 ;
        RECT 1538.770 65.660 1539.090 65.720 ;
      LAYER via ;
        RECT 1236.120 202.680 1236.380 202.940 ;
        RECT 1241.640 202.680 1241.900 202.940 ;
        RECT 1241.640 65.660 1241.900 65.920 ;
        RECT 1538.800 65.660 1539.060 65.920 ;
      LAYER met2 ;
        RECT 1236.070 216.000 1236.350 220.000 ;
        RECT 1236.180 202.970 1236.320 216.000 ;
        RECT 1236.120 202.650 1236.380 202.970 ;
        RECT 1241.640 202.650 1241.900 202.970 ;
        RECT 1241.700 65.950 1241.840 202.650 ;
        RECT 1241.640 65.630 1241.900 65.950 ;
        RECT 1538.800 65.630 1539.060 65.950 ;
        RECT 1538.860 16.730 1539.000 65.630 ;
        RECT 1538.860 16.590 1543.140 16.730 ;
        RECT 1543.000 2.400 1543.140 16.590 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 72.320 1255.730 72.380 ;
        RECT 1559.470 72.320 1559.790 72.380 ;
        RECT 1255.410 72.180 1559.790 72.320 ;
        RECT 1255.410 72.120 1255.730 72.180 ;
        RECT 1559.470 72.120 1559.790 72.180 ;
      LAYER via ;
        RECT 1255.440 72.120 1255.700 72.380 ;
        RECT 1559.500 72.120 1559.760 72.380 ;
      LAYER met2 ;
        RECT 1254.010 216.650 1254.290 220.000 ;
        RECT 1254.010 216.510 1255.640 216.650 ;
        RECT 1254.010 216.000 1254.290 216.510 ;
        RECT 1255.500 72.410 1255.640 216.510 ;
        RECT 1255.440 72.090 1255.700 72.410 ;
        RECT 1559.500 72.090 1559.760 72.410 ;
        RECT 1559.560 16.730 1559.700 72.090 ;
        RECT 1559.560 16.590 1561.080 16.730 ;
        RECT 1560.940 2.400 1561.080 16.590 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1271.970 200.500 1272.290 200.560 ;
        RECT 1276.110 200.500 1276.430 200.560 ;
        RECT 1271.970 200.360 1276.430 200.500 ;
        RECT 1271.970 200.300 1272.290 200.360 ;
        RECT 1276.110 200.300 1276.430 200.360 ;
        RECT 1276.110 24.720 1276.430 24.780 ;
        RECT 1578.790 24.720 1579.110 24.780 ;
        RECT 1276.110 24.580 1579.110 24.720 ;
        RECT 1276.110 24.520 1276.430 24.580 ;
        RECT 1578.790 24.520 1579.110 24.580 ;
      LAYER via ;
        RECT 1272.000 200.300 1272.260 200.560 ;
        RECT 1276.140 200.300 1276.400 200.560 ;
        RECT 1276.140 24.520 1276.400 24.780 ;
        RECT 1578.820 24.520 1579.080 24.780 ;
      LAYER met2 ;
        RECT 1271.950 216.000 1272.230 220.000 ;
        RECT 1272.060 200.590 1272.200 216.000 ;
        RECT 1272.000 200.270 1272.260 200.590 ;
        RECT 1276.140 200.270 1276.400 200.590 ;
        RECT 1276.200 24.810 1276.340 200.270 ;
        RECT 1276.140 24.490 1276.400 24.810 ;
        RECT 1578.820 24.490 1579.080 24.810 ;
        RECT 1578.880 2.400 1579.020 24.490 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.450 79.460 1289.770 79.520 ;
        RECT 1593.970 79.460 1594.290 79.520 ;
        RECT 1289.450 79.320 1594.290 79.460 ;
        RECT 1289.450 79.260 1289.770 79.320 ;
        RECT 1593.970 79.260 1594.290 79.320 ;
      LAYER via ;
        RECT 1289.480 79.260 1289.740 79.520 ;
        RECT 1594.000 79.260 1594.260 79.520 ;
      LAYER met2 ;
        RECT 1289.890 216.650 1290.170 220.000 ;
        RECT 1289.540 216.510 1290.170 216.650 ;
        RECT 1289.540 79.550 1289.680 216.510 ;
        RECT 1289.890 216.000 1290.170 216.510 ;
        RECT 1289.480 79.230 1289.740 79.550 ;
        RECT 1594.000 79.230 1594.260 79.550 ;
        RECT 1594.060 16.730 1594.200 79.230 ;
        RECT 1594.060 16.590 1596.500 16.730 ;
        RECT 1596.360 2.400 1596.500 16.590 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 86.260 1310.930 86.320 ;
        RECT 1608.230 86.260 1608.550 86.320 ;
        RECT 1310.610 86.120 1608.550 86.260 ;
        RECT 1310.610 86.060 1310.930 86.120 ;
        RECT 1608.230 86.060 1608.550 86.120 ;
        RECT 1608.230 17.920 1608.550 17.980 ;
        RECT 1614.210 17.920 1614.530 17.980 ;
        RECT 1608.230 17.780 1614.530 17.920 ;
        RECT 1608.230 17.720 1608.550 17.780 ;
        RECT 1614.210 17.720 1614.530 17.780 ;
      LAYER via ;
        RECT 1310.640 86.060 1310.900 86.320 ;
        RECT 1608.260 86.060 1608.520 86.320 ;
        RECT 1608.260 17.720 1608.520 17.980 ;
        RECT 1614.240 17.720 1614.500 17.980 ;
      LAYER met2 ;
        RECT 1307.830 216.650 1308.110 220.000 ;
        RECT 1307.830 216.510 1310.840 216.650 ;
        RECT 1307.830 216.000 1308.110 216.510 ;
        RECT 1310.700 86.350 1310.840 216.510 ;
        RECT 1310.640 86.030 1310.900 86.350 ;
        RECT 1608.260 86.030 1608.520 86.350 ;
        RECT 1608.320 18.010 1608.460 86.030 ;
        RECT 1608.260 17.690 1608.520 18.010 ;
        RECT 1614.240 17.690 1614.500 18.010 ;
        RECT 1614.300 2.400 1614.440 17.690 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1325.790 200.500 1326.110 200.560 ;
        RECT 1331.310 200.500 1331.630 200.560 ;
        RECT 1325.790 200.360 1331.630 200.500 ;
        RECT 1325.790 200.300 1326.110 200.360 ;
        RECT 1331.310 200.300 1331.630 200.360 ;
        RECT 1331.310 93.060 1331.630 93.120 ;
        RECT 1628.470 93.060 1628.790 93.120 ;
        RECT 1331.310 92.920 1628.790 93.060 ;
        RECT 1331.310 92.860 1331.630 92.920 ;
        RECT 1628.470 92.860 1628.790 92.920 ;
      LAYER via ;
        RECT 1325.820 200.300 1326.080 200.560 ;
        RECT 1331.340 200.300 1331.600 200.560 ;
        RECT 1331.340 92.860 1331.600 93.120 ;
        RECT 1628.500 92.860 1628.760 93.120 ;
      LAYER met2 ;
        RECT 1325.770 216.000 1326.050 220.000 ;
        RECT 1325.880 200.590 1326.020 216.000 ;
        RECT 1325.820 200.270 1326.080 200.590 ;
        RECT 1331.340 200.270 1331.600 200.590 ;
        RECT 1331.400 93.150 1331.540 200.270 ;
        RECT 1331.340 92.830 1331.600 93.150 ;
        RECT 1628.500 92.830 1628.760 93.150 ;
        RECT 1628.560 16.730 1628.700 92.830 ;
        RECT 1628.560 16.590 1632.380 16.730 ;
        RECT 1632.240 2.400 1632.380 16.590 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 107.000 1345.430 107.060 ;
        RECT 1649.170 107.000 1649.490 107.060 ;
        RECT 1345.110 106.860 1649.490 107.000 ;
        RECT 1345.110 106.800 1345.430 106.860 ;
        RECT 1649.170 106.800 1649.490 106.860 ;
      LAYER via ;
        RECT 1345.140 106.800 1345.400 107.060 ;
        RECT 1649.200 106.800 1649.460 107.060 ;
      LAYER met2 ;
        RECT 1343.250 216.650 1343.530 220.000 ;
        RECT 1343.250 216.510 1345.340 216.650 ;
        RECT 1343.250 216.000 1343.530 216.510 ;
        RECT 1345.200 107.090 1345.340 216.510 ;
        RECT 1345.140 106.770 1345.400 107.090 ;
        RECT 1649.200 106.770 1649.460 107.090 ;
        RECT 1649.260 16.730 1649.400 106.770 ;
        RECT 1649.260 16.590 1650.320 16.730 ;
        RECT 1650.180 2.400 1650.320 16.590 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.210 206.280 1361.530 206.340 ;
        RECT 1365.810 206.280 1366.130 206.340 ;
        RECT 1361.210 206.140 1366.130 206.280 ;
        RECT 1361.210 206.080 1361.530 206.140 ;
        RECT 1365.810 206.080 1366.130 206.140 ;
        RECT 1365.810 99.860 1366.130 99.920 ;
        RECT 1662.970 99.860 1663.290 99.920 ;
        RECT 1365.810 99.720 1663.290 99.860 ;
        RECT 1365.810 99.660 1366.130 99.720 ;
        RECT 1662.970 99.660 1663.290 99.720 ;
      LAYER via ;
        RECT 1361.240 206.080 1361.500 206.340 ;
        RECT 1365.840 206.080 1366.100 206.340 ;
        RECT 1365.840 99.660 1366.100 99.920 ;
        RECT 1663.000 99.660 1663.260 99.920 ;
      LAYER met2 ;
        RECT 1361.190 216.000 1361.470 220.000 ;
        RECT 1361.300 206.370 1361.440 216.000 ;
        RECT 1361.240 206.050 1361.500 206.370 ;
        RECT 1365.840 206.050 1366.100 206.370 ;
        RECT 1365.900 99.950 1366.040 206.050 ;
        RECT 1365.840 99.630 1366.100 99.950 ;
        RECT 1663.000 99.630 1663.260 99.950 ;
        RECT 1663.060 16.730 1663.200 99.630 ;
        RECT 1663.060 16.590 1668.260 16.730 ;
        RECT 1668.120 2.400 1668.260 16.590 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.610 120.600 1379.930 120.660 ;
        RECT 1683.670 120.600 1683.990 120.660 ;
        RECT 1379.610 120.460 1683.990 120.600 ;
        RECT 1379.610 120.400 1379.930 120.460 ;
        RECT 1683.670 120.400 1683.990 120.460 ;
      LAYER via ;
        RECT 1379.640 120.400 1379.900 120.660 ;
        RECT 1683.700 120.400 1683.960 120.660 ;
      LAYER met2 ;
        RECT 1379.130 216.650 1379.410 220.000 ;
        RECT 1379.130 216.510 1379.840 216.650 ;
        RECT 1379.130 216.000 1379.410 216.510 ;
        RECT 1379.700 120.690 1379.840 216.510 ;
        RECT 1379.640 120.370 1379.900 120.690 ;
        RECT 1683.700 120.370 1683.960 120.690 ;
        RECT 1683.760 17.410 1683.900 120.370 ;
        RECT 1683.760 17.270 1685.740 17.410 ;
        RECT 1685.600 2.400 1685.740 17.270 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 414.070 205.600 414.390 205.660 ;
        RECT 420.050 205.600 420.370 205.660 ;
        RECT 414.070 205.460 420.370 205.600 ;
        RECT 414.070 205.400 414.390 205.460 ;
        RECT 420.050 205.400 420.370 205.460 ;
        RECT 420.050 113.800 420.370 113.860 ;
        RECT 717.670 113.800 717.990 113.860 ;
        RECT 420.050 113.660 717.990 113.800 ;
        RECT 420.050 113.600 420.370 113.660 ;
        RECT 717.670 113.600 717.990 113.660 ;
      LAYER via ;
        RECT 414.100 205.400 414.360 205.660 ;
        RECT 420.080 205.400 420.340 205.660 ;
        RECT 420.080 113.600 420.340 113.860 ;
        RECT 717.700 113.600 717.960 113.860 ;
      LAYER met2 ;
        RECT 414.050 216.000 414.330 220.000 ;
        RECT 414.160 205.690 414.300 216.000 ;
        RECT 414.100 205.370 414.360 205.690 ;
        RECT 420.080 205.370 420.340 205.690 ;
        RECT 420.140 113.890 420.280 205.370 ;
        RECT 420.080 113.570 420.340 113.890 ;
        RECT 717.700 113.570 717.960 113.890 ;
        RECT 717.760 16.730 717.900 113.570 ;
        RECT 717.760 16.590 722.500 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 30.840 1400.630 30.900 ;
        RECT 1703.450 30.840 1703.770 30.900 ;
        RECT 1400.310 30.700 1703.770 30.840 ;
        RECT 1400.310 30.640 1400.630 30.700 ;
        RECT 1703.450 30.640 1703.770 30.700 ;
      LAYER via ;
        RECT 1400.340 30.640 1400.600 30.900 ;
        RECT 1703.480 30.640 1703.740 30.900 ;
      LAYER met2 ;
        RECT 1397.070 216.650 1397.350 220.000 ;
        RECT 1397.070 216.510 1400.540 216.650 ;
        RECT 1397.070 216.000 1397.350 216.510 ;
        RECT 1400.400 30.930 1400.540 216.510 ;
        RECT 1400.340 30.610 1400.600 30.930 ;
        RECT 1703.480 30.610 1703.740 30.930 ;
        RECT 1703.540 2.400 1703.680 30.610 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1415.030 201.860 1415.350 201.920 ;
        RECT 1421.010 201.860 1421.330 201.920 ;
        RECT 1415.030 201.720 1421.330 201.860 ;
        RECT 1415.030 201.660 1415.350 201.720 ;
        RECT 1421.010 201.660 1421.330 201.720 ;
        RECT 1421.010 37.980 1421.330 38.040 ;
        RECT 1721.390 37.980 1721.710 38.040 ;
        RECT 1421.010 37.840 1721.710 37.980 ;
        RECT 1421.010 37.780 1421.330 37.840 ;
        RECT 1721.390 37.780 1721.710 37.840 ;
      LAYER via ;
        RECT 1415.060 201.660 1415.320 201.920 ;
        RECT 1421.040 201.660 1421.300 201.920 ;
        RECT 1421.040 37.780 1421.300 38.040 ;
        RECT 1721.420 37.780 1721.680 38.040 ;
      LAYER met2 ;
        RECT 1415.010 216.000 1415.290 220.000 ;
        RECT 1415.120 201.950 1415.260 216.000 ;
        RECT 1415.060 201.630 1415.320 201.950 ;
        RECT 1421.040 201.630 1421.300 201.950 ;
        RECT 1421.100 38.070 1421.240 201.630 ;
        RECT 1421.040 37.750 1421.300 38.070 ;
        RECT 1721.420 37.750 1721.680 38.070 ;
        RECT 1721.480 2.400 1721.620 37.750 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 113.800 1435.130 113.860 ;
        RECT 1739.330 113.800 1739.650 113.860 ;
        RECT 1434.810 113.660 1739.650 113.800 ;
        RECT 1434.810 113.600 1435.130 113.660 ;
        RECT 1739.330 113.600 1739.650 113.660 ;
      LAYER via ;
        RECT 1434.840 113.600 1435.100 113.860 ;
        RECT 1739.360 113.600 1739.620 113.860 ;
      LAYER met2 ;
        RECT 1432.950 216.650 1433.230 220.000 ;
        RECT 1432.950 216.510 1435.040 216.650 ;
        RECT 1432.950 216.000 1433.230 216.510 ;
        RECT 1434.900 113.890 1435.040 216.510 ;
        RECT 1434.840 113.570 1435.100 113.890 ;
        RECT 1739.360 113.570 1739.620 113.890 ;
        RECT 1739.420 2.400 1739.560 113.570 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1450.910 202.540 1451.230 202.600 ;
        RECT 1455.510 202.540 1455.830 202.600 ;
        RECT 1450.910 202.400 1455.830 202.540 ;
        RECT 1450.910 202.340 1451.230 202.400 ;
        RECT 1455.510 202.340 1455.830 202.400 ;
        RECT 1455.510 45.120 1455.830 45.180 ;
        RECT 1756.810 45.120 1757.130 45.180 ;
        RECT 1455.510 44.980 1757.130 45.120 ;
        RECT 1455.510 44.920 1455.830 44.980 ;
        RECT 1756.810 44.920 1757.130 44.980 ;
      LAYER via ;
        RECT 1450.940 202.340 1451.200 202.600 ;
        RECT 1455.540 202.340 1455.800 202.600 ;
        RECT 1455.540 44.920 1455.800 45.180 ;
        RECT 1756.840 44.920 1757.100 45.180 ;
      LAYER met2 ;
        RECT 1450.890 216.000 1451.170 220.000 ;
        RECT 1451.000 202.630 1451.140 216.000 ;
        RECT 1450.940 202.310 1451.200 202.630 ;
        RECT 1455.540 202.310 1455.800 202.630 ;
        RECT 1455.600 45.210 1455.740 202.310 ;
        RECT 1455.540 44.890 1455.800 45.210 ;
        RECT 1756.840 44.890 1757.100 45.210 ;
        RECT 1756.900 2.400 1757.040 44.890 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1468.850 127.740 1469.170 127.800 ;
        RECT 1773.370 127.740 1773.690 127.800 ;
        RECT 1468.850 127.600 1773.690 127.740 ;
        RECT 1468.850 127.540 1469.170 127.600 ;
        RECT 1773.370 127.540 1773.690 127.600 ;
      LAYER via ;
        RECT 1468.880 127.540 1469.140 127.800 ;
        RECT 1773.400 127.540 1773.660 127.800 ;
      LAYER met2 ;
        RECT 1468.370 216.650 1468.650 220.000 ;
        RECT 1468.370 216.510 1469.080 216.650 ;
        RECT 1468.370 216.000 1468.650 216.510 ;
        RECT 1468.940 127.830 1469.080 216.510 ;
        RECT 1468.880 127.510 1469.140 127.830 ;
        RECT 1773.400 127.510 1773.660 127.830 ;
        RECT 1773.460 16.730 1773.600 127.510 ;
        RECT 1773.460 16.590 1774.980 16.730 ;
        RECT 1774.840 2.400 1774.980 16.590 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 51.920 1490.330 51.980 ;
        RECT 1787.170 51.920 1787.490 51.980 ;
        RECT 1490.010 51.780 1787.490 51.920 ;
        RECT 1490.010 51.720 1490.330 51.780 ;
        RECT 1787.170 51.720 1787.490 51.780 ;
      LAYER via ;
        RECT 1490.040 51.720 1490.300 51.980 ;
        RECT 1787.200 51.720 1787.460 51.980 ;
      LAYER met2 ;
        RECT 1486.310 216.650 1486.590 220.000 ;
        RECT 1486.310 216.510 1490.240 216.650 ;
        RECT 1486.310 216.000 1486.590 216.510 ;
        RECT 1490.100 52.010 1490.240 216.510 ;
        RECT 1490.040 51.690 1490.300 52.010 ;
        RECT 1787.200 51.690 1787.460 52.010 ;
        RECT 1787.260 16.730 1787.400 51.690 ;
        RECT 1787.260 16.590 1792.920 16.730 ;
        RECT 1792.780 2.400 1792.920 16.590 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1504.270 202.540 1504.590 202.600 ;
        RECT 1510.710 202.540 1511.030 202.600 ;
        RECT 1504.270 202.400 1511.030 202.540 ;
        RECT 1504.270 202.340 1504.590 202.400 ;
        RECT 1510.710 202.340 1511.030 202.400 ;
        RECT 1510.710 58.720 1511.030 58.780 ;
        RECT 1807.870 58.720 1808.190 58.780 ;
        RECT 1510.710 58.580 1808.190 58.720 ;
        RECT 1510.710 58.520 1511.030 58.580 ;
        RECT 1807.870 58.520 1808.190 58.580 ;
      LAYER via ;
        RECT 1504.300 202.340 1504.560 202.600 ;
        RECT 1510.740 202.340 1511.000 202.600 ;
        RECT 1510.740 58.520 1511.000 58.780 ;
        RECT 1807.900 58.520 1808.160 58.780 ;
      LAYER met2 ;
        RECT 1504.250 216.000 1504.530 220.000 ;
        RECT 1504.360 202.630 1504.500 216.000 ;
        RECT 1504.300 202.310 1504.560 202.630 ;
        RECT 1510.740 202.310 1511.000 202.630 ;
        RECT 1510.800 58.810 1510.940 202.310 ;
        RECT 1510.740 58.490 1511.000 58.810 ;
        RECT 1807.900 58.490 1808.160 58.810 ;
        RECT 1807.960 16.730 1808.100 58.490 ;
        RECT 1807.960 16.590 1810.860 16.730 ;
        RECT 1810.720 2.400 1810.860 16.590 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 65.520 1524.830 65.580 ;
        RECT 1829.030 65.520 1829.350 65.580 ;
        RECT 1524.510 65.380 1829.350 65.520 ;
        RECT 1524.510 65.320 1524.830 65.380 ;
        RECT 1829.030 65.320 1829.350 65.380 ;
      LAYER via ;
        RECT 1524.540 65.320 1524.800 65.580 ;
        RECT 1829.060 65.320 1829.320 65.580 ;
      LAYER met2 ;
        RECT 1522.190 216.650 1522.470 220.000 ;
        RECT 1522.190 216.510 1524.740 216.650 ;
        RECT 1522.190 216.000 1522.470 216.510 ;
        RECT 1524.600 65.610 1524.740 216.510 ;
        RECT 1524.540 65.290 1524.800 65.610 ;
        RECT 1829.060 65.290 1829.320 65.610 ;
        RECT 1829.120 7.210 1829.260 65.290 ;
        RECT 1828.660 7.070 1829.260 7.210 ;
        RECT 1828.660 2.400 1828.800 7.070 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1540.150 200.500 1540.470 200.560 ;
        RECT 1545.210 200.500 1545.530 200.560 ;
        RECT 1540.150 200.360 1545.530 200.500 ;
        RECT 1540.150 200.300 1540.470 200.360 ;
        RECT 1545.210 200.300 1545.530 200.360 ;
        RECT 1545.210 72.660 1545.530 72.720 ;
        RECT 1842.370 72.660 1842.690 72.720 ;
        RECT 1545.210 72.520 1842.690 72.660 ;
        RECT 1545.210 72.460 1545.530 72.520 ;
        RECT 1842.370 72.460 1842.690 72.520 ;
      LAYER via ;
        RECT 1540.180 200.300 1540.440 200.560 ;
        RECT 1545.240 200.300 1545.500 200.560 ;
        RECT 1545.240 72.460 1545.500 72.720 ;
        RECT 1842.400 72.460 1842.660 72.720 ;
      LAYER met2 ;
        RECT 1540.130 216.000 1540.410 220.000 ;
        RECT 1540.240 200.590 1540.380 216.000 ;
        RECT 1540.180 200.270 1540.440 200.590 ;
        RECT 1545.240 200.270 1545.500 200.590 ;
        RECT 1545.300 72.750 1545.440 200.270 ;
        RECT 1545.240 72.430 1545.500 72.750 ;
        RECT 1842.400 72.430 1842.660 72.750 ;
        RECT 1842.460 16.730 1842.600 72.430 ;
        RECT 1842.460 16.590 1846.280 16.730 ;
        RECT 1846.140 2.400 1846.280 16.590 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 134.540 1559.330 134.600 ;
        RECT 1863.070 134.540 1863.390 134.600 ;
        RECT 1559.010 134.400 1863.390 134.540 ;
        RECT 1559.010 134.340 1559.330 134.400 ;
        RECT 1863.070 134.340 1863.390 134.400 ;
      LAYER via ;
        RECT 1559.040 134.340 1559.300 134.600 ;
        RECT 1863.100 134.340 1863.360 134.600 ;
      LAYER met2 ;
        RECT 1558.070 216.650 1558.350 220.000 ;
        RECT 1558.070 216.510 1559.240 216.650 ;
        RECT 1558.070 216.000 1558.350 216.510 ;
        RECT 1559.100 134.630 1559.240 216.510 ;
        RECT 1559.040 134.310 1559.300 134.630 ;
        RECT 1863.100 134.310 1863.360 134.630 ;
        RECT 1863.160 16.730 1863.300 134.310 ;
        RECT 1863.160 16.590 1864.220 16.730 ;
        RECT 1864.080 2.400 1864.220 16.590 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 434.310 120.600 434.630 120.660 ;
        RECT 738.370 120.600 738.690 120.660 ;
        RECT 434.310 120.460 738.690 120.600 ;
        RECT 434.310 120.400 434.630 120.460 ;
        RECT 738.370 120.400 738.690 120.460 ;
      LAYER via ;
        RECT 434.340 120.400 434.600 120.660 ;
        RECT 738.400 120.400 738.660 120.660 ;
      LAYER met2 ;
        RECT 431.990 216.650 432.270 220.000 ;
        RECT 431.990 216.510 434.540 216.650 ;
        RECT 431.990 216.000 432.270 216.510 ;
        RECT 434.400 120.690 434.540 216.510 ;
        RECT 434.340 120.370 434.600 120.690 ;
        RECT 738.400 120.370 738.660 120.690 ;
        RECT 738.460 16.730 738.600 120.370 ;
        RECT 738.460 16.590 740.440 16.730 ;
        RECT 740.300 2.400 740.440 16.590 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1576.030 200.500 1576.350 200.560 ;
        RECT 1579.710 200.500 1580.030 200.560 ;
        RECT 1576.030 200.360 1580.030 200.500 ;
        RECT 1576.030 200.300 1576.350 200.360 ;
        RECT 1579.710 200.300 1580.030 200.360 ;
        RECT 1579.710 79.800 1580.030 79.860 ;
        RECT 1876.870 79.800 1877.190 79.860 ;
        RECT 1579.710 79.660 1877.190 79.800 ;
        RECT 1579.710 79.600 1580.030 79.660 ;
        RECT 1876.870 79.600 1877.190 79.660 ;
        RECT 1876.870 2.960 1877.190 3.020 ;
        RECT 1881.930 2.960 1882.250 3.020 ;
        RECT 1876.870 2.820 1882.250 2.960 ;
        RECT 1876.870 2.760 1877.190 2.820 ;
        RECT 1881.930 2.760 1882.250 2.820 ;
      LAYER via ;
        RECT 1576.060 200.300 1576.320 200.560 ;
        RECT 1579.740 200.300 1580.000 200.560 ;
        RECT 1579.740 79.600 1580.000 79.860 ;
        RECT 1876.900 79.600 1877.160 79.860 ;
        RECT 1876.900 2.760 1877.160 3.020 ;
        RECT 1881.960 2.760 1882.220 3.020 ;
      LAYER met2 ;
        RECT 1576.010 216.000 1576.290 220.000 ;
        RECT 1576.120 200.590 1576.260 216.000 ;
        RECT 1576.060 200.270 1576.320 200.590 ;
        RECT 1579.740 200.270 1580.000 200.590 ;
        RECT 1579.800 79.890 1579.940 200.270 ;
        RECT 1579.740 79.570 1580.000 79.890 ;
        RECT 1876.900 79.570 1877.160 79.890 ;
        RECT 1876.960 3.050 1877.100 79.570 ;
        RECT 1876.900 2.730 1877.160 3.050 ;
        RECT 1881.960 2.730 1882.220 3.050 ;
        RECT 1882.020 2.400 1882.160 2.730 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 204.240 1593.830 204.300 ;
        RECT 1728.290 204.240 1728.610 204.300 ;
        RECT 1593.510 204.100 1728.610 204.240 ;
        RECT 1593.510 204.040 1593.830 204.100 ;
        RECT 1728.290 204.040 1728.610 204.100 ;
        RECT 1728.290 30.840 1728.610 30.900 ;
        RECT 1899.870 30.840 1900.190 30.900 ;
        RECT 1728.290 30.700 1900.190 30.840 ;
        RECT 1728.290 30.640 1728.610 30.700 ;
        RECT 1899.870 30.640 1900.190 30.700 ;
      LAYER via ;
        RECT 1593.540 204.040 1593.800 204.300 ;
        RECT 1728.320 204.040 1728.580 204.300 ;
        RECT 1728.320 30.640 1728.580 30.900 ;
        RECT 1899.900 30.640 1900.160 30.900 ;
      LAYER met2 ;
        RECT 1593.490 216.000 1593.770 220.000 ;
        RECT 1593.600 204.330 1593.740 216.000 ;
        RECT 1593.540 204.010 1593.800 204.330 ;
        RECT 1728.320 204.010 1728.580 204.330 ;
        RECT 1728.380 30.930 1728.520 204.010 ;
        RECT 1728.320 30.610 1728.580 30.930 ;
        RECT 1899.900 30.610 1900.160 30.930 ;
        RECT 1899.960 2.400 1900.100 30.610 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 86.260 1614.530 86.320 ;
        RECT 1911.830 86.260 1912.150 86.320 ;
        RECT 1614.210 86.120 1912.150 86.260 ;
        RECT 1614.210 86.060 1614.530 86.120 ;
        RECT 1911.830 86.060 1912.150 86.120 ;
        RECT 1911.830 17.580 1912.150 17.640 ;
        RECT 1917.810 17.580 1918.130 17.640 ;
        RECT 1911.830 17.440 1918.130 17.580 ;
        RECT 1911.830 17.380 1912.150 17.440 ;
        RECT 1917.810 17.380 1918.130 17.440 ;
      LAYER via ;
        RECT 1614.240 86.060 1614.500 86.320 ;
        RECT 1911.860 86.060 1912.120 86.320 ;
        RECT 1911.860 17.380 1912.120 17.640 ;
        RECT 1917.840 17.380 1918.100 17.640 ;
      LAYER met2 ;
        RECT 1611.430 216.650 1611.710 220.000 ;
        RECT 1611.430 216.510 1614.440 216.650 ;
        RECT 1611.430 216.000 1611.710 216.510 ;
        RECT 1614.300 86.350 1614.440 216.510 ;
        RECT 1614.240 86.030 1614.500 86.350 ;
        RECT 1911.860 86.030 1912.120 86.350 ;
        RECT 1911.920 17.670 1912.060 86.030 ;
        RECT 1911.860 17.350 1912.120 17.670 ;
        RECT 1917.840 17.350 1918.100 17.670 ;
        RECT 1917.900 2.400 1918.040 17.350 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1629.390 200.500 1629.710 200.560 ;
        RECT 1634.910 200.500 1635.230 200.560 ;
        RECT 1629.390 200.360 1635.230 200.500 ;
        RECT 1629.390 200.300 1629.710 200.360 ;
        RECT 1634.910 200.300 1635.230 200.360 ;
        RECT 1634.910 93.060 1635.230 93.120 ;
        RECT 1932.070 93.060 1932.390 93.120 ;
        RECT 1634.910 92.920 1932.390 93.060 ;
        RECT 1634.910 92.860 1635.230 92.920 ;
        RECT 1932.070 92.860 1932.390 92.920 ;
        RECT 1932.070 2.960 1932.390 3.020 ;
        RECT 1935.290 2.960 1935.610 3.020 ;
        RECT 1932.070 2.820 1935.610 2.960 ;
        RECT 1932.070 2.760 1932.390 2.820 ;
        RECT 1935.290 2.760 1935.610 2.820 ;
      LAYER via ;
        RECT 1629.420 200.300 1629.680 200.560 ;
        RECT 1634.940 200.300 1635.200 200.560 ;
        RECT 1634.940 92.860 1635.200 93.120 ;
        RECT 1932.100 92.860 1932.360 93.120 ;
        RECT 1932.100 2.760 1932.360 3.020 ;
        RECT 1935.320 2.760 1935.580 3.020 ;
      LAYER met2 ;
        RECT 1629.370 216.000 1629.650 220.000 ;
        RECT 1629.480 200.590 1629.620 216.000 ;
        RECT 1629.420 200.270 1629.680 200.590 ;
        RECT 1634.940 200.270 1635.200 200.590 ;
        RECT 1635.000 93.150 1635.140 200.270 ;
        RECT 1634.940 92.830 1635.200 93.150 ;
        RECT 1932.100 92.830 1932.360 93.150 ;
        RECT 1932.160 3.050 1932.300 92.830 ;
        RECT 1932.100 2.730 1932.360 3.050 ;
        RECT 1935.320 2.730 1935.580 3.050 ;
        RECT 1935.380 2.400 1935.520 2.730 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1952.845 48.365 1953.015 72.675 ;
      LAYER mcon ;
        RECT 1952.845 72.505 1953.015 72.675 ;
      LAYER met1 ;
        RECT 1648.710 141.340 1649.030 141.400 ;
        RECT 1952.770 141.340 1953.090 141.400 ;
        RECT 1648.710 141.200 1953.090 141.340 ;
        RECT 1648.710 141.140 1649.030 141.200 ;
        RECT 1952.770 141.140 1953.090 141.200 ;
        RECT 1952.770 72.660 1953.090 72.720 ;
        RECT 1952.575 72.520 1953.090 72.660 ;
        RECT 1952.770 72.460 1953.090 72.520 ;
        RECT 1952.785 48.520 1953.075 48.565 ;
        RECT 1953.230 48.520 1953.550 48.580 ;
        RECT 1952.785 48.380 1953.550 48.520 ;
        RECT 1952.785 48.335 1953.075 48.380 ;
        RECT 1953.230 48.320 1953.550 48.380 ;
      LAYER via ;
        RECT 1648.740 141.140 1649.000 141.400 ;
        RECT 1952.800 141.140 1953.060 141.400 ;
        RECT 1952.800 72.460 1953.060 72.720 ;
        RECT 1953.260 48.320 1953.520 48.580 ;
      LAYER met2 ;
        RECT 1647.310 216.650 1647.590 220.000 ;
        RECT 1647.310 216.510 1648.940 216.650 ;
        RECT 1647.310 216.000 1647.590 216.510 ;
        RECT 1648.800 141.430 1648.940 216.510 ;
        RECT 1648.740 141.110 1649.000 141.430 ;
        RECT 1952.800 141.110 1953.060 141.430 ;
        RECT 1952.860 72.750 1953.000 141.110 ;
        RECT 1952.800 72.430 1953.060 72.750 ;
        RECT 1953.260 48.290 1953.520 48.610 ;
        RECT 1953.320 2.400 1953.460 48.290 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1665.270 200.500 1665.590 200.560 ;
        RECT 1669.410 200.500 1669.730 200.560 ;
        RECT 1665.270 200.360 1669.730 200.500 ;
        RECT 1665.270 200.300 1665.590 200.360 ;
        RECT 1669.410 200.300 1669.730 200.360 ;
        RECT 1669.410 99.860 1669.730 99.920 ;
        RECT 1966.570 99.860 1966.890 99.920 ;
        RECT 1669.410 99.720 1966.890 99.860 ;
        RECT 1669.410 99.660 1669.730 99.720 ;
        RECT 1966.570 99.660 1966.890 99.720 ;
        RECT 1966.570 62.120 1966.890 62.180 ;
        RECT 1971.170 62.120 1971.490 62.180 ;
        RECT 1966.570 61.980 1971.490 62.120 ;
        RECT 1966.570 61.920 1966.890 61.980 ;
        RECT 1971.170 61.920 1971.490 61.980 ;
      LAYER via ;
        RECT 1665.300 200.300 1665.560 200.560 ;
        RECT 1669.440 200.300 1669.700 200.560 ;
        RECT 1669.440 99.660 1669.700 99.920 ;
        RECT 1966.600 99.660 1966.860 99.920 ;
        RECT 1966.600 61.920 1966.860 62.180 ;
        RECT 1971.200 61.920 1971.460 62.180 ;
      LAYER met2 ;
        RECT 1665.250 216.000 1665.530 220.000 ;
        RECT 1665.360 200.590 1665.500 216.000 ;
        RECT 1665.300 200.270 1665.560 200.590 ;
        RECT 1669.440 200.270 1669.700 200.590 ;
        RECT 1669.500 99.950 1669.640 200.270 ;
        RECT 1669.440 99.630 1669.700 99.950 ;
        RECT 1966.600 99.630 1966.860 99.950 ;
        RECT 1966.660 62.210 1966.800 99.630 ;
        RECT 1966.600 61.890 1966.860 62.210 ;
        RECT 1971.200 61.890 1971.460 62.210 ;
        RECT 1971.260 2.400 1971.400 61.890 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1682.750 107.000 1683.070 107.060 ;
        RECT 1987.270 107.000 1987.590 107.060 ;
        RECT 1682.750 106.860 1987.590 107.000 ;
        RECT 1682.750 106.800 1683.070 106.860 ;
        RECT 1987.270 106.800 1987.590 106.860 ;
        RECT 1987.730 61.780 1988.050 61.840 ;
        RECT 1989.110 61.780 1989.430 61.840 ;
        RECT 1987.730 61.640 1989.430 61.780 ;
        RECT 1987.730 61.580 1988.050 61.640 ;
        RECT 1989.110 61.580 1989.430 61.640 ;
        RECT 1989.110 47.980 1989.430 48.240 ;
        RECT 1989.200 47.560 1989.340 47.980 ;
        RECT 1989.110 47.300 1989.430 47.560 ;
      LAYER via ;
        RECT 1682.780 106.800 1683.040 107.060 ;
        RECT 1987.300 106.800 1987.560 107.060 ;
        RECT 1987.760 61.580 1988.020 61.840 ;
        RECT 1989.140 61.580 1989.400 61.840 ;
        RECT 1989.140 47.980 1989.400 48.240 ;
        RECT 1989.140 47.300 1989.400 47.560 ;
      LAYER met2 ;
        RECT 1683.190 216.650 1683.470 220.000 ;
        RECT 1682.840 216.510 1683.470 216.650 ;
        RECT 1682.840 107.090 1682.980 216.510 ;
        RECT 1683.190 216.000 1683.470 216.510 ;
        RECT 1682.780 106.770 1683.040 107.090 ;
        RECT 1987.300 106.770 1987.560 107.090 ;
        RECT 1987.360 72.490 1987.500 106.770 ;
        RECT 1987.360 72.350 1987.960 72.490 ;
        RECT 1987.820 61.870 1987.960 72.350 ;
        RECT 1987.760 61.550 1988.020 61.870 ;
        RECT 1989.140 61.550 1989.400 61.870 ;
        RECT 1989.200 48.270 1989.340 61.550 ;
        RECT 1989.140 47.950 1989.400 48.270 ;
        RECT 1989.140 47.270 1989.400 47.590 ;
        RECT 1989.200 2.400 1989.340 47.270 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 38.320 1704.230 38.380 ;
        RECT 2006.590 38.320 2006.910 38.380 ;
        RECT 1703.910 38.180 2006.910 38.320 ;
        RECT 1703.910 38.120 1704.230 38.180 ;
        RECT 2006.590 38.120 2006.910 38.180 ;
      LAYER via ;
        RECT 1703.940 38.120 1704.200 38.380 ;
        RECT 2006.620 38.120 2006.880 38.380 ;
      LAYER met2 ;
        RECT 1701.130 216.650 1701.410 220.000 ;
        RECT 1701.130 216.510 1704.140 216.650 ;
        RECT 1701.130 216.000 1701.410 216.510 ;
        RECT 1704.000 38.410 1704.140 216.510 ;
        RECT 1703.940 38.090 1704.200 38.410 ;
        RECT 2006.620 38.090 2006.880 38.410 ;
        RECT 2006.680 2.400 2006.820 38.090 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1718.630 200.500 1718.950 200.560 ;
        RECT 1724.150 200.500 1724.470 200.560 ;
        RECT 1718.630 200.360 1724.470 200.500 ;
        RECT 1718.630 200.300 1718.950 200.360 ;
        RECT 1724.150 200.300 1724.470 200.360 ;
        RECT 1724.150 120.600 1724.470 120.660 ;
        RECT 2021.770 120.600 2022.090 120.660 ;
        RECT 1724.150 120.460 2022.090 120.600 ;
        RECT 1724.150 120.400 1724.470 120.460 ;
        RECT 2021.770 120.400 2022.090 120.460 ;
        RECT 2021.770 62.120 2022.090 62.180 ;
        RECT 2024.530 62.120 2024.850 62.180 ;
        RECT 2021.770 61.980 2024.850 62.120 ;
        RECT 2021.770 61.920 2022.090 61.980 ;
        RECT 2024.530 61.920 2024.850 61.980 ;
      LAYER via ;
        RECT 1718.660 200.300 1718.920 200.560 ;
        RECT 1724.180 200.300 1724.440 200.560 ;
        RECT 1724.180 120.400 1724.440 120.660 ;
        RECT 2021.800 120.400 2022.060 120.660 ;
        RECT 2021.800 61.920 2022.060 62.180 ;
        RECT 2024.560 61.920 2024.820 62.180 ;
      LAYER met2 ;
        RECT 1718.610 216.000 1718.890 220.000 ;
        RECT 1718.720 200.590 1718.860 216.000 ;
        RECT 1718.660 200.270 1718.920 200.590 ;
        RECT 1724.180 200.270 1724.440 200.590 ;
        RECT 1724.240 120.690 1724.380 200.270 ;
        RECT 1724.180 120.370 1724.440 120.690 ;
        RECT 2021.800 120.370 2022.060 120.690 ;
        RECT 2021.860 62.210 2022.000 120.370 ;
        RECT 2021.800 61.890 2022.060 62.210 ;
        RECT 2024.560 61.890 2024.820 62.210 ;
        RECT 2024.620 2.400 2024.760 61.890 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1738.410 44.780 1738.730 44.840 ;
        RECT 2043.390 44.780 2043.710 44.840 ;
        RECT 1738.410 44.640 2043.710 44.780 ;
        RECT 1738.410 44.580 1738.730 44.640 ;
        RECT 2043.390 44.580 2043.710 44.640 ;
      LAYER via ;
        RECT 1738.440 44.580 1738.700 44.840 ;
        RECT 2043.420 44.580 2043.680 44.840 ;
      LAYER met2 ;
        RECT 1736.550 216.650 1736.830 220.000 ;
        RECT 1736.550 216.510 1738.640 216.650 ;
        RECT 1736.550 216.000 1736.830 216.510 ;
        RECT 1738.500 44.870 1738.640 216.510 ;
        RECT 1738.440 44.550 1738.700 44.870 ;
        RECT 2043.420 44.550 2043.680 44.870 ;
        RECT 2043.480 37.130 2043.620 44.550 ;
        RECT 2042.560 36.990 2043.620 37.130 ;
        RECT 2042.560 2.400 2042.700 36.990 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 449.490 202.880 449.810 202.940 ;
        RECT 455.010 202.880 455.330 202.940 ;
        RECT 449.490 202.740 455.330 202.880 ;
        RECT 449.490 202.680 449.810 202.740 ;
        RECT 455.010 202.680 455.330 202.740 ;
        RECT 455.010 127.740 455.330 127.800 ;
        RECT 752.630 127.740 752.950 127.800 ;
        RECT 455.010 127.600 752.950 127.740 ;
        RECT 455.010 127.540 455.330 127.600 ;
        RECT 752.630 127.540 752.950 127.600 ;
        RECT 752.630 17.920 752.950 17.980 ;
        RECT 757.690 17.920 758.010 17.980 ;
        RECT 752.630 17.780 758.010 17.920 ;
        RECT 752.630 17.720 752.950 17.780 ;
        RECT 757.690 17.720 758.010 17.780 ;
      LAYER via ;
        RECT 449.520 202.680 449.780 202.940 ;
        RECT 455.040 202.680 455.300 202.940 ;
        RECT 455.040 127.540 455.300 127.800 ;
        RECT 752.660 127.540 752.920 127.800 ;
        RECT 752.660 17.720 752.920 17.980 ;
        RECT 757.720 17.720 757.980 17.980 ;
      LAYER met2 ;
        RECT 449.470 216.000 449.750 220.000 ;
        RECT 449.580 202.970 449.720 216.000 ;
        RECT 449.520 202.650 449.780 202.970 ;
        RECT 455.040 202.650 455.300 202.970 ;
        RECT 455.100 127.830 455.240 202.650 ;
        RECT 455.040 127.510 455.300 127.830 ;
        RECT 752.660 127.510 752.920 127.830 ;
        RECT 752.720 18.010 752.860 127.510 ;
        RECT 752.660 17.690 752.920 18.010 ;
        RECT 757.720 17.690 757.980 18.010 ;
        RECT 757.780 2.400 757.920 17.690 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.510 200.500 1754.830 200.560 ;
        RECT 1759.110 200.500 1759.430 200.560 ;
        RECT 1754.510 200.360 1759.430 200.500 ;
        RECT 1754.510 200.300 1754.830 200.360 ;
        RECT 1759.110 200.300 1759.430 200.360 ;
        RECT 1759.110 113.800 1759.430 113.860 ;
        RECT 2056.270 113.800 2056.590 113.860 ;
        RECT 1759.110 113.660 2056.590 113.800 ;
        RECT 1759.110 113.600 1759.430 113.660 ;
        RECT 2056.270 113.600 2056.590 113.660 ;
        RECT 2056.270 14.180 2056.590 14.240 ;
        RECT 2056.270 14.040 2060.640 14.180 ;
        RECT 2056.270 13.980 2056.590 14.040 ;
        RECT 2060.500 13.900 2060.640 14.040 ;
        RECT 2060.410 13.640 2060.730 13.900 ;
      LAYER via ;
        RECT 1754.540 200.300 1754.800 200.560 ;
        RECT 1759.140 200.300 1759.400 200.560 ;
        RECT 1759.140 113.600 1759.400 113.860 ;
        RECT 2056.300 113.600 2056.560 113.860 ;
        RECT 2056.300 13.980 2056.560 14.240 ;
        RECT 2060.440 13.640 2060.700 13.900 ;
      LAYER met2 ;
        RECT 1754.490 216.000 1754.770 220.000 ;
        RECT 1754.600 200.590 1754.740 216.000 ;
        RECT 1754.540 200.270 1754.800 200.590 ;
        RECT 1759.140 200.270 1759.400 200.590 ;
        RECT 1759.200 113.890 1759.340 200.270 ;
        RECT 1759.140 113.570 1759.400 113.890 ;
        RECT 2056.300 113.570 2056.560 113.890 ;
        RECT 2056.360 14.270 2056.500 113.570 ;
        RECT 2056.300 13.950 2056.560 14.270 ;
        RECT 2060.440 13.610 2060.700 13.930 ;
        RECT 2060.500 2.400 2060.640 13.610 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.450 148.140 1772.770 148.200 ;
        RECT 2076.970 148.140 2077.290 148.200 ;
        RECT 1772.450 148.000 2077.290 148.140 ;
        RECT 1772.450 147.940 1772.770 148.000 ;
        RECT 2076.970 147.940 2077.290 148.000 ;
        RECT 2076.970 14.180 2077.290 14.240 ;
        RECT 2076.970 14.040 2078.580 14.180 ;
        RECT 2076.970 13.980 2077.290 14.040 ;
        RECT 2078.440 13.900 2078.580 14.040 ;
        RECT 2078.350 13.640 2078.670 13.900 ;
      LAYER via ;
        RECT 1772.480 147.940 1772.740 148.200 ;
        RECT 2077.000 147.940 2077.260 148.200 ;
        RECT 2077.000 13.980 2077.260 14.240 ;
        RECT 2078.380 13.640 2078.640 13.900 ;
      LAYER met2 ;
        RECT 1772.430 216.000 1772.710 220.000 ;
        RECT 1772.540 148.230 1772.680 216.000 ;
        RECT 1772.480 147.910 1772.740 148.230 ;
        RECT 2077.000 147.910 2077.260 148.230 ;
        RECT 2077.060 14.270 2077.200 147.910 ;
        RECT 2077.000 13.950 2077.260 14.270 ;
        RECT 2078.380 13.610 2078.640 13.930 ;
        RECT 2078.440 2.400 2078.580 13.610 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 25.060 1793.930 25.120 ;
        RECT 2095.830 25.060 2096.150 25.120 ;
        RECT 1793.610 24.920 2096.150 25.060 ;
        RECT 1793.610 24.860 1793.930 24.920 ;
        RECT 2095.830 24.860 2096.150 24.920 ;
      LAYER via ;
        RECT 1793.640 24.860 1793.900 25.120 ;
        RECT 2095.860 24.860 2096.120 25.120 ;
      LAYER met2 ;
        RECT 1790.370 216.650 1790.650 220.000 ;
        RECT 1790.370 216.510 1793.840 216.650 ;
        RECT 1790.370 216.000 1790.650 216.510 ;
        RECT 1793.700 25.150 1793.840 216.510 ;
        RECT 1793.640 24.830 1793.900 25.150 ;
        RECT 2095.860 24.830 2096.120 25.150 ;
        RECT 2095.920 2.400 2096.060 24.830 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1808.330 200.500 1808.650 200.560 ;
        RECT 1814.310 200.500 1814.630 200.560 ;
        RECT 1808.330 200.360 1814.630 200.500 ;
        RECT 1808.330 200.300 1808.650 200.360 ;
        RECT 1814.310 200.300 1814.630 200.360 ;
        RECT 1814.310 27.440 1814.630 27.500 ;
        RECT 2113.770 27.440 2114.090 27.500 ;
        RECT 1814.310 27.300 2114.090 27.440 ;
        RECT 1814.310 27.240 1814.630 27.300 ;
        RECT 2113.770 27.240 2114.090 27.300 ;
      LAYER via ;
        RECT 1808.360 200.300 1808.620 200.560 ;
        RECT 1814.340 200.300 1814.600 200.560 ;
        RECT 1814.340 27.240 1814.600 27.500 ;
        RECT 2113.800 27.240 2114.060 27.500 ;
      LAYER met2 ;
        RECT 1808.310 216.000 1808.590 220.000 ;
        RECT 1808.420 200.590 1808.560 216.000 ;
        RECT 1808.360 200.270 1808.620 200.590 ;
        RECT 1814.340 200.270 1814.600 200.590 ;
        RECT 1814.400 27.530 1814.540 200.270 ;
        RECT 1814.340 27.210 1814.600 27.530 ;
        RECT 2113.800 27.210 2114.060 27.530 ;
        RECT 2113.860 2.400 2114.000 27.210 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.110 27.100 1828.430 27.160 ;
        RECT 2131.710 27.100 2132.030 27.160 ;
        RECT 1828.110 26.960 2132.030 27.100 ;
        RECT 1828.110 26.900 1828.430 26.960 ;
        RECT 2131.710 26.900 2132.030 26.960 ;
      LAYER via ;
        RECT 1828.140 26.900 1828.400 27.160 ;
        RECT 2131.740 26.900 2132.000 27.160 ;
      LAYER met2 ;
        RECT 1826.250 216.650 1826.530 220.000 ;
        RECT 1826.250 216.510 1828.340 216.650 ;
        RECT 1826.250 216.000 1826.530 216.510 ;
        RECT 1828.200 27.190 1828.340 216.510 ;
        RECT 1828.140 26.870 1828.400 27.190 ;
        RECT 2131.740 26.870 2132.000 27.190 ;
        RECT 2131.800 2.400 2131.940 26.870 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1844.210 200.500 1844.530 200.560 ;
        RECT 1848.810 200.500 1849.130 200.560 ;
        RECT 1844.210 200.360 1849.130 200.500 ;
        RECT 1844.210 200.300 1844.530 200.360 ;
        RECT 1848.810 200.300 1849.130 200.360 ;
        RECT 1848.810 26.420 1849.130 26.480 ;
        RECT 2149.650 26.420 2149.970 26.480 ;
        RECT 1848.810 26.280 2149.970 26.420 ;
        RECT 1848.810 26.220 1849.130 26.280 ;
        RECT 2149.650 26.220 2149.970 26.280 ;
      LAYER via ;
        RECT 1844.240 200.300 1844.500 200.560 ;
        RECT 1848.840 200.300 1849.100 200.560 ;
        RECT 1848.840 26.220 1849.100 26.480 ;
        RECT 2149.680 26.220 2149.940 26.480 ;
      LAYER met2 ;
        RECT 1844.190 216.000 1844.470 220.000 ;
        RECT 1844.300 200.590 1844.440 216.000 ;
        RECT 1844.240 200.270 1844.500 200.590 ;
        RECT 1848.840 200.270 1849.100 200.590 ;
        RECT 1848.900 26.510 1849.040 200.270 ;
        RECT 1848.840 26.190 1849.100 26.510 ;
        RECT 2149.680 26.190 2149.940 26.510 ;
        RECT 2149.740 2.400 2149.880 26.190 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 24.380 1862.930 24.440 ;
        RECT 2167.590 24.380 2167.910 24.440 ;
        RECT 1862.610 24.240 2167.910 24.380 ;
        RECT 1862.610 24.180 1862.930 24.240 ;
        RECT 2167.590 24.180 2167.910 24.240 ;
      LAYER via ;
        RECT 1862.640 24.180 1862.900 24.440 ;
        RECT 2167.620 24.180 2167.880 24.440 ;
      LAYER met2 ;
        RECT 1861.670 216.650 1861.950 220.000 ;
        RECT 1861.670 216.510 1862.840 216.650 ;
        RECT 1861.670 216.000 1861.950 216.510 ;
        RECT 1862.700 24.470 1862.840 216.510 ;
        RECT 1862.640 24.150 1862.900 24.470 ;
        RECT 2167.620 24.150 2167.880 24.470 ;
        RECT 2167.680 2.400 2167.820 24.150 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1879.630 200.500 1879.950 200.560 ;
        RECT 1883.310 200.500 1883.630 200.560 ;
        RECT 1879.630 200.360 1883.630 200.500 ;
        RECT 1879.630 200.300 1879.950 200.360 ;
        RECT 1883.310 200.300 1883.630 200.360 ;
        RECT 1883.310 25.400 1883.630 25.460 ;
        RECT 2185.070 25.400 2185.390 25.460 ;
        RECT 1883.310 25.260 2185.390 25.400 ;
        RECT 1883.310 25.200 1883.630 25.260 ;
        RECT 2185.070 25.200 2185.390 25.260 ;
      LAYER via ;
        RECT 1879.660 200.300 1879.920 200.560 ;
        RECT 1883.340 200.300 1883.600 200.560 ;
        RECT 1883.340 25.200 1883.600 25.460 ;
        RECT 2185.100 25.200 2185.360 25.460 ;
      LAYER met2 ;
        RECT 1879.610 216.000 1879.890 220.000 ;
        RECT 1879.720 200.590 1879.860 216.000 ;
        RECT 1879.660 200.270 1879.920 200.590 ;
        RECT 1883.340 200.270 1883.600 200.590 ;
        RECT 1883.400 25.490 1883.540 200.270 ;
        RECT 1883.340 25.170 1883.600 25.490 ;
        RECT 2185.100 25.170 2185.360 25.490 ;
        RECT 2185.160 2.400 2185.300 25.170 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1897.570 200.500 1897.890 200.560 ;
        RECT 1904.010 200.500 1904.330 200.560 ;
        RECT 1897.570 200.360 1904.330 200.500 ;
        RECT 1897.570 200.300 1897.890 200.360 ;
        RECT 1904.010 200.300 1904.330 200.360 ;
        RECT 1904.010 26.760 1904.330 26.820 ;
        RECT 2203.010 26.760 2203.330 26.820 ;
        RECT 1904.010 26.620 2203.330 26.760 ;
        RECT 1904.010 26.560 1904.330 26.620 ;
        RECT 2203.010 26.560 2203.330 26.620 ;
      LAYER via ;
        RECT 1897.600 200.300 1897.860 200.560 ;
        RECT 1904.040 200.300 1904.300 200.560 ;
        RECT 1904.040 26.560 1904.300 26.820 ;
        RECT 2203.040 26.560 2203.300 26.820 ;
      LAYER met2 ;
        RECT 1897.550 216.000 1897.830 220.000 ;
        RECT 1897.660 200.590 1897.800 216.000 ;
        RECT 1897.600 200.270 1897.860 200.590 ;
        RECT 1904.040 200.270 1904.300 200.590 ;
        RECT 1904.100 26.850 1904.240 200.270 ;
        RECT 1904.040 26.530 1904.300 26.850 ;
        RECT 2203.040 26.530 2203.300 26.850 ;
        RECT 2203.100 2.400 2203.240 26.530 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1942.265 24.565 1942.435 25.755 ;
      LAYER mcon ;
        RECT 1942.265 25.585 1942.435 25.755 ;
      LAYER met1 ;
        RECT 1917.810 25.740 1918.130 25.800 ;
        RECT 1942.205 25.740 1942.495 25.785 ;
        RECT 1917.810 25.600 1942.495 25.740 ;
        RECT 1917.810 25.540 1918.130 25.600 ;
        RECT 1942.205 25.555 1942.495 25.600 ;
        RECT 1942.205 24.720 1942.495 24.765 ;
        RECT 2220.950 24.720 2221.270 24.780 ;
        RECT 1942.205 24.580 2221.270 24.720 ;
        RECT 1942.205 24.535 1942.495 24.580 ;
        RECT 2220.950 24.520 2221.270 24.580 ;
      LAYER via ;
        RECT 1917.840 25.540 1918.100 25.800 ;
        RECT 2220.980 24.520 2221.240 24.780 ;
      LAYER met2 ;
        RECT 1915.490 216.650 1915.770 220.000 ;
        RECT 1915.490 216.510 1918.040 216.650 ;
        RECT 1915.490 216.000 1915.770 216.510 ;
        RECT 1917.900 25.830 1918.040 216.510 ;
        RECT 1917.840 25.510 1918.100 25.830 ;
        RECT 2220.980 24.490 2221.240 24.810 ;
        RECT 2221.040 2.400 2221.180 24.490 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 468.810 134.540 469.130 134.600 ;
        RECT 772.870 134.540 773.190 134.600 ;
        RECT 468.810 134.400 773.190 134.540 ;
        RECT 468.810 134.340 469.130 134.400 ;
        RECT 772.870 134.340 773.190 134.400 ;
      LAYER via ;
        RECT 468.840 134.340 469.100 134.600 ;
        RECT 772.900 134.340 773.160 134.600 ;
      LAYER met2 ;
        RECT 467.410 216.650 467.690 220.000 ;
        RECT 467.410 216.510 469.040 216.650 ;
        RECT 467.410 216.000 467.690 216.510 ;
        RECT 468.900 134.630 469.040 216.510 ;
        RECT 468.840 134.310 469.100 134.630 ;
        RECT 772.900 134.310 773.160 134.630 ;
        RECT 772.960 16.730 773.100 134.310 ;
        RECT 772.960 16.590 775.860 16.730 ;
        RECT 775.720 2.400 775.860 16.590 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1933.450 200.500 1933.770 200.560 ;
        RECT 1938.510 200.500 1938.830 200.560 ;
        RECT 1933.450 200.360 1938.830 200.500 ;
        RECT 1933.450 200.300 1933.770 200.360 ;
        RECT 1938.510 200.300 1938.830 200.360 ;
        RECT 1938.510 26.080 1938.830 26.140 ;
        RECT 2238.890 26.080 2239.210 26.140 ;
        RECT 1938.510 25.940 2239.210 26.080 ;
        RECT 1938.510 25.880 1938.830 25.940 ;
        RECT 2238.890 25.880 2239.210 25.940 ;
      LAYER via ;
        RECT 1933.480 200.300 1933.740 200.560 ;
        RECT 1938.540 200.300 1938.800 200.560 ;
        RECT 1938.540 25.880 1938.800 26.140 ;
        RECT 2238.920 25.880 2239.180 26.140 ;
      LAYER met2 ;
        RECT 1933.430 216.000 1933.710 220.000 ;
        RECT 1933.540 200.590 1933.680 216.000 ;
        RECT 1933.480 200.270 1933.740 200.590 ;
        RECT 1938.540 200.270 1938.800 200.590 ;
        RECT 1938.600 26.170 1938.740 200.270 ;
        RECT 1938.540 25.850 1938.800 26.170 ;
        RECT 2238.920 25.850 2239.180 26.170 ;
        RECT 2238.980 2.400 2239.120 25.850 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2069.685 23.205 2069.855 24.055 ;
        RECT 2077.045 22.525 2077.215 23.715 ;
        RECT 2168.125 22.525 2168.295 24.395 ;
        RECT 2221.945 22.865 2222.115 23.715 ;
      LAYER mcon ;
        RECT 2168.125 24.225 2168.295 24.395 ;
        RECT 2069.685 23.885 2069.855 24.055 ;
        RECT 2077.045 23.545 2077.215 23.715 ;
        RECT 2221.945 23.545 2222.115 23.715 ;
      LAYER met1 ;
        RECT 2168.065 24.380 2168.355 24.425 ;
        RECT 2168.065 24.240 2197.720 24.380 ;
        RECT 2168.065 24.195 2168.355 24.240 ;
        RECT 2069.625 24.040 2069.915 24.085 ;
        RECT 2027.840 23.900 2069.915 24.040 ;
        RECT 1952.310 23.700 1952.630 23.760 ;
        RECT 1952.310 23.560 2000.840 23.700 ;
        RECT 1952.310 23.500 1952.630 23.560 ;
        RECT 2000.700 23.360 2000.840 23.560 ;
        RECT 2027.840 23.360 2027.980 23.900 ;
        RECT 2069.625 23.855 2069.915 23.900 ;
        RECT 2076.985 23.515 2077.275 23.745 ;
        RECT 2000.700 23.220 2027.980 23.360 ;
        RECT 2069.625 23.360 2069.915 23.405 ;
        RECT 2077.060 23.360 2077.200 23.515 ;
        RECT 2069.625 23.220 2077.200 23.360 ;
        RECT 2197.580 23.360 2197.720 24.240 ;
        RECT 2221.885 23.515 2222.175 23.745 ;
        RECT 2221.960 23.360 2222.100 23.515 ;
        RECT 2197.580 23.220 2222.100 23.360 ;
        RECT 2069.625 23.175 2069.915 23.220 ;
        RECT 2221.885 23.020 2222.175 23.065 ;
        RECT 2256.370 23.020 2256.690 23.080 ;
        RECT 2221.885 22.880 2256.690 23.020 ;
        RECT 2221.885 22.835 2222.175 22.880 ;
        RECT 2256.370 22.820 2256.690 22.880 ;
        RECT 2076.985 22.680 2077.275 22.725 ;
        RECT 2168.065 22.680 2168.355 22.725 ;
        RECT 2076.985 22.540 2168.355 22.680 ;
        RECT 2076.985 22.495 2077.275 22.540 ;
        RECT 2168.065 22.495 2168.355 22.540 ;
      LAYER via ;
        RECT 1952.340 23.500 1952.600 23.760 ;
        RECT 2256.400 22.820 2256.660 23.080 ;
      LAYER met2 ;
        RECT 1951.370 216.650 1951.650 220.000 ;
        RECT 1951.370 216.510 1952.540 216.650 ;
        RECT 1951.370 216.000 1951.650 216.510 ;
        RECT 1952.400 23.790 1952.540 216.510 ;
        RECT 1952.340 23.470 1952.600 23.790 ;
        RECT 2256.400 22.790 2256.660 23.110 ;
        RECT 2256.460 2.400 2256.600 22.790 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.010 25.740 1973.330 25.800 ;
        RECT 2274.310 25.740 2274.630 25.800 ;
        RECT 1973.010 25.600 2274.630 25.740 ;
        RECT 1973.010 25.540 1973.330 25.600 ;
        RECT 2274.310 25.540 2274.630 25.600 ;
      LAYER via ;
        RECT 1973.040 25.540 1973.300 25.800 ;
        RECT 2274.340 25.540 2274.600 25.800 ;
      LAYER met2 ;
        RECT 1969.310 216.650 1969.590 220.000 ;
        RECT 1969.310 216.510 1973.240 216.650 ;
        RECT 1969.310 216.000 1969.590 216.510 ;
        RECT 1973.100 25.830 1973.240 216.510 ;
        RECT 1973.040 25.510 1973.300 25.830 ;
        RECT 2274.340 25.510 2274.600 25.830 ;
        RECT 2274.400 2.400 2274.540 25.510 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.810 79.460 1987.130 79.520 ;
        RECT 2290.870 79.460 2291.190 79.520 ;
        RECT 1986.810 79.320 2291.190 79.460 ;
        RECT 1986.810 79.260 1987.130 79.320 ;
        RECT 2290.870 79.260 2291.190 79.320 ;
      LAYER via ;
        RECT 1986.840 79.260 1987.100 79.520 ;
        RECT 2290.900 79.260 2291.160 79.520 ;
      LAYER met2 ;
        RECT 1986.790 216.000 1987.070 220.000 ;
        RECT 1986.900 79.550 1987.040 216.000 ;
        RECT 1986.840 79.230 1987.100 79.550 ;
        RECT 2290.900 79.230 2291.160 79.550 ;
        RECT 2290.960 3.130 2291.100 79.230 ;
        RECT 2290.960 2.990 2292.020 3.130 ;
        RECT 2291.880 2.960 2292.020 2.990 ;
        RECT 2291.880 2.820 2292.480 2.960 ;
        RECT 2292.340 2.400 2292.480 2.820 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.510 86.600 2007.830 86.660 ;
        RECT 2304.670 86.600 2304.990 86.660 ;
        RECT 2007.510 86.460 2304.990 86.600 ;
        RECT 2007.510 86.400 2007.830 86.460 ;
        RECT 2304.670 86.400 2304.990 86.460 ;
        RECT 2305.130 2.960 2305.450 3.020 ;
        RECT 2310.190 2.960 2310.510 3.020 ;
        RECT 2305.130 2.820 2310.510 2.960 ;
        RECT 2305.130 2.760 2305.450 2.820 ;
        RECT 2310.190 2.760 2310.510 2.820 ;
      LAYER via ;
        RECT 2007.540 86.400 2007.800 86.660 ;
        RECT 2304.700 86.400 2304.960 86.660 ;
        RECT 2305.160 2.760 2305.420 3.020 ;
        RECT 2310.220 2.760 2310.480 3.020 ;
      LAYER met2 ;
        RECT 2004.730 216.650 2005.010 220.000 ;
        RECT 2004.730 216.510 2007.740 216.650 ;
        RECT 2004.730 216.000 2005.010 216.510 ;
        RECT 2007.600 86.690 2007.740 216.510 ;
        RECT 2007.540 86.370 2007.800 86.690 ;
        RECT 2304.700 86.370 2304.960 86.690 ;
        RECT 2304.760 20.810 2304.900 86.370 ;
        RECT 2304.760 20.670 2305.360 20.810 ;
        RECT 2305.220 3.050 2305.360 20.670 ;
        RECT 2305.160 2.730 2305.420 3.050 ;
        RECT 2310.220 2.730 2310.480 3.050 ;
        RECT 2310.280 2.400 2310.420 2.730 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2022.690 200.500 2023.010 200.560 ;
        RECT 2028.210 200.500 2028.530 200.560 ;
        RECT 2022.690 200.360 2028.530 200.500 ;
        RECT 2022.690 200.300 2023.010 200.360 ;
        RECT 2028.210 200.300 2028.530 200.360 ;
        RECT 2028.210 99.860 2028.530 99.920 ;
        RECT 2325.370 99.860 2325.690 99.920 ;
        RECT 2028.210 99.720 2325.690 99.860 ;
        RECT 2028.210 99.660 2028.530 99.720 ;
        RECT 2325.370 99.660 2325.690 99.720 ;
        RECT 2325.370 2.960 2325.690 3.020 ;
        RECT 2328.130 2.960 2328.450 3.020 ;
        RECT 2325.370 2.820 2328.450 2.960 ;
        RECT 2325.370 2.760 2325.690 2.820 ;
        RECT 2328.130 2.760 2328.450 2.820 ;
      LAYER via ;
        RECT 2022.720 200.300 2022.980 200.560 ;
        RECT 2028.240 200.300 2028.500 200.560 ;
        RECT 2028.240 99.660 2028.500 99.920 ;
        RECT 2325.400 99.660 2325.660 99.920 ;
        RECT 2325.400 2.760 2325.660 3.020 ;
        RECT 2328.160 2.760 2328.420 3.020 ;
      LAYER met2 ;
        RECT 2022.670 216.000 2022.950 220.000 ;
        RECT 2022.780 200.590 2022.920 216.000 ;
        RECT 2022.720 200.270 2022.980 200.590 ;
        RECT 2028.240 200.270 2028.500 200.590 ;
        RECT 2028.300 99.950 2028.440 200.270 ;
        RECT 2028.240 99.630 2028.500 99.950 ;
        RECT 2325.400 99.630 2325.660 99.950 ;
        RECT 2325.460 3.050 2325.600 99.630 ;
        RECT 2325.400 2.730 2325.660 3.050 ;
        RECT 2328.160 2.730 2328.420 3.050 ;
        RECT 2328.220 2.400 2328.360 2.730 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 93.060 2042.330 93.120 ;
        RECT 2339.170 93.060 2339.490 93.120 ;
        RECT 2042.010 92.920 2339.490 93.060 ;
        RECT 2042.010 92.860 2042.330 92.920 ;
        RECT 2339.170 92.860 2339.490 92.920 ;
        RECT 2339.170 17.920 2339.490 17.980 ;
        RECT 2345.610 17.920 2345.930 17.980 ;
        RECT 2339.170 17.780 2345.930 17.920 ;
        RECT 2339.170 17.720 2339.490 17.780 ;
        RECT 2345.610 17.720 2345.930 17.780 ;
      LAYER via ;
        RECT 2042.040 92.860 2042.300 93.120 ;
        RECT 2339.200 92.860 2339.460 93.120 ;
        RECT 2339.200 17.720 2339.460 17.980 ;
        RECT 2345.640 17.720 2345.900 17.980 ;
      LAYER met2 ;
        RECT 2040.610 216.650 2040.890 220.000 ;
        RECT 2040.610 216.510 2042.240 216.650 ;
        RECT 2040.610 216.000 2040.890 216.510 ;
        RECT 2042.100 93.150 2042.240 216.510 ;
        RECT 2042.040 92.830 2042.300 93.150 ;
        RECT 2339.200 92.830 2339.460 93.150 ;
        RECT 2339.260 18.010 2339.400 92.830 ;
        RECT 2339.200 17.690 2339.460 18.010 ;
        RECT 2345.640 17.690 2345.900 18.010 ;
        RECT 2345.700 2.400 2345.840 17.690 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2058.570 200.500 2058.890 200.560 ;
        RECT 2062.710 200.500 2063.030 200.560 ;
        RECT 2058.570 200.360 2063.030 200.500 ;
        RECT 2058.570 200.300 2058.890 200.360 ;
        RECT 2062.710 200.300 2063.030 200.360 ;
        RECT 2062.710 113.800 2063.030 113.860 ;
        RECT 2359.870 113.800 2360.190 113.860 ;
        RECT 2062.710 113.660 2360.190 113.800 ;
        RECT 2062.710 113.600 2063.030 113.660 ;
        RECT 2359.870 113.600 2360.190 113.660 ;
        RECT 2359.870 2.960 2360.190 3.020 ;
        RECT 2363.550 2.960 2363.870 3.020 ;
        RECT 2359.870 2.820 2363.870 2.960 ;
        RECT 2359.870 2.760 2360.190 2.820 ;
        RECT 2363.550 2.760 2363.870 2.820 ;
      LAYER via ;
        RECT 2058.600 200.300 2058.860 200.560 ;
        RECT 2062.740 200.300 2063.000 200.560 ;
        RECT 2062.740 113.600 2063.000 113.860 ;
        RECT 2359.900 113.600 2360.160 113.860 ;
        RECT 2359.900 2.760 2360.160 3.020 ;
        RECT 2363.580 2.760 2363.840 3.020 ;
      LAYER met2 ;
        RECT 2058.550 216.000 2058.830 220.000 ;
        RECT 2058.660 200.590 2058.800 216.000 ;
        RECT 2058.600 200.270 2058.860 200.590 ;
        RECT 2062.740 200.270 2063.000 200.590 ;
        RECT 2062.800 113.890 2062.940 200.270 ;
        RECT 2062.740 113.570 2063.000 113.890 ;
        RECT 2359.900 113.570 2360.160 113.890 ;
        RECT 2359.960 3.050 2360.100 113.570 ;
        RECT 2359.900 2.730 2360.160 3.050 ;
        RECT 2363.580 2.730 2363.840 3.050 ;
        RECT 2363.640 2.400 2363.780 2.730 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.050 182.820 2076.370 182.880 ;
        RECT 2380.570 182.820 2380.890 182.880 ;
        RECT 2076.050 182.680 2380.890 182.820 ;
        RECT 2076.050 182.620 2076.370 182.680 ;
        RECT 2380.570 182.620 2380.890 182.680 ;
      LAYER via ;
        RECT 2076.080 182.620 2076.340 182.880 ;
        RECT 2380.600 182.620 2380.860 182.880 ;
      LAYER met2 ;
        RECT 2076.490 216.650 2076.770 220.000 ;
        RECT 2076.140 216.510 2076.770 216.650 ;
        RECT 2076.140 182.910 2076.280 216.510 ;
        RECT 2076.490 216.000 2076.770 216.510 ;
        RECT 2076.080 182.590 2076.340 182.910 ;
        RECT 2380.600 182.590 2380.860 182.910 ;
        RECT 2380.660 3.130 2380.800 182.590 ;
        RECT 2380.660 2.990 2381.260 3.130 ;
        RECT 2381.120 2.960 2381.260 2.990 ;
        RECT 2381.120 2.820 2381.720 2.960 ;
        RECT 2381.580 2.400 2381.720 2.820 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2097.210 107.000 2097.530 107.060 ;
        RECT 2394.370 107.000 2394.690 107.060 ;
        RECT 2097.210 106.860 2394.690 107.000 ;
        RECT 2097.210 106.800 2097.530 106.860 ;
        RECT 2394.370 106.800 2394.690 106.860 ;
        RECT 2394.370 2.960 2394.690 3.020 ;
        RECT 2399.430 2.960 2399.750 3.020 ;
        RECT 2394.370 2.820 2399.750 2.960 ;
        RECT 2394.370 2.760 2394.690 2.820 ;
        RECT 2399.430 2.760 2399.750 2.820 ;
      LAYER via ;
        RECT 2097.240 106.800 2097.500 107.060 ;
        RECT 2394.400 106.800 2394.660 107.060 ;
        RECT 2394.400 2.760 2394.660 3.020 ;
        RECT 2399.460 2.760 2399.720 3.020 ;
      LAYER met2 ;
        RECT 2094.430 216.650 2094.710 220.000 ;
        RECT 2094.430 216.510 2097.440 216.650 ;
        RECT 2094.430 216.000 2094.710 216.510 ;
        RECT 2097.300 107.090 2097.440 216.510 ;
        RECT 2097.240 106.770 2097.500 107.090 ;
        RECT 2394.400 106.770 2394.660 107.090 ;
        RECT 2394.460 3.050 2394.600 106.770 ;
        RECT 2394.400 2.730 2394.660 3.050 ;
        RECT 2399.460 2.730 2399.720 3.050 ;
        RECT 2399.520 2.400 2399.660 2.730 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 485.370 200.500 485.690 200.560 ;
        RECT 489.510 200.500 489.830 200.560 ;
        RECT 485.370 200.360 489.830 200.500 ;
        RECT 485.370 200.300 485.690 200.360 ;
        RECT 489.510 200.300 489.830 200.360 ;
        RECT 489.510 141.340 489.830 141.400 ;
        RECT 794.030 141.340 794.350 141.400 ;
        RECT 489.510 141.200 794.350 141.340 ;
        RECT 489.510 141.140 489.830 141.200 ;
        RECT 794.030 141.140 794.350 141.200 ;
      LAYER via ;
        RECT 485.400 200.300 485.660 200.560 ;
        RECT 489.540 200.300 489.800 200.560 ;
        RECT 489.540 141.140 489.800 141.400 ;
        RECT 794.060 141.140 794.320 141.400 ;
      LAYER met2 ;
        RECT 485.350 216.000 485.630 220.000 ;
        RECT 485.460 200.590 485.600 216.000 ;
        RECT 485.400 200.270 485.660 200.590 ;
        RECT 489.540 200.270 489.800 200.590 ;
        RECT 489.600 141.430 489.740 200.270 ;
        RECT 489.540 141.110 489.800 141.430 ;
        RECT 794.060 141.110 794.320 141.430 ;
        RECT 794.120 7.890 794.260 141.110 ;
        RECT 793.660 7.750 794.260 7.890 ;
        RECT 793.660 2.400 793.800 7.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 330.350 200.500 330.670 200.560 ;
        RECT 334.490 200.500 334.810 200.560 ;
        RECT 330.350 200.360 334.810 200.500 ;
        RECT 330.350 200.300 330.670 200.360 ;
        RECT 334.490 200.300 334.810 200.360 ;
        RECT 334.490 79.460 334.810 79.520 ;
        RECT 634.870 79.460 635.190 79.520 ;
        RECT 334.490 79.320 635.190 79.460 ;
        RECT 334.490 79.260 334.810 79.320 ;
        RECT 634.870 79.260 635.190 79.320 ;
      LAYER via ;
        RECT 330.380 200.300 330.640 200.560 ;
        RECT 334.520 200.300 334.780 200.560 ;
        RECT 334.520 79.260 334.780 79.520 ;
        RECT 634.900 79.260 635.160 79.520 ;
      LAYER met2 ;
        RECT 330.330 216.000 330.610 220.000 ;
        RECT 330.440 200.590 330.580 216.000 ;
        RECT 330.380 200.270 330.640 200.590 ;
        RECT 334.520 200.270 334.780 200.590 ;
        RECT 334.580 79.550 334.720 200.270 ;
        RECT 334.520 79.230 334.780 79.550 ;
        RECT 634.900 79.230 635.160 79.550 ;
        RECT 634.960 17.410 635.100 79.230 ;
        RECT 634.960 17.270 639.240 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2117.450 120.600 2117.770 120.660 ;
        RECT 2421.970 120.600 2422.290 120.660 ;
        RECT 2117.450 120.460 2422.290 120.600 ;
        RECT 2117.450 120.400 2117.770 120.460 ;
        RECT 2421.970 120.400 2422.290 120.460 ;
      LAYER via ;
        RECT 2117.480 120.400 2117.740 120.660 ;
        RECT 2422.000 120.400 2422.260 120.660 ;
      LAYER met2 ;
        RECT 2117.890 216.650 2118.170 220.000 ;
        RECT 2117.540 216.510 2118.170 216.650 ;
        RECT 2117.540 120.690 2117.680 216.510 ;
        RECT 2117.890 216.000 2118.170 216.510 ;
        RECT 2117.480 120.370 2117.740 120.690 ;
        RECT 2422.000 120.370 2422.260 120.690 ;
        RECT 2422.060 17.410 2422.200 120.370 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.610 128.080 2138.930 128.140 ;
        RECT 2435.770 128.080 2436.090 128.140 ;
        RECT 2138.610 127.940 2436.090 128.080 ;
        RECT 2138.610 127.880 2138.930 127.940 ;
        RECT 2435.770 127.880 2436.090 127.940 ;
      LAYER via ;
        RECT 2138.640 127.880 2138.900 128.140 ;
        RECT 2435.800 127.880 2436.060 128.140 ;
      LAYER met2 ;
        RECT 2135.830 216.650 2136.110 220.000 ;
        RECT 2135.830 216.510 2138.840 216.650 ;
        RECT 2135.830 216.000 2136.110 216.510 ;
        RECT 2138.700 128.170 2138.840 216.510 ;
        RECT 2138.640 127.850 2138.900 128.170 ;
        RECT 2435.800 127.850 2436.060 128.170 ;
        RECT 2435.860 17.410 2436.000 127.850 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2153.790 200.500 2154.110 200.560 ;
        RECT 2159.310 200.500 2159.630 200.560 ;
        RECT 2153.790 200.360 2159.630 200.500 ;
        RECT 2153.790 200.300 2154.110 200.360 ;
        RECT 2159.310 200.300 2159.630 200.360 ;
        RECT 2159.310 134.880 2159.630 134.940 ;
        RECT 2456.470 134.880 2456.790 134.940 ;
        RECT 2159.310 134.740 2456.790 134.880 ;
        RECT 2159.310 134.680 2159.630 134.740 ;
        RECT 2456.470 134.680 2456.790 134.740 ;
      LAYER via ;
        RECT 2153.820 200.300 2154.080 200.560 ;
        RECT 2159.340 200.300 2159.600 200.560 ;
        RECT 2159.340 134.680 2159.600 134.940 ;
        RECT 2456.500 134.680 2456.760 134.940 ;
      LAYER met2 ;
        RECT 2153.770 216.000 2154.050 220.000 ;
        RECT 2153.880 200.590 2154.020 216.000 ;
        RECT 2153.820 200.270 2154.080 200.590 ;
        RECT 2159.340 200.270 2159.600 200.590 ;
        RECT 2159.400 134.970 2159.540 200.270 ;
        RECT 2159.340 134.650 2159.600 134.970 ;
        RECT 2456.500 134.650 2456.760 134.970 ;
        RECT 2456.560 17.410 2456.700 134.650 ;
        RECT 2456.560 17.270 2459.000 17.410 ;
        RECT 2458.860 2.400 2459.000 17.270 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2173.110 141.340 2173.430 141.400 ;
        RECT 2470.730 141.340 2471.050 141.400 ;
        RECT 2173.110 141.200 2471.050 141.340 ;
        RECT 2173.110 141.140 2173.430 141.200 ;
        RECT 2470.730 141.140 2471.050 141.200 ;
        RECT 2470.730 18.940 2471.050 19.000 ;
        RECT 2476.710 18.940 2477.030 19.000 ;
        RECT 2470.730 18.800 2477.030 18.940 ;
        RECT 2470.730 18.740 2471.050 18.800 ;
        RECT 2476.710 18.740 2477.030 18.800 ;
      LAYER via ;
        RECT 2173.140 141.140 2173.400 141.400 ;
        RECT 2470.760 141.140 2471.020 141.400 ;
        RECT 2470.760 18.740 2471.020 19.000 ;
        RECT 2476.740 18.740 2477.000 19.000 ;
      LAYER met2 ;
        RECT 2171.710 216.650 2171.990 220.000 ;
        RECT 2171.710 216.510 2173.340 216.650 ;
        RECT 2171.710 216.000 2171.990 216.510 ;
        RECT 2173.200 141.430 2173.340 216.510 ;
        RECT 2173.140 141.110 2173.400 141.430 ;
        RECT 2470.760 141.110 2471.020 141.430 ;
        RECT 2470.820 19.030 2470.960 141.110 ;
        RECT 2470.760 18.710 2471.020 19.030 ;
        RECT 2476.740 18.710 2477.000 19.030 ;
        RECT 2476.800 2.400 2476.940 18.710 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2189.670 200.500 2189.990 200.560 ;
        RECT 2193.810 200.500 2194.130 200.560 ;
        RECT 2189.670 200.360 2194.130 200.500 ;
        RECT 2189.670 200.300 2189.990 200.360 ;
        RECT 2193.810 200.300 2194.130 200.360 ;
        RECT 2193.810 148.140 2194.130 148.200 ;
        RECT 2490.970 148.140 2491.290 148.200 ;
        RECT 2193.810 148.000 2491.290 148.140 ;
        RECT 2193.810 147.940 2194.130 148.000 ;
        RECT 2490.970 147.940 2491.290 148.000 ;
      LAYER via ;
        RECT 2189.700 200.300 2189.960 200.560 ;
        RECT 2193.840 200.300 2194.100 200.560 ;
        RECT 2193.840 147.940 2194.100 148.200 ;
        RECT 2491.000 147.940 2491.260 148.200 ;
      LAYER met2 ;
        RECT 2189.650 216.000 2189.930 220.000 ;
        RECT 2189.760 200.590 2189.900 216.000 ;
        RECT 2189.700 200.270 2189.960 200.590 ;
        RECT 2193.840 200.270 2194.100 200.590 ;
        RECT 2193.900 148.230 2194.040 200.270 ;
        RECT 2193.840 147.910 2194.100 148.230 ;
        RECT 2491.000 147.910 2491.260 148.230 ;
        RECT 2491.060 17.410 2491.200 147.910 ;
        RECT 2491.060 17.270 2494.880 17.410 ;
        RECT 2494.740 2.400 2494.880 17.270 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2207.150 155.280 2207.470 155.340 ;
        RECT 2512.130 155.280 2512.450 155.340 ;
        RECT 2207.150 155.140 2512.450 155.280 ;
        RECT 2207.150 155.080 2207.470 155.140 ;
        RECT 2512.130 155.080 2512.450 155.140 ;
      LAYER via ;
        RECT 2207.180 155.080 2207.440 155.340 ;
        RECT 2512.160 155.080 2512.420 155.340 ;
      LAYER met2 ;
        RECT 2207.590 216.650 2207.870 220.000 ;
        RECT 2207.240 216.510 2207.870 216.650 ;
        RECT 2207.240 155.370 2207.380 216.510 ;
        RECT 2207.590 216.000 2207.870 216.510 ;
        RECT 2207.180 155.050 2207.440 155.370 ;
        RECT 2512.160 155.050 2512.420 155.370 ;
        RECT 2512.220 2.400 2512.360 155.050 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2228.310 162.420 2228.630 162.480 ;
        RECT 2525.470 162.420 2525.790 162.480 ;
        RECT 2228.310 162.280 2525.790 162.420 ;
        RECT 2228.310 162.220 2228.630 162.280 ;
        RECT 2525.470 162.220 2525.790 162.280 ;
      LAYER via ;
        RECT 2228.340 162.220 2228.600 162.480 ;
        RECT 2525.500 162.220 2525.760 162.480 ;
      LAYER met2 ;
        RECT 2225.530 216.650 2225.810 220.000 ;
        RECT 2225.530 216.510 2228.540 216.650 ;
        RECT 2225.530 216.000 2225.810 216.510 ;
        RECT 2228.400 162.510 2228.540 216.510 ;
        RECT 2228.340 162.190 2228.600 162.510 ;
        RECT 2525.500 162.190 2525.760 162.510 ;
        RECT 2525.560 16.730 2525.700 162.190 ;
        RECT 2525.560 16.590 2530.300 16.730 ;
        RECT 2530.160 2.400 2530.300 16.590 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2243.030 200.500 2243.350 200.560 ;
        RECT 2248.550 200.500 2248.870 200.560 ;
        RECT 2243.030 200.360 2248.870 200.500 ;
        RECT 2243.030 200.300 2243.350 200.360 ;
        RECT 2248.550 200.300 2248.870 200.360 ;
        RECT 2248.550 169.220 2248.870 169.280 ;
        RECT 2546.170 169.220 2546.490 169.280 ;
        RECT 2248.550 169.080 2546.490 169.220 ;
        RECT 2248.550 169.020 2248.870 169.080 ;
        RECT 2546.170 169.020 2546.490 169.080 ;
      LAYER via ;
        RECT 2243.060 200.300 2243.320 200.560 ;
        RECT 2248.580 200.300 2248.840 200.560 ;
        RECT 2248.580 169.020 2248.840 169.280 ;
        RECT 2546.200 169.020 2546.460 169.280 ;
      LAYER met2 ;
        RECT 2243.010 216.000 2243.290 220.000 ;
        RECT 2243.120 200.590 2243.260 216.000 ;
        RECT 2243.060 200.270 2243.320 200.590 ;
        RECT 2248.580 200.270 2248.840 200.590 ;
        RECT 2248.640 169.310 2248.780 200.270 ;
        RECT 2248.580 168.990 2248.840 169.310 ;
        RECT 2546.200 168.990 2546.460 169.310 ;
        RECT 2546.260 16.730 2546.400 168.990 ;
        RECT 2546.260 16.590 2548.240 16.730 ;
        RECT 2548.100 2.400 2548.240 16.590 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2262.810 86.260 2263.130 86.320 ;
        RECT 2560.430 86.260 2560.750 86.320 ;
        RECT 2262.810 86.120 2560.750 86.260 ;
        RECT 2262.810 86.060 2263.130 86.120 ;
        RECT 2560.430 86.060 2560.750 86.120 ;
      LAYER via ;
        RECT 2262.840 86.060 2263.100 86.320 ;
        RECT 2560.460 86.060 2560.720 86.320 ;
      LAYER met2 ;
        RECT 2260.950 216.650 2261.230 220.000 ;
        RECT 2260.950 216.510 2263.040 216.650 ;
        RECT 2260.950 216.000 2261.230 216.510 ;
        RECT 2262.900 86.350 2263.040 216.510 ;
        RECT 2262.840 86.030 2263.100 86.350 ;
        RECT 2560.460 86.030 2560.720 86.350 ;
        RECT 2560.520 16.730 2560.660 86.030 ;
        RECT 2560.520 16.590 2566.180 16.730 ;
        RECT 2566.040 2.400 2566.180 16.590 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2278.910 200.500 2279.230 200.560 ;
        RECT 2283.510 200.500 2283.830 200.560 ;
        RECT 2278.910 200.360 2283.830 200.500 ;
        RECT 2278.910 200.300 2279.230 200.360 ;
        RECT 2283.510 200.300 2283.830 200.360 ;
        RECT 2283.510 100.200 2283.830 100.260 ;
        RECT 2580.670 100.200 2580.990 100.260 ;
        RECT 2283.510 100.060 2580.990 100.200 ;
        RECT 2283.510 100.000 2283.830 100.060 ;
        RECT 2580.670 100.000 2580.990 100.060 ;
      LAYER via ;
        RECT 2278.940 200.300 2279.200 200.560 ;
        RECT 2283.540 200.300 2283.800 200.560 ;
        RECT 2283.540 100.000 2283.800 100.260 ;
        RECT 2580.700 100.000 2580.960 100.260 ;
      LAYER met2 ;
        RECT 2278.890 216.000 2279.170 220.000 ;
        RECT 2279.000 200.590 2279.140 216.000 ;
        RECT 2278.940 200.270 2279.200 200.590 ;
        RECT 2283.540 200.270 2283.800 200.590 ;
        RECT 2283.600 100.290 2283.740 200.270 ;
        RECT 2283.540 99.970 2283.800 100.290 ;
        RECT 2580.700 99.970 2580.960 100.290 ;
        RECT 2580.760 16.730 2580.900 99.970 ;
        RECT 2580.760 16.590 2584.120 16.730 ;
        RECT 2583.980 2.400 2584.120 16.590 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 510.210 148.480 510.530 148.540 ;
        RECT 814.270 148.480 814.590 148.540 ;
        RECT 510.210 148.340 814.590 148.480 ;
        RECT 510.210 148.280 510.530 148.340 ;
        RECT 814.270 148.280 814.590 148.340 ;
      LAYER via ;
        RECT 510.240 148.280 510.500 148.540 ;
        RECT 814.300 148.280 814.560 148.540 ;
      LAYER met2 ;
        RECT 509.270 216.650 509.550 220.000 ;
        RECT 509.270 216.510 510.440 216.650 ;
        RECT 509.270 216.000 509.550 216.510 ;
        RECT 510.300 148.570 510.440 216.510 ;
        RECT 510.240 148.250 510.500 148.570 ;
        RECT 814.300 148.250 814.560 148.570 ;
        RECT 814.360 17.410 814.500 148.250 ;
        RECT 814.360 17.270 817.720 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2296.850 203.900 2297.170 203.960 ;
        RECT 2335.490 203.900 2335.810 203.960 ;
        RECT 2296.850 203.760 2335.810 203.900 ;
        RECT 2296.850 203.700 2297.170 203.760 ;
        RECT 2335.490 203.700 2335.810 203.760 ;
        RECT 2335.490 93.400 2335.810 93.460 ;
        RECT 2601.830 93.400 2602.150 93.460 ;
        RECT 2335.490 93.260 2602.150 93.400 ;
        RECT 2335.490 93.200 2335.810 93.260 ;
        RECT 2601.830 93.200 2602.150 93.260 ;
      LAYER via ;
        RECT 2296.880 203.700 2297.140 203.960 ;
        RECT 2335.520 203.700 2335.780 203.960 ;
        RECT 2335.520 93.200 2335.780 93.460 ;
        RECT 2601.860 93.200 2602.120 93.460 ;
      LAYER met2 ;
        RECT 2296.830 216.000 2297.110 220.000 ;
        RECT 2296.940 203.990 2297.080 216.000 ;
        RECT 2296.880 203.670 2297.140 203.990 ;
        RECT 2335.520 203.670 2335.780 203.990 ;
        RECT 2335.580 93.490 2335.720 203.670 ;
        RECT 2335.520 93.170 2335.780 93.490 ;
        RECT 2601.860 93.170 2602.120 93.490 ;
        RECT 2601.920 17.410 2602.060 93.170 ;
        RECT 2601.460 17.270 2602.060 17.410 ;
        RECT 2601.460 2.400 2601.600 17.270 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 25.400 2318.330 25.460 ;
        RECT 2619.310 25.400 2619.630 25.460 ;
        RECT 2318.010 25.260 2619.630 25.400 ;
        RECT 2318.010 25.200 2318.330 25.260 ;
        RECT 2619.310 25.200 2619.630 25.260 ;
      LAYER via ;
        RECT 2318.040 25.200 2318.300 25.460 ;
        RECT 2619.340 25.200 2619.600 25.460 ;
      LAYER met2 ;
        RECT 2314.770 216.650 2315.050 220.000 ;
        RECT 2314.770 216.510 2318.240 216.650 ;
        RECT 2314.770 216.000 2315.050 216.510 ;
        RECT 2318.100 25.490 2318.240 216.510 ;
        RECT 2318.040 25.170 2318.300 25.490 ;
        RECT 2619.340 25.170 2619.600 25.490 ;
        RECT 2619.400 2.400 2619.540 25.170 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2332.730 200.500 2333.050 200.560 ;
        RECT 2338.710 200.500 2339.030 200.560 ;
        RECT 2332.730 200.360 2339.030 200.500 ;
        RECT 2332.730 200.300 2333.050 200.360 ;
        RECT 2338.710 200.300 2339.030 200.360 ;
        RECT 2338.710 114.140 2339.030 114.200 ;
        RECT 2635.870 114.140 2636.190 114.200 ;
        RECT 2338.710 114.000 2636.190 114.140 ;
        RECT 2338.710 113.940 2339.030 114.000 ;
        RECT 2635.870 113.940 2636.190 114.000 ;
      LAYER via ;
        RECT 2332.760 200.300 2333.020 200.560 ;
        RECT 2338.740 200.300 2339.000 200.560 ;
        RECT 2338.740 113.940 2339.000 114.200 ;
        RECT 2635.900 113.940 2636.160 114.200 ;
      LAYER met2 ;
        RECT 2332.710 216.000 2332.990 220.000 ;
        RECT 2332.820 200.590 2332.960 216.000 ;
        RECT 2332.760 200.270 2333.020 200.590 ;
        RECT 2338.740 200.270 2339.000 200.590 ;
        RECT 2338.800 114.230 2338.940 200.270 ;
        RECT 2338.740 113.910 2339.000 114.230 ;
        RECT 2635.900 113.910 2636.160 114.230 ;
        RECT 2635.960 16.730 2636.100 113.910 ;
        RECT 2635.960 16.590 2637.480 16.730 ;
        RECT 2637.340 2.400 2637.480 16.590 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2352.510 107.340 2352.830 107.400 ;
        RECT 2649.670 107.340 2649.990 107.400 ;
        RECT 2352.510 107.200 2649.990 107.340 ;
        RECT 2352.510 107.140 2352.830 107.200 ;
        RECT 2649.670 107.140 2649.990 107.200 ;
      LAYER via ;
        RECT 2352.540 107.140 2352.800 107.400 ;
        RECT 2649.700 107.140 2649.960 107.400 ;
      LAYER met2 ;
        RECT 2350.650 216.650 2350.930 220.000 ;
        RECT 2350.650 216.510 2352.740 216.650 ;
        RECT 2350.650 216.000 2350.930 216.510 ;
        RECT 2352.600 107.430 2352.740 216.510 ;
        RECT 2352.540 107.110 2352.800 107.430 ;
        RECT 2649.700 107.110 2649.960 107.430 ;
        RECT 2649.760 17.410 2649.900 107.110 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2368.150 200.500 2368.470 200.560 ;
        RECT 2373.210 200.500 2373.530 200.560 ;
        RECT 2368.150 200.360 2373.530 200.500 ;
        RECT 2368.150 200.300 2368.470 200.360 ;
        RECT 2373.210 200.300 2373.530 200.360 ;
        RECT 2373.210 120.940 2373.530 121.000 ;
        RECT 2670.370 120.940 2670.690 121.000 ;
        RECT 2373.210 120.800 2670.690 120.940 ;
        RECT 2373.210 120.740 2373.530 120.800 ;
        RECT 2670.370 120.740 2670.690 120.800 ;
      LAYER via ;
        RECT 2368.180 200.300 2368.440 200.560 ;
        RECT 2373.240 200.300 2373.500 200.560 ;
        RECT 2373.240 120.740 2373.500 121.000 ;
        RECT 2670.400 120.740 2670.660 121.000 ;
      LAYER met2 ;
        RECT 2368.130 216.000 2368.410 220.000 ;
        RECT 2368.240 200.590 2368.380 216.000 ;
        RECT 2368.180 200.270 2368.440 200.590 ;
        RECT 2373.240 200.270 2373.500 200.590 ;
        RECT 2373.300 121.030 2373.440 200.270 ;
        RECT 2373.240 120.710 2373.500 121.030 ;
        RECT 2670.400 120.710 2670.660 121.030 ;
        RECT 2670.460 17.410 2670.600 120.710 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2387.010 127.740 2387.330 127.800 ;
        RECT 2684.170 127.740 2684.490 127.800 ;
        RECT 2387.010 127.600 2684.490 127.740 ;
        RECT 2387.010 127.540 2387.330 127.600 ;
        RECT 2684.170 127.540 2684.490 127.600 ;
        RECT 2684.170 18.260 2684.490 18.320 ;
        RECT 2690.610 18.260 2690.930 18.320 ;
        RECT 2684.170 18.120 2690.930 18.260 ;
        RECT 2684.170 18.060 2684.490 18.120 ;
        RECT 2690.610 18.060 2690.930 18.120 ;
      LAYER via ;
        RECT 2387.040 127.540 2387.300 127.800 ;
        RECT 2684.200 127.540 2684.460 127.800 ;
        RECT 2684.200 18.060 2684.460 18.320 ;
        RECT 2690.640 18.060 2690.900 18.320 ;
      LAYER met2 ;
        RECT 2386.070 216.650 2386.350 220.000 ;
        RECT 2386.070 216.510 2387.240 216.650 ;
        RECT 2386.070 216.000 2386.350 216.510 ;
        RECT 2387.100 127.830 2387.240 216.510 ;
        RECT 2387.040 127.510 2387.300 127.830 ;
        RECT 2684.200 127.510 2684.460 127.830 ;
        RECT 2684.260 18.350 2684.400 127.510 ;
        RECT 2684.200 18.030 2684.460 18.350 ;
        RECT 2690.640 18.030 2690.900 18.350 ;
        RECT 2690.700 2.400 2690.840 18.030 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2404.030 200.500 2404.350 200.560 ;
        RECT 2407.710 200.500 2408.030 200.560 ;
        RECT 2404.030 200.360 2408.030 200.500 ;
        RECT 2404.030 200.300 2404.350 200.360 ;
        RECT 2407.710 200.300 2408.030 200.360 ;
        RECT 2407.710 134.540 2408.030 134.600 ;
        RECT 2704.870 134.540 2705.190 134.600 ;
        RECT 2407.710 134.400 2705.190 134.540 ;
        RECT 2407.710 134.340 2408.030 134.400 ;
        RECT 2704.870 134.340 2705.190 134.400 ;
      LAYER via ;
        RECT 2404.060 200.300 2404.320 200.560 ;
        RECT 2407.740 200.300 2408.000 200.560 ;
        RECT 2407.740 134.340 2408.000 134.600 ;
        RECT 2704.900 134.340 2705.160 134.600 ;
      LAYER met2 ;
        RECT 2404.010 216.000 2404.290 220.000 ;
        RECT 2404.120 200.590 2404.260 216.000 ;
        RECT 2404.060 200.270 2404.320 200.590 ;
        RECT 2407.740 200.270 2408.000 200.590 ;
        RECT 2407.800 134.630 2407.940 200.270 ;
        RECT 2407.740 134.310 2408.000 134.630 ;
        RECT 2704.900 134.310 2705.160 134.630 ;
        RECT 2704.960 17.410 2705.100 134.310 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2421.970 200.500 2422.290 200.560 ;
        RECT 2427.950 200.500 2428.270 200.560 ;
        RECT 2421.970 200.360 2428.270 200.500 ;
        RECT 2421.970 200.300 2422.290 200.360 ;
        RECT 2427.950 200.300 2428.270 200.360 ;
        RECT 2427.950 141.680 2428.270 141.740 ;
        RECT 2725.570 141.680 2725.890 141.740 ;
        RECT 2427.950 141.540 2725.890 141.680 ;
        RECT 2427.950 141.480 2428.270 141.540 ;
        RECT 2725.570 141.480 2725.890 141.540 ;
      LAYER via ;
        RECT 2422.000 200.300 2422.260 200.560 ;
        RECT 2427.980 200.300 2428.240 200.560 ;
        RECT 2427.980 141.480 2428.240 141.740 ;
        RECT 2725.600 141.480 2725.860 141.740 ;
      LAYER met2 ;
        RECT 2421.950 216.000 2422.230 220.000 ;
        RECT 2422.060 200.590 2422.200 216.000 ;
        RECT 2422.000 200.270 2422.260 200.590 ;
        RECT 2427.980 200.270 2428.240 200.590 ;
        RECT 2428.040 141.770 2428.180 200.270 ;
        RECT 2427.980 141.450 2428.240 141.770 ;
        RECT 2725.600 141.450 2725.860 141.770 ;
        RECT 2725.660 17.410 2725.800 141.450 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2442.210 155.620 2442.530 155.680 ;
        RECT 2739.370 155.620 2739.690 155.680 ;
        RECT 2442.210 155.480 2739.690 155.620 ;
        RECT 2442.210 155.420 2442.530 155.480 ;
        RECT 2739.370 155.420 2739.690 155.480 ;
      LAYER via ;
        RECT 2442.240 155.420 2442.500 155.680 ;
        RECT 2739.400 155.420 2739.660 155.680 ;
      LAYER met2 ;
        RECT 2439.890 216.650 2440.170 220.000 ;
        RECT 2439.890 216.510 2442.440 216.650 ;
        RECT 2439.890 216.000 2440.170 216.510 ;
        RECT 2442.300 155.710 2442.440 216.510 ;
        RECT 2442.240 155.390 2442.500 155.710 ;
        RECT 2739.400 155.390 2739.660 155.710 ;
        RECT 2739.460 17.410 2739.600 155.390 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2457.850 200.500 2458.170 200.560 ;
        RECT 2462.910 200.500 2463.230 200.560 ;
        RECT 2457.850 200.360 2463.230 200.500 ;
        RECT 2457.850 200.300 2458.170 200.360 ;
        RECT 2462.910 200.300 2463.230 200.360 ;
        RECT 2462.910 162.080 2463.230 162.140 ;
        RECT 2760.070 162.080 2760.390 162.140 ;
        RECT 2462.910 161.940 2760.390 162.080 ;
        RECT 2462.910 161.880 2463.230 161.940 ;
        RECT 2760.070 161.880 2760.390 161.940 ;
      LAYER via ;
        RECT 2457.880 200.300 2458.140 200.560 ;
        RECT 2462.940 200.300 2463.200 200.560 ;
        RECT 2462.940 161.880 2463.200 162.140 ;
        RECT 2760.100 161.880 2760.360 162.140 ;
      LAYER met2 ;
        RECT 2457.830 216.000 2458.110 220.000 ;
        RECT 2457.940 200.590 2458.080 216.000 ;
        RECT 2457.880 200.270 2458.140 200.590 ;
        RECT 2462.940 200.270 2463.200 200.590 ;
        RECT 2463.000 162.170 2463.140 200.270 ;
        RECT 2462.940 161.850 2463.200 162.170 ;
        RECT 2760.100 161.850 2760.360 162.170 ;
        RECT 2760.160 17.410 2760.300 161.850 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 527.230 203.900 527.550 203.960 ;
        RECT 530.910 203.900 531.230 203.960 ;
        RECT 527.230 203.760 531.230 203.900 ;
        RECT 527.230 203.700 527.550 203.760 ;
        RECT 530.910 203.700 531.230 203.760 ;
        RECT 530.910 155.620 531.230 155.680 ;
        RECT 835.430 155.620 835.750 155.680 ;
        RECT 530.910 155.480 835.750 155.620 ;
        RECT 530.910 155.420 531.230 155.480 ;
        RECT 835.430 155.420 835.750 155.480 ;
      LAYER via ;
        RECT 527.260 203.700 527.520 203.960 ;
        RECT 530.940 203.700 531.200 203.960 ;
        RECT 530.940 155.420 531.200 155.680 ;
        RECT 835.460 155.420 835.720 155.680 ;
      LAYER met2 ;
        RECT 527.210 216.000 527.490 220.000 ;
        RECT 527.320 203.990 527.460 216.000 ;
        RECT 527.260 203.670 527.520 203.990 ;
        RECT 530.940 203.670 531.200 203.990 ;
        RECT 531.000 155.710 531.140 203.670 ;
        RECT 530.940 155.390 531.200 155.710 ;
        RECT 835.460 155.390 835.720 155.710 ;
        RECT 835.520 2.400 835.660 155.390 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2476.710 168.880 2477.030 168.940 ;
        RECT 2774.330 168.880 2774.650 168.940 ;
        RECT 2476.710 168.740 2774.650 168.880 ;
        RECT 2476.710 168.680 2477.030 168.740 ;
        RECT 2774.330 168.680 2774.650 168.740 ;
      LAYER via ;
        RECT 2476.740 168.680 2477.000 168.940 ;
        RECT 2774.360 168.680 2774.620 168.940 ;
      LAYER met2 ;
        RECT 2475.770 216.650 2476.050 220.000 ;
        RECT 2475.770 216.510 2476.940 216.650 ;
        RECT 2475.770 216.000 2476.050 216.510 ;
        RECT 2476.800 168.970 2476.940 216.510 ;
        RECT 2476.740 168.650 2477.000 168.970 ;
        RECT 2774.360 168.650 2774.620 168.970 ;
        RECT 2774.420 17.410 2774.560 168.650 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2493.270 200.500 2493.590 200.560 ;
        RECT 2497.410 200.500 2497.730 200.560 ;
        RECT 2493.270 200.360 2497.730 200.500 ;
        RECT 2493.270 200.300 2493.590 200.360 ;
        RECT 2497.410 200.300 2497.730 200.360 ;
        RECT 2497.410 58.720 2497.730 58.780 ;
        RECT 2794.570 58.720 2794.890 58.780 ;
        RECT 2497.410 58.580 2794.890 58.720 ;
        RECT 2497.410 58.520 2497.730 58.580 ;
        RECT 2794.570 58.520 2794.890 58.580 ;
      LAYER via ;
        RECT 2493.300 200.300 2493.560 200.560 ;
        RECT 2497.440 200.300 2497.700 200.560 ;
        RECT 2497.440 58.520 2497.700 58.780 ;
        RECT 2794.600 58.520 2794.860 58.780 ;
      LAYER met2 ;
        RECT 2493.250 216.000 2493.530 220.000 ;
        RECT 2493.360 200.590 2493.500 216.000 ;
        RECT 2493.300 200.270 2493.560 200.590 ;
        RECT 2497.440 200.270 2497.700 200.590 ;
        RECT 2497.500 58.810 2497.640 200.270 ;
        RECT 2497.440 58.490 2497.700 58.810 ;
        RECT 2794.600 58.490 2794.860 58.810 ;
        RECT 2794.660 17.410 2794.800 58.490 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2511.210 189.620 2511.530 189.680 ;
        RECT 2815.730 189.620 2816.050 189.680 ;
        RECT 2511.210 189.480 2816.050 189.620 ;
        RECT 2511.210 189.420 2511.530 189.480 ;
        RECT 2815.730 189.420 2816.050 189.480 ;
      LAYER via ;
        RECT 2511.240 189.420 2511.500 189.680 ;
        RECT 2815.760 189.420 2816.020 189.680 ;
      LAYER met2 ;
        RECT 2511.190 216.000 2511.470 220.000 ;
        RECT 2511.300 189.710 2511.440 216.000 ;
        RECT 2511.240 189.390 2511.500 189.710 ;
        RECT 2815.760 189.390 2816.020 189.710 ;
        RECT 2815.820 2.400 2815.960 189.390 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2531.910 99.860 2532.230 99.920 ;
        RECT 2829.070 99.860 2829.390 99.920 ;
        RECT 2531.910 99.720 2829.390 99.860 ;
        RECT 2531.910 99.660 2532.230 99.720 ;
        RECT 2829.070 99.660 2829.390 99.720 ;
      LAYER via ;
        RECT 2531.940 99.660 2532.200 99.920 ;
        RECT 2829.100 99.660 2829.360 99.920 ;
      LAYER met2 ;
        RECT 2529.130 216.650 2529.410 220.000 ;
        RECT 2529.130 216.510 2532.140 216.650 ;
        RECT 2529.130 216.000 2529.410 216.510 ;
        RECT 2532.000 99.950 2532.140 216.510 ;
        RECT 2531.940 99.630 2532.200 99.950 ;
        RECT 2829.100 99.630 2829.360 99.950 ;
        RECT 2829.160 17.410 2829.300 99.630 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2547.090 200.500 2547.410 200.560 ;
        RECT 2552.610 200.500 2552.930 200.560 ;
        RECT 2547.090 200.360 2552.930 200.500 ;
        RECT 2547.090 200.300 2547.410 200.360 ;
        RECT 2552.610 200.300 2552.930 200.360 ;
        RECT 2552.610 93.060 2552.930 93.120 ;
        RECT 2849.770 93.060 2850.090 93.120 ;
        RECT 2552.610 92.920 2850.090 93.060 ;
        RECT 2552.610 92.860 2552.930 92.920 ;
        RECT 2849.770 92.860 2850.090 92.920 ;
      LAYER via ;
        RECT 2547.120 200.300 2547.380 200.560 ;
        RECT 2552.640 200.300 2552.900 200.560 ;
        RECT 2552.640 92.860 2552.900 93.120 ;
        RECT 2849.800 92.860 2850.060 93.120 ;
      LAYER met2 ;
        RECT 2547.070 216.000 2547.350 220.000 ;
        RECT 2547.180 200.590 2547.320 216.000 ;
        RECT 2547.120 200.270 2547.380 200.590 ;
        RECT 2552.640 200.270 2552.900 200.590 ;
        RECT 2552.700 93.150 2552.840 200.270 ;
        RECT 2552.640 92.830 2552.900 93.150 ;
        RECT 2849.800 92.830 2850.060 93.150 ;
        RECT 2849.860 17.410 2850.000 92.830 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2566.410 16.560 2566.730 16.620 ;
        RECT 2869.090 16.560 2869.410 16.620 ;
        RECT 2566.410 16.420 2869.410 16.560 ;
        RECT 2566.410 16.360 2566.730 16.420 ;
        RECT 2869.090 16.360 2869.410 16.420 ;
      LAYER via ;
        RECT 2566.440 16.360 2566.700 16.620 ;
        RECT 2869.120 16.360 2869.380 16.620 ;
      LAYER met2 ;
        RECT 2565.010 216.650 2565.290 220.000 ;
        RECT 2565.010 216.510 2566.640 216.650 ;
        RECT 2565.010 216.000 2565.290 216.510 ;
        RECT 2566.500 16.650 2566.640 216.510 ;
        RECT 2566.440 16.330 2566.700 16.650 ;
        RECT 2869.120 16.330 2869.380 16.650 ;
        RECT 2869.180 2.400 2869.320 16.330 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2582.970 200.500 2583.290 200.560 ;
        RECT 2587.110 200.500 2587.430 200.560 ;
        RECT 2582.970 200.360 2587.430 200.500 ;
        RECT 2582.970 200.300 2583.290 200.360 ;
        RECT 2587.110 200.300 2587.430 200.360 ;
        RECT 2587.110 19.280 2587.430 19.340 ;
        RECT 2887.030 19.280 2887.350 19.340 ;
        RECT 2587.110 19.140 2887.350 19.280 ;
        RECT 2587.110 19.080 2587.430 19.140 ;
        RECT 2887.030 19.080 2887.350 19.140 ;
      LAYER via ;
        RECT 2583.000 200.300 2583.260 200.560 ;
        RECT 2587.140 200.300 2587.400 200.560 ;
        RECT 2587.140 19.080 2587.400 19.340 ;
        RECT 2887.060 19.080 2887.320 19.340 ;
      LAYER met2 ;
        RECT 2582.950 216.000 2583.230 220.000 ;
        RECT 2583.060 200.590 2583.200 216.000 ;
        RECT 2583.000 200.270 2583.260 200.590 ;
        RECT 2587.140 200.270 2587.400 200.590 ;
        RECT 2587.200 19.370 2587.340 200.270 ;
        RECT 2587.140 19.050 2587.400 19.370 ;
        RECT 2887.060 19.050 2887.320 19.370 ;
        RECT 2887.120 2.400 2887.260 19.050 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2600.890 216.000 2601.170 220.000 ;
        RECT 2601.000 16.845 2601.140 216.000 ;
        RECT 2600.930 16.475 2601.210 16.845 ;
        RECT 2904.990 16.475 2905.270 16.845 ;
        RECT 2905.060 2.400 2905.200 16.475 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2600.930 16.520 2601.210 16.800 ;
        RECT 2904.990 16.520 2905.270 16.800 ;
      LAYER met3 ;
        RECT 2600.905 16.810 2601.235 16.825 ;
        RECT 2904.965 16.810 2905.295 16.825 ;
        RECT 2600.905 16.510 2905.295 16.810 ;
        RECT 2600.905 16.495 2601.235 16.510 ;
        RECT 2904.965 16.495 2905.295 16.510 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 545.170 162.080 545.490 162.140 ;
        RECT 848.770 162.080 849.090 162.140 ;
        RECT 545.170 161.940 849.090 162.080 ;
        RECT 545.170 161.880 545.490 161.940 ;
        RECT 848.770 161.880 849.090 161.940 ;
      LAYER via ;
        RECT 545.200 161.880 545.460 162.140 ;
        RECT 848.800 161.880 849.060 162.140 ;
      LAYER met2 ;
        RECT 545.150 216.000 545.430 220.000 ;
        RECT 545.260 162.170 545.400 216.000 ;
        RECT 545.200 161.850 545.460 162.170 ;
        RECT 848.800 161.850 849.060 162.170 ;
        RECT 848.860 17.410 849.000 161.850 ;
        RECT 848.860 17.270 853.140 17.410 ;
        RECT 853.000 2.400 853.140 17.270 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 565.410 169.220 565.730 169.280 ;
        RECT 869.470 169.220 869.790 169.280 ;
        RECT 565.410 169.080 869.790 169.220 ;
        RECT 565.410 169.020 565.730 169.080 ;
        RECT 869.470 169.020 869.790 169.080 ;
      LAYER via ;
        RECT 565.440 169.020 565.700 169.280 ;
        RECT 869.500 169.020 869.760 169.280 ;
      LAYER met2 ;
        RECT 563.090 216.650 563.370 220.000 ;
        RECT 563.090 216.510 565.640 216.650 ;
        RECT 563.090 216.000 563.370 216.510 ;
        RECT 565.500 169.310 565.640 216.510 ;
        RECT 565.440 168.990 565.700 169.310 ;
        RECT 869.500 168.990 869.760 169.310 ;
        RECT 869.560 16.730 869.700 168.990 ;
        RECT 869.560 16.590 871.080 16.730 ;
        RECT 870.940 2.400 871.080 16.590 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 580.590 176.360 580.910 176.420 ;
        RECT 883.270 176.360 883.590 176.420 ;
        RECT 580.590 176.220 883.590 176.360 ;
        RECT 580.590 176.160 580.910 176.220 ;
        RECT 883.270 176.160 883.590 176.220 ;
      LAYER via ;
        RECT 580.620 176.160 580.880 176.420 ;
        RECT 883.300 176.160 883.560 176.420 ;
      LAYER met2 ;
        RECT 580.570 216.000 580.850 220.000 ;
        RECT 580.680 176.450 580.820 216.000 ;
        RECT 580.620 176.130 580.880 176.450 ;
        RECT 883.300 176.130 883.560 176.450 ;
        RECT 883.360 16.730 883.500 176.130 ;
        RECT 883.360 16.590 889.020 16.730 ;
        RECT 888.880 2.400 889.020 16.590 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 598.530 182.820 598.850 182.880 ;
        RECT 903.970 182.820 904.290 182.880 ;
        RECT 598.530 182.680 904.290 182.820 ;
        RECT 598.530 182.620 598.850 182.680 ;
        RECT 903.970 182.620 904.290 182.680 ;
      LAYER via ;
        RECT 598.560 182.620 598.820 182.880 ;
        RECT 904.000 182.620 904.260 182.880 ;
      LAYER met2 ;
        RECT 598.510 216.000 598.790 220.000 ;
        RECT 598.620 182.910 598.760 216.000 ;
        RECT 598.560 182.590 598.820 182.910 ;
        RECT 904.000 182.590 904.260 182.910 ;
        RECT 904.060 16.730 904.200 182.590 ;
        RECT 904.060 16.590 906.960 16.730 ;
        RECT 906.820 2.400 906.960 16.590 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 616.470 189.960 616.790 190.020 ;
        RECT 917.770 189.960 918.090 190.020 ;
        RECT 616.470 189.820 918.090 189.960 ;
        RECT 616.470 189.760 616.790 189.820 ;
        RECT 917.770 189.760 918.090 189.820 ;
        RECT 917.770 16.900 918.090 16.960 ;
        RECT 924.210 16.900 924.530 16.960 ;
        RECT 917.770 16.760 924.530 16.900 ;
        RECT 917.770 16.700 918.090 16.760 ;
        RECT 924.210 16.700 924.530 16.760 ;
      LAYER via ;
        RECT 616.500 189.760 616.760 190.020 ;
        RECT 917.800 189.760 918.060 190.020 ;
        RECT 917.800 16.700 918.060 16.960 ;
        RECT 924.240 16.700 924.500 16.960 ;
      LAYER met2 ;
        RECT 616.450 216.000 616.730 220.000 ;
        RECT 616.560 190.050 616.700 216.000 ;
        RECT 616.500 189.730 616.760 190.050 ;
        RECT 917.800 189.730 918.060 190.050 ;
        RECT 917.860 16.990 918.000 189.730 ;
        RECT 917.800 16.670 918.060 16.990 ;
        RECT 924.240 16.670 924.500 16.990 ;
        RECT 924.300 2.400 924.440 16.670 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 634.410 196.760 634.730 196.820 ;
        RECT 938.470 196.760 938.790 196.820 ;
        RECT 634.410 196.620 938.790 196.760 ;
        RECT 634.410 196.560 634.730 196.620 ;
        RECT 938.470 196.560 938.790 196.620 ;
      LAYER via ;
        RECT 634.440 196.560 634.700 196.820 ;
        RECT 938.500 196.560 938.760 196.820 ;
      LAYER met2 ;
        RECT 634.390 216.000 634.670 220.000 ;
        RECT 634.500 196.850 634.640 216.000 ;
        RECT 634.440 196.530 634.700 196.850 ;
        RECT 938.500 196.530 938.760 196.850 ;
        RECT 938.560 16.730 938.700 196.530 ;
        RECT 938.560 16.590 942.380 16.730 ;
        RECT 942.240 2.400 942.380 16.590 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 655.110 148.820 655.430 148.880 ;
        RECT 959.170 148.820 959.490 148.880 ;
        RECT 655.110 148.680 959.490 148.820 ;
        RECT 655.110 148.620 655.430 148.680 ;
        RECT 959.170 148.620 959.490 148.680 ;
      LAYER via ;
        RECT 655.140 148.620 655.400 148.880 ;
        RECT 959.200 148.620 959.460 148.880 ;
      LAYER met2 ;
        RECT 652.330 216.650 652.610 220.000 ;
        RECT 652.330 216.510 655.340 216.650 ;
        RECT 652.330 216.000 652.610 216.510 ;
        RECT 655.200 148.910 655.340 216.510 ;
        RECT 655.140 148.590 655.400 148.910 ;
        RECT 959.200 148.590 959.460 148.910 ;
        RECT 959.260 16.730 959.400 148.590 ;
        RECT 959.260 16.590 960.320 16.730 ;
        RECT 960.180 2.400 960.320 16.590 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 670.290 202.880 670.610 202.940 ;
        RECT 675.810 202.880 676.130 202.940 ;
        RECT 670.290 202.740 676.130 202.880 ;
        RECT 670.290 202.680 670.610 202.740 ;
        RECT 675.810 202.680 676.130 202.740 ;
        RECT 675.810 155.960 676.130 156.020 ;
        RECT 972.970 155.960 973.290 156.020 ;
        RECT 675.810 155.820 973.290 155.960 ;
        RECT 675.810 155.760 676.130 155.820 ;
        RECT 972.970 155.760 973.290 155.820 ;
      LAYER via ;
        RECT 670.320 202.680 670.580 202.940 ;
        RECT 675.840 202.680 676.100 202.940 ;
        RECT 675.840 155.760 676.100 156.020 ;
        RECT 973.000 155.760 973.260 156.020 ;
      LAYER met2 ;
        RECT 670.270 216.000 670.550 220.000 ;
        RECT 670.380 202.970 670.520 216.000 ;
        RECT 670.320 202.650 670.580 202.970 ;
        RECT 675.840 202.650 676.100 202.970 ;
        RECT 675.900 156.050 676.040 202.650 ;
        RECT 675.840 155.730 676.100 156.050 ;
        RECT 973.000 155.730 973.260 156.050 ;
        RECT 973.060 16.730 973.200 155.730 ;
        RECT 973.060 16.590 978.260 16.730 ;
        RECT 978.120 2.400 978.260 16.590 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 351.510 86.600 351.830 86.660 ;
        RECT 655.570 86.600 655.890 86.660 ;
        RECT 351.510 86.460 655.890 86.600 ;
        RECT 351.510 86.400 351.830 86.460 ;
        RECT 655.570 86.400 655.890 86.460 ;
      LAYER via ;
        RECT 351.540 86.400 351.800 86.660 ;
        RECT 655.600 86.400 655.860 86.660 ;
      LAYER met2 ;
        RECT 348.270 216.650 348.550 220.000 ;
        RECT 348.270 216.510 351.740 216.650 ;
        RECT 348.270 216.000 348.550 216.510 ;
        RECT 351.600 86.690 351.740 216.510 ;
        RECT 351.540 86.370 351.800 86.690 ;
        RECT 655.600 86.370 655.860 86.690 ;
        RECT 655.660 17.410 655.800 86.370 ;
        RECT 655.660 17.270 657.180 17.410 ;
        RECT 657.040 2.400 657.180 17.270 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.610 37.980 689.930 38.040 ;
        RECT 995.970 37.980 996.290 38.040 ;
        RECT 689.610 37.840 996.290 37.980 ;
        RECT 689.610 37.780 689.930 37.840 ;
        RECT 995.970 37.780 996.290 37.840 ;
      LAYER via ;
        RECT 689.640 37.780 689.900 38.040 ;
        RECT 996.000 37.780 996.260 38.040 ;
      LAYER met2 ;
        RECT 688.210 216.650 688.490 220.000 ;
        RECT 688.210 216.510 689.840 216.650 ;
        RECT 688.210 216.000 688.490 216.510 ;
        RECT 689.700 38.070 689.840 216.510 ;
        RECT 689.640 37.750 689.900 38.070 ;
        RECT 996.000 37.750 996.260 38.070 ;
        RECT 996.060 2.400 996.200 37.750 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 705.710 162.420 706.030 162.480 ;
        RECT 1007.470 162.420 1007.790 162.480 ;
        RECT 705.710 162.280 1007.790 162.420 ;
        RECT 705.710 162.220 706.030 162.280 ;
        RECT 1007.470 162.220 1007.790 162.280 ;
        RECT 1007.470 18.260 1007.790 18.320 ;
        RECT 1013.450 18.260 1013.770 18.320 ;
        RECT 1007.470 18.120 1013.770 18.260 ;
        RECT 1007.470 18.060 1007.790 18.120 ;
        RECT 1013.450 18.060 1013.770 18.120 ;
      LAYER via ;
        RECT 705.740 162.220 706.000 162.480 ;
        RECT 1007.500 162.220 1007.760 162.480 ;
        RECT 1007.500 18.060 1007.760 18.320 ;
        RECT 1013.480 18.060 1013.740 18.320 ;
      LAYER met2 ;
        RECT 705.690 216.000 705.970 220.000 ;
        RECT 705.800 162.510 705.940 216.000 ;
        RECT 705.740 162.190 706.000 162.510 ;
        RECT 1007.500 162.190 1007.760 162.510 ;
        RECT 1007.560 18.350 1007.700 162.190 ;
        RECT 1007.500 18.030 1007.760 18.350 ;
        RECT 1013.480 18.030 1013.740 18.350 ;
        RECT 1013.540 2.400 1013.680 18.030 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 723.650 168.880 723.970 168.940 ;
        RECT 1028.170 168.880 1028.490 168.940 ;
        RECT 723.650 168.740 1028.490 168.880 ;
        RECT 723.650 168.680 723.970 168.740 ;
        RECT 1028.170 168.680 1028.490 168.740 ;
      LAYER via ;
        RECT 723.680 168.680 723.940 168.940 ;
        RECT 1028.200 168.680 1028.460 168.940 ;
      LAYER met2 ;
        RECT 723.630 216.000 723.910 220.000 ;
        RECT 723.740 168.970 723.880 216.000 ;
        RECT 723.680 168.650 723.940 168.970 ;
        RECT 1028.200 168.650 1028.460 168.970 ;
        RECT 1028.260 16.730 1028.400 168.650 ;
        RECT 1028.260 16.590 1031.620 16.730 ;
        RECT 1031.480 2.400 1031.620 16.590 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 744.810 176.020 745.130 176.080 ;
        RECT 1049.330 176.020 1049.650 176.080 ;
        RECT 744.810 175.880 1049.650 176.020 ;
        RECT 744.810 175.820 745.130 175.880 ;
        RECT 1049.330 175.820 1049.650 175.880 ;
      LAYER via ;
        RECT 744.840 175.820 745.100 176.080 ;
        RECT 1049.360 175.820 1049.620 176.080 ;
      LAYER met2 ;
        RECT 741.570 216.650 741.850 220.000 ;
        RECT 741.570 216.510 745.040 216.650 ;
        RECT 741.570 216.000 741.850 216.510 ;
        RECT 744.900 176.110 745.040 216.510 ;
        RECT 744.840 175.790 745.100 176.110 ;
        RECT 1049.360 175.790 1049.620 176.110 ;
        RECT 1049.420 2.400 1049.560 175.790 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 759.530 183.160 759.850 183.220 ;
        RECT 1062.670 183.160 1062.990 183.220 ;
        RECT 759.530 183.020 1062.990 183.160 ;
        RECT 759.530 182.960 759.850 183.020 ;
        RECT 1062.670 182.960 1062.990 183.020 ;
      LAYER via ;
        RECT 759.560 182.960 759.820 183.220 ;
        RECT 1062.700 182.960 1062.960 183.220 ;
      LAYER met2 ;
        RECT 759.510 216.000 759.790 220.000 ;
        RECT 759.620 183.250 759.760 216.000 ;
        RECT 759.560 182.930 759.820 183.250 ;
        RECT 1062.700 182.930 1062.960 183.250 ;
        RECT 1062.760 16.730 1062.900 182.930 ;
        RECT 1062.760 16.590 1067.500 16.730 ;
        RECT 1067.360 2.400 1067.500 16.590 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 777.470 189.620 777.790 189.680 ;
        RECT 1083.370 189.620 1083.690 189.680 ;
        RECT 777.470 189.480 1083.690 189.620 ;
        RECT 777.470 189.420 777.790 189.480 ;
        RECT 1083.370 189.420 1083.690 189.480 ;
      LAYER via ;
        RECT 777.500 189.420 777.760 189.680 ;
        RECT 1083.400 189.420 1083.660 189.680 ;
      LAYER met2 ;
        RECT 777.450 216.000 777.730 220.000 ;
        RECT 777.560 189.710 777.700 216.000 ;
        RECT 777.500 189.390 777.760 189.710 ;
        RECT 1083.400 189.390 1083.660 189.710 ;
        RECT 1083.460 16.730 1083.600 189.390 ;
        RECT 1083.460 16.590 1085.440 16.730 ;
        RECT 1085.300 2.400 1085.440 16.590 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 795.410 197.100 795.730 197.160 ;
        RECT 1097.170 197.100 1097.490 197.160 ;
        RECT 795.410 196.960 1097.490 197.100 ;
        RECT 795.410 196.900 795.730 196.960 ;
        RECT 1097.170 196.900 1097.490 196.960 ;
      LAYER via ;
        RECT 795.440 196.900 795.700 197.160 ;
        RECT 1097.200 196.900 1097.460 197.160 ;
      LAYER met2 ;
        RECT 795.390 216.000 795.670 220.000 ;
        RECT 795.500 197.190 795.640 216.000 ;
        RECT 795.440 196.870 795.700 197.190 ;
        RECT 1097.200 196.870 1097.460 197.190 ;
        RECT 1097.260 16.730 1097.400 196.870 ;
        RECT 1097.260 16.590 1102.920 16.730 ;
        RECT 1102.780 2.400 1102.920 16.590 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 813.350 148.140 813.670 148.200 ;
        RECT 1117.870 148.140 1118.190 148.200 ;
        RECT 813.350 148.000 1118.190 148.140 ;
        RECT 813.350 147.940 813.670 148.000 ;
        RECT 1117.870 147.940 1118.190 148.000 ;
      LAYER via ;
        RECT 813.380 147.940 813.640 148.200 ;
        RECT 1117.900 147.940 1118.160 148.200 ;
      LAYER met2 ;
        RECT 813.330 216.000 813.610 220.000 ;
        RECT 813.440 148.230 813.580 216.000 ;
        RECT 813.380 147.910 813.640 148.230 ;
        RECT 1117.900 147.910 1118.160 148.230 ;
        RECT 1117.960 16.730 1118.100 147.910 ;
        RECT 1117.960 16.590 1120.860 16.730 ;
        RECT 1120.720 2.400 1120.860 16.590 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 830.830 200.500 831.150 200.560 ;
        RECT 834.510 200.500 834.830 200.560 ;
        RECT 830.830 200.360 834.830 200.500 ;
        RECT 830.830 200.300 831.150 200.360 ;
        RECT 834.510 200.300 834.830 200.360 ;
        RECT 834.510 155.280 834.830 155.340 ;
        RECT 1139.030 155.280 1139.350 155.340 ;
        RECT 834.510 155.140 1139.350 155.280 ;
        RECT 834.510 155.080 834.830 155.140 ;
        RECT 1139.030 155.080 1139.350 155.140 ;
      LAYER via ;
        RECT 830.860 200.300 831.120 200.560 ;
        RECT 834.540 200.300 834.800 200.560 ;
        RECT 834.540 155.080 834.800 155.340 ;
        RECT 1139.060 155.080 1139.320 155.340 ;
      LAYER met2 ;
        RECT 830.810 216.000 831.090 220.000 ;
        RECT 830.920 200.590 831.060 216.000 ;
        RECT 830.860 200.270 831.120 200.590 ;
        RECT 834.540 200.270 834.800 200.590 ;
        RECT 834.600 155.370 834.740 200.270 ;
        RECT 834.540 155.050 834.800 155.370 ;
        RECT 1139.060 155.050 1139.320 155.370 ;
        RECT 1139.120 17.410 1139.260 155.050 ;
        RECT 1138.660 17.270 1139.260 17.410 ;
        RECT 1138.660 2.400 1138.800 17.270 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 848.770 200.500 849.090 200.560 ;
        RECT 854.750 200.500 855.070 200.560 ;
        RECT 848.770 200.360 855.070 200.500 ;
        RECT 848.770 200.300 849.090 200.360 ;
        RECT 854.750 200.300 855.070 200.360 ;
        RECT 854.750 162.080 855.070 162.140 ;
        RECT 1152.370 162.080 1152.690 162.140 ;
        RECT 854.750 161.940 1152.690 162.080 ;
        RECT 854.750 161.880 855.070 161.940 ;
        RECT 1152.370 161.880 1152.690 161.940 ;
      LAYER via ;
        RECT 848.800 200.300 849.060 200.560 ;
        RECT 854.780 200.300 855.040 200.560 ;
        RECT 854.780 161.880 855.040 162.140 ;
        RECT 1152.400 161.880 1152.660 162.140 ;
      LAYER met2 ;
        RECT 848.750 216.000 849.030 220.000 ;
        RECT 848.860 200.590 849.000 216.000 ;
        RECT 848.800 200.270 849.060 200.590 ;
        RECT 854.780 200.270 855.040 200.590 ;
        RECT 854.840 162.170 854.980 200.270 ;
        RECT 854.780 161.850 855.040 162.170 ;
        RECT 1152.400 161.850 1152.660 162.170 ;
        RECT 1152.460 17.410 1152.600 161.850 ;
        RECT 1152.460 17.270 1156.740 17.410 ;
        RECT 1156.600 2.400 1156.740 17.270 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 366.230 197.100 366.550 197.160 ;
        RECT 669.370 197.100 669.690 197.160 ;
        RECT 366.230 196.960 669.690 197.100 ;
        RECT 366.230 196.900 366.550 196.960 ;
        RECT 669.370 196.900 669.690 196.960 ;
      LAYER via ;
        RECT 366.260 196.900 366.520 197.160 ;
        RECT 669.400 196.900 669.660 197.160 ;
      LAYER met2 ;
        RECT 366.210 216.000 366.490 220.000 ;
        RECT 366.320 197.190 366.460 216.000 ;
        RECT 366.260 196.870 366.520 197.190 ;
        RECT 669.400 196.870 669.660 197.190 ;
        RECT 669.460 16.730 669.600 196.870 ;
        RECT 669.460 16.590 674.660 16.730 ;
        RECT 674.520 2.400 674.660 16.590 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 869.010 24.040 869.330 24.100 ;
        RECT 1173.990 24.040 1174.310 24.100 ;
        RECT 869.010 23.900 1174.310 24.040 ;
        RECT 869.010 23.840 869.330 23.900 ;
        RECT 1173.990 23.840 1174.310 23.900 ;
      LAYER via ;
        RECT 869.040 23.840 869.300 24.100 ;
        RECT 1174.020 23.840 1174.280 24.100 ;
      LAYER met2 ;
        RECT 866.690 216.650 866.970 220.000 ;
        RECT 866.690 216.510 869.240 216.650 ;
        RECT 866.690 216.000 866.970 216.510 ;
        RECT 869.100 24.130 869.240 216.510 ;
        RECT 869.040 23.810 869.300 24.130 ;
        RECT 1174.020 23.810 1174.280 24.130 ;
        RECT 1174.080 2.400 1174.220 23.810 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 884.650 200.500 884.970 200.560 ;
        RECT 889.710 200.500 890.030 200.560 ;
        RECT 884.650 200.360 890.030 200.500 ;
        RECT 884.650 200.300 884.970 200.360 ;
        RECT 889.710 200.300 890.030 200.360 ;
        RECT 889.710 169.560 890.030 169.620 ;
        RECT 1186.870 169.560 1187.190 169.620 ;
        RECT 889.710 169.420 1187.190 169.560 ;
        RECT 889.710 169.360 890.030 169.420 ;
        RECT 1186.870 169.360 1187.190 169.420 ;
      LAYER via ;
        RECT 884.680 200.300 884.940 200.560 ;
        RECT 889.740 200.300 890.000 200.560 ;
        RECT 889.740 169.360 890.000 169.620 ;
        RECT 1186.900 169.360 1187.160 169.620 ;
      LAYER met2 ;
        RECT 884.630 216.000 884.910 220.000 ;
        RECT 884.740 200.590 884.880 216.000 ;
        RECT 884.680 200.270 884.940 200.590 ;
        RECT 889.740 200.270 890.000 200.590 ;
        RECT 889.800 169.650 889.940 200.270 ;
        RECT 889.740 169.330 890.000 169.650 ;
        RECT 1186.900 169.330 1187.160 169.650 ;
        RECT 1186.960 17.410 1187.100 169.330 ;
        RECT 1186.960 17.270 1192.160 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 903.510 176.360 903.830 176.420 ;
        RECT 1207.570 176.360 1207.890 176.420 ;
        RECT 903.510 176.220 1207.890 176.360 ;
        RECT 903.510 176.160 903.830 176.220 ;
        RECT 1207.570 176.160 1207.890 176.220 ;
      LAYER via ;
        RECT 903.540 176.160 903.800 176.420 ;
        RECT 1207.600 176.160 1207.860 176.420 ;
      LAYER met2 ;
        RECT 902.570 216.650 902.850 220.000 ;
        RECT 902.570 216.510 903.740 216.650 ;
        RECT 902.570 216.000 902.850 216.510 ;
        RECT 903.600 176.450 903.740 216.510 ;
        RECT 903.540 176.130 903.800 176.450 ;
        RECT 1207.600 176.130 1207.860 176.450 ;
        RECT 1207.660 16.730 1207.800 176.130 ;
        RECT 1207.660 16.590 1210.100 16.730 ;
        RECT 1209.960 2.400 1210.100 16.590 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 920.530 183.500 920.850 183.560 ;
        RECT 1221.370 183.500 1221.690 183.560 ;
        RECT 920.530 183.360 1221.690 183.500 ;
        RECT 920.530 183.300 920.850 183.360 ;
        RECT 1221.370 183.300 1221.690 183.360 ;
        RECT 1221.370 17.240 1221.690 17.300 ;
        RECT 1227.810 17.240 1228.130 17.300 ;
        RECT 1221.370 17.100 1228.130 17.240 ;
        RECT 1221.370 17.040 1221.690 17.100 ;
        RECT 1227.810 17.040 1228.130 17.100 ;
      LAYER via ;
        RECT 920.560 183.300 920.820 183.560 ;
        RECT 1221.400 183.300 1221.660 183.560 ;
        RECT 1221.400 17.040 1221.660 17.300 ;
        RECT 1227.840 17.040 1228.100 17.300 ;
      LAYER met2 ;
        RECT 920.510 216.000 920.790 220.000 ;
        RECT 920.620 183.590 920.760 216.000 ;
        RECT 920.560 183.270 920.820 183.590 ;
        RECT 1221.400 183.270 1221.660 183.590 ;
        RECT 1221.460 17.330 1221.600 183.270 ;
        RECT 1221.400 17.010 1221.660 17.330 ;
        RECT 1227.840 17.010 1228.100 17.330 ;
        RECT 1227.900 2.400 1228.040 17.010 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 939.850 189.960 940.170 190.020 ;
        RECT 1242.070 189.960 1242.390 190.020 ;
        RECT 939.850 189.820 1242.390 189.960 ;
        RECT 939.850 189.760 940.170 189.820 ;
        RECT 1242.070 189.760 1242.390 189.820 ;
      LAYER via ;
        RECT 939.880 189.760 940.140 190.020 ;
        RECT 1242.100 189.760 1242.360 190.020 ;
      LAYER met2 ;
        RECT 938.450 216.650 938.730 220.000 ;
        RECT 938.450 216.510 940.080 216.650 ;
        RECT 938.450 216.000 938.730 216.510 ;
        RECT 939.940 190.050 940.080 216.510 ;
        RECT 939.880 189.730 940.140 190.050 ;
        RECT 1242.100 189.730 1242.360 190.050 ;
        RECT 1242.160 16.730 1242.300 189.730 ;
        RECT 1242.160 16.590 1245.980 16.730 ;
        RECT 1245.840 2.400 1245.980 16.590 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 958.710 149.160 959.030 149.220 ;
        RECT 1263.230 149.160 1263.550 149.220 ;
        RECT 958.710 149.020 1263.550 149.160 ;
        RECT 958.710 148.960 959.030 149.020 ;
        RECT 1263.230 148.960 1263.550 149.020 ;
      LAYER via ;
        RECT 958.740 148.960 959.000 149.220 ;
        RECT 1263.260 148.960 1263.520 149.220 ;
      LAYER met2 ;
        RECT 955.930 216.650 956.210 220.000 ;
        RECT 955.930 216.510 958.940 216.650 ;
        RECT 955.930 216.000 956.210 216.510 ;
        RECT 958.800 149.250 958.940 216.510 ;
        RECT 958.740 148.930 959.000 149.250 ;
        RECT 1263.260 148.930 1263.520 149.250 ;
        RECT 1263.320 2.400 1263.460 148.930 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 973.890 196.760 974.210 196.820 ;
        RECT 1276.570 196.760 1276.890 196.820 ;
        RECT 973.890 196.620 1276.890 196.760 ;
        RECT 973.890 196.560 974.210 196.620 ;
        RECT 1276.570 196.560 1276.890 196.620 ;
      LAYER via ;
        RECT 973.920 196.560 974.180 196.820 ;
        RECT 1276.600 196.560 1276.860 196.820 ;
      LAYER met2 ;
        RECT 973.870 216.000 974.150 220.000 ;
        RECT 973.980 196.850 974.120 216.000 ;
        RECT 973.920 196.530 974.180 196.850 ;
        RECT 1276.600 196.530 1276.860 196.850 ;
        RECT 1276.660 16.730 1276.800 196.530 ;
        RECT 1276.660 16.590 1281.400 16.730 ;
        RECT 1281.260 2.400 1281.400 16.590 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 993.210 155.620 993.530 155.680 ;
        RECT 1297.270 155.620 1297.590 155.680 ;
        RECT 993.210 155.480 1297.590 155.620 ;
        RECT 993.210 155.420 993.530 155.480 ;
        RECT 1297.270 155.420 1297.590 155.480 ;
      LAYER via ;
        RECT 993.240 155.420 993.500 155.680 ;
        RECT 1297.300 155.420 1297.560 155.680 ;
      LAYER met2 ;
        RECT 991.810 216.650 992.090 220.000 ;
        RECT 991.810 216.510 993.440 216.650 ;
        RECT 991.810 216.000 992.090 216.510 ;
        RECT 993.300 155.710 993.440 216.510 ;
        RECT 993.240 155.390 993.500 155.710 ;
        RECT 1297.300 155.390 1297.560 155.710 ;
        RECT 1297.360 17.410 1297.500 155.390 ;
        RECT 1297.360 17.270 1299.340 17.410 ;
        RECT 1299.200 2.400 1299.340 17.270 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1009.770 200.500 1010.090 200.560 ;
        RECT 1013.910 200.500 1014.230 200.560 ;
        RECT 1009.770 200.360 1014.230 200.500 ;
        RECT 1009.770 200.300 1010.090 200.360 ;
        RECT 1013.910 200.300 1014.230 200.360 ;
        RECT 1013.910 162.420 1014.230 162.480 ;
        RECT 1311.070 162.420 1311.390 162.480 ;
        RECT 1013.910 162.280 1311.390 162.420 ;
        RECT 1013.910 162.220 1014.230 162.280 ;
        RECT 1311.070 162.220 1311.390 162.280 ;
        RECT 1311.070 18.940 1311.390 19.000 ;
        RECT 1317.050 18.940 1317.370 19.000 ;
        RECT 1311.070 18.800 1317.370 18.940 ;
        RECT 1311.070 18.740 1311.390 18.800 ;
        RECT 1317.050 18.740 1317.370 18.800 ;
      LAYER via ;
        RECT 1009.800 200.300 1010.060 200.560 ;
        RECT 1013.940 200.300 1014.200 200.560 ;
        RECT 1013.940 162.220 1014.200 162.480 ;
        RECT 1311.100 162.220 1311.360 162.480 ;
        RECT 1311.100 18.740 1311.360 19.000 ;
        RECT 1317.080 18.740 1317.340 19.000 ;
      LAYER met2 ;
        RECT 1009.750 216.000 1010.030 220.000 ;
        RECT 1009.860 200.590 1010.000 216.000 ;
        RECT 1009.800 200.270 1010.060 200.590 ;
        RECT 1013.940 200.270 1014.200 200.590 ;
        RECT 1014.000 162.510 1014.140 200.270 ;
        RECT 1013.940 162.190 1014.200 162.510 ;
        RECT 1311.100 162.190 1311.360 162.510 ;
        RECT 1311.160 19.030 1311.300 162.190 ;
        RECT 1311.100 18.710 1311.360 19.030 ;
        RECT 1317.080 18.710 1317.340 19.030 ;
        RECT 1317.140 2.400 1317.280 18.710 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1027.250 169.220 1027.570 169.280 ;
        RECT 1331.770 169.220 1332.090 169.280 ;
        RECT 1027.250 169.080 1332.090 169.220 ;
        RECT 1027.250 169.020 1027.570 169.080 ;
        RECT 1331.770 169.020 1332.090 169.080 ;
      LAYER via ;
        RECT 1027.280 169.020 1027.540 169.280 ;
        RECT 1331.800 169.020 1332.060 169.280 ;
      LAYER met2 ;
        RECT 1027.690 216.650 1027.970 220.000 ;
        RECT 1027.340 216.510 1027.970 216.650 ;
        RECT 1027.340 169.310 1027.480 216.510 ;
        RECT 1027.690 216.000 1027.970 216.510 ;
        RECT 1027.280 168.990 1027.540 169.310 ;
        RECT 1331.800 168.990 1332.060 169.310 ;
        RECT 1331.860 17.410 1332.000 168.990 ;
        RECT 1331.860 17.270 1335.220 17.410 ;
        RECT 1335.080 2.400 1335.220 17.270 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 384.170 189.620 384.490 189.680 ;
        RECT 690.070 189.620 690.390 189.680 ;
        RECT 384.170 189.480 690.390 189.620 ;
        RECT 384.170 189.420 384.490 189.480 ;
        RECT 690.070 189.420 690.390 189.480 ;
      LAYER via ;
        RECT 384.200 189.420 384.460 189.680 ;
        RECT 690.100 189.420 690.360 189.680 ;
      LAYER met2 ;
        RECT 384.150 216.000 384.430 220.000 ;
        RECT 384.260 189.710 384.400 216.000 ;
        RECT 384.200 189.390 384.460 189.710 ;
        RECT 690.100 189.390 690.360 189.710 ;
        RECT 690.160 16.730 690.300 189.390 ;
        RECT 690.160 16.590 692.600 16.730 ;
        RECT 692.460 2.400 692.600 16.590 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1048.410 30.840 1048.730 30.900 ;
        RECT 1352.930 30.840 1353.250 30.900 ;
        RECT 1048.410 30.700 1353.250 30.840 ;
        RECT 1048.410 30.640 1048.730 30.700 ;
        RECT 1352.930 30.640 1353.250 30.700 ;
      LAYER via ;
        RECT 1048.440 30.640 1048.700 30.900 ;
        RECT 1352.960 30.640 1353.220 30.900 ;
      LAYER met2 ;
        RECT 1045.630 216.650 1045.910 220.000 ;
        RECT 1045.630 216.510 1048.640 216.650 ;
        RECT 1045.630 216.000 1045.910 216.510 ;
        RECT 1048.500 30.930 1048.640 216.510 ;
        RECT 1048.440 30.610 1048.700 30.930 ;
        RECT 1352.960 30.610 1353.220 30.930 ;
        RECT 1353.020 16.050 1353.160 30.610 ;
        RECT 1352.560 15.910 1353.160 16.050 ;
        RECT 1352.560 2.400 1352.700 15.910 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1063.590 200.500 1063.910 200.560 ;
        RECT 1069.110 200.500 1069.430 200.560 ;
        RECT 1063.590 200.360 1069.430 200.500 ;
        RECT 1063.590 200.300 1063.910 200.360 ;
        RECT 1069.110 200.300 1069.430 200.360 ;
        RECT 1069.110 176.700 1069.430 176.760 ;
        RECT 1366.270 176.700 1366.590 176.760 ;
        RECT 1069.110 176.560 1366.590 176.700 ;
        RECT 1069.110 176.500 1069.430 176.560 ;
        RECT 1366.270 176.500 1366.590 176.560 ;
      LAYER via ;
        RECT 1063.620 200.300 1063.880 200.560 ;
        RECT 1069.140 200.300 1069.400 200.560 ;
        RECT 1069.140 176.500 1069.400 176.760 ;
        RECT 1366.300 176.500 1366.560 176.760 ;
      LAYER met2 ;
        RECT 1063.570 216.000 1063.850 220.000 ;
        RECT 1063.680 200.590 1063.820 216.000 ;
        RECT 1063.620 200.270 1063.880 200.590 ;
        RECT 1069.140 200.270 1069.400 200.590 ;
        RECT 1069.200 176.790 1069.340 200.270 ;
        RECT 1069.140 176.470 1069.400 176.790 ;
        RECT 1366.300 176.470 1366.560 176.790 ;
        RECT 1366.360 17.410 1366.500 176.470 ;
        RECT 1366.360 17.270 1370.640 17.410 ;
        RECT 1370.500 2.400 1370.640 17.270 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1081.070 182.820 1081.390 182.880 ;
        RECT 1386.970 182.820 1387.290 182.880 ;
        RECT 1081.070 182.680 1387.290 182.820 ;
        RECT 1081.070 182.620 1081.390 182.680 ;
        RECT 1386.970 182.620 1387.290 182.680 ;
      LAYER via ;
        RECT 1081.100 182.620 1081.360 182.880 ;
        RECT 1387.000 182.620 1387.260 182.880 ;
      LAYER met2 ;
        RECT 1081.050 216.000 1081.330 220.000 ;
        RECT 1081.160 182.910 1081.300 216.000 ;
        RECT 1081.100 182.590 1081.360 182.910 ;
        RECT 1387.000 182.590 1387.260 182.910 ;
        RECT 1387.060 16.730 1387.200 182.590 ;
        RECT 1387.060 16.590 1388.580 16.730 ;
        RECT 1388.440 2.400 1388.580 16.590 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1099.010 190.300 1099.330 190.360 ;
        RECT 1400.770 190.300 1401.090 190.360 ;
        RECT 1099.010 190.160 1401.090 190.300 ;
        RECT 1099.010 190.100 1099.330 190.160 ;
        RECT 1400.770 190.100 1401.090 190.160 ;
      LAYER via ;
        RECT 1099.040 190.100 1099.300 190.360 ;
        RECT 1400.800 190.100 1401.060 190.360 ;
      LAYER met2 ;
        RECT 1098.990 216.000 1099.270 220.000 ;
        RECT 1099.100 190.390 1099.240 216.000 ;
        RECT 1099.040 190.070 1099.300 190.390 ;
        RECT 1400.800 190.070 1401.060 190.390 ;
        RECT 1400.860 16.730 1401.000 190.070 ;
        RECT 1400.860 16.590 1406.520 16.730 ;
        RECT 1406.380 2.400 1406.520 16.590 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1116.950 148.480 1117.270 148.540 ;
        RECT 1421.470 148.480 1421.790 148.540 ;
        RECT 1116.950 148.340 1421.790 148.480 ;
        RECT 1116.950 148.280 1117.270 148.340 ;
        RECT 1421.470 148.280 1421.790 148.340 ;
      LAYER via ;
        RECT 1116.980 148.280 1117.240 148.540 ;
        RECT 1421.500 148.280 1421.760 148.540 ;
      LAYER met2 ;
        RECT 1116.930 216.000 1117.210 220.000 ;
        RECT 1117.040 148.570 1117.180 216.000 ;
        RECT 1116.980 148.250 1117.240 148.570 ;
        RECT 1421.500 148.250 1421.760 148.570 ;
        RECT 1421.560 16.730 1421.700 148.250 ;
        RECT 1421.560 16.590 1424.000 16.730 ;
        RECT 1423.860 2.400 1424.000 16.590 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1134.890 197.100 1135.210 197.160 ;
        RECT 1435.270 197.100 1435.590 197.160 ;
        RECT 1134.890 196.960 1435.590 197.100 ;
        RECT 1134.890 196.900 1135.210 196.960 ;
        RECT 1435.270 196.900 1435.590 196.960 ;
        RECT 1435.270 16.560 1435.590 16.620 ;
        RECT 1441.710 16.560 1442.030 16.620 ;
        RECT 1435.270 16.420 1442.030 16.560 ;
        RECT 1435.270 16.360 1435.590 16.420 ;
        RECT 1441.710 16.360 1442.030 16.420 ;
      LAYER via ;
        RECT 1134.920 196.900 1135.180 197.160 ;
        RECT 1435.300 196.900 1435.560 197.160 ;
        RECT 1435.300 16.360 1435.560 16.620 ;
        RECT 1441.740 16.360 1442.000 16.620 ;
      LAYER met2 ;
        RECT 1134.870 216.000 1135.150 220.000 ;
        RECT 1134.980 197.190 1135.120 216.000 ;
        RECT 1134.920 196.870 1135.180 197.190 ;
        RECT 1435.300 196.870 1435.560 197.190 ;
        RECT 1435.360 16.650 1435.500 196.870 ;
        RECT 1435.300 16.330 1435.560 16.650 ;
        RECT 1441.740 16.330 1442.000 16.650 ;
        RECT 1441.800 2.400 1441.940 16.330 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1152.830 200.500 1153.150 200.560 ;
        RECT 1158.350 200.500 1158.670 200.560 ;
        RECT 1152.830 200.360 1158.670 200.500 ;
        RECT 1152.830 200.300 1153.150 200.360 ;
        RECT 1158.350 200.300 1158.670 200.360 ;
        RECT 1158.350 155.280 1158.670 155.340 ;
        RECT 1455.970 155.280 1456.290 155.340 ;
        RECT 1158.350 155.140 1456.290 155.280 ;
        RECT 1158.350 155.080 1158.670 155.140 ;
        RECT 1455.970 155.080 1456.290 155.140 ;
      LAYER via ;
        RECT 1152.860 200.300 1153.120 200.560 ;
        RECT 1158.380 200.300 1158.640 200.560 ;
        RECT 1158.380 155.080 1158.640 155.340 ;
        RECT 1456.000 155.080 1456.260 155.340 ;
      LAYER met2 ;
        RECT 1152.810 216.000 1153.090 220.000 ;
        RECT 1152.920 200.590 1153.060 216.000 ;
        RECT 1152.860 200.270 1153.120 200.590 ;
        RECT 1158.380 200.270 1158.640 200.590 ;
        RECT 1158.440 155.370 1158.580 200.270 ;
        RECT 1158.380 155.050 1158.640 155.370 ;
        RECT 1456.000 155.050 1456.260 155.370 ;
        RECT 1456.060 17.410 1456.200 155.050 ;
        RECT 1456.060 17.270 1459.880 17.410 ;
        RECT 1459.740 2.400 1459.880 17.270 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1172.610 162.080 1172.930 162.140 ;
        RECT 1476.670 162.080 1476.990 162.140 ;
        RECT 1172.610 161.940 1476.990 162.080 ;
        RECT 1172.610 161.880 1172.930 161.940 ;
        RECT 1476.670 161.880 1476.990 161.940 ;
      LAYER via ;
        RECT 1172.640 161.880 1172.900 162.140 ;
        RECT 1476.700 161.880 1476.960 162.140 ;
      LAYER met2 ;
        RECT 1170.750 216.650 1171.030 220.000 ;
        RECT 1170.750 216.510 1172.840 216.650 ;
        RECT 1170.750 216.000 1171.030 216.510 ;
        RECT 1172.700 162.170 1172.840 216.510 ;
        RECT 1172.640 161.850 1172.900 162.170 ;
        RECT 1476.700 161.850 1476.960 162.170 ;
        RECT 1476.760 17.410 1476.900 161.850 ;
        RECT 1476.760 17.270 1477.820 17.410 ;
        RECT 1477.680 2.400 1477.820 17.270 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1188.710 200.500 1189.030 200.560 ;
        RECT 1193.310 200.500 1193.630 200.560 ;
        RECT 1188.710 200.360 1193.630 200.500 ;
        RECT 1188.710 200.300 1189.030 200.360 ;
        RECT 1193.310 200.300 1193.630 200.360 ;
        RECT 1193.310 169.560 1193.630 169.620 ;
        RECT 1490.470 169.560 1490.790 169.620 ;
        RECT 1193.310 169.420 1490.790 169.560 ;
        RECT 1193.310 169.360 1193.630 169.420 ;
        RECT 1490.470 169.360 1490.790 169.420 ;
      LAYER via ;
        RECT 1188.740 200.300 1189.000 200.560 ;
        RECT 1193.340 200.300 1193.600 200.560 ;
        RECT 1193.340 169.360 1193.600 169.620 ;
        RECT 1490.500 169.360 1490.760 169.620 ;
      LAYER met2 ;
        RECT 1188.690 216.000 1188.970 220.000 ;
        RECT 1188.800 200.590 1188.940 216.000 ;
        RECT 1188.740 200.270 1189.000 200.590 ;
        RECT 1193.340 200.270 1193.600 200.590 ;
        RECT 1193.400 169.650 1193.540 200.270 ;
        RECT 1193.340 169.330 1193.600 169.650 ;
        RECT 1490.500 169.330 1490.760 169.650 ;
        RECT 1490.560 16.730 1490.700 169.330 ;
        RECT 1490.560 16.590 1495.760 16.730 ;
        RECT 1495.620 2.400 1495.760 16.590 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1206.650 176.020 1206.970 176.080 ;
        RECT 1511.170 176.020 1511.490 176.080 ;
        RECT 1206.650 175.880 1511.490 176.020 ;
        RECT 1206.650 175.820 1206.970 175.880 ;
        RECT 1511.170 175.820 1511.490 175.880 ;
      LAYER via ;
        RECT 1206.680 175.820 1206.940 176.080 ;
        RECT 1511.200 175.820 1511.460 176.080 ;
      LAYER met2 ;
        RECT 1206.630 216.000 1206.910 220.000 ;
        RECT 1206.740 176.110 1206.880 216.000 ;
        RECT 1206.680 175.790 1206.940 176.110 ;
        RECT 1511.200 175.790 1511.460 176.110 ;
        RECT 1511.260 16.730 1511.400 175.790 ;
        RECT 1511.260 16.590 1513.240 16.730 ;
        RECT 1513.100 2.400 1513.240 16.590 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 402.110 202.540 402.430 202.600 ;
        RECT 406.710 202.540 407.030 202.600 ;
        RECT 402.110 202.400 407.030 202.540 ;
        RECT 402.110 202.340 402.430 202.400 ;
        RECT 406.710 202.340 407.030 202.400 ;
        RECT 406.710 72.660 407.030 72.720 ;
        RECT 704.330 72.660 704.650 72.720 ;
        RECT 406.710 72.520 704.650 72.660 ;
        RECT 406.710 72.460 407.030 72.520 ;
        RECT 704.330 72.460 704.650 72.520 ;
        RECT 704.330 17.920 704.650 17.980 ;
        RECT 710.310 17.920 710.630 17.980 ;
        RECT 704.330 17.780 710.630 17.920 ;
        RECT 704.330 17.720 704.650 17.780 ;
        RECT 710.310 17.720 710.630 17.780 ;
      LAYER via ;
        RECT 402.140 202.340 402.400 202.600 ;
        RECT 406.740 202.340 407.000 202.600 ;
        RECT 406.740 72.460 407.000 72.720 ;
        RECT 704.360 72.460 704.620 72.720 ;
        RECT 704.360 17.720 704.620 17.980 ;
        RECT 710.340 17.720 710.600 17.980 ;
      LAYER met2 ;
        RECT 402.090 216.000 402.370 220.000 ;
        RECT 402.200 202.630 402.340 216.000 ;
        RECT 402.140 202.310 402.400 202.630 ;
        RECT 406.740 202.310 407.000 202.630 ;
        RECT 406.800 72.750 406.940 202.310 ;
        RECT 406.740 72.430 407.000 72.750 ;
        RECT 704.360 72.430 704.620 72.750 ;
        RECT 704.420 18.010 704.560 72.430 ;
        RECT 704.360 17.690 704.620 18.010 ;
        RECT 710.340 17.690 710.600 18.010 ;
        RECT 710.400 2.400 710.540 17.690 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1224.130 183.500 1224.450 183.560 ;
        RECT 1524.970 183.500 1525.290 183.560 ;
        RECT 1224.130 183.360 1525.290 183.500 ;
        RECT 1224.130 183.300 1224.450 183.360 ;
        RECT 1524.970 183.300 1525.290 183.360 ;
        RECT 1524.970 17.580 1525.290 17.640 ;
        RECT 1530.950 17.580 1531.270 17.640 ;
        RECT 1524.970 17.440 1531.270 17.580 ;
        RECT 1524.970 17.380 1525.290 17.440 ;
        RECT 1530.950 17.380 1531.270 17.440 ;
      LAYER via ;
        RECT 1224.160 183.300 1224.420 183.560 ;
        RECT 1525.000 183.300 1525.260 183.560 ;
        RECT 1525.000 17.380 1525.260 17.640 ;
        RECT 1530.980 17.380 1531.240 17.640 ;
      LAYER met2 ;
        RECT 1224.110 216.000 1224.390 220.000 ;
        RECT 1224.220 183.590 1224.360 216.000 ;
        RECT 1224.160 183.270 1224.420 183.590 ;
        RECT 1525.000 183.270 1525.260 183.590 ;
        RECT 1525.060 17.670 1525.200 183.270 ;
        RECT 1525.000 17.350 1525.260 17.670 ;
        RECT 1530.980 17.350 1531.240 17.670 ;
        RECT 1531.040 2.400 1531.180 17.350 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1243.450 189.620 1243.770 189.680 ;
        RECT 1545.670 189.620 1545.990 189.680 ;
        RECT 1243.450 189.480 1545.990 189.620 ;
        RECT 1243.450 189.420 1243.770 189.480 ;
        RECT 1545.670 189.420 1545.990 189.480 ;
      LAYER via ;
        RECT 1243.480 189.420 1243.740 189.680 ;
        RECT 1545.700 189.420 1545.960 189.680 ;
      LAYER met2 ;
        RECT 1242.050 216.650 1242.330 220.000 ;
        RECT 1242.050 216.510 1243.680 216.650 ;
        RECT 1242.050 216.000 1242.330 216.510 ;
        RECT 1243.540 189.710 1243.680 216.510 ;
        RECT 1243.480 189.390 1243.740 189.710 ;
        RECT 1545.700 189.390 1545.960 189.710 ;
        RECT 1545.760 16.730 1545.900 189.390 ;
        RECT 1545.760 16.590 1549.120 16.730 ;
        RECT 1548.980 2.400 1549.120 16.590 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1262.310 24.040 1262.630 24.100 ;
        RECT 1566.830 24.040 1567.150 24.100 ;
        RECT 1262.310 23.900 1567.150 24.040 ;
        RECT 1262.310 23.840 1262.630 23.900 ;
        RECT 1566.830 23.840 1567.150 23.900 ;
      LAYER via ;
        RECT 1262.340 23.840 1262.600 24.100 ;
        RECT 1566.860 23.840 1567.120 24.100 ;
      LAYER met2 ;
        RECT 1259.990 216.650 1260.270 220.000 ;
        RECT 1259.990 216.510 1262.540 216.650 ;
        RECT 1259.990 216.000 1260.270 216.510 ;
        RECT 1262.400 24.130 1262.540 216.510 ;
        RECT 1262.340 23.810 1262.600 24.130 ;
        RECT 1566.860 23.810 1567.120 24.130 ;
        RECT 1566.920 2.400 1567.060 23.810 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1277.950 203.220 1278.270 203.280 ;
        RECT 1283.010 203.220 1283.330 203.280 ;
        RECT 1277.950 203.080 1283.330 203.220 ;
        RECT 1277.950 203.020 1278.270 203.080 ;
        RECT 1283.010 203.020 1283.330 203.080 ;
        RECT 1283.010 148.820 1283.330 148.880 ;
        RECT 1580.170 148.820 1580.490 148.880 ;
        RECT 1283.010 148.680 1580.490 148.820 ;
        RECT 1283.010 148.620 1283.330 148.680 ;
        RECT 1580.170 148.620 1580.490 148.680 ;
      LAYER via ;
        RECT 1277.980 203.020 1278.240 203.280 ;
        RECT 1283.040 203.020 1283.300 203.280 ;
        RECT 1283.040 148.620 1283.300 148.880 ;
        RECT 1580.200 148.620 1580.460 148.880 ;
      LAYER met2 ;
        RECT 1277.930 216.000 1278.210 220.000 ;
        RECT 1278.040 203.310 1278.180 216.000 ;
        RECT 1277.980 202.990 1278.240 203.310 ;
        RECT 1283.040 202.990 1283.300 203.310 ;
        RECT 1283.100 148.910 1283.240 202.990 ;
        RECT 1283.040 148.590 1283.300 148.910 ;
        RECT 1580.200 148.590 1580.460 148.910 ;
        RECT 1580.260 16.730 1580.400 148.590 ;
        RECT 1580.260 16.590 1585.000 16.730 ;
        RECT 1584.860 2.400 1585.000 16.590 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1295.890 196.760 1296.210 196.820 ;
        RECT 1600.870 196.760 1601.190 196.820 ;
        RECT 1295.890 196.620 1601.190 196.760 ;
        RECT 1295.890 196.560 1296.210 196.620 ;
        RECT 1600.870 196.560 1601.190 196.620 ;
      LAYER via ;
        RECT 1295.920 196.560 1296.180 196.820 ;
        RECT 1600.900 196.560 1601.160 196.820 ;
      LAYER met2 ;
        RECT 1295.870 216.000 1296.150 220.000 ;
        RECT 1295.980 196.850 1296.120 216.000 ;
        RECT 1295.920 196.530 1296.180 196.850 ;
        RECT 1600.900 196.530 1601.160 196.850 ;
        RECT 1600.960 16.730 1601.100 196.530 ;
        RECT 1600.960 16.590 1602.480 16.730 ;
        RECT 1602.340 2.400 1602.480 16.590 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1313.830 200.500 1314.150 200.560 ;
        RECT 1317.510 200.500 1317.830 200.560 ;
        RECT 1313.830 200.360 1317.830 200.500 ;
        RECT 1313.830 200.300 1314.150 200.360 ;
        RECT 1317.510 200.300 1317.830 200.360 ;
        RECT 1317.510 155.620 1317.830 155.680 ;
        RECT 1614.670 155.620 1614.990 155.680 ;
        RECT 1317.510 155.480 1614.990 155.620 ;
        RECT 1317.510 155.420 1317.830 155.480 ;
        RECT 1614.670 155.420 1614.990 155.480 ;
      LAYER via ;
        RECT 1313.860 200.300 1314.120 200.560 ;
        RECT 1317.540 200.300 1317.800 200.560 ;
        RECT 1317.540 155.420 1317.800 155.680 ;
        RECT 1614.700 155.420 1614.960 155.680 ;
      LAYER met2 ;
        RECT 1313.810 216.000 1314.090 220.000 ;
        RECT 1313.920 200.590 1314.060 216.000 ;
        RECT 1313.860 200.270 1314.120 200.590 ;
        RECT 1317.540 200.270 1317.800 200.590 ;
        RECT 1317.600 155.710 1317.740 200.270 ;
        RECT 1317.540 155.390 1317.800 155.710 ;
        RECT 1614.700 155.390 1614.960 155.710 ;
        RECT 1614.760 16.730 1614.900 155.390 ;
        RECT 1614.760 16.590 1620.420 16.730 ;
        RECT 1620.280 2.400 1620.420 16.590 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1332.690 162.760 1333.010 162.820 ;
        RECT 1635.370 162.760 1635.690 162.820 ;
        RECT 1332.690 162.620 1635.690 162.760 ;
        RECT 1332.690 162.560 1333.010 162.620 ;
        RECT 1635.370 162.560 1635.690 162.620 ;
      LAYER via ;
        RECT 1332.720 162.560 1332.980 162.820 ;
        RECT 1635.400 162.560 1635.660 162.820 ;
      LAYER met2 ;
        RECT 1331.750 216.000 1332.030 220.000 ;
        RECT 1331.860 184.690 1332.000 216.000 ;
        RECT 1331.860 184.550 1332.920 184.690 ;
        RECT 1332.780 162.850 1332.920 184.550 ;
        RECT 1332.720 162.530 1332.980 162.850 ;
        RECT 1635.400 162.530 1635.660 162.850 ;
        RECT 1635.460 16.730 1635.600 162.530 ;
        RECT 1635.460 16.590 1638.360 16.730 ;
        RECT 1638.220 2.400 1638.360 16.590 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.010 168.880 1352.330 168.940 ;
        RECT 1656.070 168.880 1656.390 168.940 ;
        RECT 1352.010 168.740 1656.390 168.880 ;
        RECT 1352.010 168.680 1352.330 168.740 ;
        RECT 1656.070 168.680 1656.390 168.740 ;
      LAYER via ;
        RECT 1352.040 168.680 1352.300 168.940 ;
        RECT 1656.100 168.680 1656.360 168.940 ;
      LAYER met2 ;
        RECT 1349.230 216.650 1349.510 220.000 ;
        RECT 1349.230 216.510 1352.240 216.650 ;
        RECT 1349.230 216.000 1349.510 216.510 ;
        RECT 1352.100 168.970 1352.240 216.510 ;
        RECT 1352.040 168.650 1352.300 168.970 ;
        RECT 1656.100 168.650 1656.360 168.970 ;
        RECT 1656.160 2.400 1656.300 168.650 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1367.190 176.700 1367.510 176.760 ;
        RECT 1669.870 176.700 1670.190 176.760 ;
        RECT 1367.190 176.560 1670.190 176.700 ;
        RECT 1367.190 176.500 1367.510 176.560 ;
        RECT 1669.870 176.500 1670.190 176.560 ;
      LAYER via ;
        RECT 1367.220 176.500 1367.480 176.760 ;
        RECT 1669.900 176.500 1670.160 176.760 ;
      LAYER met2 ;
        RECT 1367.170 216.000 1367.450 220.000 ;
        RECT 1367.280 176.790 1367.420 216.000 ;
        RECT 1367.220 176.470 1367.480 176.790 ;
        RECT 1669.900 176.470 1670.160 176.790 ;
        RECT 1669.960 16.730 1670.100 176.470 ;
        RECT 1669.960 16.590 1673.780 16.730 ;
        RECT 1673.640 2.400 1673.780 16.590 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1385.130 183.160 1385.450 183.220 ;
        RECT 1690.570 183.160 1690.890 183.220 ;
        RECT 1385.130 183.020 1690.890 183.160 ;
        RECT 1385.130 182.960 1385.450 183.020 ;
        RECT 1690.570 182.960 1690.890 183.020 ;
      LAYER via ;
        RECT 1385.160 182.960 1385.420 183.220 ;
        RECT 1690.600 182.960 1690.860 183.220 ;
      LAYER met2 ;
        RECT 1385.110 216.000 1385.390 220.000 ;
        RECT 1385.220 183.250 1385.360 216.000 ;
        RECT 1385.160 182.930 1385.420 183.250 ;
        RECT 1690.600 182.930 1690.860 183.250 ;
        RECT 1690.660 17.410 1690.800 182.930 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 420.510 65.860 420.830 65.920 ;
        RECT 724.570 65.860 724.890 65.920 ;
        RECT 420.510 65.720 724.890 65.860 ;
        RECT 420.510 65.660 420.830 65.720 ;
        RECT 724.570 65.660 724.890 65.720 ;
      LAYER via ;
        RECT 420.540 65.660 420.800 65.920 ;
        RECT 724.600 65.660 724.860 65.920 ;
      LAYER met2 ;
        RECT 420.030 216.650 420.310 220.000 ;
        RECT 420.030 216.510 420.740 216.650 ;
        RECT 420.030 216.000 420.310 216.510 ;
        RECT 420.600 65.950 420.740 216.510 ;
        RECT 420.540 65.630 420.800 65.950 ;
        RECT 724.600 65.630 724.860 65.950 ;
        RECT 724.660 16.730 724.800 65.630 ;
        RECT 724.660 16.590 728.480 16.730 ;
        RECT 728.340 2.400 728.480 16.590 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1403.070 189.960 1403.390 190.020 ;
        RECT 1704.370 189.960 1704.690 190.020 ;
        RECT 1403.070 189.820 1704.690 189.960 ;
        RECT 1403.070 189.760 1403.390 189.820 ;
        RECT 1704.370 189.760 1704.690 189.820 ;
      LAYER via ;
        RECT 1403.100 189.760 1403.360 190.020 ;
        RECT 1704.400 189.760 1704.660 190.020 ;
      LAYER met2 ;
        RECT 1403.050 216.000 1403.330 220.000 ;
        RECT 1403.160 190.050 1403.300 216.000 ;
        RECT 1403.100 189.730 1403.360 190.050 ;
        RECT 1704.400 189.730 1704.660 190.050 ;
        RECT 1704.460 17.410 1704.600 189.730 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1420.550 148.140 1420.870 148.200 ;
        RECT 1725.070 148.140 1725.390 148.200 ;
        RECT 1420.550 148.000 1725.390 148.140 ;
        RECT 1420.550 147.940 1420.870 148.000 ;
        RECT 1725.070 147.940 1725.390 148.000 ;
      LAYER via ;
        RECT 1420.580 147.940 1420.840 148.200 ;
        RECT 1725.100 147.940 1725.360 148.200 ;
      LAYER met2 ;
        RECT 1420.990 216.650 1421.270 220.000 ;
        RECT 1420.640 216.510 1421.270 216.650 ;
        RECT 1420.640 148.230 1420.780 216.510 ;
        RECT 1420.990 216.000 1421.270 216.510 ;
        RECT 1420.580 147.910 1420.840 148.230 ;
        RECT 1725.100 147.910 1725.360 148.230 ;
        RECT 1725.160 17.410 1725.300 147.910 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1438.950 197.440 1439.270 197.500 ;
        RECT 1738.870 197.440 1739.190 197.500 ;
        RECT 1438.950 197.300 1739.190 197.440 ;
        RECT 1438.950 197.240 1439.270 197.300 ;
        RECT 1738.870 197.240 1739.190 197.300 ;
        RECT 1738.870 17.240 1739.190 17.300 ;
        RECT 1745.310 17.240 1745.630 17.300 ;
        RECT 1738.870 17.100 1745.630 17.240 ;
        RECT 1738.870 17.040 1739.190 17.100 ;
        RECT 1745.310 17.040 1745.630 17.100 ;
      LAYER via ;
        RECT 1438.980 197.240 1439.240 197.500 ;
        RECT 1738.900 197.240 1739.160 197.500 ;
        RECT 1738.900 17.040 1739.160 17.300 ;
        RECT 1745.340 17.040 1745.600 17.300 ;
      LAYER met2 ;
        RECT 1438.930 216.000 1439.210 220.000 ;
        RECT 1439.040 197.530 1439.180 216.000 ;
        RECT 1438.980 197.210 1439.240 197.530 ;
        RECT 1738.900 197.210 1739.160 197.530 ;
        RECT 1738.960 17.330 1739.100 197.210 ;
        RECT 1738.900 17.010 1739.160 17.330 ;
        RECT 1745.340 17.010 1745.600 17.330 ;
        RECT 1745.400 2.400 1745.540 17.010 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1456.890 200.500 1457.210 200.560 ;
        RECT 1462.410 200.500 1462.730 200.560 ;
        RECT 1456.890 200.360 1462.730 200.500 ;
        RECT 1456.890 200.300 1457.210 200.360 ;
        RECT 1462.410 200.300 1462.730 200.360 ;
        RECT 1462.410 155.280 1462.730 155.340 ;
        RECT 1759.570 155.280 1759.890 155.340 ;
        RECT 1462.410 155.140 1759.890 155.280 ;
        RECT 1462.410 155.080 1462.730 155.140 ;
        RECT 1759.570 155.080 1759.890 155.140 ;
      LAYER via ;
        RECT 1456.920 200.300 1457.180 200.560 ;
        RECT 1462.440 200.300 1462.700 200.560 ;
        RECT 1462.440 155.080 1462.700 155.340 ;
        RECT 1759.600 155.080 1759.860 155.340 ;
      LAYER met2 ;
        RECT 1456.870 216.000 1457.150 220.000 ;
        RECT 1456.980 200.590 1457.120 216.000 ;
        RECT 1456.920 200.270 1457.180 200.590 ;
        RECT 1462.440 200.270 1462.700 200.590 ;
        RECT 1462.500 155.370 1462.640 200.270 ;
        RECT 1462.440 155.050 1462.700 155.370 ;
        RECT 1759.600 155.050 1759.860 155.370 ;
        RECT 1759.660 17.410 1759.800 155.050 ;
        RECT 1759.660 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1476.210 162.420 1476.530 162.480 ;
        RECT 1780.730 162.420 1781.050 162.480 ;
        RECT 1476.210 162.280 1781.050 162.420 ;
        RECT 1476.210 162.220 1476.530 162.280 ;
        RECT 1780.730 162.220 1781.050 162.280 ;
      LAYER via ;
        RECT 1476.240 162.220 1476.500 162.480 ;
        RECT 1780.760 162.220 1781.020 162.480 ;
      LAYER met2 ;
        RECT 1474.350 216.650 1474.630 220.000 ;
        RECT 1474.350 216.510 1476.440 216.650 ;
        RECT 1474.350 216.000 1474.630 216.510 ;
        RECT 1476.300 162.510 1476.440 216.510 ;
        RECT 1476.240 162.190 1476.500 162.510 ;
        RECT 1780.760 162.190 1781.020 162.510 ;
        RECT 1780.820 2.400 1780.960 162.190 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1492.310 169.220 1492.630 169.280 ;
        RECT 1794.070 169.220 1794.390 169.280 ;
        RECT 1492.310 169.080 1794.390 169.220 ;
        RECT 1492.310 169.020 1492.630 169.080 ;
        RECT 1794.070 169.020 1794.390 169.080 ;
      LAYER via ;
        RECT 1492.340 169.020 1492.600 169.280 ;
        RECT 1794.100 169.020 1794.360 169.280 ;
      LAYER met2 ;
        RECT 1492.290 216.000 1492.570 220.000 ;
        RECT 1492.400 169.310 1492.540 216.000 ;
        RECT 1492.340 168.990 1492.600 169.310 ;
        RECT 1794.100 168.990 1794.360 169.310 ;
        RECT 1794.160 16.730 1794.300 168.990 ;
        RECT 1794.160 16.590 1798.900 16.730 ;
        RECT 1798.760 2.400 1798.900 16.590 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1510.250 176.360 1510.570 176.420 ;
        RECT 1814.770 176.360 1815.090 176.420 ;
        RECT 1510.250 176.220 1815.090 176.360 ;
        RECT 1510.250 176.160 1510.570 176.220 ;
        RECT 1814.770 176.160 1815.090 176.220 ;
      LAYER via ;
        RECT 1510.280 176.160 1510.540 176.420 ;
        RECT 1814.800 176.160 1815.060 176.420 ;
      LAYER met2 ;
        RECT 1510.230 216.000 1510.510 220.000 ;
        RECT 1510.340 176.450 1510.480 216.000 ;
        RECT 1510.280 176.130 1510.540 176.450 ;
        RECT 1814.800 176.130 1815.060 176.450 ;
        RECT 1814.860 16.730 1815.000 176.130 ;
        RECT 1814.860 16.590 1816.840 16.730 ;
        RECT 1816.700 2.400 1816.840 16.590 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1528.190 183.500 1528.510 183.560 ;
        RECT 1828.570 183.500 1828.890 183.560 ;
        RECT 1528.190 183.360 1828.890 183.500 ;
        RECT 1528.190 183.300 1528.510 183.360 ;
        RECT 1828.570 183.300 1828.890 183.360 ;
        RECT 1828.570 17.580 1828.890 17.640 ;
        RECT 1834.550 17.580 1834.870 17.640 ;
        RECT 1828.570 17.440 1834.870 17.580 ;
        RECT 1828.570 17.380 1828.890 17.440 ;
        RECT 1834.550 17.380 1834.870 17.440 ;
      LAYER via ;
        RECT 1528.220 183.300 1528.480 183.560 ;
        RECT 1828.600 183.300 1828.860 183.560 ;
        RECT 1828.600 17.380 1828.860 17.640 ;
        RECT 1834.580 17.380 1834.840 17.640 ;
      LAYER met2 ;
        RECT 1528.170 216.000 1528.450 220.000 ;
        RECT 1528.280 183.590 1528.420 216.000 ;
        RECT 1528.220 183.270 1528.480 183.590 ;
        RECT 1828.600 183.270 1828.860 183.590 ;
        RECT 1828.660 17.670 1828.800 183.270 ;
        RECT 1828.600 17.350 1828.860 17.670 ;
        RECT 1834.580 17.350 1834.840 17.670 ;
        RECT 1834.640 2.400 1834.780 17.350 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1546.130 200.500 1546.450 200.560 ;
        RECT 1555.790 200.500 1556.110 200.560 ;
        RECT 1546.130 200.360 1556.110 200.500 ;
        RECT 1546.130 200.300 1546.450 200.360 ;
        RECT 1555.790 200.300 1556.110 200.360 ;
        RECT 1555.790 52.260 1556.110 52.320 ;
        RECT 1849.270 52.260 1849.590 52.320 ;
        RECT 1555.790 52.120 1849.590 52.260 ;
        RECT 1555.790 52.060 1556.110 52.120 ;
        RECT 1849.270 52.060 1849.590 52.120 ;
      LAYER via ;
        RECT 1546.160 200.300 1546.420 200.560 ;
        RECT 1555.820 200.300 1556.080 200.560 ;
        RECT 1555.820 52.060 1556.080 52.320 ;
        RECT 1849.300 52.060 1849.560 52.320 ;
      LAYER met2 ;
        RECT 1546.110 216.000 1546.390 220.000 ;
        RECT 1546.220 200.590 1546.360 216.000 ;
        RECT 1546.160 200.270 1546.420 200.590 ;
        RECT 1555.820 200.270 1556.080 200.590 ;
        RECT 1555.880 52.350 1556.020 200.270 ;
        RECT 1555.820 52.030 1556.080 52.350 ;
        RECT 1849.300 52.030 1849.560 52.350 ;
        RECT 1849.360 16.730 1849.500 52.030 ;
        RECT 1849.360 16.590 1852.260 16.730 ;
        RECT 1852.120 2.400 1852.260 16.590 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1564.070 189.620 1564.390 189.680 ;
        RECT 1870.430 189.620 1870.750 189.680 ;
        RECT 1564.070 189.480 1870.750 189.620 ;
        RECT 1564.070 189.420 1564.390 189.480 ;
        RECT 1870.430 189.420 1870.750 189.480 ;
      LAYER via ;
        RECT 1564.100 189.420 1564.360 189.680 ;
        RECT 1870.460 189.420 1870.720 189.680 ;
      LAYER met2 ;
        RECT 1564.050 216.000 1564.330 220.000 ;
        RECT 1564.160 189.710 1564.300 216.000 ;
        RECT 1564.100 189.390 1564.360 189.710 ;
        RECT 1870.460 189.390 1870.720 189.710 ;
        RECT 1870.520 17.410 1870.660 189.390 ;
        RECT 1870.060 17.270 1870.660 17.410 ;
        RECT 1870.060 2.400 1870.200 17.270 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 441.210 19.620 441.530 19.680 ;
        RECT 746.190 19.620 746.510 19.680 ;
        RECT 441.210 19.480 746.510 19.620 ;
        RECT 441.210 19.420 441.530 19.480 ;
        RECT 746.190 19.420 746.510 19.480 ;
      LAYER via ;
        RECT 441.240 19.420 441.500 19.680 ;
        RECT 746.220 19.420 746.480 19.680 ;
      LAYER met2 ;
        RECT 437.970 216.650 438.250 220.000 ;
        RECT 437.970 216.510 441.440 216.650 ;
        RECT 437.970 216.000 438.250 216.510 ;
        RECT 441.300 19.710 441.440 216.510 ;
        RECT 441.240 19.390 441.500 19.710 ;
        RECT 746.220 19.390 746.480 19.710 ;
        RECT 746.280 2.400 746.420 19.390 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1582.010 200.500 1582.330 200.560 ;
        RECT 1586.610 200.500 1586.930 200.560 ;
        RECT 1582.010 200.360 1586.930 200.500 ;
        RECT 1582.010 200.300 1582.330 200.360 ;
        RECT 1586.610 200.300 1586.930 200.360 ;
        RECT 1586.610 128.080 1586.930 128.140 ;
        RECT 1883.770 128.080 1884.090 128.140 ;
        RECT 1586.610 127.940 1884.090 128.080 ;
        RECT 1586.610 127.880 1586.930 127.940 ;
        RECT 1883.770 127.880 1884.090 127.940 ;
        RECT 1883.770 2.960 1884.090 3.020 ;
        RECT 1887.910 2.960 1888.230 3.020 ;
        RECT 1883.770 2.820 1888.230 2.960 ;
        RECT 1883.770 2.760 1884.090 2.820 ;
        RECT 1887.910 2.760 1888.230 2.820 ;
      LAYER via ;
        RECT 1582.040 200.300 1582.300 200.560 ;
        RECT 1586.640 200.300 1586.900 200.560 ;
        RECT 1586.640 127.880 1586.900 128.140 ;
        RECT 1883.800 127.880 1884.060 128.140 ;
        RECT 1883.800 2.760 1884.060 3.020 ;
        RECT 1887.940 2.760 1888.200 3.020 ;
      LAYER met2 ;
        RECT 1581.990 216.000 1582.270 220.000 ;
        RECT 1582.100 200.590 1582.240 216.000 ;
        RECT 1582.040 200.270 1582.300 200.590 ;
        RECT 1586.640 200.270 1586.900 200.590 ;
        RECT 1586.700 128.170 1586.840 200.270 ;
        RECT 1586.640 127.850 1586.900 128.170 ;
        RECT 1883.800 127.850 1884.060 128.170 ;
        RECT 1883.860 3.050 1884.000 127.850 ;
        RECT 1883.800 2.730 1884.060 3.050 ;
        RECT 1887.940 2.730 1888.200 3.050 ;
        RECT 1888.000 2.400 1888.140 2.730 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1599.490 197.100 1599.810 197.160 ;
        RECT 1904.470 197.100 1904.790 197.160 ;
        RECT 1599.490 196.960 1904.790 197.100 ;
        RECT 1599.490 196.900 1599.810 196.960 ;
        RECT 1904.470 196.900 1904.790 196.960 ;
      LAYER via ;
        RECT 1599.520 196.900 1599.780 197.160 ;
        RECT 1904.500 196.900 1904.760 197.160 ;
      LAYER met2 ;
        RECT 1599.470 216.000 1599.750 220.000 ;
        RECT 1599.580 197.190 1599.720 216.000 ;
        RECT 1599.520 196.870 1599.780 197.190 ;
        RECT 1904.500 196.870 1904.760 197.190 ;
        RECT 1904.560 3.130 1904.700 196.870 ;
        RECT 1904.560 2.990 1905.620 3.130 ;
        RECT 1905.480 2.960 1905.620 2.990 ;
        RECT 1905.480 2.820 1906.080 2.960 ;
        RECT 1905.940 2.400 1906.080 2.820 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1617.430 200.500 1617.750 200.560 ;
        RECT 1621.110 200.500 1621.430 200.560 ;
        RECT 1617.430 200.360 1621.430 200.500 ;
        RECT 1617.430 200.300 1617.750 200.360 ;
        RECT 1621.110 200.300 1621.430 200.360 ;
        RECT 1621.110 155.620 1621.430 155.680 ;
        RECT 1918.270 155.620 1918.590 155.680 ;
        RECT 1621.110 155.480 1918.590 155.620 ;
        RECT 1621.110 155.420 1621.430 155.480 ;
        RECT 1918.270 155.420 1918.590 155.480 ;
        RECT 1918.270 2.960 1918.590 3.020 ;
        RECT 1923.330 2.960 1923.650 3.020 ;
        RECT 1918.270 2.820 1923.650 2.960 ;
        RECT 1918.270 2.760 1918.590 2.820 ;
        RECT 1923.330 2.760 1923.650 2.820 ;
      LAYER via ;
        RECT 1617.460 200.300 1617.720 200.560 ;
        RECT 1621.140 200.300 1621.400 200.560 ;
        RECT 1621.140 155.420 1621.400 155.680 ;
        RECT 1918.300 155.420 1918.560 155.680 ;
        RECT 1918.300 2.760 1918.560 3.020 ;
        RECT 1923.360 2.760 1923.620 3.020 ;
      LAYER met2 ;
        RECT 1617.410 216.000 1617.690 220.000 ;
        RECT 1617.520 200.590 1617.660 216.000 ;
        RECT 1617.460 200.270 1617.720 200.590 ;
        RECT 1621.140 200.270 1621.400 200.590 ;
        RECT 1621.200 155.710 1621.340 200.270 ;
        RECT 1621.140 155.390 1621.400 155.710 ;
        RECT 1918.300 155.390 1918.560 155.710 ;
        RECT 1918.360 3.050 1918.500 155.390 ;
        RECT 1918.300 2.730 1918.560 3.050 ;
        RECT 1923.360 2.730 1923.620 3.050 ;
        RECT 1923.420 2.400 1923.560 2.730 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1635.370 200.500 1635.690 200.560 ;
        RECT 1641.350 200.500 1641.670 200.560 ;
        RECT 1635.370 200.360 1641.670 200.500 ;
        RECT 1635.370 200.300 1635.690 200.360 ;
        RECT 1641.350 200.300 1641.670 200.360 ;
        RECT 1641.350 162.080 1641.670 162.140 ;
        RECT 1938.970 162.080 1939.290 162.140 ;
        RECT 1641.350 161.940 1939.290 162.080 ;
        RECT 1641.350 161.880 1641.670 161.940 ;
        RECT 1938.970 161.880 1939.290 161.940 ;
        RECT 1938.970 2.960 1939.290 3.020 ;
        RECT 1941.270 2.960 1941.590 3.020 ;
        RECT 1938.970 2.820 1941.590 2.960 ;
        RECT 1938.970 2.760 1939.290 2.820 ;
        RECT 1941.270 2.760 1941.590 2.820 ;
      LAYER via ;
        RECT 1635.400 200.300 1635.660 200.560 ;
        RECT 1641.380 200.300 1641.640 200.560 ;
        RECT 1641.380 161.880 1641.640 162.140 ;
        RECT 1939.000 161.880 1939.260 162.140 ;
        RECT 1939.000 2.760 1939.260 3.020 ;
        RECT 1941.300 2.760 1941.560 3.020 ;
      LAYER met2 ;
        RECT 1635.350 216.000 1635.630 220.000 ;
        RECT 1635.460 200.590 1635.600 216.000 ;
        RECT 1635.400 200.270 1635.660 200.590 ;
        RECT 1641.380 200.270 1641.640 200.590 ;
        RECT 1641.440 162.170 1641.580 200.270 ;
        RECT 1641.380 161.850 1641.640 162.170 ;
        RECT 1939.000 161.850 1939.260 162.170 ;
        RECT 1939.060 3.050 1939.200 161.850 ;
        RECT 1939.000 2.730 1939.260 3.050 ;
        RECT 1941.300 2.730 1941.560 3.050 ;
        RECT 1941.360 2.400 1941.500 2.730 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.610 59.060 1655.930 59.120 ;
        RECT 1959.210 59.060 1959.530 59.120 ;
        RECT 1655.610 58.920 1959.530 59.060 ;
        RECT 1655.610 58.860 1655.930 58.920 ;
        RECT 1959.210 58.860 1959.530 58.920 ;
      LAYER via ;
        RECT 1655.640 58.860 1655.900 59.120 ;
        RECT 1959.240 58.860 1959.500 59.120 ;
      LAYER met2 ;
        RECT 1653.290 216.650 1653.570 220.000 ;
        RECT 1653.290 216.510 1655.840 216.650 ;
        RECT 1653.290 216.000 1653.570 216.510 ;
        RECT 1655.700 59.150 1655.840 216.510 ;
        RECT 1655.640 58.830 1655.900 59.150 ;
        RECT 1959.240 58.830 1959.500 59.150 ;
        RECT 1959.300 2.400 1959.440 58.830 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1977.225 48.365 1977.395 65.875 ;
      LAYER mcon ;
        RECT 1977.225 65.705 1977.395 65.875 ;
      LAYER met1 ;
        RECT 1671.250 203.900 1671.570 203.960 ;
        RECT 1838.690 203.900 1839.010 203.960 ;
        RECT 1671.250 203.760 1839.010 203.900 ;
        RECT 1671.250 203.700 1671.570 203.760 ;
        RECT 1838.690 203.700 1839.010 203.760 ;
        RECT 1838.690 65.860 1839.010 65.920 ;
        RECT 1977.165 65.860 1977.455 65.905 ;
        RECT 1838.690 65.720 1977.455 65.860 ;
        RECT 1838.690 65.660 1839.010 65.720 ;
        RECT 1977.165 65.675 1977.455 65.720 ;
        RECT 1977.150 48.520 1977.470 48.580 ;
        RECT 1976.955 48.380 1977.470 48.520 ;
        RECT 1977.150 48.320 1977.470 48.380 ;
      LAYER via ;
        RECT 1671.280 203.700 1671.540 203.960 ;
        RECT 1838.720 203.700 1838.980 203.960 ;
        RECT 1838.720 65.660 1838.980 65.920 ;
        RECT 1977.180 48.320 1977.440 48.580 ;
      LAYER met2 ;
        RECT 1671.230 216.000 1671.510 220.000 ;
        RECT 1671.340 203.990 1671.480 216.000 ;
        RECT 1671.280 203.670 1671.540 203.990 ;
        RECT 1838.720 203.670 1838.980 203.990 ;
        RECT 1838.780 65.950 1838.920 203.670 ;
        RECT 1838.720 65.630 1838.980 65.950 ;
        RECT 1977.180 48.290 1977.440 48.610 ;
        RECT 1977.240 2.400 1977.380 48.290 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1994.245 89.845 1994.415 137.955 ;
      LAYER mcon ;
        RECT 1994.245 137.785 1994.415 137.955 ;
      LAYER met1 ;
        RECT 1690.110 168.880 1690.430 168.940 ;
        RECT 1994.630 168.880 1994.950 168.940 ;
        RECT 1690.110 168.740 1994.950 168.880 ;
        RECT 1690.110 168.680 1690.430 168.740 ;
        RECT 1994.630 168.680 1994.950 168.740 ;
        RECT 1994.170 137.940 1994.490 138.000 ;
        RECT 1993.975 137.800 1994.490 137.940 ;
        RECT 1994.170 137.740 1994.490 137.800 ;
        RECT 1994.170 90.000 1994.490 90.060 ;
        RECT 1993.975 89.860 1994.490 90.000 ;
        RECT 1994.170 89.800 1994.490 89.860 ;
        RECT 1994.170 62.460 1994.490 62.520 ;
        RECT 1994.170 62.320 1995.320 62.460 ;
        RECT 1994.170 62.260 1994.490 62.320 ;
        RECT 1995.180 61.500 1995.320 62.320 ;
        RECT 1995.090 61.240 1995.410 61.500 ;
        RECT 1995.090 47.980 1995.410 48.240 ;
        RECT 1995.180 47.560 1995.320 47.980 ;
        RECT 1995.090 47.300 1995.410 47.560 ;
      LAYER via ;
        RECT 1690.140 168.680 1690.400 168.940 ;
        RECT 1994.660 168.680 1994.920 168.940 ;
        RECT 1994.200 137.740 1994.460 138.000 ;
        RECT 1994.200 89.800 1994.460 90.060 ;
        RECT 1994.200 62.260 1994.460 62.520 ;
        RECT 1995.120 61.240 1995.380 61.500 ;
        RECT 1995.120 47.980 1995.380 48.240 ;
        RECT 1995.120 47.300 1995.380 47.560 ;
      LAYER met2 ;
        RECT 1689.170 216.650 1689.450 220.000 ;
        RECT 1689.170 216.510 1690.340 216.650 ;
        RECT 1689.170 216.000 1689.450 216.510 ;
        RECT 1690.200 168.970 1690.340 216.510 ;
        RECT 1690.140 168.650 1690.400 168.970 ;
        RECT 1994.660 168.650 1994.920 168.970 ;
        RECT 1994.720 145.250 1994.860 168.650 ;
        RECT 1994.260 145.110 1994.860 145.250 ;
        RECT 1994.260 138.030 1994.400 145.110 ;
        RECT 1994.200 137.710 1994.460 138.030 ;
        RECT 1994.200 89.770 1994.460 90.090 ;
        RECT 1994.260 62.550 1994.400 89.770 ;
        RECT 1994.200 62.230 1994.460 62.550 ;
        RECT 1995.120 61.210 1995.380 61.530 ;
        RECT 1995.180 48.270 1995.320 61.210 ;
        RECT 1995.120 47.950 1995.380 48.270 ;
        RECT 1995.120 47.270 1995.380 47.590 ;
        RECT 1995.180 2.400 1995.320 47.270 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1710.810 176.020 1711.130 176.080 ;
        RECT 2007.970 176.020 2008.290 176.080 ;
        RECT 1710.810 175.880 2008.290 176.020 ;
        RECT 1710.810 175.820 1711.130 175.880 ;
        RECT 2007.970 175.820 2008.290 175.880 ;
        RECT 2007.970 62.120 2008.290 62.180 ;
        RECT 2012.570 62.120 2012.890 62.180 ;
        RECT 2007.970 61.980 2012.890 62.120 ;
        RECT 2007.970 61.920 2008.290 61.980 ;
        RECT 2012.570 61.920 2012.890 61.980 ;
      LAYER via ;
        RECT 1710.840 175.820 1711.100 176.080 ;
        RECT 2008.000 175.820 2008.260 176.080 ;
        RECT 2008.000 61.920 2008.260 62.180 ;
        RECT 2012.600 61.920 2012.860 62.180 ;
      LAYER met2 ;
        RECT 1707.110 216.650 1707.390 220.000 ;
        RECT 1707.110 216.510 1711.040 216.650 ;
        RECT 1707.110 216.000 1707.390 216.510 ;
        RECT 1710.900 176.110 1711.040 216.510 ;
        RECT 1710.840 175.790 1711.100 176.110 ;
        RECT 2008.000 175.790 2008.260 176.110 ;
        RECT 2008.060 62.210 2008.200 175.790 ;
        RECT 2008.000 61.890 2008.260 62.210 ;
        RECT 2012.600 61.890 2012.860 62.210 ;
        RECT 2012.660 2.400 2012.800 61.890 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2030.585 48.365 2030.755 72.335 ;
      LAYER mcon ;
        RECT 2030.585 72.165 2030.755 72.335 ;
      LAYER met1 ;
        RECT 1724.610 72.320 1724.930 72.380 ;
        RECT 2030.525 72.320 2030.815 72.365 ;
        RECT 1724.610 72.180 2030.815 72.320 ;
        RECT 1724.610 72.120 1724.930 72.180 ;
        RECT 2030.525 72.135 2030.815 72.180 ;
        RECT 2030.510 48.520 2030.830 48.580 ;
        RECT 2030.315 48.380 2030.830 48.520 ;
        RECT 2030.510 48.320 2030.830 48.380 ;
      LAYER via ;
        RECT 1724.640 72.120 1724.900 72.380 ;
        RECT 2030.540 48.320 2030.800 48.580 ;
      LAYER met2 ;
        RECT 1724.590 216.000 1724.870 220.000 ;
        RECT 1724.700 72.410 1724.840 216.000 ;
        RECT 1724.640 72.090 1724.900 72.410 ;
        RECT 2030.540 48.290 2030.800 48.610 ;
        RECT 2030.600 2.400 2030.740 48.290 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1742.550 182.820 1742.870 182.880 ;
        RECT 2042.470 182.820 2042.790 182.880 ;
        RECT 1742.550 182.680 2042.790 182.820 ;
        RECT 1742.550 182.620 1742.870 182.680 ;
        RECT 2042.470 182.620 2042.790 182.680 ;
        RECT 2042.470 37.980 2042.790 38.040 ;
        RECT 2048.450 37.980 2048.770 38.040 ;
        RECT 2042.470 37.840 2048.770 37.980 ;
        RECT 2042.470 37.780 2042.790 37.840 ;
        RECT 2048.450 37.780 2048.770 37.840 ;
      LAYER via ;
        RECT 1742.580 182.620 1742.840 182.880 ;
        RECT 2042.500 182.620 2042.760 182.880 ;
        RECT 2042.500 37.780 2042.760 38.040 ;
        RECT 2048.480 37.780 2048.740 38.040 ;
      LAYER met2 ;
        RECT 1742.530 216.000 1742.810 220.000 ;
        RECT 1742.640 182.910 1742.780 216.000 ;
        RECT 1742.580 182.590 1742.840 182.910 ;
        RECT 2042.500 182.590 2042.760 182.910 ;
        RECT 2042.560 38.070 2042.700 182.590 ;
        RECT 2042.500 37.750 2042.760 38.070 ;
        RECT 2048.480 37.750 2048.740 38.070 ;
        RECT 2048.540 2.400 2048.680 37.750 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 455.470 200.500 455.790 200.560 ;
        RECT 461.450 200.500 461.770 200.560 ;
        RECT 455.470 200.360 461.770 200.500 ;
        RECT 455.470 200.300 455.790 200.360 ;
        RECT 461.450 200.300 461.770 200.360 ;
        RECT 461.450 19.960 461.770 20.020 ;
        RECT 763.670 19.960 763.990 20.020 ;
        RECT 461.450 19.820 763.990 19.960 ;
        RECT 461.450 19.760 461.770 19.820 ;
        RECT 763.670 19.760 763.990 19.820 ;
      LAYER via ;
        RECT 455.500 200.300 455.760 200.560 ;
        RECT 461.480 200.300 461.740 200.560 ;
        RECT 461.480 19.760 461.740 20.020 ;
        RECT 763.700 19.760 763.960 20.020 ;
      LAYER met2 ;
        RECT 455.450 216.000 455.730 220.000 ;
        RECT 455.560 200.590 455.700 216.000 ;
        RECT 455.500 200.270 455.760 200.590 ;
        RECT 461.480 200.270 461.740 200.590 ;
        RECT 461.540 20.050 461.680 200.270 ;
        RECT 461.480 19.730 461.740 20.050 ;
        RECT 763.700 19.730 763.960 20.050 ;
        RECT 763.760 2.400 763.900 19.730 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1760.490 200.500 1760.810 200.560 ;
        RECT 1766.010 200.500 1766.330 200.560 ;
        RECT 1760.490 200.360 1766.330 200.500 ;
        RECT 1760.490 200.300 1760.810 200.360 ;
        RECT 1766.010 200.300 1766.330 200.360 ;
        RECT 1766.010 134.880 1766.330 134.940 ;
        RECT 2063.170 134.880 2063.490 134.940 ;
        RECT 1766.010 134.740 2063.490 134.880 ;
        RECT 1766.010 134.680 1766.330 134.740 ;
        RECT 2063.170 134.680 2063.490 134.740 ;
        RECT 2063.170 14.180 2063.490 14.240 ;
        RECT 2063.170 14.040 2066.620 14.180 ;
        RECT 2063.170 13.980 2063.490 14.040 ;
        RECT 2066.480 13.900 2066.620 14.040 ;
        RECT 2066.390 13.640 2066.710 13.900 ;
      LAYER via ;
        RECT 1760.520 200.300 1760.780 200.560 ;
        RECT 1766.040 200.300 1766.300 200.560 ;
        RECT 1766.040 134.680 1766.300 134.940 ;
        RECT 2063.200 134.680 2063.460 134.940 ;
        RECT 2063.200 13.980 2063.460 14.240 ;
        RECT 2066.420 13.640 2066.680 13.900 ;
      LAYER met2 ;
        RECT 1760.470 216.000 1760.750 220.000 ;
        RECT 1760.580 200.590 1760.720 216.000 ;
        RECT 1760.520 200.270 1760.780 200.590 ;
        RECT 1766.040 200.270 1766.300 200.590 ;
        RECT 1766.100 134.970 1766.240 200.270 ;
        RECT 1766.040 134.650 1766.300 134.970 ;
        RECT 2063.200 134.650 2063.460 134.970 ;
        RECT 2063.260 14.270 2063.400 134.650 ;
        RECT 2063.200 13.950 2063.460 14.270 ;
        RECT 2066.420 13.610 2066.680 13.930 ;
        RECT 2066.480 2.400 2066.620 13.610 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.810 51.580 1780.130 51.640 ;
        RECT 2084.330 51.580 2084.650 51.640 ;
        RECT 1779.810 51.440 2084.650 51.580 ;
        RECT 1779.810 51.380 1780.130 51.440 ;
        RECT 2084.330 51.380 2084.650 51.440 ;
      LAYER via ;
        RECT 1779.840 51.380 1780.100 51.640 ;
        RECT 2084.360 51.380 2084.620 51.640 ;
      LAYER met2 ;
        RECT 1778.410 216.650 1778.690 220.000 ;
        RECT 1778.410 216.510 1780.040 216.650 ;
        RECT 1778.410 216.000 1778.690 216.510 ;
        RECT 1779.900 51.670 1780.040 216.510 ;
        RECT 1779.840 51.350 1780.100 51.670 ;
        RECT 2084.360 51.350 2084.620 51.670 ;
        RECT 2084.420 2.400 2084.560 51.350 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1796.370 189.960 1796.690 190.020 ;
        RECT 2097.670 189.960 2097.990 190.020 ;
        RECT 1796.370 189.820 2097.990 189.960 ;
        RECT 1796.370 189.760 1796.690 189.820 ;
        RECT 2097.670 189.760 2097.990 189.820 ;
        RECT 2097.670 14.180 2097.990 14.240 ;
        RECT 2097.670 14.040 2102.040 14.180 ;
        RECT 2097.670 13.980 2097.990 14.040 ;
        RECT 2101.900 13.900 2102.040 14.040 ;
        RECT 2101.810 13.640 2102.130 13.900 ;
      LAYER via ;
        RECT 1796.400 189.760 1796.660 190.020 ;
        RECT 2097.700 189.760 2097.960 190.020 ;
        RECT 2097.700 13.980 2097.960 14.240 ;
        RECT 2101.840 13.640 2102.100 13.900 ;
      LAYER met2 ;
        RECT 1796.350 216.000 1796.630 220.000 ;
        RECT 1796.460 190.050 1796.600 216.000 ;
        RECT 1796.400 189.730 1796.660 190.050 ;
        RECT 2097.700 189.730 2097.960 190.050 ;
        RECT 2097.760 14.270 2097.900 189.730 ;
        RECT 2097.700 13.950 2097.960 14.270 ;
        RECT 2101.840 13.610 2102.100 13.930 ;
        RECT 2101.900 2.400 2102.040 13.610 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1813.850 127.740 1814.170 127.800 ;
        RECT 2118.370 127.740 2118.690 127.800 ;
        RECT 1813.850 127.600 2118.690 127.740 ;
        RECT 1813.850 127.540 1814.170 127.600 ;
        RECT 2118.370 127.540 2118.690 127.600 ;
      LAYER via ;
        RECT 1813.880 127.540 1814.140 127.800 ;
        RECT 2118.400 127.540 2118.660 127.800 ;
      LAYER met2 ;
        RECT 1814.290 216.650 1814.570 220.000 ;
        RECT 1813.940 216.510 1814.570 216.650 ;
        RECT 1813.940 127.830 1814.080 216.510 ;
        RECT 1814.290 216.000 1814.570 216.510 ;
        RECT 1813.880 127.510 1814.140 127.830 ;
        RECT 2118.400 127.510 2118.660 127.830 ;
        RECT 2118.460 24.210 2118.600 127.510 ;
        RECT 2118.460 24.070 2119.520 24.210 ;
        RECT 2119.380 13.330 2119.520 24.070 ;
        RECT 2119.380 13.190 2119.980 13.330 ;
        RECT 2119.840 2.400 2119.980 13.190 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1832.250 196.760 1832.570 196.820 ;
        RECT 2132.170 196.760 2132.490 196.820 ;
        RECT 1832.250 196.620 2132.490 196.760 ;
        RECT 1832.250 196.560 1832.570 196.620 ;
        RECT 2132.170 196.560 2132.490 196.620 ;
        RECT 2132.170 14.180 2132.490 14.240 ;
        RECT 2132.170 14.040 2137.920 14.180 ;
        RECT 2132.170 13.980 2132.490 14.040 ;
        RECT 2137.780 13.900 2137.920 14.040 ;
        RECT 2137.690 13.640 2138.010 13.900 ;
      LAYER via ;
        RECT 1832.280 196.560 1832.540 196.820 ;
        RECT 2132.200 196.560 2132.460 196.820 ;
        RECT 2132.200 13.980 2132.460 14.240 ;
        RECT 2137.720 13.640 2137.980 13.900 ;
      LAYER met2 ;
        RECT 1832.230 216.000 1832.510 220.000 ;
        RECT 1832.340 196.850 1832.480 216.000 ;
        RECT 1832.280 196.530 1832.540 196.850 ;
        RECT 2132.200 196.530 2132.460 196.850 ;
        RECT 2132.260 14.270 2132.400 196.530 ;
        RECT 2132.200 13.950 2132.460 14.270 ;
        RECT 2137.720 13.610 2137.980 13.930 ;
        RECT 2137.780 2.400 2137.920 13.610 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1849.730 200.500 1850.050 200.560 ;
        RECT 1855.250 200.500 1855.570 200.560 ;
        RECT 1849.730 200.360 1855.570 200.500 ;
        RECT 1849.730 200.300 1850.050 200.360 ;
        RECT 1855.250 200.300 1855.570 200.360 ;
        RECT 1855.250 155.280 1855.570 155.340 ;
        RECT 2152.870 155.280 2153.190 155.340 ;
        RECT 1855.250 155.140 2153.190 155.280 ;
        RECT 1855.250 155.080 1855.570 155.140 ;
        RECT 2152.870 155.080 2153.190 155.140 ;
        RECT 2152.410 2.960 2152.730 3.020 ;
        RECT 2155.630 2.960 2155.950 3.020 ;
        RECT 2152.410 2.820 2155.950 2.960 ;
        RECT 2152.410 2.760 2152.730 2.820 ;
        RECT 2155.630 2.760 2155.950 2.820 ;
      LAYER via ;
        RECT 1849.760 200.300 1850.020 200.560 ;
        RECT 1855.280 200.300 1855.540 200.560 ;
        RECT 1855.280 155.080 1855.540 155.340 ;
        RECT 2152.900 155.080 2153.160 155.340 ;
        RECT 2152.440 2.760 2152.700 3.020 ;
        RECT 2155.660 2.760 2155.920 3.020 ;
      LAYER met2 ;
        RECT 1849.710 216.000 1849.990 220.000 ;
        RECT 1849.820 200.590 1849.960 216.000 ;
        RECT 1849.760 200.270 1850.020 200.590 ;
        RECT 1855.280 200.270 1855.540 200.590 ;
        RECT 1855.340 155.370 1855.480 200.270 ;
        RECT 1855.280 155.050 1855.540 155.370 ;
        RECT 2152.900 155.050 2153.160 155.370 ;
        RECT 2152.960 24.380 2153.100 155.050 ;
        RECT 2152.500 24.240 2153.100 24.380 ;
        RECT 2152.500 3.050 2152.640 24.240 ;
        RECT 2152.440 2.730 2152.700 3.050 ;
        RECT 2155.660 2.730 2155.920 3.050 ;
        RECT 2155.720 2.400 2155.860 2.730 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1869.510 162.420 1869.830 162.480 ;
        RECT 2166.670 162.420 2166.990 162.480 ;
        RECT 1869.510 162.280 2166.990 162.420 ;
        RECT 1869.510 162.220 1869.830 162.280 ;
        RECT 2166.670 162.220 2166.990 162.280 ;
        RECT 2166.670 38.320 2166.990 38.380 ;
        RECT 2173.110 38.320 2173.430 38.380 ;
        RECT 2166.670 38.180 2173.430 38.320 ;
        RECT 2166.670 38.120 2166.990 38.180 ;
        RECT 2173.110 38.120 2173.430 38.180 ;
      LAYER via ;
        RECT 1869.540 162.220 1869.800 162.480 ;
        RECT 2166.700 162.220 2166.960 162.480 ;
        RECT 2166.700 38.120 2166.960 38.380 ;
        RECT 2173.140 38.120 2173.400 38.380 ;
      LAYER met2 ;
        RECT 1867.650 216.650 1867.930 220.000 ;
        RECT 1867.650 216.510 1869.740 216.650 ;
        RECT 1867.650 216.000 1867.930 216.510 ;
        RECT 1869.600 162.510 1869.740 216.510 ;
        RECT 1869.540 162.190 1869.800 162.510 ;
        RECT 2166.700 162.190 2166.960 162.510 ;
        RECT 2166.760 38.410 2166.900 162.190 ;
        RECT 2166.700 38.090 2166.960 38.410 ;
        RECT 2173.140 38.090 2173.400 38.410 ;
        RECT 2173.200 2.400 2173.340 38.090 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1885.610 200.500 1885.930 200.560 ;
        RECT 1890.210 200.500 1890.530 200.560 ;
        RECT 1885.610 200.360 1890.530 200.500 ;
        RECT 1885.610 200.300 1885.930 200.360 ;
        RECT 1890.210 200.300 1890.530 200.360 ;
        RECT 1890.210 141.680 1890.530 141.740 ;
        RECT 2187.370 141.680 2187.690 141.740 ;
        RECT 1890.210 141.540 2187.690 141.680 ;
        RECT 1890.210 141.480 1890.530 141.540 ;
        RECT 2187.370 141.480 2187.690 141.540 ;
        RECT 2187.370 14.180 2187.690 14.240 ;
        RECT 2187.370 14.040 2191.280 14.180 ;
        RECT 2187.370 13.980 2187.690 14.040 ;
        RECT 2191.140 13.900 2191.280 14.040 ;
        RECT 2191.050 13.640 2191.370 13.900 ;
      LAYER via ;
        RECT 1885.640 200.300 1885.900 200.560 ;
        RECT 1890.240 200.300 1890.500 200.560 ;
        RECT 1890.240 141.480 1890.500 141.740 ;
        RECT 2187.400 141.480 2187.660 141.740 ;
        RECT 2187.400 13.980 2187.660 14.240 ;
        RECT 2191.080 13.640 2191.340 13.900 ;
      LAYER met2 ;
        RECT 1885.590 216.000 1885.870 220.000 ;
        RECT 1885.700 200.590 1885.840 216.000 ;
        RECT 1885.640 200.270 1885.900 200.590 ;
        RECT 1890.240 200.270 1890.500 200.590 ;
        RECT 1890.300 141.770 1890.440 200.270 ;
        RECT 1890.240 141.450 1890.500 141.770 ;
        RECT 2187.400 141.450 2187.660 141.770 ;
        RECT 2187.460 14.270 2187.600 141.450 ;
        RECT 2187.400 13.950 2187.660 14.270 ;
        RECT 2191.080 13.610 2191.340 13.930 ;
        RECT 2191.140 2.400 2191.280 13.610 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1903.550 58.720 1903.870 58.780 ;
        RECT 2208.990 58.720 2209.310 58.780 ;
        RECT 1903.550 58.580 2209.310 58.720 ;
        RECT 1903.550 58.520 1903.870 58.580 ;
        RECT 2208.990 58.520 2209.310 58.580 ;
      LAYER via ;
        RECT 1903.580 58.520 1903.840 58.780 ;
        RECT 2209.020 58.520 2209.280 58.780 ;
      LAYER met2 ;
        RECT 1903.530 216.000 1903.810 220.000 ;
        RECT 1903.640 58.810 1903.780 216.000 ;
        RECT 1903.580 58.490 1903.840 58.810 ;
        RECT 2209.020 58.490 2209.280 58.810 ;
        RECT 2209.080 2.400 2209.220 58.490 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 169.220 1925.030 169.280 ;
        RECT 2221.870 169.220 2222.190 169.280 ;
        RECT 1924.710 169.080 2222.190 169.220 ;
        RECT 1924.710 169.020 1925.030 169.080 ;
        RECT 2221.870 169.020 2222.190 169.080 ;
        RECT 2221.870 14.180 2222.190 14.240 ;
        RECT 2221.870 14.040 2227.160 14.180 ;
        RECT 2221.870 13.980 2222.190 14.040 ;
        RECT 2227.020 13.900 2227.160 14.040 ;
        RECT 2226.930 13.640 2227.250 13.900 ;
      LAYER via ;
        RECT 1924.740 169.020 1925.000 169.280 ;
        RECT 2221.900 169.020 2222.160 169.280 ;
        RECT 2221.900 13.980 2222.160 14.240 ;
        RECT 2226.960 13.640 2227.220 13.900 ;
      LAYER met2 ;
        RECT 1921.470 216.650 1921.750 220.000 ;
        RECT 1921.470 216.510 1924.940 216.650 ;
        RECT 1921.470 216.000 1921.750 216.510 ;
        RECT 1924.800 169.310 1924.940 216.510 ;
        RECT 1924.740 168.990 1925.000 169.310 ;
        RECT 2221.900 168.990 2222.160 169.310 ;
        RECT 2221.960 14.270 2222.100 168.990 ;
        RECT 2221.900 13.950 2222.160 14.270 ;
        RECT 2226.960 13.610 2227.220 13.930 ;
        RECT 2227.020 2.400 2227.160 13.610 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 475.710 19.280 476.030 19.340 ;
        RECT 781.610 19.280 781.930 19.340 ;
        RECT 475.710 19.140 781.930 19.280 ;
        RECT 475.710 19.080 476.030 19.140 ;
        RECT 781.610 19.080 781.930 19.140 ;
      LAYER via ;
        RECT 475.740 19.080 476.000 19.340 ;
        RECT 781.640 19.080 781.900 19.340 ;
      LAYER met2 ;
        RECT 473.390 216.650 473.670 220.000 ;
        RECT 473.390 216.510 475.940 216.650 ;
        RECT 473.390 216.000 473.670 216.510 ;
        RECT 475.800 19.370 475.940 216.510 ;
        RECT 475.740 19.050 476.000 19.370 ;
        RECT 781.640 19.050 781.900 19.370 ;
        RECT 781.700 2.400 781.840 19.050 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1939.430 200.500 1939.750 200.560 ;
        RECT 1945.410 200.500 1945.730 200.560 ;
        RECT 1939.430 200.360 1945.730 200.500 ;
        RECT 1939.430 200.300 1939.750 200.360 ;
        RECT 1945.410 200.300 1945.730 200.360 ;
        RECT 1945.410 65.520 1945.730 65.580 ;
        RECT 2242.570 65.520 2242.890 65.580 ;
        RECT 1945.410 65.380 2242.890 65.520 ;
        RECT 1945.410 65.320 1945.730 65.380 ;
        RECT 2242.570 65.320 2242.890 65.380 ;
        RECT 2242.570 62.120 2242.890 62.180 ;
        RECT 2244.870 62.120 2245.190 62.180 ;
        RECT 2242.570 61.980 2245.190 62.120 ;
        RECT 2242.570 61.920 2242.890 61.980 ;
        RECT 2244.870 61.920 2245.190 61.980 ;
      LAYER via ;
        RECT 1939.460 200.300 1939.720 200.560 ;
        RECT 1945.440 200.300 1945.700 200.560 ;
        RECT 1945.440 65.320 1945.700 65.580 ;
        RECT 2242.600 65.320 2242.860 65.580 ;
        RECT 2242.600 61.920 2242.860 62.180 ;
        RECT 2244.900 61.920 2245.160 62.180 ;
      LAYER met2 ;
        RECT 1939.410 216.000 1939.690 220.000 ;
        RECT 1939.520 200.590 1939.660 216.000 ;
        RECT 1939.460 200.270 1939.720 200.590 ;
        RECT 1945.440 200.270 1945.700 200.590 ;
        RECT 1945.500 65.610 1945.640 200.270 ;
        RECT 1945.440 65.290 1945.700 65.610 ;
        RECT 2242.600 65.290 2242.860 65.610 ;
        RECT 2242.660 62.210 2242.800 65.290 ;
        RECT 2242.600 61.890 2242.860 62.210 ;
        RECT 2244.900 61.890 2245.160 62.210 ;
        RECT 2244.960 2.400 2245.100 61.890 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1959.210 176.360 1959.530 176.420 ;
        RECT 2256.370 176.360 2256.690 176.420 ;
        RECT 1959.210 176.220 2256.690 176.360 ;
        RECT 1959.210 176.160 1959.530 176.220 ;
        RECT 2256.370 176.160 2256.690 176.220 ;
        RECT 2256.370 38.320 2256.690 38.380 ;
        RECT 2262.350 38.320 2262.670 38.380 ;
        RECT 2256.370 38.180 2262.670 38.320 ;
        RECT 2256.370 38.120 2256.690 38.180 ;
        RECT 2262.350 38.120 2262.670 38.180 ;
      LAYER via ;
        RECT 1959.240 176.160 1959.500 176.420 ;
        RECT 2256.400 176.160 2256.660 176.420 ;
        RECT 2256.400 38.120 2256.660 38.380 ;
        RECT 2262.380 38.120 2262.640 38.380 ;
      LAYER met2 ;
        RECT 1957.350 216.650 1957.630 220.000 ;
        RECT 1957.350 216.510 1959.440 216.650 ;
        RECT 1957.350 216.000 1957.630 216.510 ;
        RECT 1959.300 176.450 1959.440 216.510 ;
        RECT 1959.240 176.130 1959.500 176.450 ;
        RECT 2256.400 176.130 2256.660 176.450 ;
        RECT 2256.460 38.410 2256.600 176.130 ;
        RECT 2256.400 38.090 2256.660 38.410 ;
        RECT 2262.380 38.090 2262.640 38.410 ;
        RECT 2262.440 2.400 2262.580 38.090 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1974.850 200.500 1975.170 200.560 ;
        RECT 1979.910 200.500 1980.230 200.560 ;
        RECT 1974.850 200.360 1980.230 200.500 ;
        RECT 1974.850 200.300 1975.170 200.360 ;
        RECT 1979.910 200.300 1980.230 200.360 ;
        RECT 1979.910 72.660 1980.230 72.720 ;
        RECT 2277.070 72.660 2277.390 72.720 ;
        RECT 1979.910 72.520 2277.390 72.660 ;
        RECT 1979.910 72.460 1980.230 72.520 ;
        RECT 2277.070 72.460 2277.390 72.520 ;
      LAYER via ;
        RECT 1974.880 200.300 1975.140 200.560 ;
        RECT 1979.940 200.300 1980.200 200.560 ;
        RECT 1979.940 72.460 1980.200 72.720 ;
        RECT 2277.100 72.460 2277.360 72.720 ;
      LAYER met2 ;
        RECT 1974.830 216.000 1975.110 220.000 ;
        RECT 1974.940 200.590 1975.080 216.000 ;
        RECT 1974.880 200.270 1975.140 200.590 ;
        RECT 1979.940 200.270 1980.200 200.590 ;
        RECT 1980.000 72.750 1980.140 200.270 ;
        RECT 1979.940 72.430 1980.200 72.750 ;
        RECT 2277.100 72.430 2277.360 72.750 ;
        RECT 2277.160 3.130 2277.300 72.430 ;
        RECT 2277.160 2.990 2280.060 3.130 ;
        RECT 2279.920 2.960 2280.060 2.990 ;
        RECT 2279.920 2.820 2280.520 2.960 ;
        RECT 2280.380 2.400 2280.520 2.820 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1993.710 30.840 1994.030 30.900 ;
        RECT 2298.230 30.840 2298.550 30.900 ;
        RECT 1993.710 30.700 2298.550 30.840 ;
        RECT 1993.710 30.640 1994.030 30.700 ;
        RECT 2298.230 30.640 2298.550 30.700 ;
      LAYER via ;
        RECT 1993.740 30.640 1994.000 30.900 ;
        RECT 2298.260 30.640 2298.520 30.900 ;
      LAYER met2 ;
        RECT 1992.770 216.650 1993.050 220.000 ;
        RECT 1992.770 216.510 1993.940 216.650 ;
        RECT 1992.770 216.000 1993.050 216.510 ;
        RECT 1993.800 30.930 1993.940 216.510 ;
        RECT 1993.740 30.610 1994.000 30.930 ;
        RECT 2298.260 30.610 2298.520 30.930 ;
        RECT 2298.320 2.400 2298.460 30.610 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2010.730 189.620 2011.050 189.680 ;
        RECT 2311.570 189.620 2311.890 189.680 ;
        RECT 2010.730 189.480 2311.890 189.620 ;
        RECT 2010.730 189.420 2011.050 189.480 ;
        RECT 2311.570 189.420 2311.890 189.480 ;
        RECT 2311.570 2.960 2311.890 3.020 ;
        RECT 2316.170 2.960 2316.490 3.020 ;
        RECT 2311.570 2.820 2316.490 2.960 ;
        RECT 2311.570 2.760 2311.890 2.820 ;
        RECT 2316.170 2.760 2316.490 2.820 ;
      LAYER via ;
        RECT 2010.760 189.420 2011.020 189.680 ;
        RECT 2311.600 189.420 2311.860 189.680 ;
        RECT 2311.600 2.760 2311.860 3.020 ;
        RECT 2316.200 2.760 2316.460 3.020 ;
      LAYER met2 ;
        RECT 2010.710 216.000 2010.990 220.000 ;
        RECT 2010.820 189.710 2010.960 216.000 ;
        RECT 2010.760 189.390 2011.020 189.710 ;
        RECT 2311.600 189.390 2311.860 189.710 ;
        RECT 2311.660 3.050 2311.800 189.390 ;
        RECT 2311.600 2.730 2311.860 3.050 ;
        RECT 2316.200 2.730 2316.460 3.050 ;
        RECT 2316.260 2.400 2316.400 2.730 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2028.670 200.500 2028.990 200.560 ;
        RECT 2034.650 200.500 2034.970 200.560 ;
        RECT 2028.670 200.360 2034.970 200.500 ;
        RECT 2028.670 200.300 2028.990 200.360 ;
        RECT 2034.650 200.300 2034.970 200.360 ;
        RECT 2034.650 148.480 2034.970 148.540 ;
        RECT 2332.270 148.480 2332.590 148.540 ;
        RECT 2034.650 148.340 2332.590 148.480 ;
        RECT 2034.650 148.280 2034.970 148.340 ;
        RECT 2332.270 148.280 2332.590 148.340 ;
        RECT 2332.270 2.960 2332.590 3.020 ;
        RECT 2334.110 2.960 2334.430 3.020 ;
        RECT 2332.270 2.820 2334.430 2.960 ;
        RECT 2332.270 2.760 2332.590 2.820 ;
        RECT 2334.110 2.760 2334.430 2.820 ;
      LAYER via ;
        RECT 2028.700 200.300 2028.960 200.560 ;
        RECT 2034.680 200.300 2034.940 200.560 ;
        RECT 2034.680 148.280 2034.940 148.540 ;
        RECT 2332.300 148.280 2332.560 148.540 ;
        RECT 2332.300 2.760 2332.560 3.020 ;
        RECT 2334.140 2.760 2334.400 3.020 ;
      LAYER met2 ;
        RECT 2028.650 216.000 2028.930 220.000 ;
        RECT 2028.760 200.590 2028.900 216.000 ;
        RECT 2028.700 200.270 2028.960 200.590 ;
        RECT 2034.680 200.270 2034.940 200.590 ;
        RECT 2034.740 148.570 2034.880 200.270 ;
        RECT 2034.680 148.250 2034.940 148.570 ;
        RECT 2332.300 148.250 2332.560 148.570 ;
        RECT 2332.360 3.050 2332.500 148.250 ;
        RECT 2332.300 2.730 2332.560 3.050 ;
        RECT 2334.140 2.730 2334.400 3.050 ;
        RECT 2334.200 2.400 2334.340 2.730 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2048.910 134.540 2049.230 134.600 ;
        RECT 2346.070 134.540 2346.390 134.600 ;
        RECT 2048.910 134.400 2346.390 134.540 ;
        RECT 2048.910 134.340 2049.230 134.400 ;
        RECT 2346.070 134.340 2346.390 134.400 ;
        RECT 2346.070 2.960 2346.390 3.020 ;
        RECT 2351.590 2.960 2351.910 3.020 ;
        RECT 2346.070 2.820 2351.910 2.960 ;
        RECT 2346.070 2.760 2346.390 2.820 ;
        RECT 2351.590 2.760 2351.910 2.820 ;
      LAYER via ;
        RECT 2048.940 134.340 2049.200 134.600 ;
        RECT 2346.100 134.340 2346.360 134.600 ;
        RECT 2346.100 2.760 2346.360 3.020 ;
        RECT 2351.620 2.760 2351.880 3.020 ;
      LAYER met2 ;
        RECT 2046.590 216.650 2046.870 220.000 ;
        RECT 2046.590 216.510 2049.140 216.650 ;
        RECT 2046.590 216.000 2046.870 216.510 ;
        RECT 2049.000 134.630 2049.140 216.510 ;
        RECT 2048.940 134.310 2049.200 134.630 ;
        RECT 2346.100 134.310 2346.360 134.630 ;
        RECT 2346.160 3.050 2346.300 134.310 ;
        RECT 2346.100 2.730 2346.360 3.050 ;
        RECT 2351.620 2.730 2351.880 3.050 ;
        RECT 2351.680 2.400 2351.820 2.730 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2064.550 200.500 2064.870 200.560 ;
        RECT 2069.610 200.500 2069.930 200.560 ;
        RECT 2064.550 200.360 2069.930 200.500 ;
        RECT 2064.550 200.300 2064.870 200.360 ;
        RECT 2069.610 200.300 2069.930 200.360 ;
        RECT 2069.610 176.020 2069.930 176.080 ;
        RECT 2366.770 176.020 2367.090 176.080 ;
        RECT 2069.610 175.880 2367.090 176.020 ;
        RECT 2069.610 175.820 2069.930 175.880 ;
        RECT 2366.770 175.820 2367.090 175.880 ;
      LAYER via ;
        RECT 2064.580 200.300 2064.840 200.560 ;
        RECT 2069.640 200.300 2069.900 200.560 ;
        RECT 2069.640 175.820 2069.900 176.080 ;
        RECT 2366.800 175.820 2367.060 176.080 ;
      LAYER met2 ;
        RECT 2064.530 216.000 2064.810 220.000 ;
        RECT 2064.640 200.590 2064.780 216.000 ;
        RECT 2064.580 200.270 2064.840 200.590 ;
        RECT 2069.640 200.270 2069.900 200.590 ;
        RECT 2069.700 176.110 2069.840 200.270 ;
        RECT 2069.640 175.790 2069.900 176.110 ;
        RECT 2366.800 175.790 2367.060 176.110 ;
        RECT 2366.860 3.130 2367.000 175.790 ;
        RECT 2366.860 2.990 2369.300 3.130 ;
        RECT 2369.160 2.960 2369.300 2.990 ;
        RECT 2369.160 2.820 2369.760 2.960 ;
        RECT 2369.620 2.400 2369.760 2.820 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2083.410 51.920 2083.730 51.980 ;
        RECT 2387.930 51.920 2388.250 51.980 ;
        RECT 2083.410 51.780 2388.250 51.920 ;
        RECT 2083.410 51.720 2083.730 51.780 ;
        RECT 2387.930 51.720 2388.250 51.780 ;
      LAYER via ;
        RECT 2083.440 51.720 2083.700 51.980 ;
        RECT 2387.960 51.720 2388.220 51.980 ;
      LAYER met2 ;
        RECT 2082.470 216.650 2082.750 220.000 ;
        RECT 2082.470 216.510 2083.640 216.650 ;
        RECT 2082.470 216.000 2082.750 216.510 ;
        RECT 2083.500 52.010 2083.640 216.510 ;
        RECT 2083.440 51.690 2083.700 52.010 ;
        RECT 2387.960 51.690 2388.220 52.010 ;
        RECT 2388.020 2.960 2388.160 51.690 ;
        RECT 2387.560 2.820 2388.160 2.960 ;
        RECT 2387.560 2.400 2387.700 2.820 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2100.430 200.500 2100.750 200.560 ;
        RECT 2104.110 200.500 2104.430 200.560 ;
        RECT 2100.430 200.360 2104.430 200.500 ;
        RECT 2100.430 200.300 2100.750 200.360 ;
        RECT 2104.110 200.300 2104.430 200.360 ;
        RECT 2104.110 162.080 2104.430 162.140 ;
        RECT 2401.270 162.080 2401.590 162.140 ;
        RECT 2104.110 161.940 2401.590 162.080 ;
        RECT 2104.110 161.880 2104.430 161.940 ;
        RECT 2401.270 161.880 2401.590 161.940 ;
      LAYER via ;
        RECT 2100.460 200.300 2100.720 200.560 ;
        RECT 2104.140 200.300 2104.400 200.560 ;
        RECT 2104.140 161.880 2104.400 162.140 ;
        RECT 2401.300 161.880 2401.560 162.140 ;
      LAYER met2 ;
        RECT 2100.410 216.000 2100.690 220.000 ;
        RECT 2100.520 200.590 2100.660 216.000 ;
        RECT 2100.460 200.270 2100.720 200.590 ;
        RECT 2104.140 200.270 2104.400 200.590 ;
        RECT 2104.200 162.170 2104.340 200.270 ;
        RECT 2104.140 161.850 2104.400 162.170 ;
        RECT 2401.300 161.850 2401.560 162.170 ;
        RECT 2401.360 17.410 2401.500 161.850 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 491.350 200.500 491.670 200.560 ;
        RECT 496.410 200.500 496.730 200.560 ;
        RECT 491.350 200.360 496.730 200.500 ;
        RECT 491.350 200.300 491.670 200.360 ;
        RECT 496.410 200.300 496.730 200.360 ;
        RECT 496.410 15.540 496.730 15.600 ;
        RECT 799.550 15.540 799.870 15.600 ;
        RECT 496.410 15.400 799.870 15.540 ;
        RECT 496.410 15.340 496.730 15.400 ;
        RECT 799.550 15.340 799.870 15.400 ;
      LAYER via ;
        RECT 491.380 200.300 491.640 200.560 ;
        RECT 496.440 200.300 496.700 200.560 ;
        RECT 496.440 15.340 496.700 15.600 ;
        RECT 799.580 15.340 799.840 15.600 ;
      LAYER met2 ;
        RECT 491.330 216.000 491.610 220.000 ;
        RECT 491.440 200.590 491.580 216.000 ;
        RECT 491.380 200.270 491.640 200.590 ;
        RECT 496.440 200.270 496.700 200.590 ;
        RECT 496.500 15.630 496.640 200.270 ;
        RECT 496.440 15.310 496.700 15.630 ;
        RECT 799.580 15.310 799.840 15.630 ;
        RECT 799.640 2.400 799.780 15.310 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 336.330 204.240 336.650 204.300 ;
        RECT 642.230 204.240 642.550 204.300 ;
        RECT 336.330 204.100 642.550 204.240 ;
        RECT 336.330 204.040 336.650 204.100 ;
        RECT 642.230 204.040 642.550 204.100 ;
      LAYER via ;
        RECT 336.360 204.040 336.620 204.300 ;
        RECT 642.260 204.040 642.520 204.300 ;
      LAYER met2 ;
        RECT 336.310 216.000 336.590 220.000 ;
        RECT 336.420 204.330 336.560 216.000 ;
        RECT 336.360 204.010 336.620 204.330 ;
        RECT 642.260 204.010 642.520 204.330 ;
        RECT 642.320 17.410 642.460 204.010 ;
        RECT 642.320 17.270 645.220 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2124.810 79.800 2125.130 79.860 ;
        RECT 2428.870 79.800 2429.190 79.860 ;
        RECT 2124.810 79.660 2429.190 79.800 ;
        RECT 2124.810 79.600 2125.130 79.660 ;
        RECT 2428.870 79.600 2429.190 79.660 ;
      LAYER via ;
        RECT 2124.840 79.600 2125.100 79.860 ;
        RECT 2428.900 79.600 2429.160 79.860 ;
      LAYER met2 ;
        RECT 2123.870 216.650 2124.150 220.000 ;
        RECT 2123.870 216.510 2125.040 216.650 ;
        RECT 2123.870 216.000 2124.150 216.510 ;
        RECT 2124.900 79.890 2125.040 216.510 ;
        RECT 2124.840 79.570 2125.100 79.890 ;
        RECT 2428.900 79.570 2429.160 79.890 ;
        RECT 2428.960 2.400 2429.100 79.570 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2141.830 200.500 2142.150 200.560 ;
        RECT 2145.510 200.500 2145.830 200.560 ;
        RECT 2141.830 200.360 2145.830 200.500 ;
        RECT 2141.830 200.300 2142.150 200.360 ;
        RECT 2145.510 200.300 2145.830 200.360 ;
        RECT 2145.510 17.580 2145.830 17.640 ;
        RECT 2446.810 17.580 2447.130 17.640 ;
        RECT 2145.510 17.440 2447.130 17.580 ;
        RECT 2145.510 17.380 2145.830 17.440 ;
        RECT 2446.810 17.380 2447.130 17.440 ;
      LAYER via ;
        RECT 2141.860 200.300 2142.120 200.560 ;
        RECT 2145.540 200.300 2145.800 200.560 ;
        RECT 2145.540 17.380 2145.800 17.640 ;
        RECT 2446.840 17.380 2447.100 17.640 ;
      LAYER met2 ;
        RECT 2141.810 216.000 2142.090 220.000 ;
        RECT 2141.920 200.590 2142.060 216.000 ;
        RECT 2141.860 200.270 2142.120 200.590 ;
        RECT 2145.540 200.270 2145.800 200.590 ;
        RECT 2145.600 17.670 2145.740 200.270 ;
        RECT 2145.540 17.350 2145.800 17.670 ;
        RECT 2446.840 17.350 2447.100 17.670 ;
        RECT 2446.900 2.400 2447.040 17.350 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2159.770 200.500 2160.090 200.560 ;
        RECT 2165.750 200.500 2166.070 200.560 ;
        RECT 2159.770 200.360 2166.070 200.500 ;
        RECT 2159.770 200.300 2160.090 200.360 ;
        RECT 2165.750 200.300 2166.070 200.360 ;
        RECT 2165.750 16.220 2166.070 16.280 ;
        RECT 2464.750 16.220 2465.070 16.280 ;
        RECT 2165.750 16.080 2465.070 16.220 ;
        RECT 2165.750 16.020 2166.070 16.080 ;
        RECT 2464.750 16.020 2465.070 16.080 ;
      LAYER via ;
        RECT 2159.800 200.300 2160.060 200.560 ;
        RECT 2165.780 200.300 2166.040 200.560 ;
        RECT 2165.780 16.020 2166.040 16.280 ;
        RECT 2464.780 16.020 2465.040 16.280 ;
      LAYER met2 ;
        RECT 2159.750 216.000 2160.030 220.000 ;
        RECT 2159.860 200.590 2160.000 216.000 ;
        RECT 2159.800 200.270 2160.060 200.590 ;
        RECT 2165.780 200.270 2166.040 200.590 ;
        RECT 2165.840 16.310 2165.980 200.270 ;
        RECT 2165.780 15.990 2166.040 16.310 ;
        RECT 2464.780 15.990 2465.040 16.310 ;
        RECT 2464.840 2.400 2464.980 15.990 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 17.240 2180.330 17.300 ;
        RECT 2482.690 17.240 2483.010 17.300 ;
        RECT 2180.010 17.100 2483.010 17.240 ;
        RECT 2180.010 17.040 2180.330 17.100 ;
        RECT 2482.690 17.040 2483.010 17.100 ;
      LAYER via ;
        RECT 2180.040 17.040 2180.300 17.300 ;
        RECT 2482.720 17.040 2482.980 17.300 ;
      LAYER met2 ;
        RECT 2177.690 216.650 2177.970 220.000 ;
        RECT 2177.690 216.510 2180.240 216.650 ;
        RECT 2177.690 216.000 2177.970 216.510 ;
        RECT 2180.100 17.330 2180.240 216.510 ;
        RECT 2180.040 17.010 2180.300 17.330 ;
        RECT 2482.720 17.010 2482.980 17.330 ;
        RECT 2482.780 2.400 2482.920 17.010 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2195.650 200.500 2195.970 200.560 ;
        RECT 2200.710 200.500 2201.030 200.560 ;
        RECT 2195.650 200.360 2201.030 200.500 ;
        RECT 2195.650 200.300 2195.970 200.360 ;
        RECT 2200.710 200.300 2201.030 200.360 ;
        RECT 2200.710 16.900 2201.030 16.960 ;
        RECT 2500.630 16.900 2500.950 16.960 ;
        RECT 2200.710 16.760 2500.950 16.900 ;
        RECT 2200.710 16.700 2201.030 16.760 ;
        RECT 2500.630 16.700 2500.950 16.760 ;
      LAYER via ;
        RECT 2195.680 200.300 2195.940 200.560 ;
        RECT 2200.740 200.300 2201.000 200.560 ;
        RECT 2200.740 16.700 2201.000 16.960 ;
        RECT 2500.660 16.700 2500.920 16.960 ;
      LAYER met2 ;
        RECT 2195.630 216.000 2195.910 220.000 ;
        RECT 2195.740 200.590 2195.880 216.000 ;
        RECT 2195.680 200.270 2195.940 200.590 ;
        RECT 2200.740 200.270 2201.000 200.590 ;
        RECT 2200.800 16.990 2200.940 200.270 ;
        RECT 2200.740 16.670 2201.000 16.990 ;
        RECT 2500.660 16.670 2500.920 16.990 ;
        RECT 2500.720 2.400 2500.860 16.670 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.510 20.640 2214.830 20.700 ;
        RECT 2517.650 20.640 2517.970 20.700 ;
        RECT 2214.510 20.500 2517.970 20.640 ;
        RECT 2214.510 20.440 2214.830 20.500 ;
        RECT 2517.650 20.440 2517.970 20.500 ;
      LAYER via ;
        RECT 2214.540 20.440 2214.800 20.700 ;
        RECT 2517.680 20.440 2517.940 20.700 ;
      LAYER met2 ;
        RECT 2213.570 216.650 2213.850 220.000 ;
        RECT 2213.570 216.510 2214.740 216.650 ;
        RECT 2213.570 216.000 2213.850 216.510 ;
        RECT 2214.600 20.730 2214.740 216.510 ;
        RECT 2214.540 20.410 2214.800 20.730 ;
        RECT 2517.680 20.410 2517.940 20.730 ;
        RECT 2517.740 19.450 2517.880 20.410 ;
        RECT 2517.740 19.310 2518.340 19.450 ;
        RECT 2518.200 2.400 2518.340 19.310 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2231.070 200.500 2231.390 200.560 ;
        RECT 2235.210 200.500 2235.530 200.560 ;
        RECT 2231.070 200.360 2235.530 200.500 ;
        RECT 2231.070 200.300 2231.390 200.360 ;
        RECT 2235.210 200.300 2235.530 200.360 ;
        RECT 2235.210 16.560 2235.530 16.620 ;
        RECT 2536.050 16.560 2536.370 16.620 ;
        RECT 2235.210 16.420 2536.370 16.560 ;
        RECT 2235.210 16.360 2235.530 16.420 ;
        RECT 2536.050 16.360 2536.370 16.420 ;
      LAYER via ;
        RECT 2231.100 200.300 2231.360 200.560 ;
        RECT 2235.240 200.300 2235.500 200.560 ;
        RECT 2235.240 16.360 2235.500 16.620 ;
        RECT 2536.080 16.360 2536.340 16.620 ;
      LAYER met2 ;
        RECT 2231.050 216.000 2231.330 220.000 ;
        RECT 2231.160 200.590 2231.300 216.000 ;
        RECT 2231.100 200.270 2231.360 200.590 ;
        RECT 2235.240 200.270 2235.500 200.590 ;
        RECT 2235.300 16.650 2235.440 200.270 ;
        RECT 2235.240 16.330 2235.500 16.650 ;
        RECT 2536.080 16.330 2536.340 16.650 ;
        RECT 2536.140 2.400 2536.280 16.330 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2248.990 216.000 2249.270 220.000 ;
        RECT 2249.100 17.525 2249.240 216.000 ;
        RECT 2249.030 17.155 2249.310 17.525 ;
        RECT 2554.010 17.155 2554.290 17.525 ;
        RECT 2554.080 2.400 2554.220 17.155 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
      LAYER via2 ;
        RECT 2249.030 17.200 2249.310 17.480 ;
        RECT 2554.010 17.200 2554.290 17.480 ;
      LAYER met3 ;
        RECT 2249.005 17.490 2249.335 17.505 ;
        RECT 2553.985 17.490 2554.315 17.505 ;
        RECT 2249.005 17.190 2554.315 17.490 ;
        RECT 2249.005 17.175 2249.335 17.190 ;
        RECT 2553.985 17.175 2554.315 17.190 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 15.880 2270.030 15.940 ;
        RECT 2571.930 15.880 2572.250 15.940 ;
        RECT 2269.710 15.740 2572.250 15.880 ;
        RECT 2269.710 15.680 2270.030 15.740 ;
        RECT 2571.930 15.680 2572.250 15.740 ;
      LAYER via ;
        RECT 2269.740 15.680 2270.000 15.940 ;
        RECT 2571.960 15.680 2572.220 15.940 ;
      LAYER met2 ;
        RECT 2266.930 216.650 2267.210 220.000 ;
        RECT 2266.930 216.510 2269.940 216.650 ;
        RECT 2266.930 216.000 2267.210 216.510 ;
        RECT 2269.800 15.970 2269.940 216.510 ;
        RECT 2269.740 15.650 2270.000 15.970 ;
        RECT 2571.960 15.650 2572.220 15.970 ;
        RECT 2572.020 2.400 2572.160 15.650 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2284.890 200.500 2285.210 200.560 ;
        RECT 2290.410 200.500 2290.730 200.560 ;
        RECT 2284.890 200.360 2290.730 200.500 ;
        RECT 2284.890 200.300 2285.210 200.360 ;
        RECT 2290.410 200.300 2290.730 200.360 ;
        RECT 2290.410 19.620 2290.730 19.680 ;
        RECT 2589.410 19.620 2589.730 19.680 ;
        RECT 2290.410 19.480 2589.730 19.620 ;
        RECT 2290.410 19.420 2290.730 19.480 ;
        RECT 2589.410 19.420 2589.730 19.480 ;
      LAYER via ;
        RECT 2284.920 200.300 2285.180 200.560 ;
        RECT 2290.440 200.300 2290.700 200.560 ;
        RECT 2290.440 19.420 2290.700 19.680 ;
        RECT 2589.440 19.420 2589.700 19.680 ;
      LAYER met2 ;
        RECT 2284.870 216.000 2285.150 220.000 ;
        RECT 2284.980 200.590 2285.120 216.000 ;
        RECT 2284.920 200.270 2285.180 200.590 ;
        RECT 2290.440 200.270 2290.700 200.590 ;
        RECT 2290.500 19.710 2290.640 200.270 ;
        RECT 2290.440 19.390 2290.700 19.710 ;
        RECT 2589.440 19.390 2589.700 19.710 ;
        RECT 2589.500 2.400 2589.640 19.390 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 531.445 203.745 531.615 204.595 ;
      LAYER mcon ;
        RECT 531.445 204.425 531.615 204.595 ;
      LAYER met1 ;
        RECT 515.270 204.580 515.590 204.640 ;
        RECT 531.385 204.580 531.675 204.625 ;
        RECT 515.270 204.440 531.675 204.580 ;
        RECT 515.270 204.380 515.590 204.440 ;
        RECT 531.385 204.395 531.675 204.440 ;
        RECT 531.385 203.900 531.675 203.945 ;
        RECT 821.630 203.900 821.950 203.960 ;
        RECT 531.385 203.760 821.950 203.900 ;
        RECT 531.385 203.715 531.675 203.760 ;
        RECT 821.630 203.700 821.950 203.760 ;
      LAYER via ;
        RECT 515.300 204.380 515.560 204.640 ;
        RECT 821.660 203.700 821.920 203.960 ;
      LAYER met2 ;
        RECT 515.250 216.000 515.530 220.000 ;
        RECT 515.360 204.670 515.500 216.000 ;
        RECT 515.300 204.350 515.560 204.670 ;
        RECT 821.660 203.670 821.920 203.990 ;
        RECT 821.720 17.410 821.860 203.670 ;
        RECT 821.720 17.270 823.700 17.410 ;
        RECT 823.560 2.400 823.700 17.270 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2346.145 17.765 2346.315 19.975 ;
      LAYER mcon ;
        RECT 2346.145 19.805 2346.315 19.975 ;
      LAYER met1 ;
        RECT 2304.670 19.960 2304.990 20.020 ;
        RECT 2346.085 19.960 2346.375 20.005 ;
        RECT 2304.670 19.820 2346.375 19.960 ;
        RECT 2304.670 19.760 2304.990 19.820 ;
        RECT 2346.085 19.775 2346.375 19.820 ;
        RECT 2346.085 17.920 2346.375 17.965 ;
        RECT 2607.350 17.920 2607.670 17.980 ;
        RECT 2346.085 17.780 2607.670 17.920 ;
        RECT 2346.085 17.735 2346.375 17.780 ;
        RECT 2607.350 17.720 2607.670 17.780 ;
      LAYER via ;
        RECT 2304.700 19.760 2304.960 20.020 ;
        RECT 2607.380 17.720 2607.640 17.980 ;
      LAYER met2 ;
        RECT 2302.810 216.650 2303.090 220.000 ;
        RECT 2302.810 216.510 2304.440 216.650 ;
        RECT 2302.810 216.000 2303.090 216.510 ;
        RECT 2304.300 18.770 2304.440 216.510 ;
        RECT 2304.700 19.730 2304.960 20.050 ;
        RECT 2304.760 18.770 2304.900 19.730 ;
        RECT 2304.300 18.630 2304.900 18.770 ;
        RECT 2607.380 17.690 2607.640 18.010 ;
        RECT 2607.440 2.400 2607.580 17.690 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2320.770 200.500 2321.090 200.560 ;
        RECT 2324.910 200.500 2325.230 200.560 ;
        RECT 2320.770 200.360 2325.230 200.500 ;
        RECT 2320.770 200.300 2321.090 200.360 ;
        RECT 2324.910 200.300 2325.230 200.360 ;
        RECT 2324.910 20.300 2325.230 20.360 ;
        RECT 2324.910 20.160 2346.760 20.300 ;
        RECT 2324.910 20.100 2325.230 20.160 ;
        RECT 2346.620 19.960 2346.760 20.160 ;
        RECT 2625.290 19.960 2625.610 20.020 ;
        RECT 2346.620 19.820 2625.610 19.960 ;
        RECT 2625.290 19.760 2625.610 19.820 ;
      LAYER via ;
        RECT 2320.800 200.300 2321.060 200.560 ;
        RECT 2324.940 200.300 2325.200 200.560 ;
        RECT 2324.940 20.100 2325.200 20.360 ;
        RECT 2625.320 19.760 2625.580 20.020 ;
      LAYER met2 ;
        RECT 2320.750 216.000 2321.030 220.000 ;
        RECT 2320.860 200.590 2321.000 216.000 ;
        RECT 2320.800 200.270 2321.060 200.590 ;
        RECT 2324.940 200.270 2325.200 200.590 ;
        RECT 2325.000 20.390 2325.140 200.270 ;
        RECT 2324.940 20.070 2325.200 20.390 ;
        RECT 2625.320 19.730 2625.580 20.050 ;
        RECT 2625.380 2.400 2625.520 19.730 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2338.710 203.560 2339.030 203.620 ;
        RECT 2642.770 203.560 2643.090 203.620 ;
        RECT 2338.710 203.420 2643.090 203.560 ;
        RECT 2338.710 203.360 2339.030 203.420 ;
        RECT 2642.770 203.360 2643.090 203.420 ;
      LAYER via ;
        RECT 2338.740 203.360 2339.000 203.620 ;
        RECT 2642.800 203.360 2643.060 203.620 ;
      LAYER met2 ;
        RECT 2338.690 216.000 2338.970 220.000 ;
        RECT 2338.800 203.650 2338.940 216.000 ;
        RECT 2338.740 203.330 2339.000 203.650 ;
        RECT 2642.800 203.330 2643.060 203.650 ;
        RECT 2642.860 17.410 2643.000 203.330 ;
        RECT 2642.860 17.270 2643.460 17.410 ;
        RECT 2643.320 2.400 2643.460 17.270 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2642.845 15.385 2643.015 18.275 ;
      LAYER mcon ;
        RECT 2642.845 18.105 2643.015 18.275 ;
      LAYER met1 ;
        RECT 2359.410 18.260 2359.730 18.320 ;
        RECT 2642.785 18.260 2643.075 18.305 ;
        RECT 2359.410 18.120 2643.075 18.260 ;
        RECT 2359.410 18.060 2359.730 18.120 ;
        RECT 2642.785 18.075 2643.075 18.120 ;
        RECT 2642.785 15.540 2643.075 15.585 ;
        RECT 2661.170 15.540 2661.490 15.600 ;
        RECT 2642.785 15.400 2661.490 15.540 ;
        RECT 2642.785 15.355 2643.075 15.400 ;
        RECT 2661.170 15.340 2661.490 15.400 ;
      LAYER via ;
        RECT 2359.440 18.060 2359.700 18.320 ;
        RECT 2661.200 15.340 2661.460 15.600 ;
      LAYER met2 ;
        RECT 2356.630 216.650 2356.910 220.000 ;
        RECT 2356.630 216.510 2359.640 216.650 ;
        RECT 2356.630 216.000 2356.910 216.510 ;
        RECT 2359.500 18.350 2359.640 216.510 ;
        RECT 2359.440 18.030 2359.700 18.350 ;
        RECT 2661.200 15.310 2661.460 15.630 ;
        RECT 2661.260 2.400 2661.400 15.310 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2374.130 204.580 2374.450 204.640 ;
        RECT 2677.270 204.580 2677.590 204.640 ;
        RECT 2374.130 204.440 2677.590 204.580 ;
        RECT 2374.130 204.380 2374.450 204.440 ;
        RECT 2677.270 204.380 2677.590 204.440 ;
      LAYER via ;
        RECT 2374.160 204.380 2374.420 204.640 ;
        RECT 2677.300 204.380 2677.560 204.640 ;
      LAYER met2 ;
        RECT 2374.110 216.000 2374.390 220.000 ;
        RECT 2374.220 204.670 2374.360 216.000 ;
        RECT 2374.160 204.350 2374.420 204.670 ;
        RECT 2677.300 204.350 2677.560 204.670 ;
        RECT 2677.360 17.410 2677.500 204.350 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2393.910 18.600 2394.230 18.660 ;
        RECT 2696.590 18.600 2696.910 18.660 ;
        RECT 2393.910 18.460 2696.910 18.600 ;
        RECT 2393.910 18.400 2394.230 18.460 ;
        RECT 2696.590 18.400 2696.910 18.460 ;
      LAYER via ;
        RECT 2393.940 18.400 2394.200 18.660 ;
        RECT 2696.620 18.400 2696.880 18.660 ;
      LAYER met2 ;
        RECT 2392.050 216.650 2392.330 220.000 ;
        RECT 2392.050 216.510 2394.140 216.650 ;
        RECT 2392.050 216.000 2392.330 216.510 ;
        RECT 2394.000 18.690 2394.140 216.510 ;
        RECT 2393.940 18.370 2394.200 18.690 ;
        RECT 2696.620 18.370 2696.880 18.690 ;
        RECT 2696.680 2.400 2696.820 18.370 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2410.010 204.240 2410.330 204.300 ;
        RECT 2711.770 204.240 2712.090 204.300 ;
        RECT 2410.010 204.100 2712.090 204.240 ;
        RECT 2410.010 204.040 2410.330 204.100 ;
        RECT 2711.770 204.040 2712.090 204.100 ;
      LAYER via ;
        RECT 2410.040 204.040 2410.300 204.300 ;
        RECT 2711.800 204.040 2712.060 204.300 ;
      LAYER met2 ;
        RECT 2409.990 216.000 2410.270 220.000 ;
        RECT 2410.100 204.330 2410.240 216.000 ;
        RECT 2410.040 204.010 2410.300 204.330 ;
        RECT 2711.800 204.010 2712.060 204.330 ;
        RECT 2711.860 17.410 2712.000 204.010 ;
        RECT 2711.860 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2427.930 216.650 2428.210 220.000 ;
        RECT 2427.930 216.510 2428.640 216.650 ;
        RECT 2427.930 216.000 2428.210 216.510 ;
        RECT 2428.500 18.205 2428.640 216.510 ;
        RECT 2428.430 17.835 2428.710 18.205 ;
        RECT 2732.490 17.835 2732.770 18.205 ;
        RECT 2732.560 2.400 2732.700 17.835 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 2428.430 17.880 2428.710 18.160 ;
        RECT 2732.490 17.880 2732.770 18.160 ;
      LAYER met3 ;
        RECT 2428.405 18.170 2428.735 18.185 ;
        RECT 2732.465 18.170 2732.795 18.185 ;
        RECT 2428.405 17.870 2732.795 18.170 ;
        RECT 2428.405 17.855 2428.735 17.870 ;
        RECT 2732.465 17.855 2732.795 17.870 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2445.890 203.900 2446.210 203.960 ;
        RECT 2746.270 203.900 2746.590 203.960 ;
        RECT 2445.890 203.760 2746.590 203.900 ;
        RECT 2445.890 203.700 2446.210 203.760 ;
        RECT 2746.270 203.700 2746.590 203.760 ;
      LAYER via ;
        RECT 2445.920 203.700 2446.180 203.960 ;
        RECT 2746.300 203.700 2746.560 203.960 ;
      LAYER met2 ;
        RECT 2445.870 216.000 2446.150 220.000 ;
        RECT 2445.980 203.990 2446.120 216.000 ;
        RECT 2445.920 203.670 2446.180 203.990 ;
        RECT 2746.300 203.670 2746.560 203.990 ;
        RECT 2746.360 17.410 2746.500 203.670 ;
        RECT 2746.360 17.270 2750.640 17.410 ;
        RECT 2750.500 2.400 2750.640 17.270 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2463.830 200.500 2464.150 200.560 ;
        RECT 2469.810 200.500 2470.130 200.560 ;
        RECT 2463.830 200.360 2470.130 200.500 ;
        RECT 2463.830 200.300 2464.150 200.360 ;
        RECT 2469.810 200.300 2470.130 200.360 ;
        RECT 2469.810 17.580 2470.130 17.640 ;
        RECT 2767.890 17.580 2768.210 17.640 ;
        RECT 2469.810 17.440 2768.210 17.580 ;
        RECT 2469.810 17.380 2470.130 17.440 ;
        RECT 2767.890 17.380 2768.210 17.440 ;
      LAYER via ;
        RECT 2463.860 200.300 2464.120 200.560 ;
        RECT 2469.840 200.300 2470.100 200.560 ;
        RECT 2469.840 17.380 2470.100 17.640 ;
        RECT 2767.920 17.380 2768.180 17.640 ;
      LAYER met2 ;
        RECT 2463.810 216.000 2464.090 220.000 ;
        RECT 2463.920 200.590 2464.060 216.000 ;
        RECT 2463.860 200.270 2464.120 200.590 ;
        RECT 2469.840 200.270 2470.100 200.590 ;
        RECT 2469.900 17.670 2470.040 200.270 ;
        RECT 2469.840 17.350 2470.100 17.670 ;
        RECT 2767.920 17.350 2768.180 17.670 ;
        RECT 2767.980 2.400 2768.120 17.350 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 533.210 200.500 533.530 200.560 ;
        RECT 537.810 200.500 538.130 200.560 ;
        RECT 533.210 200.360 538.130 200.500 ;
        RECT 533.210 200.300 533.530 200.360 ;
        RECT 537.810 200.300 538.130 200.360 ;
        RECT 537.810 16.220 538.130 16.280 ;
        RECT 840.950 16.220 841.270 16.280 ;
        RECT 537.810 16.080 841.270 16.220 ;
        RECT 537.810 16.020 538.130 16.080 ;
        RECT 840.950 16.020 841.270 16.080 ;
      LAYER via ;
        RECT 533.240 200.300 533.500 200.560 ;
        RECT 537.840 200.300 538.100 200.560 ;
        RECT 537.840 16.020 538.100 16.280 ;
        RECT 840.980 16.020 841.240 16.280 ;
      LAYER met2 ;
        RECT 533.190 216.000 533.470 220.000 ;
        RECT 533.300 200.590 533.440 216.000 ;
        RECT 533.240 200.270 533.500 200.590 ;
        RECT 537.840 200.270 538.100 200.590 ;
        RECT 537.900 16.310 538.040 200.270 ;
        RECT 537.840 15.990 538.100 16.310 ;
        RECT 840.980 15.990 841.240 16.310 ;
        RECT 841.040 2.400 841.180 15.990 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2483.610 18.940 2483.930 19.000 ;
        RECT 2785.830 18.940 2786.150 19.000 ;
        RECT 2483.610 18.800 2786.150 18.940 ;
        RECT 2483.610 18.740 2483.930 18.800 ;
        RECT 2785.830 18.740 2786.150 18.800 ;
      LAYER via ;
        RECT 2483.640 18.740 2483.900 19.000 ;
        RECT 2785.860 18.740 2786.120 19.000 ;
      LAYER met2 ;
        RECT 2481.750 216.650 2482.030 220.000 ;
        RECT 2481.750 216.510 2483.840 216.650 ;
        RECT 2481.750 216.000 2482.030 216.510 ;
        RECT 2483.700 19.030 2483.840 216.510 ;
        RECT 2483.640 18.710 2483.900 19.030 ;
        RECT 2785.860 18.710 2786.120 19.030 ;
        RECT 2785.920 2.400 2786.060 18.710 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2499.250 200.500 2499.570 200.560 ;
        RECT 2504.310 200.500 2504.630 200.560 ;
        RECT 2499.250 200.360 2504.630 200.500 ;
        RECT 2499.250 200.300 2499.570 200.360 ;
        RECT 2504.310 200.300 2504.630 200.360 ;
        RECT 2504.310 16.900 2504.630 16.960 ;
        RECT 2803.770 16.900 2804.090 16.960 ;
        RECT 2504.310 16.760 2804.090 16.900 ;
        RECT 2504.310 16.700 2504.630 16.760 ;
        RECT 2803.770 16.700 2804.090 16.760 ;
      LAYER via ;
        RECT 2499.280 200.300 2499.540 200.560 ;
        RECT 2504.340 200.300 2504.600 200.560 ;
        RECT 2504.340 16.700 2504.600 16.960 ;
        RECT 2803.800 16.700 2804.060 16.960 ;
      LAYER met2 ;
        RECT 2499.230 216.000 2499.510 220.000 ;
        RECT 2499.340 200.590 2499.480 216.000 ;
        RECT 2499.280 200.270 2499.540 200.590 ;
        RECT 2504.340 200.270 2504.600 200.590 ;
        RECT 2504.400 16.990 2504.540 200.270 ;
        RECT 2504.340 16.670 2504.600 16.990 ;
        RECT 2803.800 16.670 2804.060 16.990 ;
        RECT 2803.860 2.400 2804.000 16.670 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2518.110 20.300 2518.430 20.360 ;
        RECT 2821.710 20.300 2822.030 20.360 ;
        RECT 2518.110 20.160 2822.030 20.300 ;
        RECT 2518.110 20.100 2518.430 20.160 ;
        RECT 2821.710 20.100 2822.030 20.160 ;
      LAYER via ;
        RECT 2518.140 20.100 2518.400 20.360 ;
        RECT 2821.740 20.100 2822.000 20.360 ;
      LAYER met2 ;
        RECT 2517.170 216.650 2517.450 220.000 ;
        RECT 2517.170 216.510 2518.340 216.650 ;
        RECT 2517.170 216.000 2517.450 216.510 ;
        RECT 2518.200 20.390 2518.340 216.510 ;
        RECT 2518.140 20.070 2518.400 20.390 ;
        RECT 2821.740 20.070 2822.000 20.390 ;
        RECT 2821.800 2.400 2821.940 20.070 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2538.810 20.640 2539.130 20.700 ;
        RECT 2839.190 20.640 2839.510 20.700 ;
        RECT 2538.810 20.500 2839.510 20.640 ;
        RECT 2538.810 20.440 2539.130 20.500 ;
        RECT 2839.190 20.440 2839.510 20.500 ;
      LAYER via ;
        RECT 2538.840 20.440 2539.100 20.700 ;
        RECT 2839.220 20.440 2839.480 20.700 ;
      LAYER met2 ;
        RECT 2535.110 216.650 2535.390 220.000 ;
        RECT 2535.110 216.510 2539.040 216.650 ;
        RECT 2535.110 216.000 2535.390 216.510 ;
        RECT 2538.900 20.730 2539.040 216.510 ;
        RECT 2538.840 20.410 2539.100 20.730 ;
        RECT 2839.220 20.410 2839.480 20.730 ;
        RECT 2839.280 2.400 2839.420 20.410 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2553.070 200.500 2553.390 200.560 ;
        RECT 2559.510 200.500 2559.830 200.560 ;
        RECT 2553.070 200.360 2559.830 200.500 ;
        RECT 2553.070 200.300 2553.390 200.360 ;
        RECT 2559.510 200.300 2559.830 200.360 ;
        RECT 2559.510 16.220 2559.830 16.280 ;
        RECT 2857.130 16.220 2857.450 16.280 ;
        RECT 2559.510 16.080 2857.450 16.220 ;
        RECT 2559.510 16.020 2559.830 16.080 ;
        RECT 2857.130 16.020 2857.450 16.080 ;
      LAYER via ;
        RECT 2553.100 200.300 2553.360 200.560 ;
        RECT 2559.540 200.300 2559.800 200.560 ;
        RECT 2559.540 16.020 2559.800 16.280 ;
        RECT 2857.160 16.020 2857.420 16.280 ;
      LAYER met2 ;
        RECT 2553.050 216.000 2553.330 220.000 ;
        RECT 2553.160 200.590 2553.300 216.000 ;
        RECT 2553.100 200.270 2553.360 200.590 ;
        RECT 2559.540 200.270 2559.800 200.590 ;
        RECT 2559.600 16.310 2559.740 200.270 ;
        RECT 2559.540 15.990 2559.800 16.310 ;
        RECT 2857.160 15.990 2857.420 16.310 ;
        RECT 2857.220 2.400 2857.360 15.990 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 15.880 2573.630 15.940 ;
        RECT 2875.070 15.880 2875.390 15.940 ;
        RECT 2573.310 15.740 2875.390 15.880 ;
        RECT 2573.310 15.680 2573.630 15.740 ;
        RECT 2875.070 15.680 2875.390 15.740 ;
      LAYER via ;
        RECT 2573.340 15.680 2573.600 15.940 ;
        RECT 2875.100 15.680 2875.360 15.940 ;
      LAYER met2 ;
        RECT 2570.990 216.650 2571.270 220.000 ;
        RECT 2570.990 216.510 2573.540 216.650 ;
        RECT 2570.990 216.000 2571.270 216.510 ;
        RECT 2573.400 15.970 2573.540 216.510 ;
        RECT 2573.340 15.650 2573.600 15.970 ;
        RECT 2875.100 15.650 2875.360 15.970 ;
        RECT 2875.160 2.400 2875.300 15.650 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2588.950 200.500 2589.270 200.560 ;
        RECT 2594.010 200.500 2594.330 200.560 ;
        RECT 2588.950 200.360 2594.330 200.500 ;
        RECT 2588.950 200.300 2589.270 200.360 ;
        RECT 2594.010 200.300 2594.330 200.360 ;
        RECT 2594.010 17.240 2594.330 17.300 ;
        RECT 2893.010 17.240 2893.330 17.300 ;
        RECT 2594.010 17.100 2893.330 17.240 ;
        RECT 2594.010 17.040 2594.330 17.100 ;
        RECT 2893.010 17.040 2893.330 17.100 ;
      LAYER via ;
        RECT 2588.980 200.300 2589.240 200.560 ;
        RECT 2594.040 200.300 2594.300 200.560 ;
        RECT 2594.040 17.040 2594.300 17.300 ;
        RECT 2893.040 17.040 2893.300 17.300 ;
      LAYER met2 ;
        RECT 2588.930 216.000 2589.210 220.000 ;
        RECT 2589.040 200.590 2589.180 216.000 ;
        RECT 2588.980 200.270 2589.240 200.590 ;
        RECT 2594.040 200.270 2594.300 200.590 ;
        RECT 2594.100 17.330 2594.240 200.270 ;
        RECT 2594.040 17.010 2594.300 17.330 ;
        RECT 2893.040 17.010 2893.300 17.330 ;
        RECT 2893.100 2.400 2893.240 17.010 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2607.810 17.920 2608.130 17.980 ;
        RECT 2910.950 17.920 2911.270 17.980 ;
        RECT 2607.810 17.780 2911.270 17.920 ;
        RECT 2607.810 17.720 2608.130 17.780 ;
        RECT 2910.950 17.720 2911.270 17.780 ;
      LAYER via ;
        RECT 2607.840 17.720 2608.100 17.980 ;
        RECT 2910.980 17.720 2911.240 17.980 ;
      LAYER met2 ;
        RECT 2606.870 216.650 2607.150 220.000 ;
        RECT 2606.870 216.510 2608.040 216.650 ;
        RECT 2606.870 216.000 2607.150 216.510 ;
        RECT 2607.900 18.010 2608.040 216.510 ;
        RECT 2607.840 17.690 2608.100 18.010 ;
        RECT 2910.980 17.690 2911.240 18.010 ;
        RECT 2911.040 2.400 2911.180 17.690 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.150 205.600 551.470 205.660 ;
        RECT 856.130 205.600 856.450 205.660 ;
        RECT 551.150 205.460 856.450 205.600 ;
        RECT 551.150 205.400 551.470 205.460 ;
        RECT 856.130 205.400 856.450 205.460 ;
      LAYER via ;
        RECT 551.180 205.400 551.440 205.660 ;
        RECT 856.160 205.400 856.420 205.660 ;
      LAYER met2 ;
        RECT 551.130 216.000 551.410 220.000 ;
        RECT 551.240 205.690 551.380 216.000 ;
        RECT 551.180 205.370 551.440 205.690 ;
        RECT 856.160 205.370 856.420 205.690 ;
        RECT 856.220 16.730 856.360 205.370 ;
        RECT 856.220 16.590 859.120 16.730 ;
        RECT 858.980 2.400 859.120 16.590 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 568.630 204.580 568.950 204.640 ;
        RECT 572.310 204.580 572.630 204.640 ;
        RECT 568.630 204.440 572.630 204.580 ;
        RECT 568.630 204.380 568.950 204.440 ;
        RECT 572.310 204.380 572.630 204.440 ;
        RECT 572.310 18.940 572.630 19.000 ;
        RECT 876.370 18.940 876.690 19.000 ;
        RECT 572.310 18.800 876.690 18.940 ;
        RECT 572.310 18.740 572.630 18.800 ;
        RECT 876.370 18.740 876.690 18.800 ;
      LAYER via ;
        RECT 568.660 204.380 568.920 204.640 ;
        RECT 572.340 204.380 572.600 204.640 ;
        RECT 572.340 18.740 572.600 19.000 ;
        RECT 876.400 18.740 876.660 19.000 ;
      LAYER met2 ;
        RECT 568.610 216.000 568.890 220.000 ;
        RECT 568.720 204.670 568.860 216.000 ;
        RECT 568.660 204.350 568.920 204.670 ;
        RECT 572.340 204.350 572.600 204.670 ;
        RECT 572.400 19.030 572.540 204.350 ;
        RECT 572.340 18.710 572.600 19.030 ;
        RECT 876.400 18.710 876.660 19.030 ;
        RECT 876.460 16.050 876.600 18.710 ;
        RECT 876.460 15.910 877.060 16.050 ;
        RECT 876.920 2.400 877.060 15.910 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.570 202.540 586.890 202.600 ;
        RECT 593.010 202.540 593.330 202.600 ;
        RECT 586.570 202.400 593.330 202.540 ;
        RECT 586.570 202.340 586.890 202.400 ;
        RECT 593.010 202.340 593.330 202.400 ;
        RECT 593.010 16.560 593.330 16.620 ;
        RECT 593.010 16.420 865.100 16.560 ;
        RECT 593.010 16.360 593.330 16.420 ;
        RECT 864.960 16.220 865.100 16.420 ;
        RECT 894.770 16.220 895.090 16.280 ;
        RECT 864.960 16.080 895.090 16.220 ;
        RECT 894.770 16.020 895.090 16.080 ;
      LAYER via ;
        RECT 586.600 202.340 586.860 202.600 ;
        RECT 593.040 202.340 593.300 202.600 ;
        RECT 593.040 16.360 593.300 16.620 ;
        RECT 894.800 16.020 895.060 16.280 ;
      LAYER met2 ;
        RECT 586.550 216.000 586.830 220.000 ;
        RECT 586.660 202.630 586.800 216.000 ;
        RECT 586.600 202.310 586.860 202.630 ;
        RECT 593.040 202.310 593.300 202.630 ;
        RECT 593.100 16.650 593.240 202.310 ;
        RECT 593.040 16.330 593.300 16.650 ;
        RECT 894.800 15.990 895.060 16.310 ;
        RECT 894.860 2.400 895.000 15.990 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 18.600 607.130 18.660 ;
        RECT 912.710 18.600 913.030 18.660 ;
        RECT 606.810 18.460 913.030 18.600 ;
        RECT 606.810 18.400 607.130 18.460 ;
        RECT 912.710 18.400 913.030 18.460 ;
      LAYER via ;
        RECT 606.840 18.400 607.100 18.660 ;
        RECT 912.740 18.400 913.000 18.660 ;
      LAYER met2 ;
        RECT 604.490 216.650 604.770 220.000 ;
        RECT 604.490 216.510 607.040 216.650 ;
        RECT 604.490 216.000 604.770 216.510 ;
        RECT 606.900 18.690 607.040 216.510 ;
        RECT 606.840 18.370 607.100 18.690 ;
        RECT 912.740 18.370 913.000 18.690 ;
        RECT 912.800 2.400 912.940 18.370 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 905.425 16.065 905.595 16.915 ;
      LAYER mcon ;
        RECT 905.425 16.745 905.595 16.915 ;
      LAYER met1 ;
        RECT 622.450 200.500 622.770 200.560 ;
        RECT 627.510 200.500 627.830 200.560 ;
        RECT 622.450 200.360 627.830 200.500 ;
        RECT 622.450 200.300 622.770 200.360 ;
        RECT 627.510 200.300 627.830 200.360 ;
        RECT 627.510 16.900 627.830 16.960 ;
        RECT 905.365 16.900 905.655 16.945 ;
        RECT 627.510 16.760 905.655 16.900 ;
        RECT 627.510 16.700 627.830 16.760 ;
        RECT 905.365 16.715 905.655 16.760 ;
        RECT 905.365 16.220 905.655 16.265 ;
        RECT 930.190 16.220 930.510 16.280 ;
        RECT 905.365 16.080 930.510 16.220 ;
        RECT 905.365 16.035 905.655 16.080 ;
        RECT 930.190 16.020 930.510 16.080 ;
      LAYER via ;
        RECT 622.480 200.300 622.740 200.560 ;
        RECT 627.540 200.300 627.800 200.560 ;
        RECT 627.540 16.700 627.800 16.960 ;
        RECT 930.220 16.020 930.480 16.280 ;
      LAYER met2 ;
        RECT 622.430 216.000 622.710 220.000 ;
        RECT 622.540 200.590 622.680 216.000 ;
        RECT 622.480 200.270 622.740 200.590 ;
        RECT 627.540 200.270 627.800 200.590 ;
        RECT 627.600 16.990 627.740 200.270 ;
        RECT 627.540 16.670 627.800 16.990 ;
        RECT 930.220 15.990 930.480 16.310 ;
        RECT 930.280 2.400 930.420 15.990 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 641.310 18.260 641.630 18.320 ;
        RECT 948.130 18.260 948.450 18.320 ;
        RECT 641.310 18.120 948.450 18.260 ;
        RECT 641.310 18.060 641.630 18.120 ;
        RECT 948.130 18.060 948.450 18.120 ;
      LAYER via ;
        RECT 641.340 18.060 641.600 18.320 ;
        RECT 948.160 18.060 948.420 18.320 ;
      LAYER met2 ;
        RECT 640.370 216.650 640.650 220.000 ;
        RECT 640.370 216.510 641.540 216.650 ;
        RECT 640.370 216.000 640.650 216.510 ;
        RECT 641.400 18.350 641.540 216.510 ;
        RECT 641.340 18.030 641.600 18.350 ;
        RECT 948.160 18.030 948.420 18.350 ;
        RECT 948.220 2.400 948.360 18.030 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 658.330 205.260 658.650 205.320 ;
        RECT 966.990 205.260 967.310 205.320 ;
        RECT 658.330 205.120 967.310 205.260 ;
        RECT 658.330 205.060 658.650 205.120 ;
        RECT 966.990 205.060 967.310 205.120 ;
      LAYER via ;
        RECT 658.360 205.060 658.620 205.320 ;
        RECT 967.020 205.060 967.280 205.320 ;
      LAYER met2 ;
        RECT 658.310 216.000 658.590 220.000 ;
        RECT 658.420 205.350 658.560 216.000 ;
        RECT 658.360 205.030 658.620 205.350 ;
        RECT 967.020 205.030 967.280 205.350 ;
        RECT 967.080 16.730 967.220 205.030 ;
        RECT 966.160 16.590 967.220 16.730 ;
        RECT 966.160 2.400 966.300 16.590 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 676.270 200.500 676.590 200.560 ;
        RECT 682.710 200.500 683.030 200.560 ;
        RECT 676.270 200.360 683.030 200.500 ;
        RECT 676.270 200.300 676.590 200.360 ;
        RECT 682.710 200.300 683.030 200.360 ;
        RECT 682.710 20.640 683.030 20.700 ;
        RECT 984.010 20.640 984.330 20.700 ;
        RECT 682.710 20.500 984.330 20.640 ;
        RECT 682.710 20.440 683.030 20.500 ;
        RECT 984.010 20.440 984.330 20.500 ;
      LAYER via ;
        RECT 676.300 200.300 676.560 200.560 ;
        RECT 682.740 200.300 683.000 200.560 ;
        RECT 682.740 20.440 683.000 20.700 ;
        RECT 984.040 20.440 984.300 20.700 ;
      LAYER met2 ;
        RECT 676.250 216.000 676.530 220.000 ;
        RECT 676.360 200.590 676.500 216.000 ;
        RECT 676.300 200.270 676.560 200.590 ;
        RECT 682.740 200.270 683.000 200.590 ;
        RECT 682.800 20.730 682.940 200.270 ;
        RECT 682.740 20.410 683.000 20.730 ;
        RECT 984.040 20.410 984.300 20.730 ;
        RECT 984.100 2.400 984.240 20.410 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 354.270 200.500 354.590 200.560 ;
        RECT 358.410 200.500 358.730 200.560 ;
        RECT 354.270 200.360 358.730 200.500 ;
        RECT 354.270 200.300 354.590 200.360 ;
        RECT 358.410 200.300 358.730 200.360 ;
        RECT 358.410 17.920 358.730 17.980 ;
        RECT 662.470 17.920 662.790 17.980 ;
        RECT 358.410 17.780 662.790 17.920 ;
        RECT 358.410 17.720 358.730 17.780 ;
        RECT 662.470 17.720 662.790 17.780 ;
      LAYER via ;
        RECT 354.300 200.300 354.560 200.560 ;
        RECT 358.440 200.300 358.700 200.560 ;
        RECT 358.440 17.720 358.700 17.980 ;
        RECT 662.500 17.720 662.760 17.980 ;
      LAYER met2 ;
        RECT 354.250 216.000 354.530 220.000 ;
        RECT 354.360 200.590 354.500 216.000 ;
        RECT 354.300 200.270 354.560 200.590 ;
        RECT 358.440 200.270 358.700 200.590 ;
        RECT 358.500 18.010 358.640 200.270 ;
        RECT 358.440 17.690 358.700 18.010 ;
        RECT 662.500 17.690 662.760 18.010 ;
        RECT 662.560 16.730 662.700 17.690 ;
        RECT 662.560 16.590 663.160 16.730 ;
        RECT 663.020 2.400 663.160 16.590 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 753.625 203.065 753.795 204.935 ;
        RECT 952.345 203.745 952.515 204.935 ;
        RECT 976.265 203.745 976.435 205.275 ;
      LAYER mcon ;
        RECT 976.265 205.105 976.435 205.275 ;
        RECT 753.625 204.765 753.795 204.935 ;
        RECT 952.345 204.765 952.515 204.935 ;
      LAYER met1 ;
        RECT 976.205 205.260 976.495 205.305 ;
        RECT 1001.030 205.260 1001.350 205.320 ;
        RECT 976.205 205.120 1001.350 205.260 ;
        RECT 976.205 205.075 976.495 205.120 ;
        RECT 1001.030 205.060 1001.350 205.120 ;
        RECT 753.565 204.920 753.855 204.965 ;
        RECT 952.285 204.920 952.575 204.965 ;
        RECT 753.565 204.780 952.575 204.920 ;
        RECT 753.565 204.735 753.855 204.780 ;
        RECT 952.285 204.735 952.575 204.780 ;
        RECT 952.285 203.900 952.575 203.945 ;
        RECT 976.205 203.900 976.495 203.945 ;
        RECT 952.285 203.760 976.495 203.900 ;
        RECT 952.285 203.715 952.575 203.760 ;
        RECT 976.205 203.715 976.495 203.760 ;
        RECT 694.210 203.220 694.530 203.280 ;
        RECT 753.565 203.220 753.855 203.265 ;
        RECT 694.210 203.080 753.855 203.220 ;
        RECT 694.210 203.020 694.530 203.080 ;
        RECT 753.565 203.035 753.855 203.080 ;
      LAYER via ;
        RECT 1001.060 205.060 1001.320 205.320 ;
        RECT 694.240 203.020 694.500 203.280 ;
      LAYER met2 ;
        RECT 694.190 216.000 694.470 220.000 ;
        RECT 694.300 203.310 694.440 216.000 ;
        RECT 1001.060 205.030 1001.320 205.350 ;
        RECT 694.240 202.990 694.500 203.310 ;
        RECT 1001.120 16.730 1001.260 205.030 ;
        RECT 1001.120 16.590 1002.180 16.730 ;
        RECT 1002.040 2.400 1002.180 16.590 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 711.690 202.880 712.010 202.940 ;
        RECT 717.210 202.880 717.530 202.940 ;
        RECT 711.690 202.740 717.530 202.880 ;
        RECT 711.690 202.680 712.010 202.740 ;
        RECT 717.210 202.680 717.530 202.740 ;
        RECT 717.210 20.300 717.530 20.360 ;
        RECT 1019.430 20.300 1019.750 20.360 ;
        RECT 717.210 20.160 1019.750 20.300 ;
        RECT 717.210 20.100 717.530 20.160 ;
        RECT 1019.430 20.100 1019.750 20.160 ;
      LAYER via ;
        RECT 711.720 202.680 711.980 202.940 ;
        RECT 717.240 202.680 717.500 202.940 ;
        RECT 717.240 20.100 717.500 20.360 ;
        RECT 1019.460 20.100 1019.720 20.360 ;
      LAYER met2 ;
        RECT 711.670 216.000 711.950 220.000 ;
        RECT 711.780 202.970 711.920 216.000 ;
        RECT 711.720 202.650 711.980 202.970 ;
        RECT 717.240 202.650 717.500 202.970 ;
        RECT 717.300 20.390 717.440 202.650 ;
        RECT 717.240 20.070 717.500 20.390 ;
        RECT 1019.460 20.070 1019.720 20.390 ;
        RECT 1019.520 2.400 1019.660 20.070 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 729.630 204.240 729.950 204.300 ;
        RECT 1035.530 204.240 1035.850 204.300 ;
        RECT 729.630 204.100 1035.850 204.240 ;
        RECT 729.630 204.040 729.950 204.100 ;
        RECT 1035.530 204.040 1035.850 204.100 ;
      LAYER via ;
        RECT 729.660 204.040 729.920 204.300 ;
        RECT 1035.560 204.040 1035.820 204.300 ;
      LAYER met2 ;
        RECT 729.610 216.000 729.890 220.000 ;
        RECT 729.720 204.330 729.860 216.000 ;
        RECT 729.660 204.010 729.920 204.330 ;
        RECT 1035.560 204.010 1035.820 204.330 ;
        RECT 1035.620 16.730 1035.760 204.010 ;
        RECT 1035.620 16.590 1037.600 16.730 ;
        RECT 1037.460 2.400 1037.600 16.590 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 747.570 200.500 747.890 200.560 ;
        RECT 751.710 200.500 752.030 200.560 ;
        RECT 747.570 200.360 752.030 200.500 ;
        RECT 747.570 200.300 747.890 200.360 ;
        RECT 751.710 200.300 752.030 200.360 ;
        RECT 751.710 19.620 752.030 19.680 ;
        RECT 1055.310 19.620 1055.630 19.680 ;
        RECT 751.710 19.480 1055.630 19.620 ;
        RECT 751.710 19.420 752.030 19.480 ;
        RECT 1055.310 19.420 1055.630 19.480 ;
      LAYER via ;
        RECT 747.600 200.300 747.860 200.560 ;
        RECT 751.740 200.300 752.000 200.560 ;
        RECT 751.740 19.420 752.000 19.680 ;
        RECT 1055.340 19.420 1055.600 19.680 ;
      LAYER met2 ;
        RECT 747.550 216.000 747.830 220.000 ;
        RECT 747.660 200.590 747.800 216.000 ;
        RECT 747.600 200.270 747.860 200.590 ;
        RECT 751.740 200.270 752.000 200.590 ;
        RECT 751.800 19.710 751.940 200.270 ;
        RECT 751.740 19.390 752.000 19.710 ;
        RECT 1055.340 19.390 1055.600 19.710 ;
        RECT 1055.400 2.400 1055.540 19.390 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 765.510 17.580 765.830 17.640 ;
        RECT 1073.250 17.580 1073.570 17.640 ;
        RECT 765.510 17.440 1073.570 17.580 ;
        RECT 765.510 17.380 765.830 17.440 ;
        RECT 1073.250 17.380 1073.570 17.440 ;
      LAYER via ;
        RECT 765.540 17.380 765.800 17.640 ;
        RECT 1073.280 17.380 1073.540 17.640 ;
      LAYER met2 ;
        RECT 765.490 216.000 765.770 220.000 ;
        RECT 765.600 17.670 765.740 216.000 ;
        RECT 765.540 17.350 765.800 17.670 ;
        RECT 1073.280 17.350 1073.540 17.670 ;
        RECT 1073.340 2.400 1073.480 17.350 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 786.210 17.920 786.530 17.980 ;
        RECT 1090.270 17.920 1090.590 17.980 ;
        RECT 786.210 17.780 1090.590 17.920 ;
        RECT 786.210 17.720 786.530 17.780 ;
        RECT 1090.270 17.720 1090.590 17.780 ;
      LAYER via ;
        RECT 786.240 17.720 786.500 17.980 ;
        RECT 1090.300 17.720 1090.560 17.980 ;
      LAYER met2 ;
        RECT 783.430 216.650 783.710 220.000 ;
        RECT 783.430 216.510 786.440 216.650 ;
        RECT 783.430 216.000 783.710 216.510 ;
        RECT 786.300 18.010 786.440 216.510 ;
        RECT 786.240 17.690 786.500 18.010 ;
        RECT 1090.300 17.690 1090.560 18.010 ;
        RECT 1090.360 16.730 1090.500 17.690 ;
        RECT 1090.360 16.590 1090.960 16.730 ;
        RECT 1090.820 2.400 1090.960 16.590 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 801.390 200.500 801.710 200.560 ;
        RECT 806.910 200.500 807.230 200.560 ;
        RECT 801.390 200.360 807.230 200.500 ;
        RECT 801.390 200.300 801.710 200.360 ;
        RECT 806.910 200.300 807.230 200.360 ;
        RECT 806.910 19.960 807.230 20.020 ;
        RECT 1108.670 19.960 1108.990 20.020 ;
        RECT 806.910 19.820 1108.990 19.960 ;
        RECT 806.910 19.760 807.230 19.820 ;
        RECT 1108.670 19.760 1108.990 19.820 ;
      LAYER via ;
        RECT 801.420 200.300 801.680 200.560 ;
        RECT 806.940 200.300 807.200 200.560 ;
        RECT 806.940 19.760 807.200 20.020 ;
        RECT 1108.700 19.760 1108.960 20.020 ;
      LAYER met2 ;
        RECT 801.370 216.000 801.650 220.000 ;
        RECT 801.480 200.590 801.620 216.000 ;
        RECT 801.420 200.270 801.680 200.590 ;
        RECT 806.940 200.270 807.200 200.590 ;
        RECT 807.000 20.050 807.140 200.270 ;
        RECT 806.940 19.730 807.200 20.050 ;
        RECT 1108.700 19.730 1108.960 20.050 ;
        RECT 1108.760 2.400 1108.900 19.730 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 820.710 19.280 821.030 19.340 ;
        RECT 1126.610 19.280 1126.930 19.340 ;
        RECT 820.710 19.140 1126.930 19.280 ;
        RECT 820.710 19.080 821.030 19.140 ;
        RECT 1126.610 19.080 1126.930 19.140 ;
      LAYER via ;
        RECT 820.740 19.080 821.000 19.340 ;
        RECT 1126.640 19.080 1126.900 19.340 ;
      LAYER met2 ;
        RECT 819.310 216.650 819.590 220.000 ;
        RECT 819.310 216.510 820.940 216.650 ;
        RECT 819.310 216.000 819.590 216.510 ;
        RECT 820.800 19.370 820.940 216.510 ;
        RECT 820.740 19.050 821.000 19.370 ;
        RECT 1126.640 19.050 1126.900 19.370 ;
        RECT 1126.700 2.400 1126.840 19.050 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 836.810 205.940 837.130 206.000 ;
        RECT 1139.490 205.940 1139.810 206.000 ;
        RECT 836.810 205.800 1139.810 205.940 ;
        RECT 836.810 205.740 837.130 205.800 ;
        RECT 1139.490 205.740 1139.810 205.800 ;
      LAYER via ;
        RECT 836.840 205.740 837.100 206.000 ;
        RECT 1139.520 205.740 1139.780 206.000 ;
      LAYER met2 ;
        RECT 836.790 216.000 837.070 220.000 ;
        RECT 836.900 206.030 837.040 216.000 ;
        RECT 836.840 205.710 837.100 206.030 ;
        RECT 1139.520 205.710 1139.780 206.030 ;
        RECT 1139.580 16.730 1139.720 205.710 ;
        RECT 1139.580 16.590 1144.780 16.730 ;
        RECT 1144.640 2.400 1144.780 16.590 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 855.210 17.240 855.530 17.300 ;
        RECT 1162.490 17.240 1162.810 17.300 ;
        RECT 855.210 17.100 1162.810 17.240 ;
        RECT 855.210 17.040 855.530 17.100 ;
        RECT 1162.490 17.040 1162.810 17.100 ;
      LAYER via ;
        RECT 855.240 17.040 855.500 17.300 ;
        RECT 1162.520 17.040 1162.780 17.300 ;
      LAYER met2 ;
        RECT 854.730 216.650 855.010 220.000 ;
        RECT 854.730 216.510 855.440 216.650 ;
        RECT 854.730 216.000 855.010 216.510 ;
        RECT 855.300 17.330 855.440 216.510 ;
        RECT 855.240 17.010 855.500 17.330 ;
        RECT 1162.520 17.010 1162.780 17.330 ;
        RECT 1162.580 2.400 1162.720 17.010 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 371.750 17.240 372.070 17.300 ;
        RECT 680.410 17.240 680.730 17.300 ;
        RECT 371.750 17.100 680.730 17.240 ;
        RECT 371.750 17.040 372.070 17.100 ;
        RECT 680.410 17.040 680.730 17.100 ;
      LAYER via ;
        RECT 371.780 17.040 372.040 17.300 ;
        RECT 680.440 17.040 680.700 17.300 ;
      LAYER met2 ;
        RECT 372.190 216.650 372.470 220.000 ;
        RECT 371.840 216.510 372.470 216.650 ;
        RECT 371.840 17.330 371.980 216.510 ;
        RECT 372.190 216.000 372.470 216.510 ;
        RECT 371.780 17.010 372.040 17.330 ;
        RECT 680.440 17.010 680.700 17.330 ;
        RECT 680.500 2.400 680.640 17.010 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 872.690 204.580 873.010 204.640 ;
        RECT 1180.890 204.580 1181.210 204.640 ;
        RECT 872.690 204.440 1181.210 204.580 ;
        RECT 872.690 204.380 873.010 204.440 ;
        RECT 1180.890 204.380 1181.210 204.440 ;
      LAYER via ;
        RECT 872.720 204.380 872.980 204.640 ;
        RECT 1180.920 204.380 1181.180 204.640 ;
      LAYER met2 ;
        RECT 872.670 216.000 872.950 220.000 ;
        RECT 872.780 204.670 872.920 216.000 ;
        RECT 872.720 204.350 872.980 204.670 ;
        RECT 1180.920 204.350 1181.180 204.670 ;
        RECT 1180.980 17.410 1181.120 204.350 ;
        RECT 1180.060 17.270 1181.120 17.410 ;
        RECT 1180.060 2.400 1180.200 17.270 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 890.630 200.500 890.950 200.560 ;
        RECT 896.610 200.500 896.930 200.560 ;
        RECT 890.630 200.360 896.930 200.500 ;
        RECT 890.630 200.300 890.950 200.360 ;
        RECT 896.610 200.300 896.930 200.360 ;
        RECT 896.610 16.560 896.930 16.620 ;
        RECT 1197.910 16.560 1198.230 16.620 ;
        RECT 896.610 16.420 1198.230 16.560 ;
        RECT 896.610 16.360 896.930 16.420 ;
        RECT 1197.910 16.360 1198.230 16.420 ;
      LAYER via ;
        RECT 890.660 200.300 890.920 200.560 ;
        RECT 896.640 200.300 896.900 200.560 ;
        RECT 896.640 16.360 896.900 16.620 ;
        RECT 1197.940 16.360 1198.200 16.620 ;
      LAYER met2 ;
        RECT 890.610 216.000 890.890 220.000 ;
        RECT 890.720 200.590 890.860 216.000 ;
        RECT 890.660 200.270 890.920 200.590 ;
        RECT 896.640 200.270 896.900 200.590 ;
        RECT 896.700 16.650 896.840 200.270 ;
        RECT 896.640 16.330 896.900 16.650 ;
        RECT 1197.940 16.330 1198.200 16.650 ;
        RECT 1198.000 2.400 1198.140 16.330 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 908.570 203.560 908.890 203.620 ;
        RECT 1214.930 203.560 1215.250 203.620 ;
        RECT 908.570 203.420 1215.250 203.560 ;
        RECT 908.570 203.360 908.890 203.420 ;
        RECT 1214.930 203.360 1215.250 203.420 ;
      LAYER via ;
        RECT 908.600 203.360 908.860 203.620 ;
        RECT 1214.960 203.360 1215.220 203.620 ;
      LAYER met2 ;
        RECT 908.550 216.000 908.830 220.000 ;
        RECT 908.660 203.650 908.800 216.000 ;
        RECT 908.600 203.330 908.860 203.650 ;
        RECT 1214.960 203.330 1215.220 203.650 ;
        RECT 1215.020 16.730 1215.160 203.330 ;
        RECT 1215.020 16.590 1216.080 16.730 ;
        RECT 1215.940 2.400 1216.080 16.590 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 926.510 200.500 926.830 200.560 ;
        RECT 931.110 200.500 931.430 200.560 ;
        RECT 926.510 200.360 931.430 200.500 ;
        RECT 926.510 200.300 926.830 200.360 ;
        RECT 931.110 200.300 931.430 200.360 ;
        RECT 931.110 16.900 931.430 16.960 ;
        RECT 1233.790 16.900 1234.110 16.960 ;
        RECT 931.110 16.760 1234.110 16.900 ;
        RECT 931.110 16.700 931.430 16.760 ;
        RECT 1233.790 16.700 1234.110 16.760 ;
      LAYER via ;
        RECT 926.540 200.300 926.800 200.560 ;
        RECT 931.140 200.300 931.400 200.560 ;
        RECT 931.140 16.700 931.400 16.960 ;
        RECT 1233.820 16.700 1234.080 16.960 ;
      LAYER met2 ;
        RECT 926.490 216.000 926.770 220.000 ;
        RECT 926.600 200.590 926.740 216.000 ;
        RECT 926.540 200.270 926.800 200.590 ;
        RECT 931.140 200.270 931.400 200.590 ;
        RECT 931.200 16.990 931.340 200.270 ;
        RECT 931.140 16.670 931.400 16.990 ;
        RECT 1233.820 16.670 1234.080 16.990 ;
        RECT 1233.880 2.400 1234.020 16.670 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 944.450 205.600 944.770 205.660 ;
        RECT 1249.430 205.600 1249.750 205.660 ;
        RECT 944.450 205.460 1249.750 205.600 ;
        RECT 944.450 205.400 944.770 205.460 ;
        RECT 1249.430 205.400 1249.750 205.460 ;
      LAYER via ;
        RECT 944.480 205.400 944.740 205.660 ;
        RECT 1249.460 205.400 1249.720 205.660 ;
      LAYER met2 ;
        RECT 944.430 216.000 944.710 220.000 ;
        RECT 944.540 205.690 944.680 216.000 ;
        RECT 944.480 205.370 944.740 205.690 ;
        RECT 1249.460 205.370 1249.720 205.690 ;
        RECT 1249.520 16.730 1249.660 205.370 ;
        RECT 1249.520 16.590 1251.960 16.730 ;
        RECT 1251.820 2.400 1251.960 16.590 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 965.610 15.880 965.930 15.940 ;
        RECT 1269.210 15.880 1269.530 15.940 ;
        RECT 965.610 15.740 1269.530 15.880 ;
        RECT 965.610 15.680 965.930 15.740 ;
        RECT 1269.210 15.680 1269.530 15.740 ;
      LAYER via ;
        RECT 965.640 15.680 965.900 15.940 ;
        RECT 1269.240 15.680 1269.500 15.940 ;
      LAYER met2 ;
        RECT 961.910 216.650 962.190 220.000 ;
        RECT 961.910 216.510 965.840 216.650 ;
        RECT 961.910 216.000 962.190 216.510 ;
        RECT 965.700 15.970 965.840 216.510 ;
        RECT 965.640 15.650 965.900 15.970 ;
        RECT 1269.240 15.650 1269.500 15.970 ;
        RECT 1269.300 2.400 1269.440 15.650 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 979.870 200.500 980.190 200.560 ;
        RECT 986.310 200.500 986.630 200.560 ;
        RECT 979.870 200.360 986.630 200.500 ;
        RECT 979.870 200.300 980.190 200.360 ;
        RECT 986.310 200.300 986.630 200.360 ;
        RECT 986.310 20.640 986.630 20.700 ;
        RECT 1287.150 20.640 1287.470 20.700 ;
        RECT 986.310 20.500 1287.470 20.640 ;
        RECT 986.310 20.440 986.630 20.500 ;
        RECT 1287.150 20.440 1287.470 20.500 ;
      LAYER via ;
        RECT 979.900 200.300 980.160 200.560 ;
        RECT 986.340 200.300 986.600 200.560 ;
        RECT 986.340 20.440 986.600 20.700 ;
        RECT 1287.180 20.440 1287.440 20.700 ;
      LAYER met2 ;
        RECT 979.850 216.000 980.130 220.000 ;
        RECT 979.960 200.590 980.100 216.000 ;
        RECT 979.900 200.270 980.160 200.590 ;
        RECT 986.340 200.270 986.600 200.590 ;
        RECT 986.400 20.730 986.540 200.270 ;
        RECT 986.340 20.410 986.600 20.730 ;
        RECT 1287.180 20.410 1287.440 20.730 ;
        RECT 1287.240 2.400 1287.380 20.410 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1000.110 18.940 1000.430 19.000 ;
        RECT 1305.090 18.940 1305.410 19.000 ;
        RECT 1000.110 18.800 1305.410 18.940 ;
        RECT 1000.110 18.740 1000.430 18.800 ;
        RECT 1305.090 18.740 1305.410 18.800 ;
      LAYER via ;
        RECT 1000.140 18.740 1000.400 19.000 ;
        RECT 1305.120 18.740 1305.380 19.000 ;
      LAYER met2 ;
        RECT 997.790 216.650 998.070 220.000 ;
        RECT 997.790 216.510 1000.340 216.650 ;
        RECT 997.790 216.000 998.070 216.510 ;
        RECT 1000.200 19.030 1000.340 216.510 ;
        RECT 1000.140 18.710 1000.400 19.030 ;
        RECT 1305.120 18.710 1305.380 19.030 ;
        RECT 1305.180 2.400 1305.320 18.710 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1015.750 200.500 1016.070 200.560 ;
        RECT 1020.810 200.500 1021.130 200.560 ;
        RECT 1015.750 200.360 1021.130 200.500 ;
        RECT 1015.750 200.300 1016.070 200.360 ;
        RECT 1020.810 200.300 1021.130 200.360 ;
        RECT 1020.810 20.300 1021.130 20.360 ;
        RECT 1323.030 20.300 1323.350 20.360 ;
        RECT 1020.810 20.160 1323.350 20.300 ;
        RECT 1020.810 20.100 1021.130 20.160 ;
        RECT 1323.030 20.100 1323.350 20.160 ;
      LAYER via ;
        RECT 1015.780 200.300 1016.040 200.560 ;
        RECT 1020.840 200.300 1021.100 200.560 ;
        RECT 1020.840 20.100 1021.100 20.360 ;
        RECT 1323.060 20.100 1323.320 20.360 ;
      LAYER met2 ;
        RECT 1015.730 216.000 1016.010 220.000 ;
        RECT 1015.840 200.590 1015.980 216.000 ;
        RECT 1015.780 200.270 1016.040 200.590 ;
        RECT 1020.840 200.270 1021.100 200.590 ;
        RECT 1020.900 20.390 1021.040 200.270 ;
        RECT 1020.840 20.070 1021.100 20.390 ;
        RECT 1323.060 20.070 1323.320 20.390 ;
        RECT 1323.120 2.400 1323.260 20.070 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1034.610 18.600 1034.930 18.660 ;
        RECT 1340.510 18.600 1340.830 18.660 ;
        RECT 1034.610 18.460 1340.830 18.600 ;
        RECT 1034.610 18.400 1034.930 18.460 ;
        RECT 1340.510 18.400 1340.830 18.460 ;
      LAYER via ;
        RECT 1034.640 18.400 1034.900 18.660 ;
        RECT 1340.540 18.400 1340.800 18.660 ;
      LAYER met2 ;
        RECT 1033.670 216.650 1033.950 220.000 ;
        RECT 1033.670 216.510 1034.840 216.650 ;
        RECT 1033.670 216.000 1033.950 216.510 ;
        RECT 1034.700 18.690 1034.840 216.510 ;
        RECT 1034.640 18.370 1034.900 18.690 ;
        RECT 1340.540 18.370 1340.800 18.690 ;
        RECT 1340.600 2.400 1340.740 18.370 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 17.920 698.670 17.980 ;
        RECT 663.020 17.780 698.670 17.920 ;
        RECT 392.910 17.580 393.230 17.640 ;
        RECT 663.020 17.580 663.160 17.780 ;
        RECT 698.350 17.720 698.670 17.780 ;
        RECT 392.910 17.440 663.160 17.580 ;
        RECT 392.910 17.380 393.230 17.440 ;
      LAYER via ;
        RECT 392.940 17.380 393.200 17.640 ;
        RECT 698.380 17.720 698.640 17.980 ;
      LAYER met2 ;
        RECT 390.130 216.650 390.410 220.000 ;
        RECT 390.130 216.510 393.140 216.650 ;
        RECT 390.130 216.000 390.410 216.510 ;
        RECT 393.000 17.670 393.140 216.510 ;
        RECT 698.380 17.690 698.640 18.010 ;
        RECT 392.940 17.350 393.200 17.670 ;
        RECT 698.440 2.400 698.580 17.690 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1051.630 204.920 1051.950 204.980 ;
        RECT 1352.470 204.920 1352.790 204.980 ;
        RECT 1051.630 204.780 1352.790 204.920 ;
        RECT 1051.630 204.720 1051.950 204.780 ;
        RECT 1352.470 204.720 1352.790 204.780 ;
        RECT 1352.470 16.560 1352.790 16.620 ;
        RECT 1358.450 16.560 1358.770 16.620 ;
        RECT 1352.470 16.420 1358.770 16.560 ;
        RECT 1352.470 16.360 1352.790 16.420 ;
        RECT 1358.450 16.360 1358.770 16.420 ;
      LAYER via ;
        RECT 1051.660 204.720 1051.920 204.980 ;
        RECT 1352.500 204.720 1352.760 204.980 ;
        RECT 1352.500 16.360 1352.760 16.620 ;
        RECT 1358.480 16.360 1358.740 16.620 ;
      LAYER met2 ;
        RECT 1051.610 216.000 1051.890 220.000 ;
        RECT 1051.720 205.010 1051.860 216.000 ;
        RECT 1051.660 204.690 1051.920 205.010 ;
        RECT 1352.500 204.690 1352.760 205.010 ;
        RECT 1352.560 16.650 1352.700 204.690 ;
        RECT 1352.500 16.330 1352.760 16.650 ;
        RECT 1358.480 16.330 1358.740 16.650 ;
        RECT 1358.540 2.400 1358.680 16.330 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1069.570 200.500 1069.890 200.560 ;
        RECT 1076.010 200.500 1076.330 200.560 ;
        RECT 1069.570 200.360 1076.330 200.500 ;
        RECT 1069.570 200.300 1069.890 200.360 ;
        RECT 1076.010 200.300 1076.330 200.360 ;
        RECT 1076.010 19.620 1076.330 19.680 ;
        RECT 1376.390 19.620 1376.710 19.680 ;
        RECT 1076.010 19.480 1376.710 19.620 ;
        RECT 1076.010 19.420 1076.330 19.480 ;
        RECT 1376.390 19.420 1376.710 19.480 ;
      LAYER via ;
        RECT 1069.600 200.300 1069.860 200.560 ;
        RECT 1076.040 200.300 1076.300 200.560 ;
        RECT 1076.040 19.420 1076.300 19.680 ;
        RECT 1376.420 19.420 1376.680 19.680 ;
      LAYER met2 ;
        RECT 1069.550 216.000 1069.830 220.000 ;
        RECT 1069.660 200.590 1069.800 216.000 ;
        RECT 1069.600 200.270 1069.860 200.590 ;
        RECT 1076.040 200.270 1076.300 200.590 ;
        RECT 1076.100 19.710 1076.240 200.270 ;
        RECT 1076.040 19.390 1076.300 19.710 ;
        RECT 1376.420 19.390 1376.680 19.710 ;
        RECT 1376.480 2.400 1376.620 19.390 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1087.050 204.240 1087.370 204.300 ;
        RECT 1394.790 204.240 1395.110 204.300 ;
        RECT 1087.050 204.100 1395.110 204.240 ;
        RECT 1087.050 204.040 1087.370 204.100 ;
        RECT 1394.790 204.040 1395.110 204.100 ;
      LAYER via ;
        RECT 1087.080 204.040 1087.340 204.300 ;
        RECT 1394.820 204.040 1395.080 204.300 ;
      LAYER met2 ;
        RECT 1087.030 216.000 1087.310 220.000 ;
        RECT 1087.140 204.330 1087.280 216.000 ;
        RECT 1087.080 204.010 1087.340 204.330 ;
        RECT 1394.820 204.010 1395.080 204.330 ;
        RECT 1394.880 17.410 1395.020 204.010 ;
        RECT 1394.420 17.270 1395.020 17.410 ;
        RECT 1394.420 2.400 1394.560 17.270 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1104.990 200.500 1105.310 200.560 ;
        RECT 1110.510 200.500 1110.830 200.560 ;
        RECT 1104.990 200.360 1110.830 200.500 ;
        RECT 1104.990 200.300 1105.310 200.360 ;
        RECT 1110.510 200.300 1110.830 200.360 ;
        RECT 1110.510 16.220 1110.830 16.280 ;
        RECT 1412.270 16.220 1412.590 16.280 ;
        RECT 1110.510 16.080 1412.590 16.220 ;
        RECT 1110.510 16.020 1110.830 16.080 ;
        RECT 1412.270 16.020 1412.590 16.080 ;
      LAYER via ;
        RECT 1105.020 200.300 1105.280 200.560 ;
        RECT 1110.540 200.300 1110.800 200.560 ;
        RECT 1110.540 16.020 1110.800 16.280 ;
        RECT 1412.300 16.020 1412.560 16.280 ;
      LAYER met2 ;
        RECT 1104.970 216.000 1105.250 220.000 ;
        RECT 1105.080 200.590 1105.220 216.000 ;
        RECT 1105.020 200.270 1105.280 200.590 ;
        RECT 1110.540 200.270 1110.800 200.590 ;
        RECT 1110.600 16.310 1110.740 200.270 ;
        RECT 1110.540 15.990 1110.800 16.310 ;
        RECT 1412.300 15.990 1412.560 16.310 ;
        RECT 1412.360 2.400 1412.500 15.990 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1122.930 203.900 1123.250 203.960 ;
        RECT 1428.830 203.900 1429.150 203.960 ;
        RECT 1122.930 203.760 1429.150 203.900 ;
        RECT 1122.930 203.700 1123.250 203.760 ;
        RECT 1428.830 203.700 1429.150 203.760 ;
      LAYER via ;
        RECT 1122.960 203.700 1123.220 203.960 ;
        RECT 1428.860 203.700 1429.120 203.960 ;
      LAYER met2 ;
        RECT 1122.910 216.000 1123.190 220.000 ;
        RECT 1123.020 203.990 1123.160 216.000 ;
        RECT 1122.960 203.670 1123.220 203.990 ;
        RECT 1428.860 203.670 1429.120 203.990 ;
        RECT 1428.920 16.730 1429.060 203.670 ;
        RECT 1428.920 16.590 1429.980 16.730 ;
        RECT 1429.840 2.400 1429.980 16.590 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1140.870 200.500 1141.190 200.560 ;
        RECT 1145.010 200.500 1145.330 200.560 ;
        RECT 1140.870 200.360 1145.330 200.500 ;
        RECT 1140.870 200.300 1141.190 200.360 ;
        RECT 1145.010 200.300 1145.330 200.360 ;
        RECT 1145.010 19.280 1145.330 19.340 ;
        RECT 1447.690 19.280 1448.010 19.340 ;
        RECT 1145.010 19.140 1448.010 19.280 ;
        RECT 1145.010 19.080 1145.330 19.140 ;
        RECT 1447.690 19.080 1448.010 19.140 ;
      LAYER via ;
        RECT 1140.900 200.300 1141.160 200.560 ;
        RECT 1145.040 200.300 1145.300 200.560 ;
        RECT 1145.040 19.080 1145.300 19.340 ;
        RECT 1447.720 19.080 1447.980 19.340 ;
      LAYER met2 ;
        RECT 1140.850 216.000 1141.130 220.000 ;
        RECT 1140.960 200.590 1141.100 216.000 ;
        RECT 1140.900 200.270 1141.160 200.590 ;
        RECT 1145.040 200.270 1145.300 200.590 ;
        RECT 1145.100 19.370 1145.240 200.270 ;
        RECT 1145.040 19.050 1145.300 19.370 ;
        RECT 1447.720 19.050 1447.980 19.370 ;
        RECT 1447.780 2.400 1447.920 19.050 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1158.810 17.580 1159.130 17.640 ;
        RECT 1465.630 17.580 1465.950 17.640 ;
        RECT 1158.810 17.440 1465.950 17.580 ;
        RECT 1158.810 17.380 1159.130 17.440 ;
        RECT 1465.630 17.380 1465.950 17.440 ;
      LAYER via ;
        RECT 1158.840 17.380 1159.100 17.640 ;
        RECT 1465.660 17.380 1465.920 17.640 ;
      LAYER met2 ;
        RECT 1158.790 216.000 1159.070 220.000 ;
        RECT 1158.900 17.670 1159.040 216.000 ;
        RECT 1158.840 17.350 1159.100 17.670 ;
        RECT 1465.660 17.350 1465.920 17.670 ;
        RECT 1465.720 2.400 1465.860 17.350 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.510 18.260 1179.830 18.320 ;
        RECT 1483.570 18.260 1483.890 18.320 ;
        RECT 1179.510 18.120 1483.890 18.260 ;
        RECT 1179.510 18.060 1179.830 18.120 ;
        RECT 1483.570 18.060 1483.890 18.120 ;
      LAYER via ;
        RECT 1179.540 18.060 1179.800 18.320 ;
        RECT 1483.600 18.060 1483.860 18.320 ;
      LAYER met2 ;
        RECT 1176.730 216.650 1177.010 220.000 ;
        RECT 1176.730 216.510 1179.740 216.650 ;
        RECT 1176.730 216.000 1177.010 216.510 ;
        RECT 1179.600 18.350 1179.740 216.510 ;
        RECT 1179.540 18.030 1179.800 18.350 ;
        RECT 1483.600 18.030 1483.860 18.350 ;
        RECT 1483.660 2.400 1483.800 18.030 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.690 200.500 1195.010 200.560 ;
        RECT 1200.210 200.500 1200.530 200.560 ;
        RECT 1194.690 200.360 1200.530 200.500 ;
        RECT 1194.690 200.300 1195.010 200.360 ;
        RECT 1200.210 200.300 1200.530 200.360 ;
        RECT 1200.210 19.960 1200.530 20.020 ;
        RECT 1501.510 19.960 1501.830 20.020 ;
        RECT 1200.210 19.820 1501.830 19.960 ;
        RECT 1200.210 19.760 1200.530 19.820 ;
        RECT 1501.510 19.760 1501.830 19.820 ;
      LAYER via ;
        RECT 1194.720 200.300 1194.980 200.560 ;
        RECT 1200.240 200.300 1200.500 200.560 ;
        RECT 1200.240 19.760 1200.500 20.020 ;
        RECT 1501.540 19.760 1501.800 20.020 ;
      LAYER met2 ;
        RECT 1194.670 216.000 1194.950 220.000 ;
        RECT 1194.780 200.590 1194.920 216.000 ;
        RECT 1194.720 200.270 1194.980 200.590 ;
        RECT 1200.240 200.270 1200.500 200.590 ;
        RECT 1200.300 20.050 1200.440 200.270 ;
        RECT 1200.240 19.730 1200.500 20.050 ;
        RECT 1501.540 19.730 1501.800 20.050 ;
        RECT 1501.600 2.400 1501.740 19.730 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.010 17.920 1214.330 17.980 ;
        RECT 1518.990 17.920 1519.310 17.980 ;
        RECT 1214.010 17.780 1519.310 17.920 ;
        RECT 1214.010 17.720 1214.330 17.780 ;
        RECT 1518.990 17.720 1519.310 17.780 ;
      LAYER via ;
        RECT 1214.040 17.720 1214.300 17.980 ;
        RECT 1519.020 17.720 1519.280 17.980 ;
      LAYER met2 ;
        RECT 1212.150 216.650 1212.430 220.000 ;
        RECT 1212.150 216.510 1214.240 216.650 ;
        RECT 1212.150 216.000 1212.430 216.510 ;
        RECT 1214.100 18.010 1214.240 216.510 ;
        RECT 1214.040 17.690 1214.300 18.010 ;
        RECT 1519.020 17.690 1519.280 18.010 ;
        RECT 1519.080 2.400 1519.220 17.690 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 408.090 205.940 408.410 206.000 ;
        RECT 711.230 205.940 711.550 206.000 ;
        RECT 408.090 205.800 711.550 205.940 ;
        RECT 408.090 205.740 408.410 205.800 ;
        RECT 711.230 205.740 711.550 205.800 ;
      LAYER via ;
        RECT 408.120 205.740 408.380 206.000 ;
        RECT 711.260 205.740 711.520 206.000 ;
      LAYER met2 ;
        RECT 408.070 216.000 408.350 220.000 ;
        RECT 408.180 206.030 408.320 216.000 ;
        RECT 408.120 205.710 408.380 206.030 ;
        RECT 711.260 205.710 711.520 206.030 ;
        RECT 711.320 16.730 711.460 205.710 ;
        RECT 711.320 16.590 716.520 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1230.110 200.500 1230.430 200.560 ;
        RECT 1234.710 200.500 1235.030 200.560 ;
        RECT 1230.110 200.360 1235.030 200.500 ;
        RECT 1230.110 200.300 1230.430 200.360 ;
        RECT 1234.710 200.300 1235.030 200.360 ;
        RECT 1234.710 16.900 1235.030 16.960 ;
        RECT 1536.930 16.900 1537.250 16.960 ;
        RECT 1234.710 16.760 1537.250 16.900 ;
        RECT 1234.710 16.700 1235.030 16.760 ;
        RECT 1536.930 16.700 1537.250 16.760 ;
      LAYER via ;
        RECT 1230.140 200.300 1230.400 200.560 ;
        RECT 1234.740 200.300 1235.000 200.560 ;
        RECT 1234.740 16.700 1235.000 16.960 ;
        RECT 1536.960 16.700 1537.220 16.960 ;
      LAYER met2 ;
        RECT 1230.090 216.000 1230.370 220.000 ;
        RECT 1230.200 200.590 1230.340 216.000 ;
        RECT 1230.140 200.270 1230.400 200.590 ;
        RECT 1234.740 200.270 1235.000 200.590 ;
        RECT 1234.800 16.990 1234.940 200.270 ;
        RECT 1234.740 16.670 1235.000 16.990 ;
        RECT 1536.960 16.670 1537.220 16.990 ;
        RECT 1537.020 2.400 1537.160 16.670 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.510 17.240 1248.830 17.300 ;
        RECT 1554.870 17.240 1555.190 17.300 ;
        RECT 1248.510 17.100 1555.190 17.240 ;
        RECT 1248.510 17.040 1248.830 17.100 ;
        RECT 1554.870 17.040 1555.190 17.100 ;
      LAYER via ;
        RECT 1248.540 17.040 1248.800 17.300 ;
        RECT 1554.900 17.040 1555.160 17.300 ;
      LAYER met2 ;
        RECT 1248.030 216.650 1248.310 220.000 ;
        RECT 1248.030 216.510 1248.740 216.650 ;
        RECT 1248.030 216.000 1248.310 216.510 ;
        RECT 1248.600 17.330 1248.740 216.510 ;
        RECT 1248.540 17.010 1248.800 17.330 ;
        RECT 1554.900 17.010 1555.160 17.330 ;
        RECT 1554.960 2.400 1555.100 17.010 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1352.545 205.445 1352.715 206.635 ;
        RECT 1373.705 205.105 1373.875 206.635 ;
        RECT 1400.845 205.105 1401.015 205.955 ;
        RECT 1448.685 205.105 1448.855 205.955 ;
        RECT 1449.145 204.765 1449.775 204.935 ;
        RECT 1545.745 204.085 1545.915 204.935 ;
      LAYER mcon ;
        RECT 1352.545 206.465 1352.715 206.635 ;
        RECT 1373.705 206.465 1373.875 206.635 ;
        RECT 1400.845 205.785 1401.015 205.955 ;
        RECT 1448.685 205.785 1448.855 205.955 ;
        RECT 1449.605 204.765 1449.775 204.935 ;
        RECT 1545.745 204.765 1545.915 204.935 ;
      LAYER met1 ;
        RECT 1352.485 206.620 1352.775 206.665 ;
        RECT 1373.645 206.620 1373.935 206.665 ;
        RECT 1352.485 206.480 1373.935 206.620 ;
        RECT 1352.485 206.435 1352.775 206.480 ;
        RECT 1373.645 206.435 1373.935 206.480 ;
        RECT 1265.990 205.940 1266.310 206.000 ;
        RECT 1400.785 205.940 1401.075 205.985 ;
        RECT 1448.625 205.940 1448.915 205.985 ;
        RECT 1265.990 205.800 1269.900 205.940 ;
        RECT 1265.990 205.740 1266.310 205.800 ;
        RECT 1269.760 205.600 1269.900 205.800 ;
        RECT 1400.785 205.800 1448.915 205.940 ;
        RECT 1400.785 205.755 1401.075 205.800 ;
        RECT 1448.625 205.755 1448.915 205.800 ;
        RECT 1352.485 205.600 1352.775 205.645 ;
        RECT 1269.760 205.460 1352.775 205.600 ;
        RECT 1352.485 205.415 1352.775 205.460 ;
        RECT 1373.645 205.260 1373.935 205.305 ;
        RECT 1400.785 205.260 1401.075 205.305 ;
        RECT 1373.645 205.120 1401.075 205.260 ;
        RECT 1373.645 205.075 1373.935 205.120 ;
        RECT 1400.785 205.075 1401.075 205.120 ;
        RECT 1448.625 205.260 1448.915 205.305 ;
        RECT 1448.625 205.120 1449.300 205.260 ;
        RECT 1448.625 205.075 1448.915 205.120 ;
        RECT 1449.160 204.965 1449.300 205.120 ;
        RECT 1449.085 204.735 1449.375 204.965 ;
        RECT 1449.545 204.920 1449.835 204.965 ;
        RECT 1545.685 204.920 1545.975 204.965 ;
        RECT 1449.545 204.780 1545.975 204.920 ;
        RECT 1449.545 204.735 1449.835 204.780 ;
        RECT 1545.685 204.735 1545.975 204.780 ;
        RECT 1545.685 204.240 1545.975 204.285 ;
        RECT 1567.290 204.240 1567.610 204.300 ;
        RECT 1545.685 204.100 1567.610 204.240 ;
        RECT 1545.685 204.055 1545.975 204.100 ;
        RECT 1567.290 204.040 1567.610 204.100 ;
      LAYER via ;
        RECT 1266.020 205.740 1266.280 206.000 ;
        RECT 1567.320 204.040 1567.580 204.300 ;
      LAYER met2 ;
        RECT 1265.970 216.000 1266.250 220.000 ;
        RECT 1266.080 206.030 1266.220 216.000 ;
        RECT 1266.020 205.710 1266.280 206.030 ;
        RECT 1567.320 204.010 1567.580 204.330 ;
        RECT 1567.380 16.730 1567.520 204.010 ;
        RECT 1567.380 16.590 1573.040 16.730 ;
        RECT 1572.900 2.400 1573.040 16.590 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.930 200.500 1284.250 200.560 ;
        RECT 1289.910 200.500 1290.230 200.560 ;
        RECT 1283.930 200.360 1290.230 200.500 ;
        RECT 1283.930 200.300 1284.250 200.360 ;
        RECT 1289.910 200.300 1290.230 200.360 ;
        RECT 1289.910 20.640 1290.230 20.700 ;
        RECT 1590.290 20.640 1590.610 20.700 ;
        RECT 1289.910 20.500 1590.610 20.640 ;
        RECT 1289.910 20.440 1290.230 20.500 ;
        RECT 1590.290 20.440 1590.610 20.500 ;
      LAYER via ;
        RECT 1283.960 200.300 1284.220 200.560 ;
        RECT 1289.940 200.300 1290.200 200.560 ;
        RECT 1289.940 20.440 1290.200 20.700 ;
        RECT 1590.320 20.440 1590.580 20.700 ;
      LAYER met2 ;
        RECT 1283.910 216.000 1284.190 220.000 ;
        RECT 1284.020 200.590 1284.160 216.000 ;
        RECT 1283.960 200.270 1284.220 200.590 ;
        RECT 1289.940 200.270 1290.200 200.590 ;
        RECT 1290.000 20.730 1290.140 200.270 ;
        RECT 1289.940 20.410 1290.200 20.730 ;
        RECT 1590.320 20.410 1590.580 20.730 ;
        RECT 1590.380 2.400 1590.520 20.410 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1301.870 203.560 1302.190 203.620 ;
        RECT 1608.690 203.560 1609.010 203.620 ;
        RECT 1301.870 203.420 1609.010 203.560 ;
        RECT 1301.870 203.360 1302.190 203.420 ;
        RECT 1608.690 203.360 1609.010 203.420 ;
      LAYER via ;
        RECT 1301.900 203.360 1302.160 203.620 ;
        RECT 1608.720 203.360 1608.980 203.620 ;
      LAYER met2 ;
        RECT 1301.850 216.000 1302.130 220.000 ;
        RECT 1301.960 203.650 1302.100 216.000 ;
        RECT 1301.900 203.330 1302.160 203.650 ;
        RECT 1608.720 203.330 1608.980 203.650 ;
        RECT 1608.780 17.410 1608.920 203.330 ;
        RECT 1608.320 17.270 1608.920 17.410 ;
        RECT 1608.320 2.400 1608.460 17.270 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1319.810 200.500 1320.130 200.560 ;
        RECT 1324.410 200.500 1324.730 200.560 ;
        RECT 1319.810 200.360 1324.730 200.500 ;
        RECT 1319.810 200.300 1320.130 200.360 ;
        RECT 1324.410 200.300 1324.730 200.360 ;
        RECT 1324.410 20.300 1324.730 20.360 ;
        RECT 1626.170 20.300 1626.490 20.360 ;
        RECT 1324.410 20.160 1626.490 20.300 ;
        RECT 1324.410 20.100 1324.730 20.160 ;
        RECT 1626.170 20.100 1626.490 20.160 ;
      LAYER via ;
        RECT 1319.840 200.300 1320.100 200.560 ;
        RECT 1324.440 200.300 1324.700 200.560 ;
        RECT 1324.440 20.100 1324.700 20.360 ;
        RECT 1626.200 20.100 1626.460 20.360 ;
      LAYER met2 ;
        RECT 1319.790 216.000 1320.070 220.000 ;
        RECT 1319.900 200.590 1320.040 216.000 ;
        RECT 1319.840 200.270 1320.100 200.590 ;
        RECT 1324.440 200.270 1324.700 200.590 ;
        RECT 1324.500 20.390 1324.640 200.270 ;
        RECT 1324.440 20.070 1324.700 20.390 ;
        RECT 1626.200 20.070 1626.460 20.390 ;
        RECT 1626.260 2.400 1626.400 20.070 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1338.210 204.580 1338.530 204.640 ;
        RECT 1642.730 204.580 1643.050 204.640 ;
        RECT 1338.210 204.440 1643.050 204.580 ;
        RECT 1338.210 204.380 1338.530 204.440 ;
        RECT 1642.730 204.380 1643.050 204.440 ;
      LAYER via ;
        RECT 1338.240 204.380 1338.500 204.640 ;
        RECT 1642.760 204.380 1643.020 204.640 ;
      LAYER met2 ;
        RECT 1337.270 216.650 1337.550 220.000 ;
        RECT 1337.270 216.510 1338.440 216.650 ;
        RECT 1337.270 216.000 1337.550 216.510 ;
        RECT 1338.300 204.670 1338.440 216.510 ;
        RECT 1338.240 204.350 1338.500 204.670 ;
        RECT 1642.760 204.350 1643.020 204.670 ;
        RECT 1642.820 16.730 1642.960 204.350 ;
        RECT 1642.820 16.590 1644.340 16.730 ;
        RECT 1644.200 2.400 1644.340 16.590 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1355.230 200.500 1355.550 200.560 ;
        RECT 1362.590 200.500 1362.910 200.560 ;
        RECT 1355.230 200.360 1362.910 200.500 ;
        RECT 1355.230 200.300 1355.550 200.360 ;
        RECT 1362.590 200.300 1362.910 200.360 ;
        RECT 1362.590 141.680 1362.910 141.740 ;
        RECT 1656.530 141.680 1656.850 141.740 ;
        RECT 1362.590 141.540 1656.850 141.680 ;
        RECT 1362.590 141.480 1362.910 141.540 ;
        RECT 1656.530 141.480 1656.850 141.540 ;
      LAYER via ;
        RECT 1355.260 200.300 1355.520 200.560 ;
        RECT 1362.620 200.300 1362.880 200.560 ;
        RECT 1362.620 141.480 1362.880 141.740 ;
        RECT 1656.560 141.480 1656.820 141.740 ;
      LAYER met2 ;
        RECT 1355.210 216.000 1355.490 220.000 ;
        RECT 1355.320 200.590 1355.460 216.000 ;
        RECT 1355.260 200.270 1355.520 200.590 ;
        RECT 1362.620 200.270 1362.880 200.590 ;
        RECT 1362.680 141.770 1362.820 200.270 ;
        RECT 1362.620 141.450 1362.880 141.770 ;
        RECT 1656.560 141.450 1656.820 141.770 ;
        RECT 1656.620 16.730 1656.760 141.450 ;
        RECT 1656.620 16.590 1662.280 16.730 ;
        RECT 1662.140 2.400 1662.280 16.590 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1373.170 200.500 1373.490 200.560 ;
        RECT 1379.150 200.500 1379.470 200.560 ;
        RECT 1373.170 200.360 1379.470 200.500 ;
        RECT 1373.170 200.300 1373.490 200.360 ;
        RECT 1379.150 200.300 1379.470 200.360 ;
        RECT 1379.150 134.880 1379.470 134.940 ;
        RECT 1676.770 134.880 1677.090 134.940 ;
        RECT 1379.150 134.740 1677.090 134.880 ;
        RECT 1379.150 134.680 1379.470 134.740 ;
        RECT 1676.770 134.680 1677.090 134.740 ;
      LAYER via ;
        RECT 1373.200 200.300 1373.460 200.560 ;
        RECT 1379.180 200.300 1379.440 200.560 ;
        RECT 1379.180 134.680 1379.440 134.940 ;
        RECT 1676.800 134.680 1677.060 134.940 ;
      LAYER met2 ;
        RECT 1373.150 216.000 1373.430 220.000 ;
        RECT 1373.260 200.590 1373.400 216.000 ;
        RECT 1373.200 200.270 1373.460 200.590 ;
        RECT 1379.180 200.270 1379.440 200.590 ;
        RECT 1379.240 134.970 1379.380 200.270 ;
        RECT 1379.180 134.650 1379.440 134.970 ;
        RECT 1676.800 134.650 1677.060 134.970 ;
        RECT 1676.860 17.410 1677.000 134.650 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1393.410 114.140 1393.730 114.200 ;
        RECT 1697.470 114.140 1697.790 114.200 ;
        RECT 1393.410 114.000 1697.790 114.140 ;
        RECT 1393.410 113.940 1393.730 114.000 ;
        RECT 1697.470 113.940 1697.790 114.000 ;
      LAYER via ;
        RECT 1393.440 113.940 1393.700 114.200 ;
        RECT 1697.500 113.940 1697.760 114.200 ;
      LAYER met2 ;
        RECT 1391.090 216.650 1391.370 220.000 ;
        RECT 1391.090 216.510 1393.640 216.650 ;
        RECT 1391.090 216.000 1391.370 216.510 ;
        RECT 1393.500 114.230 1393.640 216.510 ;
        RECT 1393.440 113.910 1393.700 114.230 ;
        RECT 1697.500 113.910 1697.760 114.230 ;
        RECT 1697.560 2.400 1697.700 113.910 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.010 216.650 426.290 220.000 ;
        RECT 426.010 216.510 427.640 216.650 ;
        RECT 426.010 216.000 426.290 216.510 ;
        RECT 427.500 16.845 427.640 216.510 ;
        RECT 427.430 16.475 427.710 16.845 ;
        RECT 734.250 16.475 734.530 16.845 ;
        RECT 734.320 2.400 734.460 16.475 ;
        RECT 734.110 -4.800 734.670 2.400 ;
      LAYER via2 ;
        RECT 427.430 16.520 427.710 16.800 ;
        RECT 734.250 16.520 734.530 16.800 ;
      LAYER met3 ;
        RECT 427.405 16.810 427.735 16.825 ;
        RECT 734.225 16.810 734.555 16.825 ;
        RECT 427.405 16.510 734.555 16.810 ;
        RECT 427.405 16.495 427.735 16.510 ;
        RECT 734.225 16.495 734.555 16.510 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.050 200.500 1409.370 200.560 ;
        RECT 1414.110 200.500 1414.430 200.560 ;
        RECT 1409.050 200.360 1414.430 200.500 ;
        RECT 1409.050 200.300 1409.370 200.360 ;
        RECT 1414.110 200.300 1414.430 200.360 ;
        RECT 1414.110 31.180 1414.430 31.240 ;
        RECT 1715.410 31.180 1715.730 31.240 ;
        RECT 1414.110 31.040 1715.730 31.180 ;
        RECT 1414.110 30.980 1414.430 31.040 ;
        RECT 1715.410 30.980 1715.730 31.040 ;
      LAYER via ;
        RECT 1409.080 200.300 1409.340 200.560 ;
        RECT 1414.140 200.300 1414.400 200.560 ;
        RECT 1414.140 30.980 1414.400 31.240 ;
        RECT 1715.440 30.980 1715.700 31.240 ;
      LAYER met2 ;
        RECT 1409.030 216.000 1409.310 220.000 ;
        RECT 1409.140 200.590 1409.280 216.000 ;
        RECT 1409.080 200.270 1409.340 200.590 ;
        RECT 1414.140 200.270 1414.400 200.590 ;
        RECT 1414.200 31.270 1414.340 200.270 ;
        RECT 1414.140 30.950 1414.400 31.270 ;
        RECT 1715.440 30.950 1715.700 31.270 ;
        RECT 1715.500 2.400 1715.640 30.950 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.910 120.940 1428.230 121.000 ;
        RECT 1731.970 120.940 1732.290 121.000 ;
        RECT 1427.910 120.800 1732.290 120.940 ;
        RECT 1427.910 120.740 1428.230 120.800 ;
        RECT 1731.970 120.740 1732.290 120.800 ;
      LAYER via ;
        RECT 1427.940 120.740 1428.200 121.000 ;
        RECT 1732.000 120.740 1732.260 121.000 ;
      LAYER met2 ;
        RECT 1426.970 216.650 1427.250 220.000 ;
        RECT 1426.970 216.510 1428.140 216.650 ;
        RECT 1426.970 216.000 1427.250 216.510 ;
        RECT 1428.000 121.030 1428.140 216.510 ;
        RECT 1427.940 120.710 1428.200 121.030 ;
        RECT 1732.000 120.710 1732.260 121.030 ;
        RECT 1732.060 17.410 1732.200 120.710 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.610 18.940 1448.930 19.000 ;
        RECT 1751.290 18.940 1751.610 19.000 ;
        RECT 1448.610 18.800 1751.610 18.940 ;
        RECT 1448.610 18.740 1448.930 18.800 ;
        RECT 1751.290 18.740 1751.610 18.800 ;
      LAYER via ;
        RECT 1448.640 18.740 1448.900 19.000 ;
        RECT 1751.320 18.740 1751.580 19.000 ;
      LAYER met2 ;
        RECT 1444.910 216.650 1445.190 220.000 ;
        RECT 1444.910 216.510 1448.840 216.650 ;
        RECT 1444.910 216.000 1445.190 216.510 ;
        RECT 1448.700 19.030 1448.840 216.510 ;
        RECT 1448.640 18.710 1448.900 19.030 ;
        RECT 1751.320 18.710 1751.580 19.030 ;
        RECT 1751.380 2.400 1751.520 18.710 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.870 200.500 1463.190 200.560 ;
        RECT 1469.310 200.500 1469.630 200.560 ;
        RECT 1462.870 200.360 1469.630 200.500 ;
        RECT 1462.870 200.300 1463.190 200.360 ;
        RECT 1469.310 200.300 1469.630 200.360 ;
        RECT 1469.310 19.280 1469.630 19.340 ;
        RECT 1768.770 19.280 1769.090 19.340 ;
        RECT 1469.310 19.140 1769.090 19.280 ;
        RECT 1469.310 19.080 1469.630 19.140 ;
        RECT 1768.770 19.080 1769.090 19.140 ;
      LAYER via ;
        RECT 1462.900 200.300 1463.160 200.560 ;
        RECT 1469.340 200.300 1469.600 200.560 ;
        RECT 1469.340 19.080 1469.600 19.340 ;
        RECT 1768.800 19.080 1769.060 19.340 ;
      LAYER met2 ;
        RECT 1462.850 216.000 1463.130 220.000 ;
        RECT 1462.960 200.590 1463.100 216.000 ;
        RECT 1462.900 200.270 1463.160 200.590 ;
        RECT 1469.340 200.270 1469.600 200.590 ;
        RECT 1469.400 19.370 1469.540 200.270 ;
        RECT 1469.340 19.050 1469.600 19.370 ;
        RECT 1768.800 19.050 1769.060 19.370 ;
        RECT 1768.860 2.400 1769.000 19.050 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.110 19.620 1483.430 19.680 ;
        RECT 1786.710 19.620 1787.030 19.680 ;
        RECT 1483.110 19.480 1787.030 19.620 ;
        RECT 1483.110 19.420 1483.430 19.480 ;
        RECT 1786.710 19.420 1787.030 19.480 ;
      LAYER via ;
        RECT 1483.140 19.420 1483.400 19.680 ;
        RECT 1786.740 19.420 1787.000 19.680 ;
      LAYER met2 ;
        RECT 1480.330 216.650 1480.610 220.000 ;
        RECT 1480.330 216.510 1483.340 216.650 ;
        RECT 1480.330 216.000 1480.610 216.510 ;
        RECT 1483.200 19.710 1483.340 216.510 ;
        RECT 1483.140 19.390 1483.400 19.710 ;
        RECT 1786.740 19.390 1787.000 19.710 ;
        RECT 1786.800 2.400 1786.940 19.390 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1498.290 202.880 1498.610 202.940 ;
        RECT 1503.810 202.880 1504.130 202.940 ;
        RECT 1498.290 202.740 1504.130 202.880 ;
        RECT 1498.290 202.680 1498.610 202.740 ;
        RECT 1503.810 202.680 1504.130 202.740 ;
        RECT 1503.810 19.960 1504.130 20.020 ;
        RECT 1804.650 19.960 1804.970 20.020 ;
        RECT 1503.810 19.820 1804.970 19.960 ;
        RECT 1503.810 19.760 1504.130 19.820 ;
        RECT 1804.650 19.760 1804.970 19.820 ;
      LAYER via ;
        RECT 1498.320 202.680 1498.580 202.940 ;
        RECT 1503.840 202.680 1504.100 202.940 ;
        RECT 1503.840 19.760 1504.100 20.020 ;
        RECT 1804.680 19.760 1804.940 20.020 ;
      LAYER met2 ;
        RECT 1498.270 216.000 1498.550 220.000 ;
        RECT 1498.380 202.970 1498.520 216.000 ;
        RECT 1498.320 202.650 1498.580 202.970 ;
        RECT 1503.840 202.650 1504.100 202.970 ;
        RECT 1503.900 20.050 1504.040 202.650 ;
        RECT 1503.840 19.730 1504.100 20.050 ;
        RECT 1804.680 19.730 1804.940 20.050 ;
        RECT 1804.740 2.400 1804.880 19.730 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.610 24.380 1517.930 24.440 ;
        RECT 1822.590 24.380 1822.910 24.440 ;
        RECT 1517.610 24.240 1822.910 24.380 ;
        RECT 1517.610 24.180 1517.930 24.240 ;
        RECT 1822.590 24.180 1822.910 24.240 ;
      LAYER via ;
        RECT 1517.640 24.180 1517.900 24.440 ;
        RECT 1822.620 24.180 1822.880 24.440 ;
      LAYER met2 ;
        RECT 1516.210 216.650 1516.490 220.000 ;
        RECT 1516.210 216.510 1517.840 216.650 ;
        RECT 1516.210 216.000 1516.490 216.510 ;
        RECT 1517.700 24.470 1517.840 216.510 ;
        RECT 1517.640 24.150 1517.900 24.470 ;
        RECT 1822.620 24.150 1822.880 24.470 ;
        RECT 1822.680 2.400 1822.820 24.150 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1534.170 200.500 1534.490 200.560 ;
        RECT 1538.310 200.500 1538.630 200.560 ;
        RECT 1534.170 200.360 1538.630 200.500 ;
        RECT 1534.170 200.300 1534.490 200.360 ;
        RECT 1538.310 200.300 1538.630 200.360 ;
        RECT 1538.310 18.600 1538.630 18.660 ;
        RECT 1840.070 18.600 1840.390 18.660 ;
        RECT 1538.310 18.460 1840.390 18.600 ;
        RECT 1538.310 18.400 1538.630 18.460 ;
        RECT 1840.070 18.400 1840.390 18.460 ;
      LAYER via ;
        RECT 1534.200 200.300 1534.460 200.560 ;
        RECT 1538.340 200.300 1538.600 200.560 ;
        RECT 1538.340 18.400 1538.600 18.660 ;
        RECT 1840.100 18.400 1840.360 18.660 ;
      LAYER met2 ;
        RECT 1534.150 216.000 1534.430 220.000 ;
        RECT 1534.260 200.590 1534.400 216.000 ;
        RECT 1534.200 200.270 1534.460 200.590 ;
        RECT 1538.340 200.270 1538.600 200.590 ;
        RECT 1538.400 18.690 1538.540 200.270 ;
        RECT 1538.340 18.370 1538.600 18.690 ;
        RECT 1840.100 18.370 1840.360 18.690 ;
        RECT 1840.160 2.400 1840.300 18.370 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1828.185 14.705 1828.355 17.595 ;
      LAYER mcon ;
        RECT 1828.185 17.425 1828.355 17.595 ;
      LAYER met1 ;
        RECT 1552.110 18.260 1552.430 18.320 ;
        RECT 1552.110 18.120 1573.500 18.260 ;
        RECT 1552.110 18.060 1552.430 18.120 ;
        RECT 1573.360 17.580 1573.500 18.120 ;
        RECT 1828.125 17.580 1828.415 17.625 ;
        RECT 1573.360 17.440 1828.415 17.580 ;
        RECT 1828.125 17.395 1828.415 17.440 ;
        RECT 1828.125 14.860 1828.415 14.905 ;
        RECT 1858.010 14.860 1858.330 14.920 ;
        RECT 1828.125 14.720 1858.330 14.860 ;
        RECT 1828.125 14.675 1828.415 14.720 ;
        RECT 1858.010 14.660 1858.330 14.720 ;
      LAYER via ;
        RECT 1552.140 18.060 1552.400 18.320 ;
        RECT 1858.040 14.660 1858.300 14.920 ;
      LAYER met2 ;
        RECT 1552.090 216.000 1552.370 220.000 ;
        RECT 1552.200 18.350 1552.340 216.000 ;
        RECT 1552.140 18.030 1552.400 18.350 ;
        RECT 1858.040 14.630 1858.300 14.950 ;
        RECT 1858.100 2.400 1858.240 14.630 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 17.720 1573.130 17.980 ;
        RECT 1572.900 16.900 1573.040 17.720 ;
        RECT 1875.950 16.900 1876.270 16.960 ;
        RECT 1572.900 16.760 1876.270 16.900 ;
        RECT 1875.950 16.700 1876.270 16.760 ;
      LAYER via ;
        RECT 1572.840 17.720 1573.100 17.980 ;
        RECT 1875.980 16.700 1876.240 16.960 ;
      LAYER met2 ;
        RECT 1570.030 216.650 1570.310 220.000 ;
        RECT 1570.030 216.510 1573.040 216.650 ;
        RECT 1570.030 216.000 1570.310 216.510 ;
        RECT 1572.900 18.010 1573.040 216.510 ;
        RECT 1572.840 17.690 1573.100 18.010 ;
        RECT 1875.980 16.670 1876.240 16.990 ;
        RECT 1876.040 2.400 1876.180 16.670 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 482.685 204.765 482.855 205.615 ;
        RECT 496.945 204.765 497.115 206.295 ;
        RECT 530.985 205.105 531.155 206.295 ;
        RECT 724.185 202.045 724.355 204.935 ;
        RECT 724.645 198.305 724.815 202.215 ;
      LAYER mcon ;
        RECT 496.945 206.125 497.115 206.295 ;
        RECT 482.685 205.445 482.855 205.615 ;
        RECT 530.985 206.125 531.155 206.295 ;
        RECT 724.185 204.765 724.355 204.935 ;
        RECT 724.645 202.045 724.815 202.215 ;
      LAYER met1 ;
        RECT 496.885 206.280 497.175 206.325 ;
        RECT 530.925 206.280 531.215 206.325 ;
        RECT 496.885 206.140 531.215 206.280 ;
        RECT 496.885 206.095 497.175 206.140 ;
        RECT 530.925 206.095 531.215 206.140 ;
        RECT 443.510 205.600 443.830 205.660 ;
        RECT 482.625 205.600 482.915 205.645 ;
        RECT 443.510 205.460 482.915 205.600 ;
        RECT 443.510 205.400 443.830 205.460 ;
        RECT 482.625 205.415 482.915 205.460 ;
        RECT 530.925 205.260 531.215 205.305 ;
        RECT 530.925 205.120 545.400 205.260 ;
        RECT 530.925 205.075 531.215 205.120 ;
        RECT 482.625 204.920 482.915 204.965 ;
        RECT 496.885 204.920 497.175 204.965 ;
        RECT 482.625 204.780 497.175 204.920 ;
        RECT 545.260 204.920 545.400 205.120 ;
        RECT 724.125 204.920 724.415 204.965 ;
        RECT 545.260 204.780 724.415 204.920 ;
        RECT 482.625 204.735 482.915 204.780 ;
        RECT 496.885 204.735 497.175 204.780 ;
        RECT 724.125 204.735 724.415 204.780 ;
        RECT 724.200 202.400 724.800 202.540 ;
        RECT 724.200 202.245 724.340 202.400 ;
        RECT 724.660 202.245 724.800 202.400 ;
        RECT 724.125 202.015 724.415 202.245 ;
        RECT 724.585 202.015 724.875 202.245 ;
        RECT 724.585 198.460 724.875 198.505 ;
        RECT 753.090 198.460 753.410 198.520 ;
        RECT 724.585 198.320 753.410 198.460 ;
        RECT 724.585 198.275 724.875 198.320 ;
        RECT 753.090 198.260 753.410 198.320 ;
      LAYER via ;
        RECT 443.540 205.400 443.800 205.660 ;
        RECT 753.120 198.260 753.380 198.520 ;
      LAYER met2 ;
        RECT 443.490 216.000 443.770 220.000 ;
        RECT 443.600 205.690 443.740 216.000 ;
        RECT 443.540 205.370 443.800 205.690 ;
        RECT 753.120 198.230 753.380 198.550 ;
        RECT 753.180 17.410 753.320 198.230 ;
        RECT 752.260 17.270 753.320 17.410 ;
        RECT 752.260 2.400 752.400 17.270 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.990 200.500 1588.310 200.560 ;
        RECT 1593.510 200.500 1593.830 200.560 ;
        RECT 1587.990 200.360 1593.830 200.500 ;
        RECT 1587.990 200.300 1588.310 200.360 ;
        RECT 1593.510 200.300 1593.830 200.360 ;
        RECT 1593.510 16.220 1593.830 16.280 ;
        RECT 1893.890 16.220 1894.210 16.280 ;
        RECT 1593.510 16.080 1894.210 16.220 ;
        RECT 1593.510 16.020 1593.830 16.080 ;
        RECT 1893.890 16.020 1894.210 16.080 ;
      LAYER via ;
        RECT 1588.020 200.300 1588.280 200.560 ;
        RECT 1593.540 200.300 1593.800 200.560 ;
        RECT 1593.540 16.020 1593.800 16.280 ;
        RECT 1893.920 16.020 1894.180 16.280 ;
      LAYER met2 ;
        RECT 1587.970 216.000 1588.250 220.000 ;
        RECT 1588.080 200.590 1588.220 216.000 ;
        RECT 1588.020 200.270 1588.280 200.590 ;
        RECT 1593.540 200.270 1593.800 200.590 ;
        RECT 1593.600 16.310 1593.740 200.270 ;
        RECT 1593.540 15.990 1593.800 16.310 ;
        RECT 1893.920 15.990 1894.180 16.310 ;
        RECT 1893.980 2.400 1894.120 15.990 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1607.310 18.260 1607.630 18.320 ;
        RECT 1911.370 18.260 1911.690 18.320 ;
        RECT 1607.310 18.120 1911.690 18.260 ;
        RECT 1607.310 18.060 1607.630 18.120 ;
        RECT 1911.370 18.060 1911.690 18.120 ;
      LAYER via ;
        RECT 1607.340 18.060 1607.600 18.320 ;
        RECT 1911.400 18.060 1911.660 18.320 ;
      LAYER met2 ;
        RECT 1605.450 216.650 1605.730 220.000 ;
        RECT 1605.450 216.510 1607.540 216.650 ;
        RECT 1605.450 216.000 1605.730 216.510 ;
        RECT 1607.400 18.350 1607.540 216.510 ;
        RECT 1607.340 18.030 1607.600 18.350 ;
        RECT 1911.400 18.030 1911.660 18.350 ;
        RECT 1911.460 16.730 1911.600 18.030 ;
        RECT 1911.460 16.590 1912.060 16.730 ;
        RECT 1911.920 2.400 1912.060 16.590 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1623.410 200.500 1623.730 200.560 ;
        RECT 1628.010 200.500 1628.330 200.560 ;
        RECT 1623.410 200.360 1628.330 200.500 ;
        RECT 1623.410 200.300 1623.730 200.360 ;
        RECT 1628.010 200.300 1628.330 200.360 ;
        RECT 1628.010 20.300 1628.330 20.360 ;
        RECT 1929.310 20.300 1929.630 20.360 ;
        RECT 1628.010 20.160 1929.630 20.300 ;
        RECT 1628.010 20.100 1628.330 20.160 ;
        RECT 1929.310 20.100 1929.630 20.160 ;
      LAYER via ;
        RECT 1623.440 200.300 1623.700 200.560 ;
        RECT 1628.040 200.300 1628.300 200.560 ;
        RECT 1628.040 20.100 1628.300 20.360 ;
        RECT 1929.340 20.100 1929.600 20.360 ;
      LAYER met2 ;
        RECT 1623.390 216.000 1623.670 220.000 ;
        RECT 1623.500 200.590 1623.640 216.000 ;
        RECT 1623.440 200.270 1623.700 200.590 ;
        RECT 1628.040 200.270 1628.300 200.590 ;
        RECT 1628.100 20.390 1628.240 200.270 ;
        RECT 1628.040 20.070 1628.300 20.390 ;
        RECT 1929.340 20.070 1929.600 20.390 ;
        RECT 1929.400 2.400 1929.540 20.070 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1641.810 17.920 1642.130 17.980 ;
        RECT 1947.250 17.920 1947.570 17.980 ;
        RECT 1641.810 17.780 1947.570 17.920 ;
        RECT 1641.810 17.720 1642.130 17.780 ;
        RECT 1947.250 17.720 1947.570 17.780 ;
      LAYER via ;
        RECT 1641.840 17.720 1642.100 17.980 ;
        RECT 1947.280 17.720 1947.540 17.980 ;
      LAYER met2 ;
        RECT 1641.330 216.650 1641.610 220.000 ;
        RECT 1641.330 216.510 1642.040 216.650 ;
        RECT 1641.330 216.000 1641.610 216.510 ;
        RECT 1641.900 18.010 1642.040 216.510 ;
        RECT 1641.840 17.690 1642.100 18.010 ;
        RECT 1947.280 17.690 1947.540 18.010 ;
        RECT 1947.340 2.400 1947.480 17.690 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.510 15.200 1662.830 15.260 ;
        RECT 1965.190 15.200 1965.510 15.260 ;
        RECT 1662.510 15.060 1965.510 15.200 ;
        RECT 1662.510 15.000 1662.830 15.060 ;
        RECT 1965.190 15.000 1965.510 15.060 ;
      LAYER via ;
        RECT 1662.540 15.000 1662.800 15.260 ;
        RECT 1965.220 15.000 1965.480 15.260 ;
      LAYER met2 ;
        RECT 1659.270 216.650 1659.550 220.000 ;
        RECT 1659.270 216.510 1662.740 216.650 ;
        RECT 1659.270 216.000 1659.550 216.510 ;
        RECT 1662.600 15.290 1662.740 216.510 ;
        RECT 1662.540 14.970 1662.800 15.290 ;
        RECT 1965.220 14.970 1965.480 15.290 ;
        RECT 1965.280 2.400 1965.420 14.970 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1677.230 200.500 1677.550 200.560 ;
        RECT 1683.210 200.500 1683.530 200.560 ;
        RECT 1677.230 200.360 1683.530 200.500 ;
        RECT 1677.230 200.300 1677.550 200.360 ;
        RECT 1683.210 200.300 1683.530 200.360 ;
        RECT 1683.210 15.540 1683.530 15.600 ;
        RECT 1983.130 15.540 1983.450 15.600 ;
        RECT 1683.210 15.400 1983.450 15.540 ;
        RECT 1683.210 15.340 1683.530 15.400 ;
        RECT 1983.130 15.340 1983.450 15.400 ;
      LAYER via ;
        RECT 1677.260 200.300 1677.520 200.560 ;
        RECT 1683.240 200.300 1683.500 200.560 ;
        RECT 1683.240 15.340 1683.500 15.600 ;
        RECT 1983.160 15.340 1983.420 15.600 ;
      LAYER met2 ;
        RECT 1677.210 216.000 1677.490 220.000 ;
        RECT 1677.320 200.590 1677.460 216.000 ;
        RECT 1677.260 200.270 1677.520 200.590 ;
        RECT 1683.240 200.270 1683.500 200.590 ;
        RECT 1683.300 15.630 1683.440 200.270 ;
        RECT 1683.240 15.310 1683.500 15.630 ;
        RECT 1983.160 15.310 1983.420 15.630 ;
        RECT 1983.220 2.400 1983.360 15.310 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1695.150 216.650 1695.430 220.000 ;
        RECT 1695.150 216.510 1697.240 216.650 ;
        RECT 1695.150 216.000 1695.430 216.510 ;
        RECT 1697.100 16.845 1697.240 216.510 ;
        RECT 1697.030 16.475 1697.310 16.845 ;
        RECT 2001.090 16.475 2001.370 16.845 ;
        RECT 2001.160 2.400 2001.300 16.475 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
      LAYER via2 ;
        RECT 1697.030 16.520 1697.310 16.800 ;
        RECT 2001.090 16.520 2001.370 16.800 ;
      LAYER met3 ;
        RECT 1697.005 16.810 1697.335 16.825 ;
        RECT 2001.065 16.810 2001.395 16.825 ;
        RECT 1697.005 16.510 2001.395 16.810 ;
        RECT 1697.005 16.495 1697.335 16.510 ;
        RECT 2001.065 16.495 2001.395 16.510 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1713.110 200.500 1713.430 200.560 ;
        RECT 1717.710 200.500 1718.030 200.560 ;
        RECT 1713.110 200.360 1718.030 200.500 ;
        RECT 1713.110 200.300 1713.430 200.360 ;
        RECT 1717.710 200.300 1718.030 200.360 ;
        RECT 1717.710 15.880 1718.030 15.940 ;
        RECT 2018.550 15.880 2018.870 15.940 ;
        RECT 1717.710 15.740 2018.870 15.880 ;
        RECT 1717.710 15.680 1718.030 15.740 ;
        RECT 2018.550 15.680 2018.870 15.740 ;
      LAYER via ;
        RECT 1713.140 200.300 1713.400 200.560 ;
        RECT 1717.740 200.300 1718.000 200.560 ;
        RECT 1717.740 15.680 1718.000 15.940 ;
        RECT 2018.580 15.680 2018.840 15.940 ;
      LAYER met2 ;
        RECT 1713.090 216.000 1713.370 220.000 ;
        RECT 1713.200 200.590 1713.340 216.000 ;
        RECT 1713.140 200.270 1713.400 200.590 ;
        RECT 1717.740 200.270 1718.000 200.590 ;
        RECT 1717.800 15.970 1717.940 200.270 ;
        RECT 1717.740 15.650 1718.000 15.970 ;
        RECT 2018.580 15.650 2018.840 15.970 ;
        RECT 2018.640 2.400 2018.780 15.650 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2036.105 89.845 2036.275 137.955 ;
      LAYER mcon ;
        RECT 2036.105 137.785 2036.275 137.955 ;
      LAYER met1 ;
        RECT 1730.590 203.560 1730.910 203.620 ;
        RECT 2036.030 203.560 2036.350 203.620 ;
        RECT 1730.590 203.420 2036.350 203.560 ;
        RECT 1730.590 203.360 1730.910 203.420 ;
        RECT 2036.030 203.360 2036.350 203.420 ;
        RECT 2036.030 137.940 2036.350 138.000 ;
        RECT 2035.835 137.800 2036.350 137.940 ;
        RECT 2036.030 137.740 2036.350 137.800 ;
        RECT 2036.030 90.000 2036.350 90.060 ;
        RECT 2035.835 89.860 2036.350 90.000 ;
        RECT 2036.030 89.800 2036.350 89.860 ;
        RECT 2036.030 62.260 2036.350 62.520 ;
        RECT 2036.120 61.780 2036.260 62.260 ;
        RECT 2036.490 61.780 2036.810 61.840 ;
        RECT 2036.120 61.640 2036.810 61.780 ;
        RECT 2036.490 61.580 2036.810 61.640 ;
      LAYER via ;
        RECT 1730.620 203.360 1730.880 203.620 ;
        RECT 2036.060 203.360 2036.320 203.620 ;
        RECT 2036.060 137.740 2036.320 138.000 ;
        RECT 2036.060 89.800 2036.320 90.060 ;
        RECT 2036.060 62.260 2036.320 62.520 ;
        RECT 2036.520 61.580 2036.780 61.840 ;
      LAYER met2 ;
        RECT 1730.570 216.000 1730.850 220.000 ;
        RECT 1730.680 203.650 1730.820 216.000 ;
        RECT 1730.620 203.330 1730.880 203.650 ;
        RECT 2036.060 203.330 2036.320 203.650 ;
        RECT 2036.120 146.045 2036.260 203.330 ;
        RECT 2036.050 145.675 2036.330 146.045 ;
        RECT 2036.050 144.995 2036.330 145.365 ;
        RECT 2036.120 138.030 2036.260 144.995 ;
        RECT 2036.060 137.710 2036.320 138.030 ;
        RECT 2036.060 89.770 2036.320 90.090 ;
        RECT 2036.120 62.550 2036.260 89.770 ;
        RECT 2036.060 62.230 2036.320 62.550 ;
        RECT 2036.520 61.550 2036.780 61.870 ;
        RECT 2036.580 2.400 2036.720 61.550 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
      LAYER via2 ;
        RECT 2036.050 145.720 2036.330 146.000 ;
        RECT 2036.050 145.040 2036.330 145.320 ;
      LAYER met3 ;
        RECT 2036.025 146.010 2036.355 146.025 ;
        RECT 2035.350 145.710 2036.355 146.010 ;
        RECT 2035.350 145.330 2035.650 145.710 ;
        RECT 2036.025 145.695 2036.355 145.710 ;
        RECT 2036.025 145.330 2036.355 145.345 ;
        RECT 2035.350 145.030 2036.355 145.330 ;
        RECT 2036.025 145.015 2036.355 145.030 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1752.210 20.640 1752.530 20.700 ;
        RECT 2054.430 20.640 2054.750 20.700 ;
        RECT 1752.210 20.500 2054.750 20.640 ;
        RECT 1752.210 20.440 1752.530 20.500 ;
        RECT 2054.430 20.440 2054.750 20.500 ;
      LAYER via ;
        RECT 1752.240 20.440 1752.500 20.700 ;
        RECT 2054.460 20.440 2054.720 20.700 ;
      LAYER met2 ;
        RECT 1748.510 216.650 1748.790 220.000 ;
        RECT 1748.510 216.510 1752.440 216.650 ;
        RECT 1748.510 216.000 1748.790 216.510 ;
        RECT 1752.300 20.730 1752.440 216.510 ;
        RECT 1752.240 20.410 1752.500 20.730 ;
        RECT 2054.460 20.410 2054.720 20.730 ;
        RECT 2054.520 2.400 2054.660 20.410 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.430 216.650 461.710 220.000 ;
        RECT 461.430 216.510 462.140 216.650 ;
        RECT 461.430 216.000 461.710 216.510 ;
        RECT 462.000 17.525 462.140 216.510 ;
        RECT 461.930 17.155 462.210 17.525 ;
        RECT 769.670 17.155 769.950 17.525 ;
        RECT 769.740 2.400 769.880 17.155 ;
        RECT 769.530 -4.800 770.090 2.400 ;
      LAYER via2 ;
        RECT 461.930 17.200 462.210 17.480 ;
        RECT 769.670 17.200 769.950 17.480 ;
      LAYER met3 ;
        RECT 461.905 17.490 462.235 17.505 ;
        RECT 769.645 17.490 769.975 17.505 ;
        RECT 461.905 17.190 769.975 17.490 ;
        RECT 461.905 17.175 462.235 17.190 ;
        RECT 769.645 17.175 769.975 17.190 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.470 200.500 1766.790 200.560 ;
        RECT 1772.910 200.500 1773.230 200.560 ;
        RECT 1766.470 200.360 1773.230 200.500 ;
        RECT 1766.470 200.300 1766.790 200.360 ;
        RECT 1772.910 200.300 1773.230 200.360 ;
        RECT 1772.910 18.940 1773.230 19.000 ;
        RECT 2072.370 18.940 2072.690 19.000 ;
        RECT 1772.910 18.800 2072.690 18.940 ;
        RECT 1772.910 18.740 1773.230 18.800 ;
        RECT 2072.370 18.740 2072.690 18.800 ;
      LAYER via ;
        RECT 1766.500 200.300 1766.760 200.560 ;
        RECT 1772.940 200.300 1773.200 200.560 ;
        RECT 1772.940 18.740 1773.200 19.000 ;
        RECT 2072.400 18.740 2072.660 19.000 ;
      LAYER met2 ;
        RECT 1766.450 216.000 1766.730 220.000 ;
        RECT 1766.560 200.590 1766.700 216.000 ;
        RECT 1766.500 200.270 1766.760 200.590 ;
        RECT 1772.940 200.270 1773.200 200.590 ;
        RECT 1773.000 19.030 1773.140 200.270 ;
        RECT 1772.940 18.710 1773.200 19.030 ;
        RECT 2072.400 18.710 2072.660 19.030 ;
        RECT 2072.460 2.400 2072.600 18.710 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1785.790 16.560 1786.110 16.620 ;
        RECT 2089.850 16.560 2090.170 16.620 ;
        RECT 1785.790 16.420 2090.170 16.560 ;
        RECT 1785.790 16.360 1786.110 16.420 ;
        RECT 2089.850 16.360 2090.170 16.420 ;
      LAYER via ;
        RECT 1785.820 16.360 1786.080 16.620 ;
        RECT 2089.880 16.360 2090.140 16.620 ;
      LAYER met2 ;
        RECT 1784.390 216.650 1784.670 220.000 ;
        RECT 1784.390 216.510 1786.940 216.650 ;
        RECT 1784.390 216.000 1784.670 216.510 ;
        RECT 1786.800 34.410 1786.940 216.510 ;
        RECT 1785.880 34.270 1786.940 34.410 ;
        RECT 1785.880 16.650 1786.020 34.270 ;
        RECT 1785.820 16.330 1786.080 16.650 ;
        RECT 2089.880 16.330 2090.140 16.650 ;
        RECT 2089.940 2.400 2090.080 16.330 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1802.350 200.500 1802.670 200.560 ;
        RECT 1807.410 200.500 1807.730 200.560 ;
        RECT 1802.350 200.360 1807.730 200.500 ;
        RECT 1802.350 200.300 1802.670 200.360 ;
        RECT 1807.410 200.300 1807.730 200.360 ;
        RECT 1807.410 19.280 1807.730 19.340 ;
        RECT 2107.790 19.280 2108.110 19.340 ;
        RECT 1807.410 19.140 2108.110 19.280 ;
        RECT 1807.410 19.080 1807.730 19.140 ;
        RECT 2107.790 19.080 2108.110 19.140 ;
      LAYER via ;
        RECT 1802.380 200.300 1802.640 200.560 ;
        RECT 1807.440 200.300 1807.700 200.560 ;
        RECT 1807.440 19.080 1807.700 19.340 ;
        RECT 2107.820 19.080 2108.080 19.340 ;
      LAYER met2 ;
        RECT 1802.330 216.000 1802.610 220.000 ;
        RECT 1802.440 200.590 1802.580 216.000 ;
        RECT 1802.380 200.270 1802.640 200.590 ;
        RECT 1807.440 200.270 1807.700 200.590 ;
        RECT 1807.500 19.370 1807.640 200.270 ;
        RECT 1807.440 19.050 1807.700 19.370 ;
        RECT 2107.820 19.050 2108.080 19.370 ;
        RECT 2107.880 2.400 2108.020 19.050 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1820.270 216.650 1820.550 220.000 ;
        RECT 1820.270 216.510 1821.440 216.650 ;
        RECT 1820.270 216.000 1820.550 216.510 ;
        RECT 1821.300 17.525 1821.440 216.510 ;
        RECT 1821.230 17.155 1821.510 17.525 ;
        RECT 2125.750 17.155 2126.030 17.525 ;
        RECT 2125.820 2.400 2125.960 17.155 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
      LAYER via2 ;
        RECT 1821.230 17.200 1821.510 17.480 ;
        RECT 2125.750 17.200 2126.030 17.480 ;
      LAYER met3 ;
        RECT 1821.205 17.490 1821.535 17.505 ;
        RECT 2125.725 17.490 2126.055 17.505 ;
        RECT 1821.205 17.190 2126.055 17.490 ;
        RECT 1821.205 17.175 1821.535 17.190 ;
        RECT 2125.725 17.175 2126.055 17.190 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2143.745 2.805 2143.915 14.195 ;
      LAYER mcon ;
        RECT 2143.745 14.025 2143.915 14.195 ;
      LAYER met1 ;
        RECT 1838.230 204.580 1838.550 204.640 ;
        RECT 2139.530 204.580 2139.850 204.640 ;
        RECT 1838.230 204.440 2139.850 204.580 ;
        RECT 1838.230 204.380 1838.550 204.440 ;
        RECT 2139.530 204.380 2139.850 204.440 ;
        RECT 2139.530 14.180 2139.850 14.240 ;
        RECT 2143.685 14.180 2143.975 14.225 ;
        RECT 2139.530 14.040 2143.975 14.180 ;
        RECT 2139.530 13.980 2139.850 14.040 ;
        RECT 2143.685 13.995 2143.975 14.040 ;
        RECT 2143.670 2.960 2143.990 3.020 ;
        RECT 2143.475 2.820 2143.990 2.960 ;
        RECT 2143.670 2.760 2143.990 2.820 ;
      LAYER via ;
        RECT 1838.260 204.380 1838.520 204.640 ;
        RECT 2139.560 204.380 2139.820 204.640 ;
        RECT 2139.560 13.980 2139.820 14.240 ;
        RECT 2143.700 2.760 2143.960 3.020 ;
      LAYER met2 ;
        RECT 1838.210 216.000 1838.490 220.000 ;
        RECT 1838.320 204.670 1838.460 216.000 ;
        RECT 1838.260 204.350 1838.520 204.670 ;
        RECT 2139.560 204.350 2139.820 204.670 ;
        RECT 2139.620 14.270 2139.760 204.350 ;
        RECT 2139.560 13.950 2139.820 14.270 ;
        RECT 2143.700 2.730 2143.960 3.050 ;
        RECT 2143.760 2.400 2143.900 2.730 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1855.710 17.240 1856.030 17.300 ;
        RECT 2161.610 17.240 2161.930 17.300 ;
        RECT 1855.710 17.100 2161.930 17.240 ;
        RECT 1855.710 17.040 1856.030 17.100 ;
        RECT 2161.610 17.040 2161.930 17.100 ;
      LAYER via ;
        RECT 1855.740 17.040 1856.000 17.300 ;
        RECT 2161.640 17.040 2161.900 17.300 ;
      LAYER met2 ;
        RECT 1855.690 216.000 1855.970 220.000 ;
        RECT 1855.800 17.330 1855.940 216.000 ;
        RECT 1855.740 17.010 1856.000 17.330 ;
        RECT 2161.640 17.010 2161.900 17.330 ;
        RECT 2161.700 2.400 2161.840 17.010 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2179.165 2.805 2179.335 14.195 ;
      LAYER mcon ;
        RECT 2179.165 14.025 2179.335 14.195 ;
      LAYER met1 ;
        RECT 1873.650 204.920 1873.970 204.980 ;
        RECT 2174.030 204.920 2174.350 204.980 ;
        RECT 1873.650 204.780 2174.350 204.920 ;
        RECT 1873.650 204.720 1873.970 204.780 ;
        RECT 2174.030 204.720 2174.350 204.780 ;
        RECT 2174.030 14.180 2174.350 14.240 ;
        RECT 2179.105 14.180 2179.395 14.225 ;
        RECT 2174.030 14.040 2179.395 14.180 ;
        RECT 2174.030 13.980 2174.350 14.040 ;
        RECT 2179.105 13.995 2179.395 14.040 ;
        RECT 2179.090 2.960 2179.410 3.020 ;
        RECT 2178.895 2.820 2179.410 2.960 ;
        RECT 2179.090 2.760 2179.410 2.820 ;
      LAYER via ;
        RECT 1873.680 204.720 1873.940 204.980 ;
        RECT 2174.060 204.720 2174.320 204.980 ;
        RECT 2174.060 13.980 2174.320 14.240 ;
        RECT 2179.120 2.760 2179.380 3.020 ;
      LAYER met2 ;
        RECT 1873.630 216.000 1873.910 220.000 ;
        RECT 1873.740 205.010 1873.880 216.000 ;
        RECT 1873.680 204.690 1873.940 205.010 ;
        RECT 2174.060 204.690 2174.320 205.010 ;
        RECT 2174.120 14.270 2174.260 204.690 ;
        RECT 2174.060 13.950 2174.320 14.270 ;
        RECT 2179.120 2.730 2179.380 3.050 ;
        RECT 2179.180 2.400 2179.320 2.730 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.590 200.500 1891.910 200.560 ;
        RECT 1897.110 200.500 1897.430 200.560 ;
        RECT 1891.590 200.360 1897.430 200.500 ;
        RECT 1891.590 200.300 1891.910 200.360 ;
        RECT 1897.110 200.300 1897.430 200.360 ;
        RECT 1897.110 19.960 1897.430 20.020 ;
        RECT 2197.030 19.960 2197.350 20.020 ;
        RECT 1897.110 19.820 2197.350 19.960 ;
        RECT 1897.110 19.760 1897.430 19.820 ;
        RECT 2197.030 19.760 2197.350 19.820 ;
      LAYER via ;
        RECT 1891.620 200.300 1891.880 200.560 ;
        RECT 1897.140 200.300 1897.400 200.560 ;
        RECT 1897.140 19.760 1897.400 20.020 ;
        RECT 2197.060 19.760 2197.320 20.020 ;
      LAYER met2 ;
        RECT 1891.570 216.000 1891.850 220.000 ;
        RECT 1891.680 200.590 1891.820 216.000 ;
        RECT 1891.620 200.270 1891.880 200.590 ;
        RECT 1897.140 200.270 1897.400 200.590 ;
        RECT 1897.200 20.050 1897.340 200.270 ;
        RECT 1897.140 19.730 1897.400 20.050 ;
        RECT 2197.060 19.730 2197.320 20.050 ;
        RECT 2197.120 2.400 2197.260 19.730 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2215.965 186.405 2216.135 203.915 ;
        RECT 2215.965 48.365 2216.135 137.955 ;
      LAYER mcon ;
        RECT 2215.965 203.745 2216.135 203.915 ;
        RECT 2215.965 137.785 2216.135 137.955 ;
      LAYER met1 ;
        RECT 1909.530 203.900 1909.850 203.960 ;
        RECT 2215.905 203.900 2216.195 203.945 ;
        RECT 1909.530 203.760 2216.195 203.900 ;
        RECT 1909.530 203.700 1909.850 203.760 ;
        RECT 2215.905 203.715 2216.195 203.760 ;
        RECT 2215.890 186.560 2216.210 186.620 ;
        RECT 2215.695 186.420 2216.210 186.560 ;
        RECT 2215.890 186.360 2216.210 186.420 ;
        RECT 2215.890 137.940 2216.210 138.000 ;
        RECT 2215.695 137.800 2216.210 137.940 ;
        RECT 2215.890 137.740 2216.210 137.800 ;
        RECT 2215.890 48.520 2216.210 48.580 ;
        RECT 2215.695 48.380 2216.210 48.520 ;
        RECT 2215.890 48.320 2216.210 48.380 ;
        RECT 2214.970 2.960 2215.290 3.020 ;
        RECT 2215.890 2.960 2216.210 3.020 ;
        RECT 2214.970 2.820 2216.210 2.960 ;
        RECT 2214.970 2.760 2215.290 2.820 ;
        RECT 2215.890 2.760 2216.210 2.820 ;
      LAYER via ;
        RECT 1909.560 203.700 1909.820 203.960 ;
        RECT 2215.920 186.360 2216.180 186.620 ;
        RECT 2215.920 137.740 2216.180 138.000 ;
        RECT 2215.920 48.320 2216.180 48.580 ;
        RECT 2215.000 2.760 2215.260 3.020 ;
        RECT 2215.920 2.760 2216.180 3.020 ;
      LAYER met2 ;
        RECT 1909.510 216.000 1909.790 220.000 ;
        RECT 1909.620 203.990 1909.760 216.000 ;
        RECT 1909.560 203.670 1909.820 203.990 ;
        RECT 2215.920 186.330 2216.180 186.650 ;
        RECT 2215.980 138.030 2216.120 186.330 ;
        RECT 2215.920 137.710 2216.180 138.030 ;
        RECT 2215.920 48.290 2216.180 48.610 ;
        RECT 2215.980 3.050 2216.120 48.290 ;
        RECT 2215.000 2.730 2215.260 3.050 ;
        RECT 2215.920 2.730 2216.180 3.050 ;
        RECT 2215.060 2.400 2215.200 2.730 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1927.470 200.500 1927.790 200.560 ;
        RECT 1931.610 200.500 1931.930 200.560 ;
        RECT 1927.470 200.360 1931.930 200.500 ;
        RECT 1927.470 200.300 1927.790 200.360 ;
        RECT 1931.610 200.300 1931.930 200.360 ;
        RECT 1931.610 19.620 1931.930 19.680 ;
        RECT 2232.910 19.620 2233.230 19.680 ;
        RECT 1931.610 19.480 2233.230 19.620 ;
        RECT 1931.610 19.420 1931.930 19.480 ;
        RECT 2232.910 19.420 2233.230 19.480 ;
      LAYER via ;
        RECT 1927.500 200.300 1927.760 200.560 ;
        RECT 1931.640 200.300 1931.900 200.560 ;
        RECT 1931.640 19.420 1931.900 19.680 ;
        RECT 2232.940 19.420 2233.200 19.680 ;
      LAYER met2 ;
        RECT 1927.450 216.000 1927.730 220.000 ;
        RECT 1927.560 200.590 1927.700 216.000 ;
        RECT 1927.500 200.270 1927.760 200.590 ;
        RECT 1931.640 200.270 1931.900 200.590 ;
        RECT 1931.700 19.710 1931.840 200.270 ;
        RECT 1931.640 19.390 1931.900 19.710 ;
        RECT 2232.940 19.390 2233.200 19.710 ;
        RECT 2233.000 2.400 2233.140 19.390 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 479.390 203.560 479.710 203.620 ;
        RECT 787.130 203.560 787.450 203.620 ;
        RECT 479.390 203.420 787.450 203.560 ;
        RECT 479.390 203.360 479.710 203.420 ;
        RECT 787.130 203.360 787.450 203.420 ;
      LAYER via ;
        RECT 479.420 203.360 479.680 203.620 ;
        RECT 787.160 203.360 787.420 203.620 ;
      LAYER met2 ;
        RECT 479.370 216.000 479.650 220.000 ;
        RECT 479.480 203.650 479.620 216.000 ;
        RECT 479.420 203.330 479.680 203.650 ;
        RECT 787.160 203.330 787.420 203.650 ;
        RECT 787.220 7.890 787.360 203.330 ;
        RECT 787.220 7.750 787.820 7.890 ;
        RECT 787.680 2.400 787.820 7.750 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2250.005 186.405 2250.175 204.255 ;
      LAYER mcon ;
        RECT 2250.005 204.085 2250.175 204.255 ;
      LAYER met1 ;
        RECT 1945.410 204.240 1945.730 204.300 ;
        RECT 2249.945 204.240 2250.235 204.285 ;
        RECT 1945.410 204.100 2250.235 204.240 ;
        RECT 1945.410 204.040 1945.730 204.100 ;
        RECT 2249.945 204.055 2250.235 204.100 ;
        RECT 2249.930 186.560 2250.250 186.620 ;
        RECT 2249.735 186.420 2250.250 186.560 ;
        RECT 2249.930 186.360 2250.250 186.420 ;
        RECT 2249.930 137.940 2250.250 138.000 ;
        RECT 2251.770 137.940 2252.090 138.000 ;
        RECT 2249.930 137.800 2252.090 137.940 ;
        RECT 2249.930 137.740 2250.250 137.800 ;
        RECT 2251.770 137.740 2252.090 137.800 ;
        RECT 2250.850 2.960 2251.170 3.020 ;
        RECT 2251.770 2.960 2252.090 3.020 ;
        RECT 2250.850 2.820 2252.090 2.960 ;
        RECT 2250.850 2.760 2251.170 2.820 ;
        RECT 2251.770 2.760 2252.090 2.820 ;
      LAYER via ;
        RECT 1945.440 204.040 1945.700 204.300 ;
        RECT 2249.960 186.360 2250.220 186.620 ;
        RECT 2249.960 137.740 2250.220 138.000 ;
        RECT 2251.800 137.740 2252.060 138.000 ;
        RECT 2250.880 2.760 2251.140 3.020 ;
        RECT 2251.800 2.760 2252.060 3.020 ;
      LAYER met2 ;
        RECT 1945.390 216.000 1945.670 220.000 ;
        RECT 1945.500 204.330 1945.640 216.000 ;
        RECT 1945.440 204.010 1945.700 204.330 ;
        RECT 2249.960 186.330 2250.220 186.650 ;
        RECT 2250.020 138.030 2250.160 186.330 ;
        RECT 2249.960 137.710 2250.220 138.030 ;
        RECT 2251.800 137.710 2252.060 138.030 ;
        RECT 2251.860 3.050 2252.000 137.710 ;
        RECT 2250.880 2.730 2251.140 3.050 ;
        RECT 2251.800 2.730 2252.060 3.050 ;
        RECT 2250.940 2.400 2251.080 2.730 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 20.300 1966.430 20.360 ;
        RECT 2268.330 20.300 2268.650 20.360 ;
        RECT 1966.110 20.160 2268.650 20.300 ;
        RECT 1966.110 20.100 1966.430 20.160 ;
        RECT 2268.330 20.100 2268.650 20.160 ;
      LAYER via ;
        RECT 1966.140 20.100 1966.400 20.360 ;
        RECT 2268.360 20.100 2268.620 20.360 ;
      LAYER met2 ;
        RECT 1963.330 216.650 1963.610 220.000 ;
        RECT 1963.330 216.510 1966.340 216.650 ;
        RECT 1963.330 216.000 1963.610 216.510 ;
        RECT 1966.200 20.390 1966.340 216.510 ;
        RECT 1966.140 20.070 1966.400 20.390 ;
        RECT 2268.360 20.070 2268.620 20.390 ;
        RECT 2268.420 2.400 2268.560 20.070 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1980.830 205.600 1981.150 205.660 ;
        RECT 2284.430 205.600 2284.750 205.660 ;
        RECT 1980.830 205.460 2284.750 205.600 ;
        RECT 1980.830 205.400 1981.150 205.460 ;
        RECT 2284.430 205.400 2284.750 205.460 ;
      LAYER via ;
        RECT 1980.860 205.400 1981.120 205.660 ;
        RECT 2284.460 205.400 2284.720 205.660 ;
      LAYER met2 ;
        RECT 1980.810 216.000 1981.090 220.000 ;
        RECT 1980.920 205.690 1981.060 216.000 ;
        RECT 1980.860 205.370 1981.120 205.690 ;
        RECT 2284.460 205.370 2284.720 205.690 ;
        RECT 2284.520 3.130 2284.660 205.370 ;
        RECT 2284.520 2.990 2286.040 3.130 ;
        RECT 2285.900 2.960 2286.040 2.990 ;
        RECT 2285.900 2.820 2286.500 2.960 ;
        RECT 2286.360 2.400 2286.500 2.820 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2000.610 17.920 2000.930 17.980 ;
        RECT 2304.210 17.920 2304.530 17.980 ;
        RECT 2000.610 17.780 2304.530 17.920 ;
        RECT 2000.610 17.720 2000.930 17.780 ;
        RECT 2304.210 17.720 2304.530 17.780 ;
      LAYER via ;
        RECT 2000.640 17.720 2000.900 17.980 ;
        RECT 2304.240 17.720 2304.500 17.980 ;
      LAYER met2 ;
        RECT 1998.750 216.650 1999.030 220.000 ;
        RECT 1998.750 216.510 2000.840 216.650 ;
        RECT 1998.750 216.000 1999.030 216.510 ;
        RECT 2000.700 18.010 2000.840 216.510 ;
        RECT 2000.640 17.690 2000.900 18.010 ;
        RECT 2304.240 17.690 2304.500 18.010 ;
        RECT 2304.300 2.400 2304.440 17.690 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2016.710 205.260 2017.030 205.320 ;
        RECT 2318.930 205.260 2319.250 205.320 ;
        RECT 2016.710 205.120 2319.250 205.260 ;
        RECT 2016.710 205.060 2017.030 205.120 ;
        RECT 2318.930 205.060 2319.250 205.120 ;
        RECT 2318.930 2.960 2319.250 3.020 ;
        RECT 2322.150 2.960 2322.470 3.020 ;
        RECT 2318.930 2.820 2322.470 2.960 ;
        RECT 2318.930 2.760 2319.250 2.820 ;
        RECT 2322.150 2.760 2322.470 2.820 ;
      LAYER via ;
        RECT 2016.740 205.060 2017.000 205.320 ;
        RECT 2318.960 205.060 2319.220 205.320 ;
        RECT 2318.960 2.760 2319.220 3.020 ;
        RECT 2322.180 2.760 2322.440 3.020 ;
      LAYER met2 ;
        RECT 2016.690 216.000 2016.970 220.000 ;
        RECT 2016.800 205.350 2016.940 216.000 ;
        RECT 2016.740 205.030 2017.000 205.350 ;
        RECT 2318.960 205.030 2319.220 205.350 ;
        RECT 2319.020 3.050 2319.160 205.030 ;
        RECT 2318.960 2.730 2319.220 3.050 ;
        RECT 2322.180 2.730 2322.440 3.050 ;
        RECT 2322.240 2.400 2322.380 2.730 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2034.630 216.650 2034.910 220.000 ;
        RECT 2034.630 216.510 2035.340 216.650 ;
        RECT 2034.630 216.000 2034.910 216.510 ;
        RECT 2035.200 16.845 2035.340 216.510 ;
        RECT 2035.130 16.475 2035.410 16.845 ;
        RECT 2339.650 16.475 2339.930 16.845 ;
        RECT 2339.720 2.400 2339.860 16.475 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
      LAYER via2 ;
        RECT 2035.130 16.520 2035.410 16.800 ;
        RECT 2339.650 16.520 2339.930 16.800 ;
      LAYER met3 ;
        RECT 2035.105 16.810 2035.435 16.825 ;
        RECT 2339.625 16.810 2339.955 16.825 ;
        RECT 2035.105 16.510 2339.955 16.810 ;
        RECT 2035.105 16.495 2035.435 16.510 ;
        RECT 2339.625 16.495 2339.955 16.510 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 18.260 2056.130 18.320 ;
        RECT 2357.570 18.260 2357.890 18.320 ;
        RECT 2055.810 18.120 2357.890 18.260 ;
        RECT 2055.810 18.060 2056.130 18.120 ;
        RECT 2357.570 18.060 2357.890 18.120 ;
      LAYER via ;
        RECT 2055.840 18.060 2056.100 18.320 ;
        RECT 2357.600 18.060 2357.860 18.320 ;
      LAYER met2 ;
        RECT 2052.570 216.650 2052.850 220.000 ;
        RECT 2052.570 216.510 2056.040 216.650 ;
        RECT 2052.570 216.000 2052.850 216.510 ;
        RECT 2055.900 18.350 2056.040 216.510 ;
        RECT 2055.840 18.030 2056.100 18.350 ;
        RECT 2357.600 18.030 2357.860 18.350 ;
        RECT 2357.660 2.400 2357.800 18.030 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2070.530 200.500 2070.850 200.560 ;
        RECT 2076.510 200.500 2076.830 200.560 ;
        RECT 2070.530 200.360 2076.830 200.500 ;
        RECT 2070.530 200.300 2070.850 200.360 ;
        RECT 2076.510 200.300 2076.830 200.360 ;
        RECT 2076.510 18.600 2076.830 18.660 ;
        RECT 2375.510 18.600 2375.830 18.660 ;
        RECT 2076.510 18.460 2375.830 18.600 ;
        RECT 2076.510 18.400 2076.830 18.460 ;
        RECT 2375.510 18.400 2375.830 18.460 ;
      LAYER via ;
        RECT 2070.560 200.300 2070.820 200.560 ;
        RECT 2076.540 200.300 2076.800 200.560 ;
        RECT 2076.540 18.400 2076.800 18.660 ;
        RECT 2375.540 18.400 2375.800 18.660 ;
      LAYER met2 ;
        RECT 2070.510 216.000 2070.790 220.000 ;
        RECT 2070.620 200.590 2070.760 216.000 ;
        RECT 2070.560 200.270 2070.820 200.590 ;
        RECT 2076.540 200.270 2076.800 200.590 ;
        RECT 2076.600 18.690 2076.740 200.270 ;
        RECT 2076.540 18.370 2076.800 18.690 ;
        RECT 2375.540 18.370 2375.800 18.690 ;
        RECT 2375.600 2.400 2375.740 18.370 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 18.940 2090.630 19.000 ;
        RECT 2393.450 18.940 2393.770 19.000 ;
        RECT 2090.310 18.800 2393.770 18.940 ;
        RECT 2090.310 18.740 2090.630 18.800 ;
        RECT 2393.450 18.740 2393.770 18.800 ;
      LAYER via ;
        RECT 2090.340 18.740 2090.600 19.000 ;
        RECT 2393.480 18.740 2393.740 19.000 ;
      LAYER met2 ;
        RECT 2088.450 216.650 2088.730 220.000 ;
        RECT 2088.450 216.510 2090.540 216.650 ;
        RECT 2088.450 216.000 2088.730 216.510 ;
        RECT 2090.400 19.030 2090.540 216.510 ;
        RECT 2090.340 18.710 2090.600 19.030 ;
        RECT 2393.480 18.710 2393.740 19.030 ;
        RECT 2393.540 2.400 2393.680 18.710 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2105.950 200.500 2106.270 200.560 ;
        RECT 2111.010 200.500 2111.330 200.560 ;
        RECT 2105.950 200.360 2111.330 200.500 ;
        RECT 2105.950 200.300 2106.270 200.360 ;
        RECT 2111.010 200.300 2111.330 200.360 ;
        RECT 2111.010 19.280 2111.330 19.340 ;
        RECT 2411.390 19.280 2411.710 19.340 ;
        RECT 2111.010 19.140 2411.710 19.280 ;
        RECT 2111.010 19.080 2111.330 19.140 ;
        RECT 2411.390 19.080 2411.710 19.140 ;
      LAYER via ;
        RECT 2105.980 200.300 2106.240 200.560 ;
        RECT 2111.040 200.300 2111.300 200.560 ;
        RECT 2111.040 19.080 2111.300 19.340 ;
        RECT 2411.420 19.080 2411.680 19.340 ;
      LAYER met2 ;
        RECT 2105.930 216.000 2106.210 220.000 ;
        RECT 2106.040 200.590 2106.180 216.000 ;
        RECT 2105.980 200.270 2106.240 200.590 ;
        RECT 2111.040 200.270 2111.300 200.590 ;
        RECT 2111.100 19.370 2111.240 200.270 ;
        RECT 2111.040 19.050 2111.300 19.370 ;
        RECT 2411.420 19.050 2411.680 19.370 ;
        RECT 2411.480 2.400 2411.620 19.050 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 497.330 200.500 497.650 200.560 ;
        RECT 503.310 200.500 503.630 200.560 ;
        RECT 497.330 200.360 503.630 200.500 ;
        RECT 497.330 200.300 497.650 200.360 ;
        RECT 503.310 200.300 503.630 200.360 ;
        RECT 503.310 15.880 503.630 15.940 ;
        RECT 805.530 15.880 805.850 15.940 ;
        RECT 503.310 15.740 805.850 15.880 ;
        RECT 503.310 15.680 503.630 15.740 ;
        RECT 805.530 15.680 805.850 15.740 ;
      LAYER via ;
        RECT 497.360 200.300 497.620 200.560 ;
        RECT 503.340 200.300 503.600 200.560 ;
        RECT 503.340 15.680 503.600 15.940 ;
        RECT 805.560 15.680 805.820 15.940 ;
      LAYER met2 ;
        RECT 497.310 216.000 497.590 220.000 ;
        RECT 497.420 200.590 497.560 216.000 ;
        RECT 497.360 200.270 497.620 200.590 ;
        RECT 503.340 200.270 503.600 200.590 ;
        RECT 503.400 15.970 503.540 200.270 ;
        RECT 503.340 15.650 503.600 15.970 ;
        RECT 805.560 15.650 805.820 15.970 ;
        RECT 805.620 2.400 805.760 15.650 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 310.570 17.240 310.890 17.300 ;
        RECT 2.830 17.100 310.890 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 310.570 17.040 310.890 17.100 ;
      LAYER via ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 310.600 17.040 310.860 17.300 ;
      LAYER met2 ;
        RECT 312.850 216.650 313.130 220.000 ;
        RECT 310.660 216.510 313.130 216.650 ;
        RECT 310.660 17.330 310.800 216.510 ;
        RECT 312.850 216.000 313.130 216.510 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 310.600 17.010 310.860 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 317.470 17.580 317.790 17.640 ;
        RECT 8.350 17.440 317.790 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 317.470 17.380 317.790 17.440 ;
      LAYER via ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 317.500 17.380 317.760 17.640 ;
      LAYER met2 ;
        RECT 318.370 216.650 318.650 220.000 ;
        RECT 317.560 216.510 318.650 216.650 ;
        RECT 317.560 17.670 317.700 216.510 ;
        RECT 318.370 216.000 318.650 216.510 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 317.500 17.350 317.760 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 3226.000 367.020 3529.000 ;
        RECT 544.020 3226.000 547.020 3529.000 ;
        RECT 724.020 3226.000 727.020 3529.000 ;
        RECT 904.020 3226.000 907.020 3529.000 ;
        RECT 1084.020 3226.000 1087.020 3529.000 ;
        RECT 1264.020 3226.000 1267.020 3529.000 ;
        RECT 1444.020 3226.000 1447.020 3529.000 ;
        RECT 1624.020 3226.000 1627.020 3529.000 ;
        RECT 1804.020 3226.000 1807.020 3529.000 ;
        RECT 1984.020 3226.000 1987.020 3529.000 ;
        RECT 2164.020 3226.000 2167.020 3529.000 ;
        RECT 2344.020 3226.000 2347.020 3529.000 ;
        RECT 2524.020 3226.000 2527.020 3529.000 ;
        RECT 331.040 226.640 332.640 3202.800 ;
        RECT 364.020 -9.320 367.020 206.000 ;
        RECT 544.020 -9.320 547.020 206.000 ;
        RECT 724.020 -9.320 727.020 206.000 ;
        RECT 904.020 -9.320 907.020 206.000 ;
        RECT 1084.020 -9.320 1087.020 206.000 ;
        RECT 1264.020 -9.320 1267.020 206.000 ;
        RECT 1444.020 -9.320 1447.020 206.000 ;
        RECT 1624.020 -9.320 1627.020 206.000 ;
        RECT 1804.020 -9.320 1807.020 206.000 ;
        RECT 1984.020 -9.320 1987.020 206.000 ;
        RECT 2164.020 -9.320 2167.020 206.000 ;
        RECT 2344.020 -9.320 2347.020 206.000 ;
        RECT 2524.020 -9.320 2527.020 206.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 331.250 3071.090 332.430 3072.270 ;
        RECT 331.250 3069.490 332.430 3070.670 ;
        RECT 331.250 2891.090 332.430 2892.270 ;
        RECT 331.250 2889.490 332.430 2890.670 ;
        RECT 331.250 2711.090 332.430 2712.270 ;
        RECT 331.250 2709.490 332.430 2710.670 ;
        RECT 331.250 2531.090 332.430 2532.270 ;
        RECT 331.250 2529.490 332.430 2530.670 ;
        RECT 331.250 2351.090 332.430 2352.270 ;
        RECT 331.250 2349.490 332.430 2350.670 ;
        RECT 331.250 2171.090 332.430 2172.270 ;
        RECT 331.250 2169.490 332.430 2170.670 ;
        RECT 331.250 1991.090 332.430 1992.270 ;
        RECT 331.250 1989.490 332.430 1990.670 ;
        RECT 331.250 1811.090 332.430 1812.270 ;
        RECT 331.250 1809.490 332.430 1810.670 ;
        RECT 331.250 1631.090 332.430 1632.270 ;
        RECT 331.250 1629.490 332.430 1630.670 ;
        RECT 331.250 1451.090 332.430 1452.270 ;
        RECT 331.250 1449.490 332.430 1450.670 ;
        RECT 331.250 1271.090 332.430 1272.270 ;
        RECT 331.250 1269.490 332.430 1270.670 ;
        RECT 331.250 1091.090 332.430 1092.270 ;
        RECT 331.250 1089.490 332.430 1090.670 ;
        RECT 331.250 911.090 332.430 912.270 ;
        RECT 331.250 909.490 332.430 910.670 ;
        RECT 331.250 731.090 332.430 732.270 ;
        RECT 331.250 729.490 332.430 730.670 ;
        RECT 331.250 551.090 332.430 552.270 ;
        RECT 331.250 549.490 332.430 550.670 ;
        RECT 331.250 371.090 332.430 372.270 ;
        RECT 331.250 369.490 332.430 370.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 331.040 3072.380 332.640 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 331.040 3069.370 332.640 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 331.040 2892.380 332.640 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 331.040 2889.370 332.640 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 331.040 2712.380 332.640 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 331.040 2709.370 332.640 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 331.040 2532.380 332.640 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 331.040 2529.370 332.640 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 331.040 2352.380 332.640 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 331.040 2349.370 332.640 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 331.040 2172.380 332.640 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 331.040 2169.370 332.640 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 331.040 1992.380 332.640 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 331.040 1989.370 332.640 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 331.040 1812.380 332.640 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 331.040 1809.370 332.640 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 331.040 1632.380 332.640 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 331.040 1629.370 332.640 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 331.040 1452.380 332.640 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 331.040 1449.370 332.640 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 331.040 1272.380 332.640 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 331.040 1269.370 332.640 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 331.040 1092.380 332.640 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 331.040 1089.370 332.640 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 331.040 912.380 332.640 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 331.040 909.370 332.640 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 331.040 732.380 332.640 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 331.040 729.370 332.640 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 331.040 552.380 332.640 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 331.040 549.370 332.640 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 331.040 372.380 332.640 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 331.040 369.370 332.640 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 3226.000 457.020 3529.000 ;
        RECT 634.020 3226.000 637.020 3529.000 ;
        RECT 814.020 3226.000 817.020 3529.000 ;
        RECT 994.020 3226.000 997.020 3529.000 ;
        RECT 1174.020 3226.000 1177.020 3529.000 ;
        RECT 1354.020 3226.000 1357.020 3529.000 ;
        RECT 1534.020 3226.000 1537.020 3529.000 ;
        RECT 1714.020 3226.000 1717.020 3529.000 ;
        RECT 1894.020 3226.000 1897.020 3529.000 ;
        RECT 2074.020 3226.000 2077.020 3529.000 ;
        RECT 2254.020 3226.000 2257.020 3529.000 ;
        RECT 2434.020 3226.000 2437.020 3529.000 ;
        RECT 2614.020 3226.000 2617.020 3529.000 ;
        RECT 407.840 226.640 409.440 3202.800 ;
        RECT 454.020 -9.320 457.020 206.000 ;
        RECT 634.020 -9.320 637.020 206.000 ;
        RECT 814.020 -9.320 817.020 206.000 ;
        RECT 994.020 -9.320 997.020 206.000 ;
        RECT 1174.020 -9.320 1177.020 206.000 ;
        RECT 1354.020 -9.320 1357.020 206.000 ;
        RECT 1534.020 -9.320 1537.020 206.000 ;
        RECT 1714.020 -9.320 1717.020 206.000 ;
        RECT 1894.020 -9.320 1897.020 206.000 ;
        RECT 2074.020 -9.320 2077.020 206.000 ;
        RECT 2254.020 -9.320 2257.020 206.000 ;
        RECT 2434.020 -9.320 2437.020 206.000 ;
        RECT 2614.020 -9.320 2617.020 206.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 408.050 3161.090 409.230 3162.270 ;
        RECT 408.050 3159.490 409.230 3160.670 ;
        RECT 408.050 2981.090 409.230 2982.270 ;
        RECT 408.050 2979.490 409.230 2980.670 ;
        RECT 408.050 2801.090 409.230 2802.270 ;
        RECT 408.050 2799.490 409.230 2800.670 ;
        RECT 408.050 2621.090 409.230 2622.270 ;
        RECT 408.050 2619.490 409.230 2620.670 ;
        RECT 408.050 2441.090 409.230 2442.270 ;
        RECT 408.050 2439.490 409.230 2440.670 ;
        RECT 408.050 2261.090 409.230 2262.270 ;
        RECT 408.050 2259.490 409.230 2260.670 ;
        RECT 408.050 2081.090 409.230 2082.270 ;
        RECT 408.050 2079.490 409.230 2080.670 ;
        RECT 408.050 1901.090 409.230 1902.270 ;
        RECT 408.050 1899.490 409.230 1900.670 ;
        RECT 408.050 1721.090 409.230 1722.270 ;
        RECT 408.050 1719.490 409.230 1720.670 ;
        RECT 408.050 1541.090 409.230 1542.270 ;
        RECT 408.050 1539.490 409.230 1540.670 ;
        RECT 408.050 1361.090 409.230 1362.270 ;
        RECT 408.050 1359.490 409.230 1360.670 ;
        RECT 408.050 1181.090 409.230 1182.270 ;
        RECT 408.050 1179.490 409.230 1180.670 ;
        RECT 408.050 1001.090 409.230 1002.270 ;
        RECT 408.050 999.490 409.230 1000.670 ;
        RECT 408.050 821.090 409.230 822.270 ;
        RECT 408.050 819.490 409.230 820.670 ;
        RECT 408.050 641.090 409.230 642.270 ;
        RECT 408.050 639.490 409.230 640.670 ;
        RECT 408.050 461.090 409.230 462.270 ;
        RECT 408.050 459.490 409.230 460.670 ;
        RECT 408.050 281.090 409.230 282.270 ;
        RECT 408.050 279.490 409.230 280.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 407.840 3162.380 409.440 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 407.840 3159.370 409.440 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 407.840 2982.380 409.440 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 407.840 2979.370 409.440 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 407.840 2802.380 409.440 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 407.840 2799.370 409.440 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 407.840 2622.380 409.440 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 407.840 2619.370 409.440 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 407.840 2442.380 409.440 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 407.840 2439.370 409.440 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 407.840 2262.380 409.440 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 407.840 2259.370 409.440 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 407.840 2082.380 409.440 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 407.840 2079.370 409.440 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 407.840 1902.380 409.440 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 407.840 1899.370 409.440 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 407.840 1722.380 409.440 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 407.840 1719.370 409.440 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 407.840 1542.380 409.440 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 407.840 1539.370 409.440 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 407.840 1362.380 409.440 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 407.840 1359.370 409.440 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 407.840 1182.380 409.440 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 407.840 1179.370 409.440 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 407.840 1002.380 409.440 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 407.840 999.370 409.440 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 407.840 822.380 409.440 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 407.840 819.370 409.440 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 407.840 642.380 409.440 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 407.840 639.370 409.440 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 407.840 462.380 409.440 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 407.840 459.370 409.440 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 407.840 282.380 409.440 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 407.840 279.370 409.440 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 315.520 226.795 2604.480 3202.645 ;
      LAYER met1 ;
        RECT 315.520 224.540 2604.480 3202.800 ;
      LAYER met2 ;
        RECT 312.850 3211.720 352.130 3212.000 ;
        RECT 352.970 3211.720 437.230 3212.000 ;
        RECT 438.070 3211.720 522.330 3212.000 ;
        RECT 523.170 3211.720 607.430 3212.000 ;
        RECT 608.270 3211.720 692.530 3212.000 ;
        RECT 693.370 3211.720 777.630 3212.000 ;
        RECT 778.470 3211.720 863.190 3212.000 ;
        RECT 864.030 3211.720 948.290 3212.000 ;
        RECT 949.130 3211.720 1033.390 3212.000 ;
        RECT 1034.230 3211.720 1118.490 3212.000 ;
        RECT 1119.330 3211.720 1203.590 3212.000 ;
        RECT 1204.430 3211.720 1289.150 3212.000 ;
        RECT 1289.990 3211.720 1374.250 3212.000 ;
        RECT 1375.090 3211.720 1459.350 3212.000 ;
        RECT 1460.190 3211.720 1544.450 3212.000 ;
        RECT 1545.290 3211.720 1629.550 3212.000 ;
        RECT 1630.390 3211.720 1714.650 3212.000 ;
        RECT 1715.490 3211.720 1800.210 3212.000 ;
        RECT 1801.050 3211.720 1885.310 3212.000 ;
        RECT 1886.150 3211.720 1970.410 3212.000 ;
        RECT 1971.250 3211.720 2055.510 3212.000 ;
        RECT 2056.350 3211.720 2140.610 3212.000 ;
        RECT 2141.450 3211.720 2226.170 3212.000 ;
        RECT 2227.010 3211.720 2311.270 3212.000 ;
        RECT 2312.110 3211.720 2396.370 3212.000 ;
        RECT 2397.210 3211.720 2481.470 3212.000 ;
        RECT 2482.310 3211.720 2566.570 3212.000 ;
        RECT 2567.410 3211.720 2602.540 3212.000 ;
        RECT 312.850 220.280 2602.540 3211.720 ;
        RECT 313.410 220.000 318.090 220.280 ;
        RECT 318.930 220.000 324.070 220.280 ;
        RECT 324.910 220.000 330.050 220.280 ;
        RECT 330.890 220.000 336.030 220.280 ;
        RECT 336.870 220.000 342.010 220.280 ;
        RECT 342.850 220.000 347.990 220.280 ;
        RECT 348.830 220.000 353.970 220.280 ;
        RECT 354.810 220.000 359.950 220.280 ;
        RECT 360.790 220.000 365.930 220.280 ;
        RECT 366.770 220.000 371.910 220.280 ;
        RECT 372.750 220.000 377.890 220.280 ;
        RECT 378.730 220.000 383.870 220.280 ;
        RECT 384.710 220.000 389.850 220.280 ;
        RECT 390.690 220.000 395.830 220.280 ;
        RECT 396.670 220.000 401.810 220.280 ;
        RECT 402.650 220.000 407.790 220.280 ;
        RECT 408.630 220.000 413.770 220.280 ;
        RECT 414.610 220.000 419.750 220.280 ;
        RECT 420.590 220.000 425.730 220.280 ;
        RECT 426.570 220.000 431.710 220.280 ;
        RECT 432.550 220.000 437.690 220.280 ;
        RECT 438.530 220.000 443.210 220.280 ;
        RECT 444.050 220.000 449.190 220.280 ;
        RECT 450.030 220.000 455.170 220.280 ;
        RECT 456.010 220.000 461.150 220.280 ;
        RECT 461.990 220.000 467.130 220.280 ;
        RECT 467.970 220.000 473.110 220.280 ;
        RECT 473.950 220.000 479.090 220.280 ;
        RECT 479.930 220.000 485.070 220.280 ;
        RECT 485.910 220.000 491.050 220.280 ;
        RECT 491.890 220.000 497.030 220.280 ;
        RECT 497.870 220.000 503.010 220.280 ;
        RECT 503.850 220.000 508.990 220.280 ;
        RECT 509.830 220.000 514.970 220.280 ;
        RECT 515.810 220.000 520.950 220.280 ;
        RECT 521.790 220.000 526.930 220.280 ;
        RECT 527.770 220.000 532.910 220.280 ;
        RECT 533.750 220.000 538.890 220.280 ;
        RECT 539.730 220.000 544.870 220.280 ;
        RECT 545.710 220.000 550.850 220.280 ;
        RECT 551.690 220.000 556.830 220.280 ;
        RECT 557.670 220.000 562.810 220.280 ;
        RECT 563.650 220.000 568.330 220.280 ;
        RECT 569.170 220.000 574.310 220.280 ;
        RECT 575.150 220.000 580.290 220.280 ;
        RECT 581.130 220.000 586.270 220.280 ;
        RECT 587.110 220.000 592.250 220.280 ;
        RECT 593.090 220.000 598.230 220.280 ;
        RECT 599.070 220.000 604.210 220.280 ;
        RECT 605.050 220.000 610.190 220.280 ;
        RECT 611.030 220.000 616.170 220.280 ;
        RECT 617.010 220.000 622.150 220.280 ;
        RECT 622.990 220.000 628.130 220.280 ;
        RECT 628.970 220.000 634.110 220.280 ;
        RECT 634.950 220.000 640.090 220.280 ;
        RECT 640.930 220.000 646.070 220.280 ;
        RECT 646.910 220.000 652.050 220.280 ;
        RECT 652.890 220.000 658.030 220.280 ;
        RECT 658.870 220.000 664.010 220.280 ;
        RECT 664.850 220.000 669.990 220.280 ;
        RECT 670.830 220.000 675.970 220.280 ;
        RECT 676.810 220.000 681.950 220.280 ;
        RECT 682.790 220.000 687.930 220.280 ;
        RECT 688.770 220.000 693.910 220.280 ;
        RECT 694.750 220.000 699.430 220.280 ;
        RECT 700.270 220.000 705.410 220.280 ;
        RECT 706.250 220.000 711.390 220.280 ;
        RECT 712.230 220.000 717.370 220.280 ;
        RECT 718.210 220.000 723.350 220.280 ;
        RECT 724.190 220.000 729.330 220.280 ;
        RECT 730.170 220.000 735.310 220.280 ;
        RECT 736.150 220.000 741.290 220.280 ;
        RECT 742.130 220.000 747.270 220.280 ;
        RECT 748.110 220.000 753.250 220.280 ;
        RECT 754.090 220.000 759.230 220.280 ;
        RECT 760.070 220.000 765.210 220.280 ;
        RECT 766.050 220.000 771.190 220.280 ;
        RECT 772.030 220.000 777.170 220.280 ;
        RECT 778.010 220.000 783.150 220.280 ;
        RECT 783.990 220.000 789.130 220.280 ;
        RECT 789.970 220.000 795.110 220.280 ;
        RECT 795.950 220.000 801.090 220.280 ;
        RECT 801.930 220.000 807.070 220.280 ;
        RECT 807.910 220.000 813.050 220.280 ;
        RECT 813.890 220.000 819.030 220.280 ;
        RECT 819.870 220.000 824.550 220.280 ;
        RECT 825.390 220.000 830.530 220.280 ;
        RECT 831.370 220.000 836.510 220.280 ;
        RECT 837.350 220.000 842.490 220.280 ;
        RECT 843.330 220.000 848.470 220.280 ;
        RECT 849.310 220.000 854.450 220.280 ;
        RECT 855.290 220.000 860.430 220.280 ;
        RECT 861.270 220.000 866.410 220.280 ;
        RECT 867.250 220.000 872.390 220.280 ;
        RECT 873.230 220.000 878.370 220.280 ;
        RECT 879.210 220.000 884.350 220.280 ;
        RECT 885.190 220.000 890.330 220.280 ;
        RECT 891.170 220.000 896.310 220.280 ;
        RECT 897.150 220.000 902.290 220.280 ;
        RECT 903.130 220.000 908.270 220.280 ;
        RECT 909.110 220.000 914.250 220.280 ;
        RECT 915.090 220.000 920.230 220.280 ;
        RECT 921.070 220.000 926.210 220.280 ;
        RECT 927.050 220.000 932.190 220.280 ;
        RECT 933.030 220.000 938.170 220.280 ;
        RECT 939.010 220.000 944.150 220.280 ;
        RECT 944.990 220.000 950.130 220.280 ;
        RECT 950.970 220.000 955.650 220.280 ;
        RECT 956.490 220.000 961.630 220.280 ;
        RECT 962.470 220.000 967.610 220.280 ;
        RECT 968.450 220.000 973.590 220.280 ;
        RECT 974.430 220.000 979.570 220.280 ;
        RECT 980.410 220.000 985.550 220.280 ;
        RECT 986.390 220.000 991.530 220.280 ;
        RECT 992.370 220.000 997.510 220.280 ;
        RECT 998.350 220.000 1003.490 220.280 ;
        RECT 1004.330 220.000 1009.470 220.280 ;
        RECT 1010.310 220.000 1015.450 220.280 ;
        RECT 1016.290 220.000 1021.430 220.280 ;
        RECT 1022.270 220.000 1027.410 220.280 ;
        RECT 1028.250 220.000 1033.390 220.280 ;
        RECT 1034.230 220.000 1039.370 220.280 ;
        RECT 1040.210 220.000 1045.350 220.280 ;
        RECT 1046.190 220.000 1051.330 220.280 ;
        RECT 1052.170 220.000 1057.310 220.280 ;
        RECT 1058.150 220.000 1063.290 220.280 ;
        RECT 1064.130 220.000 1069.270 220.280 ;
        RECT 1070.110 220.000 1075.250 220.280 ;
        RECT 1076.090 220.000 1080.770 220.280 ;
        RECT 1081.610 220.000 1086.750 220.280 ;
        RECT 1087.590 220.000 1092.730 220.280 ;
        RECT 1093.570 220.000 1098.710 220.280 ;
        RECT 1099.550 220.000 1104.690 220.280 ;
        RECT 1105.530 220.000 1110.670 220.280 ;
        RECT 1111.510 220.000 1116.650 220.280 ;
        RECT 1117.490 220.000 1122.630 220.280 ;
        RECT 1123.470 220.000 1128.610 220.280 ;
        RECT 1129.450 220.000 1134.590 220.280 ;
        RECT 1135.430 220.000 1140.570 220.280 ;
        RECT 1141.410 220.000 1146.550 220.280 ;
        RECT 1147.390 220.000 1152.530 220.280 ;
        RECT 1153.370 220.000 1158.510 220.280 ;
        RECT 1159.350 220.000 1164.490 220.280 ;
        RECT 1165.330 220.000 1170.470 220.280 ;
        RECT 1171.310 220.000 1176.450 220.280 ;
        RECT 1177.290 220.000 1182.430 220.280 ;
        RECT 1183.270 220.000 1188.410 220.280 ;
        RECT 1189.250 220.000 1194.390 220.280 ;
        RECT 1195.230 220.000 1200.370 220.280 ;
        RECT 1201.210 220.000 1206.350 220.280 ;
        RECT 1207.190 220.000 1211.870 220.280 ;
        RECT 1212.710 220.000 1217.850 220.280 ;
        RECT 1218.690 220.000 1223.830 220.280 ;
        RECT 1224.670 220.000 1229.810 220.280 ;
        RECT 1230.650 220.000 1235.790 220.280 ;
        RECT 1236.630 220.000 1241.770 220.280 ;
        RECT 1242.610 220.000 1247.750 220.280 ;
        RECT 1248.590 220.000 1253.730 220.280 ;
        RECT 1254.570 220.000 1259.710 220.280 ;
        RECT 1260.550 220.000 1265.690 220.280 ;
        RECT 1266.530 220.000 1271.670 220.280 ;
        RECT 1272.510 220.000 1277.650 220.280 ;
        RECT 1278.490 220.000 1283.630 220.280 ;
        RECT 1284.470 220.000 1289.610 220.280 ;
        RECT 1290.450 220.000 1295.590 220.280 ;
        RECT 1296.430 220.000 1301.570 220.280 ;
        RECT 1302.410 220.000 1307.550 220.280 ;
        RECT 1308.390 220.000 1313.530 220.280 ;
        RECT 1314.370 220.000 1319.510 220.280 ;
        RECT 1320.350 220.000 1325.490 220.280 ;
        RECT 1326.330 220.000 1331.470 220.280 ;
        RECT 1332.310 220.000 1336.990 220.280 ;
        RECT 1337.830 220.000 1342.970 220.280 ;
        RECT 1343.810 220.000 1348.950 220.280 ;
        RECT 1349.790 220.000 1354.930 220.280 ;
        RECT 1355.770 220.000 1360.910 220.280 ;
        RECT 1361.750 220.000 1366.890 220.280 ;
        RECT 1367.730 220.000 1372.870 220.280 ;
        RECT 1373.710 220.000 1378.850 220.280 ;
        RECT 1379.690 220.000 1384.830 220.280 ;
        RECT 1385.670 220.000 1390.810 220.280 ;
        RECT 1391.650 220.000 1396.790 220.280 ;
        RECT 1397.630 220.000 1402.770 220.280 ;
        RECT 1403.610 220.000 1408.750 220.280 ;
        RECT 1409.590 220.000 1414.730 220.280 ;
        RECT 1415.570 220.000 1420.710 220.280 ;
        RECT 1421.550 220.000 1426.690 220.280 ;
        RECT 1427.530 220.000 1432.670 220.280 ;
        RECT 1433.510 220.000 1438.650 220.280 ;
        RECT 1439.490 220.000 1444.630 220.280 ;
        RECT 1445.470 220.000 1450.610 220.280 ;
        RECT 1451.450 220.000 1456.590 220.280 ;
        RECT 1457.430 220.000 1462.570 220.280 ;
        RECT 1463.410 220.000 1468.090 220.280 ;
        RECT 1468.930 220.000 1474.070 220.280 ;
        RECT 1474.910 220.000 1480.050 220.280 ;
        RECT 1480.890 220.000 1486.030 220.280 ;
        RECT 1486.870 220.000 1492.010 220.280 ;
        RECT 1492.850 220.000 1497.990 220.280 ;
        RECT 1498.830 220.000 1503.970 220.280 ;
        RECT 1504.810 220.000 1509.950 220.280 ;
        RECT 1510.790 220.000 1515.930 220.280 ;
        RECT 1516.770 220.000 1521.910 220.280 ;
        RECT 1522.750 220.000 1527.890 220.280 ;
        RECT 1528.730 220.000 1533.870 220.280 ;
        RECT 1534.710 220.000 1539.850 220.280 ;
        RECT 1540.690 220.000 1545.830 220.280 ;
        RECT 1546.670 220.000 1551.810 220.280 ;
        RECT 1552.650 220.000 1557.790 220.280 ;
        RECT 1558.630 220.000 1563.770 220.280 ;
        RECT 1564.610 220.000 1569.750 220.280 ;
        RECT 1570.590 220.000 1575.730 220.280 ;
        RECT 1576.570 220.000 1581.710 220.280 ;
        RECT 1582.550 220.000 1587.690 220.280 ;
        RECT 1588.530 220.000 1593.210 220.280 ;
        RECT 1594.050 220.000 1599.190 220.280 ;
        RECT 1600.030 220.000 1605.170 220.280 ;
        RECT 1606.010 220.000 1611.150 220.280 ;
        RECT 1611.990 220.000 1617.130 220.280 ;
        RECT 1617.970 220.000 1623.110 220.280 ;
        RECT 1623.950 220.000 1629.090 220.280 ;
        RECT 1629.930 220.000 1635.070 220.280 ;
        RECT 1635.910 220.000 1641.050 220.280 ;
        RECT 1641.890 220.000 1647.030 220.280 ;
        RECT 1647.870 220.000 1653.010 220.280 ;
        RECT 1653.850 220.000 1658.990 220.280 ;
        RECT 1659.830 220.000 1664.970 220.280 ;
        RECT 1665.810 220.000 1670.950 220.280 ;
        RECT 1671.790 220.000 1676.930 220.280 ;
        RECT 1677.770 220.000 1682.910 220.280 ;
        RECT 1683.750 220.000 1688.890 220.280 ;
        RECT 1689.730 220.000 1694.870 220.280 ;
        RECT 1695.710 220.000 1700.850 220.280 ;
        RECT 1701.690 220.000 1706.830 220.280 ;
        RECT 1707.670 220.000 1712.810 220.280 ;
        RECT 1713.650 220.000 1718.330 220.280 ;
        RECT 1719.170 220.000 1724.310 220.280 ;
        RECT 1725.150 220.000 1730.290 220.280 ;
        RECT 1731.130 220.000 1736.270 220.280 ;
        RECT 1737.110 220.000 1742.250 220.280 ;
        RECT 1743.090 220.000 1748.230 220.280 ;
        RECT 1749.070 220.000 1754.210 220.280 ;
        RECT 1755.050 220.000 1760.190 220.280 ;
        RECT 1761.030 220.000 1766.170 220.280 ;
        RECT 1767.010 220.000 1772.150 220.280 ;
        RECT 1772.990 220.000 1778.130 220.280 ;
        RECT 1778.970 220.000 1784.110 220.280 ;
        RECT 1784.950 220.000 1790.090 220.280 ;
        RECT 1790.930 220.000 1796.070 220.280 ;
        RECT 1796.910 220.000 1802.050 220.280 ;
        RECT 1802.890 220.000 1808.030 220.280 ;
        RECT 1808.870 220.000 1814.010 220.280 ;
        RECT 1814.850 220.000 1819.990 220.280 ;
        RECT 1820.830 220.000 1825.970 220.280 ;
        RECT 1826.810 220.000 1831.950 220.280 ;
        RECT 1832.790 220.000 1837.930 220.280 ;
        RECT 1838.770 220.000 1843.910 220.280 ;
        RECT 1844.750 220.000 1849.430 220.280 ;
        RECT 1850.270 220.000 1855.410 220.280 ;
        RECT 1856.250 220.000 1861.390 220.280 ;
        RECT 1862.230 220.000 1867.370 220.280 ;
        RECT 1868.210 220.000 1873.350 220.280 ;
        RECT 1874.190 220.000 1879.330 220.280 ;
        RECT 1880.170 220.000 1885.310 220.280 ;
        RECT 1886.150 220.000 1891.290 220.280 ;
        RECT 1892.130 220.000 1897.270 220.280 ;
        RECT 1898.110 220.000 1903.250 220.280 ;
        RECT 1904.090 220.000 1909.230 220.280 ;
        RECT 1910.070 220.000 1915.210 220.280 ;
        RECT 1916.050 220.000 1921.190 220.280 ;
        RECT 1922.030 220.000 1927.170 220.280 ;
        RECT 1928.010 220.000 1933.150 220.280 ;
        RECT 1933.990 220.000 1939.130 220.280 ;
        RECT 1939.970 220.000 1945.110 220.280 ;
        RECT 1945.950 220.000 1951.090 220.280 ;
        RECT 1951.930 220.000 1957.070 220.280 ;
        RECT 1957.910 220.000 1963.050 220.280 ;
        RECT 1963.890 220.000 1969.030 220.280 ;
        RECT 1969.870 220.000 1974.550 220.280 ;
        RECT 1975.390 220.000 1980.530 220.280 ;
        RECT 1981.370 220.000 1986.510 220.280 ;
        RECT 1987.350 220.000 1992.490 220.280 ;
        RECT 1993.330 220.000 1998.470 220.280 ;
        RECT 1999.310 220.000 2004.450 220.280 ;
        RECT 2005.290 220.000 2010.430 220.280 ;
        RECT 2011.270 220.000 2016.410 220.280 ;
        RECT 2017.250 220.000 2022.390 220.280 ;
        RECT 2023.230 220.000 2028.370 220.280 ;
        RECT 2029.210 220.000 2034.350 220.280 ;
        RECT 2035.190 220.000 2040.330 220.280 ;
        RECT 2041.170 220.000 2046.310 220.280 ;
        RECT 2047.150 220.000 2052.290 220.280 ;
        RECT 2053.130 220.000 2058.270 220.280 ;
        RECT 2059.110 220.000 2064.250 220.280 ;
        RECT 2065.090 220.000 2070.230 220.280 ;
        RECT 2071.070 220.000 2076.210 220.280 ;
        RECT 2077.050 220.000 2082.190 220.280 ;
        RECT 2083.030 220.000 2088.170 220.280 ;
        RECT 2089.010 220.000 2094.150 220.280 ;
        RECT 2094.990 220.000 2100.130 220.280 ;
        RECT 2100.970 220.000 2105.650 220.280 ;
        RECT 2106.490 220.000 2111.630 220.280 ;
        RECT 2112.470 220.000 2117.610 220.280 ;
        RECT 2118.450 220.000 2123.590 220.280 ;
        RECT 2124.430 220.000 2129.570 220.280 ;
        RECT 2130.410 220.000 2135.550 220.280 ;
        RECT 2136.390 220.000 2141.530 220.280 ;
        RECT 2142.370 220.000 2147.510 220.280 ;
        RECT 2148.350 220.000 2153.490 220.280 ;
        RECT 2154.330 220.000 2159.470 220.280 ;
        RECT 2160.310 220.000 2165.450 220.280 ;
        RECT 2166.290 220.000 2171.430 220.280 ;
        RECT 2172.270 220.000 2177.410 220.280 ;
        RECT 2178.250 220.000 2183.390 220.280 ;
        RECT 2184.230 220.000 2189.370 220.280 ;
        RECT 2190.210 220.000 2195.350 220.280 ;
        RECT 2196.190 220.000 2201.330 220.280 ;
        RECT 2202.170 220.000 2207.310 220.280 ;
        RECT 2208.150 220.000 2213.290 220.280 ;
        RECT 2214.130 220.000 2219.270 220.280 ;
        RECT 2220.110 220.000 2225.250 220.280 ;
        RECT 2226.090 220.000 2230.770 220.280 ;
        RECT 2231.610 220.000 2236.750 220.280 ;
        RECT 2237.590 220.000 2242.730 220.280 ;
        RECT 2243.570 220.000 2248.710 220.280 ;
        RECT 2249.550 220.000 2254.690 220.280 ;
        RECT 2255.530 220.000 2260.670 220.280 ;
        RECT 2261.510 220.000 2266.650 220.280 ;
        RECT 2267.490 220.000 2272.630 220.280 ;
        RECT 2273.470 220.000 2278.610 220.280 ;
        RECT 2279.450 220.000 2284.590 220.280 ;
        RECT 2285.430 220.000 2290.570 220.280 ;
        RECT 2291.410 220.000 2296.550 220.280 ;
        RECT 2297.390 220.000 2302.530 220.280 ;
        RECT 2303.370 220.000 2308.510 220.280 ;
        RECT 2309.350 220.000 2314.490 220.280 ;
        RECT 2315.330 220.000 2320.470 220.280 ;
        RECT 2321.310 220.000 2326.450 220.280 ;
        RECT 2327.290 220.000 2332.430 220.280 ;
        RECT 2333.270 220.000 2338.410 220.280 ;
        RECT 2339.250 220.000 2344.390 220.280 ;
        RECT 2345.230 220.000 2350.370 220.280 ;
        RECT 2351.210 220.000 2356.350 220.280 ;
        RECT 2357.190 220.000 2361.870 220.280 ;
        RECT 2362.710 220.000 2367.850 220.280 ;
        RECT 2368.690 220.000 2373.830 220.280 ;
        RECT 2374.670 220.000 2379.810 220.280 ;
        RECT 2380.650 220.000 2385.790 220.280 ;
        RECT 2386.630 220.000 2391.770 220.280 ;
        RECT 2392.610 220.000 2397.750 220.280 ;
        RECT 2398.590 220.000 2403.730 220.280 ;
        RECT 2404.570 220.000 2409.710 220.280 ;
        RECT 2410.550 220.000 2415.690 220.280 ;
        RECT 2416.530 220.000 2421.670 220.280 ;
        RECT 2422.510 220.000 2427.650 220.280 ;
        RECT 2428.490 220.000 2433.630 220.280 ;
        RECT 2434.470 220.000 2439.610 220.280 ;
        RECT 2440.450 220.000 2445.590 220.280 ;
        RECT 2446.430 220.000 2451.570 220.280 ;
        RECT 2452.410 220.000 2457.550 220.280 ;
        RECT 2458.390 220.000 2463.530 220.280 ;
        RECT 2464.370 220.000 2469.510 220.280 ;
        RECT 2470.350 220.000 2475.490 220.280 ;
        RECT 2476.330 220.000 2481.470 220.280 ;
        RECT 2482.310 220.000 2486.990 220.280 ;
        RECT 2487.830 220.000 2492.970 220.280 ;
        RECT 2493.810 220.000 2498.950 220.280 ;
        RECT 2499.790 220.000 2504.930 220.280 ;
        RECT 2505.770 220.000 2510.910 220.280 ;
        RECT 2511.750 220.000 2516.890 220.280 ;
        RECT 2517.730 220.000 2522.870 220.280 ;
        RECT 2523.710 220.000 2528.850 220.280 ;
        RECT 2529.690 220.000 2534.830 220.280 ;
        RECT 2535.670 220.000 2540.810 220.280 ;
        RECT 2541.650 220.000 2546.790 220.280 ;
        RECT 2547.630 220.000 2552.770 220.280 ;
        RECT 2553.610 220.000 2558.750 220.280 ;
        RECT 2559.590 220.000 2564.730 220.280 ;
        RECT 2565.570 220.000 2570.710 220.280 ;
        RECT 2571.550 220.000 2576.690 220.280 ;
        RECT 2577.530 220.000 2582.670 220.280 ;
        RECT 2583.510 220.000 2588.650 220.280 ;
        RECT 2589.490 220.000 2594.630 220.280 ;
        RECT 2595.470 220.000 2600.610 220.280 ;
        RECT 2601.450 220.000 2602.540 220.280 ;
      LAYER met3 ;
        RECT 312.825 3183.200 2606.010 3202.725 ;
        RECT 312.825 3181.800 2605.600 3183.200 ;
        RECT 312.825 3180.480 2606.010 3181.800 ;
        RECT 314.400 3179.080 2606.010 3180.480 ;
        RECT 312.825 3116.560 2606.010 3179.080 ;
        RECT 312.825 3115.160 2605.600 3116.560 ;
        RECT 312.825 3109.080 2606.010 3115.160 ;
        RECT 314.400 3107.680 2606.010 3109.080 ;
        RECT 312.825 3049.920 2606.010 3107.680 ;
        RECT 312.825 3048.520 2605.600 3049.920 ;
        RECT 312.825 3037.680 2606.010 3048.520 ;
        RECT 314.400 3036.280 2606.010 3037.680 ;
        RECT 312.825 2983.280 2606.010 3036.280 ;
        RECT 312.825 2981.880 2605.600 2983.280 ;
        RECT 312.825 2966.280 2606.010 2981.880 ;
        RECT 314.400 2964.880 2606.010 2966.280 ;
        RECT 312.825 2916.640 2606.010 2964.880 ;
        RECT 312.825 2915.240 2605.600 2916.640 ;
        RECT 312.825 2894.880 2606.010 2915.240 ;
        RECT 314.400 2893.480 2606.010 2894.880 ;
        RECT 312.825 2850.000 2606.010 2893.480 ;
        RECT 312.825 2848.600 2605.600 2850.000 ;
        RECT 312.825 2823.480 2606.010 2848.600 ;
        RECT 314.400 2822.080 2606.010 2823.480 ;
        RECT 312.825 2783.360 2606.010 2822.080 ;
        RECT 312.825 2781.960 2605.600 2783.360 ;
        RECT 312.825 2752.080 2606.010 2781.960 ;
        RECT 314.400 2750.680 2606.010 2752.080 ;
        RECT 312.825 2716.720 2606.010 2750.680 ;
        RECT 312.825 2715.320 2605.600 2716.720 ;
        RECT 312.825 2680.680 2606.010 2715.320 ;
        RECT 314.400 2679.280 2606.010 2680.680 ;
        RECT 312.825 2650.080 2606.010 2679.280 ;
        RECT 312.825 2648.680 2605.600 2650.080 ;
        RECT 312.825 2609.280 2606.010 2648.680 ;
        RECT 314.400 2607.880 2606.010 2609.280 ;
        RECT 312.825 2583.440 2606.010 2607.880 ;
        RECT 312.825 2582.040 2605.600 2583.440 ;
        RECT 312.825 2537.880 2606.010 2582.040 ;
        RECT 314.400 2536.480 2606.010 2537.880 ;
        RECT 312.825 2516.800 2606.010 2536.480 ;
        RECT 312.825 2515.400 2605.600 2516.800 ;
        RECT 312.825 2466.480 2606.010 2515.400 ;
        RECT 314.400 2465.080 2606.010 2466.480 ;
        RECT 312.825 2450.160 2606.010 2465.080 ;
        RECT 312.825 2448.760 2605.600 2450.160 ;
        RECT 312.825 2395.080 2606.010 2448.760 ;
        RECT 314.400 2393.680 2606.010 2395.080 ;
        RECT 312.825 2383.520 2606.010 2393.680 ;
        RECT 312.825 2382.120 2605.600 2383.520 ;
        RECT 312.825 2323.680 2606.010 2382.120 ;
        RECT 314.400 2322.280 2606.010 2323.680 ;
        RECT 312.825 2316.880 2606.010 2322.280 ;
        RECT 312.825 2315.480 2605.600 2316.880 ;
        RECT 312.825 2252.280 2606.010 2315.480 ;
        RECT 314.400 2250.880 2606.010 2252.280 ;
        RECT 312.825 2250.240 2606.010 2250.880 ;
        RECT 312.825 2248.840 2605.600 2250.240 ;
        RECT 312.825 2183.600 2606.010 2248.840 ;
        RECT 312.825 2182.200 2605.600 2183.600 ;
        RECT 312.825 2180.880 2606.010 2182.200 ;
        RECT 314.400 2179.480 2606.010 2180.880 ;
        RECT 312.825 2116.960 2606.010 2179.480 ;
        RECT 312.825 2115.560 2605.600 2116.960 ;
        RECT 312.825 2109.480 2606.010 2115.560 ;
        RECT 314.400 2108.080 2606.010 2109.480 ;
        RECT 312.825 2050.320 2606.010 2108.080 ;
        RECT 312.825 2048.920 2605.600 2050.320 ;
        RECT 312.825 2038.080 2606.010 2048.920 ;
        RECT 314.400 2036.680 2606.010 2038.080 ;
        RECT 312.825 1983.680 2606.010 2036.680 ;
        RECT 312.825 1982.280 2605.600 1983.680 ;
        RECT 312.825 1966.680 2606.010 1982.280 ;
        RECT 314.400 1965.280 2606.010 1966.680 ;
        RECT 312.825 1917.040 2606.010 1965.280 ;
        RECT 312.825 1915.640 2605.600 1917.040 ;
        RECT 312.825 1895.280 2606.010 1915.640 ;
        RECT 314.400 1893.880 2606.010 1895.280 ;
        RECT 312.825 1850.400 2606.010 1893.880 ;
        RECT 312.825 1849.000 2605.600 1850.400 ;
        RECT 312.825 1823.880 2606.010 1849.000 ;
        RECT 314.400 1822.480 2606.010 1823.880 ;
        RECT 312.825 1783.760 2606.010 1822.480 ;
        RECT 312.825 1782.360 2605.600 1783.760 ;
        RECT 312.825 1752.480 2606.010 1782.360 ;
        RECT 314.400 1751.080 2606.010 1752.480 ;
        RECT 312.825 1716.440 2606.010 1751.080 ;
        RECT 312.825 1715.040 2605.600 1716.440 ;
        RECT 312.825 1680.400 2606.010 1715.040 ;
        RECT 314.400 1679.000 2606.010 1680.400 ;
        RECT 312.825 1649.800 2606.010 1679.000 ;
        RECT 312.825 1648.400 2605.600 1649.800 ;
        RECT 312.825 1609.000 2606.010 1648.400 ;
        RECT 314.400 1607.600 2606.010 1609.000 ;
        RECT 312.825 1583.160 2606.010 1607.600 ;
        RECT 312.825 1581.760 2605.600 1583.160 ;
        RECT 312.825 1537.600 2606.010 1581.760 ;
        RECT 314.400 1536.200 2606.010 1537.600 ;
        RECT 312.825 1516.520 2606.010 1536.200 ;
        RECT 312.825 1515.120 2605.600 1516.520 ;
        RECT 312.825 1466.200 2606.010 1515.120 ;
        RECT 314.400 1464.800 2606.010 1466.200 ;
        RECT 312.825 1449.880 2606.010 1464.800 ;
        RECT 312.825 1448.480 2605.600 1449.880 ;
        RECT 312.825 1394.800 2606.010 1448.480 ;
        RECT 314.400 1393.400 2606.010 1394.800 ;
        RECT 312.825 1383.240 2606.010 1393.400 ;
        RECT 312.825 1381.840 2605.600 1383.240 ;
        RECT 312.825 1323.400 2606.010 1381.840 ;
        RECT 314.400 1322.000 2606.010 1323.400 ;
        RECT 312.825 1316.600 2606.010 1322.000 ;
        RECT 312.825 1315.200 2605.600 1316.600 ;
        RECT 312.825 1252.000 2606.010 1315.200 ;
        RECT 314.400 1250.600 2606.010 1252.000 ;
        RECT 312.825 1249.960 2606.010 1250.600 ;
        RECT 312.825 1248.560 2605.600 1249.960 ;
        RECT 312.825 1183.320 2606.010 1248.560 ;
        RECT 312.825 1181.920 2605.600 1183.320 ;
        RECT 312.825 1180.600 2606.010 1181.920 ;
        RECT 314.400 1179.200 2606.010 1180.600 ;
        RECT 312.825 1116.680 2606.010 1179.200 ;
        RECT 312.825 1115.280 2605.600 1116.680 ;
        RECT 312.825 1109.200 2606.010 1115.280 ;
        RECT 314.400 1107.800 2606.010 1109.200 ;
        RECT 312.825 1050.040 2606.010 1107.800 ;
        RECT 312.825 1048.640 2605.600 1050.040 ;
        RECT 312.825 1037.800 2606.010 1048.640 ;
        RECT 314.400 1036.400 2606.010 1037.800 ;
        RECT 312.825 983.400 2606.010 1036.400 ;
        RECT 312.825 982.000 2605.600 983.400 ;
        RECT 312.825 966.400 2606.010 982.000 ;
        RECT 314.400 965.000 2606.010 966.400 ;
        RECT 312.825 916.760 2606.010 965.000 ;
        RECT 312.825 915.360 2605.600 916.760 ;
        RECT 312.825 895.000 2606.010 915.360 ;
        RECT 314.400 893.600 2606.010 895.000 ;
        RECT 312.825 850.120 2606.010 893.600 ;
        RECT 312.825 848.720 2605.600 850.120 ;
        RECT 312.825 823.600 2606.010 848.720 ;
        RECT 314.400 822.200 2606.010 823.600 ;
        RECT 312.825 783.480 2606.010 822.200 ;
        RECT 312.825 782.080 2605.600 783.480 ;
        RECT 312.825 752.200 2606.010 782.080 ;
        RECT 314.400 750.800 2606.010 752.200 ;
        RECT 312.825 716.840 2606.010 750.800 ;
        RECT 312.825 715.440 2605.600 716.840 ;
        RECT 312.825 680.800 2606.010 715.440 ;
        RECT 314.400 679.400 2606.010 680.800 ;
        RECT 312.825 650.200 2606.010 679.400 ;
        RECT 312.825 648.800 2605.600 650.200 ;
        RECT 312.825 609.400 2606.010 648.800 ;
        RECT 314.400 608.000 2606.010 609.400 ;
        RECT 312.825 583.560 2606.010 608.000 ;
        RECT 312.825 582.160 2605.600 583.560 ;
        RECT 312.825 538.000 2606.010 582.160 ;
        RECT 314.400 536.600 2606.010 538.000 ;
        RECT 312.825 516.920 2606.010 536.600 ;
        RECT 312.825 515.520 2605.600 516.920 ;
        RECT 312.825 466.600 2606.010 515.520 ;
        RECT 314.400 465.200 2606.010 466.600 ;
        RECT 312.825 450.280 2606.010 465.200 ;
        RECT 312.825 448.880 2605.600 450.280 ;
        RECT 312.825 395.200 2606.010 448.880 ;
        RECT 314.400 393.800 2606.010 395.200 ;
        RECT 312.825 383.640 2606.010 393.800 ;
        RECT 312.825 382.240 2605.600 383.640 ;
        RECT 312.825 323.800 2606.010 382.240 ;
        RECT 314.400 322.400 2606.010 323.800 ;
        RECT 312.825 317.000 2606.010 322.400 ;
        RECT 312.825 315.600 2605.600 317.000 ;
        RECT 312.825 252.400 2606.010 315.600 ;
        RECT 314.400 251.000 2606.010 252.400 ;
        RECT 312.825 250.360 2606.010 251.000 ;
        RECT 312.825 248.960 2605.600 250.360 ;
        RECT 312.825 226.715 2606.010 248.960 ;
      LAYER met4 ;
        RECT 326.855 226.640 330.640 3202.800 ;
        RECT 333.040 226.640 407.440 3202.800 ;
        RECT 409.840 226.640 2592.225 3202.800 ;
  END
END user_project_wrapper
END LIBRARY

