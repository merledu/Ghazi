magic
tech sky130A
magscale 1 2
timestamp 1608008999
<< locali >>
rect 8125 685899 8159 695453
rect 72525 683247 72559 692733
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72709 678895 72743 683077
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 72801 656931 72835 666485
rect 219081 656931 219115 666485
rect 427921 48331 427955 49181
rect 434821 48331 434855 49249
rect 427921 29019 427955 38573
rect 434821 29019 434855 38573
rect 328469 9707 328503 19261
rect 330033 9707 330067 18649
rect 394709 9707 394743 19261
rect 397469 9707 397503 19261
rect 427921 9707 427955 19261
rect 434821 9775 434855 19261
rect 376769 4811 376803 4913
rect 386337 4743 386371 4913
rect 422309 4879 422343 4981
rect 402989 4675 403023 4845
rect 386463 4641 386613 4675
rect 428197 4879 428231 4981
rect 406393 4675 406427 4845
rect 415409 4539 415443 4641
rect 424977 4539 425011 4709
rect 347513 3859 347547 4097
rect 326295 3553 326445 3587
rect 425069 2363 425103 4641
rect 431141 595 431175 9605
rect 435833 595 435867 9605
rect 442951 3689 443193 3723
rect 528569 3179 528603 3757
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 692733 72559 692767
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 72525 683213 72559 683247
rect 154313 685797 154347 685831
rect 72709 683077 72743 683111
rect 72709 678861 72743 678895
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 284033 676209 284067 676243
rect 72801 666485 72835 666519
rect 72801 656897 72835 656931
rect 219081 666485 219115 666519
rect 219081 656897 219115 656931
rect 434821 49249 434855 49283
rect 427921 49181 427955 49215
rect 427921 48297 427955 48331
rect 434821 48297 434855 48331
rect 427921 38573 427955 38607
rect 427921 28985 427955 29019
rect 434821 38573 434855 38607
rect 434821 28985 434855 29019
rect 328469 19261 328503 19295
rect 394709 19261 394743 19295
rect 328469 9673 328503 9707
rect 330033 18649 330067 18683
rect 330033 9673 330067 9707
rect 394709 9673 394743 9707
rect 397469 19261 397503 19295
rect 397469 9673 397503 9707
rect 427921 19261 427955 19295
rect 434821 19261 434855 19295
rect 434821 9741 434855 9775
rect 427921 9673 427955 9707
rect 431141 9605 431175 9639
rect 422309 4981 422343 5015
rect 376769 4913 376803 4947
rect 376769 4777 376803 4811
rect 386337 4913 386371 4947
rect 386337 4709 386371 4743
rect 402989 4845 403023 4879
rect 386429 4641 386463 4675
rect 386613 4641 386647 4675
rect 402989 4641 403023 4675
rect 406393 4845 406427 4879
rect 422309 4845 422343 4879
rect 428197 4981 428231 5015
rect 428197 4845 428231 4879
rect 424977 4709 425011 4743
rect 406393 4641 406427 4675
rect 415409 4641 415443 4675
rect 415409 4505 415443 4539
rect 424977 4505 425011 4539
rect 425069 4641 425103 4675
rect 347513 4097 347547 4131
rect 347513 3825 347547 3859
rect 326261 3553 326295 3587
rect 326445 3553 326479 3587
rect 425069 2329 425103 2363
rect 431141 561 431175 595
rect 435833 9605 435867 9639
rect 528569 3757 528603 3791
rect 442917 3689 442951 3723
rect 443193 3689 443227 3723
rect 528569 3145 528603 3179
rect 435833 561 435867 595
<< metal1 >>
rect 411162 700408 411168 700460
rect 411220 700448 411226 700460
rect 429838 700448 429844 700460
rect 411220 700420 429844 700448
rect 411220 700408 411226 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 463602 700408 463608 700460
rect 463660 700448 463666 700460
rect 494790 700448 494796 700460
rect 463660 700420 494796 700448
rect 463660 700408 463666 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 514662 700408 514668 700460
rect 514720 700448 514726 700460
rect 559650 700448 559656 700460
rect 514720 700420 559656 700448
rect 514720 700408 514726 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 394602 700340 394608 700392
rect 394660 700380 394666 700392
rect 413646 700380 413652 700392
rect 394660 700352 413652 700380
rect 394660 700340 394666 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 445662 700340 445668 700392
rect 445720 700380 445726 700392
rect 478506 700380 478512 700392
rect 445720 700352 478512 700380
rect 445720 700340 445726 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 496722 700340 496728 700392
rect 496780 700380 496786 700392
rect 543458 700380 543464 700392
rect 496780 700352 543464 700380
rect 496780 700340 496786 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 343542 700272 343548 700324
rect 343600 700312 343606 700324
rect 348786 700312 348792 700324
rect 343600 700284 348792 700312
rect 343600 700272 343606 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 378042 700272 378048 700324
rect 378100 700312 378106 700324
rect 397454 700312 397460 700324
rect 378100 700284 397460 700312
rect 378100 700272 378106 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 429102 700272 429108 700324
rect 429160 700312 429166 700324
rect 462314 700312 462320 700324
rect 429160 700284 462320 700312
rect 429160 700272 429166 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 480162 700272 480168 700324
rect 480220 700312 480226 700324
rect 527174 700312 527180 700324
rect 480220 700284 527180 700312
rect 480220 700272 480226 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 326982 699660 326988 699712
rect 327040 699700 327046 699712
rect 332502 699700 332508 699712
rect 327040 699672 332508 699700
rect 327040 699660 327046 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 360102 699660 360108 699712
rect 360160 699700 360166 699712
rect 364978 699700 364984 699712
rect 360160 699672 364984 699700
rect 360160 699660 360166 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 523770 696940 523776 696992
rect 523828 696980 523834 696992
rect 580166 696980 580172 696992
rect 523828 696952 580172 696980
rect 523828 696940 523834 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 692767 72571 692773
rect 72513 692733 72525 692767
rect 72559 692764 72571 692767
rect 72694 692764 72700 692776
rect 72559 692736 72700 692764
rect 72559 692733 72571 692736
rect 72513 692727 72571 692733
rect 72694 692724 72700 692736
rect 72752 692724 72758 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 523678 685856 523684 685908
rect 523736 685896 523742 685908
rect 580166 685896 580172 685908
rect 523736 685868 580172 685896
rect 523736 685856 523742 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 683244 72516 683256
rect 72471 683216 72516 683244
rect 72510 683204 72516 683216
rect 72568 683204 72574 683256
rect 72510 683068 72516 683120
rect 72568 683108 72574 683120
rect 72697 683111 72755 683117
rect 72697 683108 72709 683111
rect 72568 683080 72709 683108
rect 72568 683068 72574 683080
rect 72697 683077 72709 683080
rect 72743 683077 72755 683111
rect 72697 683071 72755 683077
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 219066 679028 219072 679040
rect 218992 679000 219072 679028
rect 218992 678972 219020 679000
rect 219066 678988 219072 679000
rect 219124 678988 219130 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 218974 678920 218980 678972
rect 219032 678920 219038 678972
rect 72694 678892 72700 678904
rect 72655 678864 72700 678892
rect 72694 678852 72700 678864
rect 72752 678852 72758 678904
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 72694 669264 72700 669316
rect 72752 669304 72758 669316
rect 72878 669304 72884 669316
rect 72752 669276 72884 669304
rect 72752 669264 72758 669276
rect 72878 669264 72884 669276
rect 72936 669264 72942 669316
rect 218974 669264 218980 669316
rect 219032 669304 219038 669316
rect 219158 669304 219164 669316
rect 219032 669276 219164 669304
rect 219032 669264 219038 669276
rect 219158 669264 219164 669276
rect 219216 669264 219222 669316
rect 72789 666519 72847 666525
rect 72789 666485 72801 666519
rect 72835 666516 72847 666519
rect 72878 666516 72884 666528
rect 72835 666488 72884 666516
rect 72835 666485 72847 666488
rect 72789 666479 72847 666485
rect 72878 666476 72884 666488
rect 72936 666476 72942 666528
rect 219069 666519 219127 666525
rect 219069 666485 219081 666519
rect 219115 666516 219127 666519
rect 219158 666516 219164 666528
rect 219115 666488 219164 666516
rect 219115 666485 219127 666488
rect 219069 666479 219127 666485
rect 219158 666476 219164 666488
rect 219216 666476 219222 666528
rect 72786 656928 72792 656940
rect 72747 656900 72792 656928
rect 72786 656888 72792 656900
rect 72844 656888 72850 656940
rect 219066 656928 219072 656940
rect 219027 656900 219072 656928
rect 219066 656888 219072 656900
rect 219124 656888 219130 656940
rect 377122 655460 377128 655512
rect 377180 655500 377186 655512
rect 378042 655500 378048 655512
rect 377180 655472 378048 655500
rect 377180 655460 377186 655472
rect 378042 655460 378048 655472
rect 378100 655460 378106 655512
rect 428182 655460 428188 655512
rect 428240 655500 428246 655512
rect 429102 655500 429108 655512
rect 428240 655472 429108 655500
rect 428240 655460 428246 655472
rect 429102 655460 429108 655472
rect 429160 655460 429166 655512
rect 462314 655460 462320 655512
rect 462372 655500 462378 655512
rect 463602 655500 463608 655512
rect 462372 655472 463608 655500
rect 462372 655460 462378 655472
rect 463602 655460 463608 655472
rect 463660 655460 463666 655512
rect 479334 655460 479340 655512
rect 479392 655500 479398 655512
rect 480162 655500 480168 655512
rect 479392 655472 480168 655500
rect 479392 655460 479398 655472
rect 480162 655460 480168 655472
rect 480220 655460 480226 655512
rect 513374 655256 513380 655308
rect 513432 655296 513438 655308
rect 514662 655296 514668 655308
rect 513432 655268 514668 655296
rect 513432 655256 513438 655268
rect 514662 655256 514668 655268
rect 514720 655256 514726 655308
rect 325970 655120 325976 655172
rect 326028 655160 326034 655172
rect 326982 655160 326988 655172
rect 326028 655132 326988 655160
rect 326028 655120 326034 655132
rect 326982 655120 326988 655132
rect 327040 655120 327046 655172
rect 8018 654916 8024 654968
rect 8076 654956 8082 654968
rect 70486 654956 70492 654968
rect 8076 654928 70492 654956
rect 8076 654916 8082 654928
rect 70486 654916 70492 654928
rect 70544 654916 70550 654968
rect 72786 654916 72792 654968
rect 72844 654956 72850 654968
rect 121546 654956 121552 654968
rect 72844 654928 121552 654956
rect 72844 654916 72850 654928
rect 121546 654916 121552 654928
rect 121604 654916 121610 654968
rect 137738 654916 137744 654968
rect 137796 654956 137802 654968
rect 172698 654956 172704 654968
rect 137796 654928 172704 654956
rect 137796 654916 137802 654928
rect 172698 654916 172704 654928
rect 172756 654916 172762 654968
rect 41322 654848 41328 654900
rect 41380 654888 41386 654900
rect 104526 654888 104532 654900
rect 41380 654860 104532 654888
rect 41380 654848 41386 654860
rect 104526 654848 104532 654860
rect 104584 654848 104590 654900
rect 106182 654848 106188 654900
rect 106240 654888 106246 654900
rect 155586 654888 155592 654900
rect 106240 654860 155592 654888
rect 106240 654848 106246 654860
rect 155586 654848 155592 654860
rect 155644 654848 155650 654900
rect 171042 654848 171048 654900
rect 171100 654888 171106 654900
rect 206738 654888 206744 654900
rect 171100 654860 206744 654888
rect 171100 654848 171106 654860
rect 206738 654848 206744 654860
rect 206796 654848 206802 654900
rect 219066 654848 219072 654900
rect 219124 654888 219130 654900
rect 240778 654888 240784 654900
rect 219124 654860 240784 654888
rect 219124 654848 219130 654860
rect 240778 654848 240784 654860
rect 240836 654848 240842 654900
rect 24762 654780 24768 654832
rect 24820 654820 24826 654832
rect 87506 654820 87512 654832
rect 24820 654792 87512 654820
rect 24820 654780 24826 654792
rect 87506 654780 87512 654792
rect 87564 654780 87570 654832
rect 89622 654780 89628 654832
rect 89680 654820 89686 654832
rect 138566 654820 138572 654832
rect 89680 654792 138572 654820
rect 89680 654780 89686 654792
rect 138566 654780 138572 654792
rect 138624 654780 138630 654832
rect 154298 654780 154304 654832
rect 154356 654820 154362 654832
rect 189718 654820 189724 654832
rect 154356 654792 189724 654820
rect 154356 654780 154362 654792
rect 189718 654780 189724 654792
rect 189776 654780 189782 654832
rect 202782 654780 202788 654832
rect 202840 654820 202846 654832
rect 223758 654820 223764 654832
rect 202840 654792 223764 654820
rect 202840 654780 202846 654792
rect 223758 654780 223764 654792
rect 223816 654780 223822 654832
rect 235902 654780 235908 654832
rect 235960 654820 235966 654832
rect 257890 654820 257896 654832
rect 235960 654792 257896 654820
rect 235960 654780 235966 654792
rect 257890 654780 257896 654792
rect 257948 654780 257954 654832
rect 267642 654780 267648 654832
rect 267700 654820 267706 654832
rect 274910 654820 274916 654832
rect 267700 654792 274916 654820
rect 267700 654780 267706 654792
rect 274910 654780 274916 654792
rect 274968 654780 274974 654832
rect 284018 654780 284024 654832
rect 284076 654820 284082 654832
rect 291930 654820 291936 654832
rect 284076 654792 291936 654820
rect 284076 654780 284082 654792
rect 291930 654780 291936 654792
rect 291988 654780 291994 654832
rect 300762 654100 300768 654152
rect 300820 654140 300826 654152
rect 308950 654140 308956 654152
rect 300820 654112 308956 654140
rect 300820 654100 300826 654112
rect 308950 654100 308956 654112
rect 309008 654100 309014 654152
rect 3602 645804 3608 645856
rect 3660 645844 3666 645856
rect 59354 645844 59360 645856
rect 3660 645816 59360 645844
rect 3660 645804 3666 645816
rect 59354 645804 59360 645816
rect 59412 645804 59418 645856
rect 523770 638936 523776 638988
rect 523828 638976 523834 638988
rect 580166 638976 580172 638988
rect 523828 638948 580172 638976
rect 523828 638936 523834 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 3418 630572 3424 630624
rect 3476 630612 3482 630624
rect 59354 630612 59360 630624
rect 3476 630584 59360 630612
rect 3476 630572 3482 630584
rect 59354 630572 59360 630584
rect 59412 630572 59418 630624
rect 524322 619556 524328 619608
rect 524380 619596 524386 619608
rect 580258 619596 580264 619608
rect 524380 619568 580264 619596
rect 524380 619556 524386 619568
rect 580258 619556 580264 619568
rect 580316 619556 580322 619608
rect 3510 616768 3516 616820
rect 3568 616808 3574 616820
rect 59354 616808 59360 616820
rect 3568 616780 59360 616808
rect 3568 616768 3574 616780
rect 59354 616768 59360 616780
rect 59412 616768 59418 616820
rect 523126 605752 523132 605804
rect 523184 605792 523190 605804
rect 580442 605792 580448 605804
rect 523184 605764 580448 605792
rect 523184 605752 523190 605764
rect 580442 605752 580448 605764
rect 580500 605752 580506 605804
rect 3602 603032 3608 603084
rect 3660 603072 3666 603084
rect 59354 603072 59360 603084
rect 3660 603044 59360 603072
rect 3660 603032 3666 603044
rect 59354 603032 59360 603044
rect 59412 603032 59418 603084
rect 523678 592016 523684 592068
rect 523736 592056 523742 592068
rect 579798 592056 579804 592068
rect 523736 592028 579804 592056
rect 523736 592016 523742 592028
rect 579798 592016 579804 592028
rect 579856 592016 579862 592068
rect 3418 587800 3424 587852
rect 3476 587840 3482 587852
rect 59354 587840 59360 587852
rect 3476 587812 59360 587840
rect 3476 587800 3482 587812
rect 59354 587800 59360 587812
rect 59412 587800 59418 587852
rect 524322 579572 524328 579624
rect 524380 579612 524386 579624
rect 580350 579612 580356 579624
rect 524380 579584 580356 579612
rect 524380 579572 524386 579584
rect 580350 579572 580356 579584
rect 580408 579572 580414 579624
rect 3510 573996 3516 574048
rect 3568 574036 3574 574048
rect 59354 574036 59360 574048
rect 3568 574008 59360 574036
rect 3568 573996 3574 574008
rect 59354 573996 59360 574008
rect 59412 573996 59418 574048
rect 523126 565768 523132 565820
rect 523184 565808 523190 565820
rect 580442 565808 580448 565820
rect 523184 565780 580448 565808
rect 523184 565768 523190 565780
rect 580442 565768 580448 565780
rect 580500 565768 580506 565820
rect 3418 560192 3424 560244
rect 3476 560232 3482 560244
rect 59354 560232 59360 560244
rect 3476 560204 59360 560232
rect 3476 560192 3482 560204
rect 59354 560192 59360 560204
rect 59412 560192 59418 560244
rect 523770 556180 523776 556232
rect 523828 556220 523834 556232
rect 580166 556220 580172 556232
rect 523828 556192 580172 556220
rect 523828 556180 523834 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 523494 545096 523500 545148
rect 523552 545136 523558 545148
rect 580166 545136 580172 545148
rect 523552 545108 580172 545136
rect 523552 545096 523558 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 3418 545028 3424 545080
rect 3476 545068 3482 545080
rect 59354 545068 59360 545080
rect 3476 545040 59360 545068
rect 3476 545028 3482 545040
rect 59354 545028 59360 545040
rect 59412 545028 59418 545080
rect 523678 539520 523684 539572
rect 523736 539560 523742 539572
rect 580258 539560 580264 539572
rect 523736 539532 580264 539560
rect 523736 539520 523742 539532
rect 580258 539520 580264 539532
rect 580316 539520 580322 539572
rect 3418 531224 3424 531276
rect 3476 531264 3482 531276
rect 59354 531264 59360 531276
rect 3476 531236 59360 531264
rect 3476 531224 3482 531236
rect 59354 531224 59360 531236
rect 59412 531224 59418 531276
rect 3418 516128 3424 516180
rect 3476 516168 3482 516180
rect 59354 516168 59360 516180
rect 3476 516140 59360 516168
rect 3476 516128 3482 516140
rect 59354 516128 59360 516140
rect 59412 516128 59418 516180
rect 523770 509260 523776 509312
rect 523828 509300 523834 509312
rect 580166 509300 580172 509312
rect 523828 509272 580172 509300
rect 523828 509260 523834 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 59354 501004 59360 501016
rect 3384 500976 59360 501004
rect 3384 500964 3390 500976
rect 59354 500964 59360 500976
rect 59412 500964 59418 501016
rect 523678 499468 523684 499520
rect 523736 499508 523742 499520
rect 580258 499508 580264 499520
rect 523736 499480 580264 499508
rect 523736 499468 523742 499480
rect 580258 499468 580264 499480
rect 580316 499468 580322 499520
rect 523678 498176 523684 498228
rect 523736 498216 523742 498228
rect 580166 498216 580172 498228
rect 523736 498188 580172 498216
rect 523736 498176 523742 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3418 487160 3424 487212
rect 3476 487200 3482 487212
rect 59354 487200 59360 487212
rect 3476 487172 59360 487200
rect 3476 487160 3482 487172
rect 59354 487160 59360 487172
rect 59412 487160 59418 487212
rect 3418 473356 3424 473408
rect 3476 473396 3482 473408
rect 59354 473396 59360 473408
rect 3476 473368 59360 473396
rect 3476 473356 3482 473368
rect 59354 473356 59360 473368
rect 59412 473356 59418 473408
rect 523678 462340 523684 462392
rect 523736 462380 523742 462392
rect 580166 462380 580172 462392
rect 523736 462352 580172 462380
rect 523736 462340 523742 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 524322 459484 524328 459536
rect 524380 459524 524386 459536
rect 580258 459524 580264 459536
rect 524380 459496 580264 459524
rect 524380 459484 524386 459496
rect 580258 459484 580264 459496
rect 580316 459484 580322 459536
rect 3510 458192 3516 458244
rect 3568 458232 3574 458244
rect 59354 458232 59360 458244
rect 3568 458204 59360 458232
rect 3568 458192 3574 458204
rect 59354 458192 59360 458204
rect 59412 458192 59418 458244
rect 523770 451256 523776 451308
rect 523828 451296 523834 451308
rect 580166 451296 580172 451308
rect 523828 451268 580172 451296
rect 523828 451256 523834 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 3418 444388 3424 444440
rect 3476 444428 3482 444440
rect 59354 444428 59360 444440
rect 3476 444400 59360 444428
rect 3476 444388 3482 444400
rect 59354 444388 59360 444400
rect 59412 444388 59418 444440
rect 523678 438880 523684 438932
rect 523736 438920 523742 438932
rect 580166 438920 580172 438932
rect 523736 438892 580172 438920
rect 523736 438880 523742 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3510 429156 3516 429208
rect 3568 429196 3574 429208
rect 59354 429196 59360 429208
rect 3568 429168 59360 429196
rect 3568 429156 3574 429168
rect 59354 429156 59360 429168
rect 59412 429156 59418 429208
rect 3418 415420 3424 415472
rect 3476 415460 3482 415472
rect 59354 415460 59360 415472
rect 3476 415432 59360 415460
rect 3476 415420 3482 415432
rect 59354 415420 59360 415432
rect 59412 415420 59418 415472
rect 523678 415420 523684 415472
rect 523736 415460 523742 415472
rect 580166 415460 580172 415472
rect 523736 415432 580172 415460
rect 523736 415420 523742 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 523770 404336 523776 404388
rect 523828 404376 523834 404388
rect 580166 404376 580172 404388
rect 523828 404348 580172 404376
rect 523828 404336 523834 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3602 401616 3608 401668
rect 3660 401656 3666 401668
rect 59354 401656 59360 401668
rect 3660 401628 59360 401656
rect 3660 401616 3666 401628
rect 59354 401616 59360 401628
rect 59412 401616 59418 401668
rect 523678 391960 523684 392012
rect 523736 392000 523742 392012
rect 580166 392000 580172 392012
rect 523736 391972 580172 392000
rect 523736 391960 523742 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 3510 372580 3516 372632
rect 3568 372620 3574 372632
rect 59354 372620 59360 372632
rect 3568 372592 59360 372620
rect 3568 372580 3574 372592
rect 59354 372580 59360 372592
rect 59412 372580 59418 372632
rect 524230 368500 524236 368552
rect 524288 368540 524294 368552
rect 580166 368540 580172 368552
rect 524288 368512 580172 368540
rect 524288 368500 524294 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 3418 358776 3424 358828
rect 3476 358816 3482 358828
rect 59354 358816 59360 358828
rect 3476 358788 59360 358816
rect 3476 358776 3482 358788
rect 59354 358776 59360 358788
rect 59412 358776 59418 358828
rect 523678 357416 523684 357468
rect 523736 357456 523742 357468
rect 580166 357456 580172 357468
rect 523736 357428 580172 357456
rect 523736 357416 523742 357428
rect 580166 357416 580172 357428
rect 580224 357416 580230 357468
rect 523770 345040 523776 345092
rect 523828 345080 523834 345092
rect 580166 345080 580172 345092
rect 523828 345052 580172 345080
rect 523828 345040 523834 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 3602 338036 3608 338088
rect 3660 338076 3666 338088
rect 59998 338076 60004 338088
rect 3660 338048 60004 338076
rect 3660 338036 3666 338048
rect 59998 338036 60004 338048
rect 60056 338036 60062 338088
rect 3602 329808 3608 329860
rect 3660 329848 3666 329860
rect 59354 329848 59360 329860
rect 3660 329820 59360 329848
rect 3660 329808 3666 329820
rect 59354 329808 59360 329820
rect 59412 329808 59418 329860
rect 524322 322872 524328 322924
rect 524380 322912 524386 322924
rect 580166 322912 580172 322924
rect 524380 322884 580172 322912
rect 524380 322872 524386 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 3694 316004 3700 316056
rect 3752 316044 3758 316056
rect 59354 316044 59360 316056
rect 3752 316016 59360 316044
rect 3752 316004 3758 316016
rect 59354 316004 59360 316016
rect 59412 316004 59418 316056
rect 524322 311788 524328 311840
rect 524380 311828 524386 311840
rect 580166 311828 580172 311840
rect 524380 311800 580172 311828
rect 524380 311788 524386 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 524322 298732 524328 298784
rect 524380 298772 524386 298784
rect 580166 298772 580172 298784
rect 524380 298744 580172 298772
rect 524380 298732 524386 298744
rect 580166 298732 580172 298744
rect 580224 298732 580230 298784
rect 3050 295264 3056 295316
rect 3108 295304 3114 295316
rect 60182 295304 60188 295316
rect 3108 295276 60188 295304
rect 3108 295264 3114 295276
rect 60182 295264 60188 295276
rect 60240 295264 60246 295316
rect 3510 287036 3516 287088
rect 3568 287076 3574 287088
rect 59354 287076 59360 287088
rect 3568 287048 59360 287076
rect 3568 287036 3574 287048
rect 59354 287036 59360 287048
rect 59412 287036 59418 287088
rect 523678 275952 523684 276004
rect 523736 275992 523742 276004
rect 580166 275992 580172 276004
rect 523736 275964 580172 275992
rect 523736 275952 523742 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 3602 273232 3608 273284
rect 3660 273272 3666 273284
rect 59354 273272 59360 273284
rect 3660 273244 59360 273272
rect 3660 273232 3666 273244
rect 59354 273232 59360 273244
rect 59412 273232 59418 273284
rect 523678 264868 523684 264920
rect 523736 264908 523742 264920
rect 580166 264908 580172 264920
rect 523736 264880 580172 264908
rect 523736 264868 523742 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 3142 252492 3148 252544
rect 3200 252532 3206 252544
rect 60090 252532 60096 252544
rect 3200 252504 60096 252532
rect 3200 252492 3206 252504
rect 60090 252492 60096 252504
rect 60148 252492 60154 252544
rect 523678 252492 523684 252544
rect 523736 252532 523742 252544
rect 579798 252532 579804 252544
rect 523736 252504 579804 252532
rect 523736 252492 523742 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 3418 244264 3424 244316
rect 3476 244304 3482 244316
rect 59354 244304 59360 244316
rect 3476 244276 59360 244304
rect 3476 244264 3482 244276
rect 59354 244264 59360 244276
rect 59412 244264 59418 244316
rect 3694 229100 3700 229152
rect 3752 229140 3758 229152
rect 59354 229140 59360 229152
rect 3752 229112 59360 229140
rect 3752 229100 3758 229112
rect 59354 229100 59360 229112
rect 59412 229100 59418 229152
rect 523678 229032 523684 229084
rect 523736 229072 523742 229084
rect 580166 229072 580172 229084
rect 523736 229044 580172 229072
rect 523736 229032 523742 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 523770 217948 523776 218000
rect 523828 217988 523834 218000
rect 580166 217988 580172 218000
rect 523828 217960 580172 217988
rect 523828 217948 523834 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 3142 208292 3148 208344
rect 3200 208332 3206 208344
rect 59998 208332 60004 208344
rect 3200 208304 60004 208332
rect 3200 208292 3206 208304
rect 59998 208292 60004 208304
rect 60056 208292 60062 208344
rect 523862 205572 523868 205624
rect 523920 205612 523926 205624
rect 579798 205612 579804 205624
rect 523920 205584 579804 205612
rect 523920 205572 523926 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 3510 201492 3516 201544
rect 3568 201532 3574 201544
rect 59354 201532 59360 201544
rect 3568 201504 59360 201532
rect 3568 201492 3574 201504
rect 59354 201492 59360 201504
rect 59412 201492 59418 201544
rect 3602 186328 3608 186380
rect 3660 186368 3666 186380
rect 59354 186368 59360 186380
rect 3660 186340 59360 186368
rect 3660 186328 3666 186340
rect 59354 186328 59360 186340
rect 59412 186328 59418 186380
rect 523678 182112 523684 182164
rect 523736 182152 523742 182164
rect 580166 182152 580172 182164
rect 523736 182124 580172 182152
rect 523736 182112 523742 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 523770 171028 523776 171080
rect 523828 171068 523834 171080
rect 580166 171068 580172 171080
rect 523828 171040 580172 171068
rect 523828 171028 523834 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 3418 165520 3424 165572
rect 3476 165560 3482 165572
rect 60090 165560 60096 165572
rect 3476 165532 60096 165560
rect 3476 165520 3482 165532
rect 60090 165520 60096 165532
rect 60148 165520 60154 165572
rect 3418 158720 3424 158772
rect 3476 158760 3482 158772
rect 59354 158760 59360 158772
rect 3476 158732 59360 158760
rect 3476 158720 3482 158732
rect 59354 158720 59360 158732
rect 59412 158720 59418 158772
rect 523862 158652 523868 158704
rect 523920 158692 523926 158704
rect 579798 158692 579804 158704
rect 523920 158664 579804 158692
rect 523920 158652 523926 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 3694 143556 3700 143608
rect 3752 143596 3758 143608
rect 59354 143596 59360 143608
rect 3752 143568 59360 143596
rect 3752 143556 3758 143568
rect 59354 143556 59360 143568
rect 59412 143556 59418 143608
rect 523678 135192 523684 135244
rect 523736 135232 523742 135244
rect 580166 135232 580172 135244
rect 523736 135204 580172 135232
rect 523736 135192 523742 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 523770 124108 523776 124160
rect 523828 124148 523834 124160
rect 580166 124148 580172 124160
rect 523828 124120 580172 124148
rect 523828 124108 523834 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 2958 122748 2964 122800
rect 3016 122788 3022 122800
rect 59998 122788 60004 122800
rect 3016 122760 60004 122788
rect 3016 122748 3022 122760
rect 59998 122748 60004 122760
rect 60056 122748 60062 122800
rect 3510 115948 3516 116000
rect 3568 115988 3574 116000
rect 59354 115988 59360 116000
rect 3568 115960 59360 115988
rect 3568 115948 3574 115960
rect 59354 115948 59360 115960
rect 59412 115948 59418 116000
rect 523862 111732 523868 111784
rect 523920 111772 523926 111784
rect 579798 111772 579804 111784
rect 523920 111744 579804 111772
rect 523920 111732 523926 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3602 100716 3608 100768
rect 3660 100756 3666 100768
rect 59354 100756 59360 100768
rect 3660 100728 59360 100756
rect 3660 100716 3666 100728
rect 59354 100716 59360 100728
rect 59412 100716 59418 100768
rect 523678 88272 523684 88324
rect 523736 88312 523742 88324
rect 580166 88312 580172 88324
rect 523736 88284 580172 88312
rect 523736 88272 523742 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 3050 79976 3056 80028
rect 3108 80016 3114 80028
rect 60090 80016 60096 80028
rect 3108 79988 60096 80016
rect 3108 79976 3114 79988
rect 60090 79976 60096 79988
rect 60148 79976 60154 80028
rect 523770 77188 523776 77240
rect 523828 77228 523834 77240
rect 580166 77228 580172 77240
rect 523828 77200 580172 77228
rect 523828 77188 523834 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 3418 73176 3424 73228
rect 3476 73216 3482 73228
rect 59354 73216 59360 73228
rect 3476 73188 59360 73216
rect 3476 73176 3482 73188
rect 59354 73176 59360 73188
rect 59412 73176 59418 73228
rect 523862 64812 523868 64864
rect 523920 64852 523926 64864
rect 579798 64852 579804 64864
rect 523920 64824 579804 64852
rect 523920 64812 523926 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 3510 57944 3516 57996
rect 3568 57984 3574 57996
rect 59354 57984 59360 57996
rect 3568 57956 59360 57984
rect 3568 57944 3574 57956
rect 59354 57944 59360 57956
rect 59412 57944 59418 57996
rect 477218 49648 477224 49700
rect 477276 49688 477282 49700
rect 482278 49688 482284 49700
rect 477276 49660 482284 49688
rect 477276 49648 477282 49660
rect 482278 49648 482284 49660
rect 482336 49648 482342 49700
rect 167362 49444 167368 49496
rect 167420 49484 167426 49496
rect 227898 49484 227904 49496
rect 167420 49456 227904 49484
rect 167420 49444 167426 49456
rect 227898 49444 227904 49456
rect 227956 49444 227962 49496
rect 110230 49376 110236 49428
rect 110288 49416 110294 49428
rect 171226 49416 171232 49428
rect 110288 49388 171232 49416
rect 110288 49376 110294 49388
rect 171226 49376 171232 49388
rect 171284 49376 171290 49428
rect 396166 49376 396172 49428
rect 396224 49416 396230 49428
rect 456886 49416 456892 49428
rect 396224 49388 456892 49416
rect 396224 49376 396230 49388
rect 456886 49376 456892 49388
rect 456944 49376 456950 49428
rect 88702 49308 88708 49360
rect 88760 49348 88766 49360
rect 150618 49348 150624 49360
rect 88760 49320 150624 49348
rect 88760 49308 88766 49320
rect 150618 49308 150624 49320
rect 150676 49308 150682 49360
rect 188890 49308 188896 49360
rect 188948 49348 188954 49360
rect 249886 49348 249892 49360
rect 188948 49320 249892 49348
rect 188948 49308 188954 49320
rect 249886 49308 249892 49320
rect 249944 49308 249950 49360
rect 403342 49308 403348 49360
rect 403400 49348 403406 49360
rect 463786 49348 463792 49360
rect 403400 49320 463792 49348
rect 403400 49308 403406 49320
rect 463786 49308 463792 49320
rect 463844 49308 463850 49360
rect 103054 49240 103060 49292
rect 103112 49280 103118 49292
rect 164326 49280 164332 49292
rect 103112 49252 164332 49280
rect 103112 49240 103118 49252
rect 164326 49240 164332 49252
rect 164384 49240 164390 49292
rect 174538 49240 174544 49292
rect 174596 49280 174602 49292
rect 236178 49280 236184 49292
rect 174596 49252 236184 49280
rect 174596 49240 174602 49252
rect 236178 49240 236184 49252
rect 236236 49240 236242 49292
rect 253198 49240 253204 49292
rect 253256 49280 253262 49292
rect 313458 49280 313464 49292
rect 253256 49252 313464 49280
rect 253256 49240 253262 49252
rect 313458 49240 313464 49252
rect 313516 49240 313522 49292
rect 374730 49240 374736 49292
rect 374788 49280 374794 49292
rect 434809 49283 434867 49289
rect 434809 49280 434821 49283
rect 374788 49252 434821 49280
rect 374788 49240 374794 49252
rect 434809 49249 434821 49252
rect 434855 49249 434867 49283
rect 434809 49243 434867 49249
rect 81618 49172 81624 49224
rect 81676 49212 81682 49224
rect 142246 49212 142252 49224
rect 81676 49184 142252 49212
rect 81676 49172 81682 49184
rect 142246 49172 142252 49184
rect 142304 49172 142310 49224
rect 145926 49172 145932 49224
rect 145984 49212 145990 49224
rect 207106 49212 207112 49224
rect 145984 49184 207112 49212
rect 145984 49172 145990 49184
rect 207106 49172 207112 49184
rect 207164 49172 207170 49224
rect 210326 49172 210332 49224
rect 210384 49212 210390 49224
rect 270494 49212 270500 49224
rect 210384 49184 270500 49212
rect 210384 49172 210390 49184
rect 270494 49172 270500 49184
rect 270552 49172 270558 49224
rect 367646 49172 367652 49224
rect 367704 49212 367710 49224
rect 427909 49215 427967 49221
rect 427909 49212 427921 49215
rect 367704 49184 427921 49212
rect 367704 49172 367710 49184
rect 427909 49181 427921 49184
rect 427955 49181 427967 49215
rect 427909 49175 427967 49181
rect 474826 49172 474832 49224
rect 474884 49212 474890 49224
rect 535454 49212 535460 49224
rect 474884 49184 535460 49212
rect 474884 49172 474890 49184
rect 535454 49172 535460 49184
rect 535512 49172 535518 49224
rect 74442 49104 74448 49156
rect 74500 49144 74506 49156
rect 135438 49144 135444 49156
rect 74500 49116 135444 49144
rect 74500 49104 74506 49116
rect 135438 49104 135444 49116
rect 135496 49104 135502 49156
rect 138842 49104 138848 49156
rect 138900 49144 138906 49156
rect 200206 49144 200212 49156
rect 138900 49116 200212 49144
rect 138900 49104 138906 49116
rect 200206 49104 200212 49116
rect 200264 49104 200270 49156
rect 224586 49104 224592 49156
rect 224644 49144 224650 49156
rect 285766 49144 285772 49156
rect 224644 49116 285772 49144
rect 224644 49104 224650 49116
rect 285766 49104 285772 49116
rect 285824 49104 285830 49156
rect 311618 49104 311624 49156
rect 311676 49144 311682 49156
rect 345658 49144 345664 49156
rect 311676 49116 345664 49144
rect 311676 49104 311682 49116
rect 345658 49104 345664 49116
rect 345716 49104 345722 49156
rect 389082 49104 389088 49156
rect 389140 49144 389146 49156
rect 449986 49144 449992 49156
rect 389140 49116 449992 49144
rect 389140 49104 389146 49116
rect 449986 49104 449992 49116
rect 450044 49104 450050 49156
rect 482002 49104 482008 49156
rect 482060 49144 482066 49156
rect 542354 49144 542360 49156
rect 482060 49116 542360 49144
rect 482060 49104 482066 49116
rect 542354 49104 542360 49116
rect 542412 49104 542418 49156
rect 67266 49036 67272 49088
rect 67324 49076 67330 49088
rect 128446 49076 128452 49088
rect 67324 49048 128452 49076
rect 67324 49036 67330 49048
rect 128446 49036 128452 49048
rect 128504 49036 128510 49088
rect 131666 49036 131672 49088
rect 131724 49076 131730 49088
rect 193398 49076 193404 49088
rect 131724 49048 193404 49076
rect 131724 49036 131730 49048
rect 193398 49036 193404 49048
rect 193456 49036 193462 49088
rect 217410 49036 217416 49088
rect 217468 49076 217474 49088
rect 278958 49076 278964 49088
rect 217468 49048 278964 49076
rect 217468 49036 217474 49048
rect 278958 49036 278964 49048
rect 279016 49036 279022 49088
rect 346118 49036 346124 49088
rect 346176 49076 346182 49088
rect 407206 49076 407212 49088
rect 346176 49048 407212 49076
rect 346176 49036 346182 49048
rect 407206 49036 407212 49048
rect 407264 49036 407270 49088
rect 489178 49036 489184 49088
rect 489236 49076 489242 49088
rect 549254 49076 549260 49088
rect 489236 49048 549260 49076
rect 489236 49036 489242 49048
rect 549254 49036 549260 49048
rect 549312 49036 549318 49088
rect 95878 48968 95884 49020
rect 95936 49008 95942 49020
rect 157426 49008 157432 49020
rect 95936 48980 157432 49008
rect 95936 48968 95942 48980
rect 157426 48968 157432 48980
rect 157484 48968 157490 49020
rect 181714 48968 181720 49020
rect 181772 49008 181778 49020
rect 242986 49008 242992 49020
rect 181772 48980 242992 49008
rect 181772 48968 181778 48980
rect 242986 48968 242992 48980
rect 243044 48968 243050 49020
rect 260374 48968 260380 49020
rect 260432 49008 260438 49020
rect 321738 49008 321744 49020
rect 260432 48980 321744 49008
rect 260432 48968 260438 48980
rect 321738 48968 321744 48980
rect 321796 48968 321802 49020
rect 354490 48968 354496 49020
rect 354548 49008 354554 49020
rect 367738 49008 367744 49020
rect 354548 48980 367744 49008
rect 354548 48968 354554 48980
rect 367738 48968 367744 48980
rect 367796 48968 367802 49020
rect 381906 48968 381912 49020
rect 381964 49008 381970 49020
rect 443178 49008 443184 49020
rect 381964 48980 443184 49008
rect 381964 48968 381970 48980
rect 443178 48968 443184 48980
rect 443236 48968 443242 49020
rect 467742 48968 467748 49020
rect 467800 49008 467806 49020
rect 528554 49008 528560 49020
rect 467800 48980 528560 49008
rect 467800 48968 467806 48980
rect 528554 48968 528560 48980
rect 528612 48968 528618 49020
rect 66070 48764 66076 48816
rect 66128 48804 66134 48816
rect 66898 48804 66904 48816
rect 66128 48776 66904 48804
rect 66128 48764 66134 48776
rect 66898 48764 66904 48776
rect 66956 48764 66962 48816
rect 70854 48764 70860 48816
rect 70912 48804 70918 48816
rect 71682 48804 71688 48816
rect 70912 48776 71688 48804
rect 70912 48764 70918 48776
rect 71682 48764 71688 48776
rect 71740 48764 71746 48816
rect 72050 48764 72056 48816
rect 72108 48804 72114 48816
rect 73062 48804 73068 48816
rect 72108 48776 73068 48804
rect 72108 48764 72114 48776
rect 73062 48764 73068 48776
rect 73120 48764 73126 48816
rect 73246 48764 73252 48816
rect 73304 48804 73310 48816
rect 74442 48804 74448 48816
rect 73304 48776 74448 48804
rect 73304 48764 73310 48776
rect 74442 48764 74448 48776
rect 74500 48764 74506 48816
rect 80422 48764 80428 48816
rect 80480 48804 80486 48816
rect 81342 48804 81348 48816
rect 80480 48776 81348 48804
rect 80480 48764 80486 48776
rect 81342 48764 81348 48776
rect 81400 48764 81406 48816
rect 89898 48764 89904 48816
rect 89956 48804 89962 48816
rect 91002 48804 91008 48816
rect 89956 48776 91008 48804
rect 89956 48764 89962 48776
rect 91002 48764 91008 48776
rect 91060 48764 91066 48816
rect 91094 48764 91100 48816
rect 91152 48804 91158 48816
rect 92290 48804 92296 48816
rect 91152 48776 92296 48804
rect 91152 48764 91158 48776
rect 92290 48764 92296 48776
rect 92348 48764 92354 48816
rect 97074 48764 97080 48816
rect 97132 48804 97138 48816
rect 97902 48804 97908 48816
rect 97132 48776 97908 48804
rect 97132 48764 97138 48776
rect 97902 48764 97908 48776
rect 97960 48764 97966 48816
rect 98270 48764 98276 48816
rect 98328 48804 98334 48816
rect 99282 48804 99288 48816
rect 98328 48776 99288 48804
rect 98328 48764 98334 48776
rect 99282 48764 99288 48776
rect 99340 48764 99346 48816
rect 99466 48764 99472 48816
rect 99524 48804 99530 48816
rect 100662 48804 100668 48816
rect 99524 48776 100668 48804
rect 99524 48764 99530 48776
rect 100662 48764 100668 48776
rect 100720 48764 100726 48816
rect 105446 48764 105452 48816
rect 105504 48804 105510 48816
rect 106182 48804 106188 48816
rect 105504 48776 106188 48804
rect 105504 48764 105510 48776
rect 106182 48764 106188 48776
rect 106240 48764 106246 48816
rect 106642 48764 106648 48816
rect 106700 48804 106706 48816
rect 107562 48804 107568 48816
rect 106700 48776 107568 48804
rect 106700 48764 106706 48776
rect 107562 48764 107568 48776
rect 107620 48764 107626 48816
rect 107838 48764 107844 48816
rect 107896 48804 107902 48816
rect 108942 48804 108948 48816
rect 107896 48776 108948 48804
rect 107896 48764 107902 48776
rect 108942 48764 108948 48776
rect 109000 48764 109006 48816
rect 109034 48764 109040 48816
rect 109092 48804 109098 48816
rect 110322 48804 110328 48816
rect 109092 48776 110328 48804
rect 109092 48764 109098 48776
rect 110322 48764 110328 48776
rect 110380 48764 110386 48816
rect 113726 48764 113732 48816
rect 113784 48804 113790 48816
rect 114462 48804 114468 48816
rect 113784 48776 114468 48804
rect 113784 48764 113790 48776
rect 114462 48764 114468 48776
rect 114520 48764 114526 48816
rect 114922 48764 114928 48816
rect 114980 48804 114986 48816
rect 115842 48804 115848 48816
rect 114980 48776 115848 48804
rect 114980 48764 114986 48776
rect 115842 48764 115848 48776
rect 115900 48764 115906 48816
rect 116118 48764 116124 48816
rect 116176 48804 116182 48816
rect 117222 48804 117228 48816
rect 116176 48776 117228 48804
rect 116176 48764 116182 48776
rect 117222 48764 117228 48776
rect 117280 48764 117286 48816
rect 117314 48764 117320 48816
rect 117372 48804 117378 48816
rect 118602 48804 118608 48816
rect 117372 48776 118608 48804
rect 117372 48764 117378 48776
rect 118602 48764 118608 48776
rect 118660 48764 118666 48816
rect 123294 48764 123300 48816
rect 123352 48804 123358 48816
rect 124122 48804 124128 48816
rect 123352 48776 124128 48804
rect 123352 48764 123358 48776
rect 124122 48764 124128 48776
rect 124180 48764 124186 48816
rect 124490 48764 124496 48816
rect 124548 48804 124554 48816
rect 125502 48804 125508 48816
rect 124548 48776 125508 48804
rect 124548 48764 124554 48776
rect 125502 48764 125508 48776
rect 125560 48764 125566 48816
rect 132862 48764 132868 48816
rect 132920 48804 132926 48816
rect 133782 48804 133788 48816
rect 132920 48776 133788 48804
rect 132920 48764 132926 48776
rect 133782 48764 133788 48776
rect 133840 48764 133846 48816
rect 134058 48764 134064 48816
rect 134116 48804 134122 48816
rect 135162 48804 135168 48816
rect 134116 48776 135168 48804
rect 134116 48764 134122 48776
rect 135162 48764 135168 48776
rect 135220 48764 135226 48816
rect 141142 48764 141148 48816
rect 141200 48804 141206 48816
rect 142062 48804 142068 48816
rect 141200 48776 142068 48804
rect 141200 48764 141206 48776
rect 142062 48764 142068 48776
rect 142120 48764 142126 48816
rect 142338 48764 142344 48816
rect 142396 48804 142402 48816
rect 143442 48804 143448 48816
rect 142396 48776 143448 48804
rect 142396 48764 142402 48776
rect 143442 48764 143448 48776
rect 143500 48764 143506 48816
rect 149514 48764 149520 48816
rect 149572 48804 149578 48816
rect 150342 48804 150348 48816
rect 149572 48776 150348 48804
rect 149572 48764 149578 48776
rect 150342 48764 150348 48776
rect 150400 48764 150406 48816
rect 150710 48764 150716 48816
rect 150768 48804 150774 48816
rect 151722 48804 151728 48816
rect 150768 48776 151728 48804
rect 150768 48764 150774 48776
rect 151722 48764 151728 48776
rect 151780 48764 151786 48816
rect 151906 48764 151912 48816
rect 151964 48804 151970 48816
rect 153010 48804 153016 48816
rect 151964 48776 153016 48804
rect 151964 48764 151970 48776
rect 153010 48764 153016 48776
rect 153068 48764 153074 48816
rect 157886 48764 157892 48816
rect 157944 48804 157950 48816
rect 158622 48804 158628 48816
rect 157944 48776 158628 48804
rect 157944 48764 157950 48776
rect 158622 48764 158628 48776
rect 158680 48764 158686 48816
rect 159082 48764 159088 48816
rect 159140 48804 159146 48816
rect 160002 48804 160008 48816
rect 159140 48776 160008 48804
rect 159140 48764 159146 48776
rect 160002 48764 160008 48776
rect 160060 48764 160066 48816
rect 160278 48764 160284 48816
rect 160336 48804 160342 48816
rect 161382 48804 161388 48816
rect 160336 48776 161388 48804
rect 160336 48764 160342 48776
rect 161382 48764 161388 48776
rect 161440 48764 161446 48816
rect 161474 48764 161480 48816
rect 161532 48804 161538 48816
rect 162762 48804 162768 48816
rect 161532 48776 162768 48804
rect 161532 48764 161538 48776
rect 162762 48764 162768 48776
rect 162820 48764 162826 48816
rect 168558 48764 168564 48816
rect 168616 48804 168622 48816
rect 169662 48804 169668 48816
rect 168616 48776 169668 48804
rect 168616 48764 168622 48776
rect 169662 48764 169668 48776
rect 169720 48764 169726 48816
rect 169754 48764 169760 48816
rect 169812 48804 169818 48816
rect 170950 48804 170956 48816
rect 169812 48776 170956 48804
rect 169812 48764 169818 48776
rect 170950 48764 170956 48776
rect 171008 48764 171014 48816
rect 175734 48764 175740 48816
rect 175792 48804 175798 48816
rect 176562 48804 176568 48816
rect 175792 48776 176568 48804
rect 175792 48764 175798 48776
rect 176562 48764 176568 48776
rect 176620 48764 176626 48816
rect 176930 48764 176936 48816
rect 176988 48804 176994 48816
rect 177942 48804 177948 48816
rect 176988 48776 177948 48804
rect 176988 48764 176994 48776
rect 177942 48764 177948 48776
rect 178000 48764 178006 48816
rect 178126 48764 178132 48816
rect 178184 48804 178190 48816
rect 179322 48804 179328 48816
rect 178184 48776 179328 48804
rect 178184 48764 178190 48776
rect 179322 48764 179328 48776
rect 179380 48764 179386 48816
rect 185302 48764 185308 48816
rect 185360 48804 185366 48816
rect 186222 48804 186228 48816
rect 185360 48776 186228 48804
rect 185360 48764 185366 48776
rect 186222 48764 186228 48776
rect 186280 48764 186286 48816
rect 186498 48764 186504 48816
rect 186556 48804 186562 48816
rect 187602 48804 187608 48816
rect 186556 48776 187608 48804
rect 186556 48764 186562 48776
rect 187602 48764 187608 48776
rect 187660 48764 187666 48816
rect 187694 48764 187700 48816
rect 187752 48804 187758 48816
rect 188982 48804 188988 48816
rect 187752 48776 188988 48804
rect 187752 48764 187758 48776
rect 188982 48764 188988 48776
rect 189040 48764 189046 48816
rect 193582 48764 193588 48816
rect 193640 48804 193646 48816
rect 194502 48804 194508 48816
rect 193640 48776 194508 48804
rect 193640 48764 193646 48776
rect 194502 48764 194508 48776
rect 194560 48764 194566 48816
rect 201954 48764 201960 48816
rect 202012 48804 202018 48816
rect 202782 48804 202788 48816
rect 202012 48776 202788 48804
rect 202012 48764 202018 48776
rect 202782 48764 202788 48776
rect 202840 48764 202846 48816
rect 203150 48764 203156 48816
rect 203208 48804 203214 48816
rect 204162 48804 204168 48816
rect 203208 48776 204168 48804
rect 203208 48764 203214 48776
rect 204162 48764 204168 48776
rect 204220 48764 204226 48816
rect 204346 48764 204352 48816
rect 204404 48804 204410 48816
rect 205542 48804 205548 48816
rect 204404 48776 205548 48804
rect 204404 48764 204410 48776
rect 205542 48764 205548 48776
rect 205600 48764 205606 48816
rect 211522 48764 211528 48816
rect 211580 48804 211586 48816
rect 212442 48804 212448 48816
rect 211580 48776 212448 48804
rect 211580 48764 211586 48776
rect 212442 48764 212448 48776
rect 212500 48764 212506 48816
rect 212718 48764 212724 48816
rect 212776 48804 212782 48816
rect 213822 48804 213828 48816
rect 212776 48776 213828 48804
rect 212776 48764 212782 48776
rect 213822 48764 213828 48776
rect 213880 48764 213886 48816
rect 213914 48764 213920 48816
rect 213972 48804 213978 48816
rect 215202 48804 215208 48816
rect 213972 48776 215208 48804
rect 213972 48764 213978 48776
rect 215202 48764 215208 48776
rect 215260 48764 215266 48816
rect 218606 48764 218612 48816
rect 218664 48804 218670 48816
rect 219342 48804 219348 48816
rect 218664 48776 219348 48804
rect 218664 48764 218670 48776
rect 219342 48764 219348 48776
rect 219400 48764 219406 48816
rect 220998 48764 221004 48816
rect 221056 48804 221062 48816
rect 222102 48804 222108 48816
rect 221056 48776 222108 48804
rect 221056 48764 221062 48776
rect 222102 48764 222108 48776
rect 222160 48764 222166 48816
rect 222194 48764 222200 48816
rect 222252 48804 222258 48816
rect 223482 48804 223488 48816
rect 222252 48776 223488 48804
rect 222252 48764 222258 48776
rect 223482 48764 223488 48776
rect 223540 48764 223546 48816
rect 228174 48764 228180 48816
rect 228232 48804 228238 48816
rect 229002 48804 229008 48816
rect 228232 48776 229008 48804
rect 228232 48764 228238 48776
rect 229002 48764 229008 48776
rect 229060 48764 229066 48816
rect 229370 48764 229376 48816
rect 229428 48804 229434 48816
rect 230382 48804 230388 48816
rect 229428 48776 230388 48804
rect 229428 48764 229434 48776
rect 230382 48764 230388 48776
rect 230440 48764 230446 48816
rect 237742 48764 237748 48816
rect 237800 48804 237806 48816
rect 238662 48804 238668 48816
rect 237800 48776 238668 48804
rect 237800 48764 237806 48776
rect 238662 48764 238668 48776
rect 238720 48764 238726 48816
rect 246022 48764 246028 48816
rect 246080 48804 246086 48816
rect 246942 48804 246948 48816
rect 246080 48776 246948 48804
rect 246080 48764 246086 48776
rect 246942 48764 246948 48776
rect 247000 48764 247006 48816
rect 247218 48764 247224 48816
rect 247276 48804 247282 48816
rect 248322 48804 248328 48816
rect 247276 48776 248328 48804
rect 247276 48764 247282 48776
rect 248322 48764 248328 48776
rect 248380 48764 248386 48816
rect 248414 48764 248420 48816
rect 248472 48804 248478 48816
rect 249610 48804 249616 48816
rect 248472 48776 249616 48804
rect 248472 48764 248478 48776
rect 249610 48764 249616 48776
rect 249668 48764 249674 48816
rect 254394 48764 254400 48816
rect 254452 48804 254458 48816
rect 255222 48804 255228 48816
rect 254452 48776 255228 48804
rect 254452 48764 254458 48776
rect 255222 48764 255228 48776
rect 255280 48764 255286 48816
rect 255590 48764 255596 48816
rect 255648 48804 255654 48816
rect 256602 48804 256608 48816
rect 255648 48776 256608 48804
rect 255648 48764 255654 48776
rect 256602 48764 256608 48776
rect 256660 48764 256666 48816
rect 256786 48764 256792 48816
rect 256844 48804 256850 48816
rect 257982 48804 257988 48816
rect 256844 48776 257988 48804
rect 256844 48764 256850 48776
rect 257982 48764 257988 48776
rect 258040 48764 258046 48816
rect 263962 48764 263968 48816
rect 264020 48804 264026 48816
rect 264882 48804 264888 48816
rect 264020 48776 264888 48804
rect 264020 48764 264026 48776
rect 264882 48764 264888 48776
rect 264940 48764 264946 48816
rect 265158 48764 265164 48816
rect 265216 48804 265222 48816
rect 266262 48804 266268 48816
rect 265216 48776 266268 48804
rect 265216 48764 265222 48776
rect 266262 48764 266268 48776
rect 266320 48764 266326 48816
rect 266354 48764 266360 48816
rect 266412 48804 266418 48816
rect 267550 48804 267556 48816
rect 266412 48776 267556 48804
rect 266412 48764 266418 48776
rect 267550 48764 267556 48776
rect 267608 48764 267614 48816
rect 272242 48764 272248 48816
rect 272300 48804 272306 48816
rect 273162 48804 273168 48816
rect 272300 48776 273168 48804
rect 272300 48764 272306 48776
rect 273162 48764 273168 48776
rect 273220 48764 273226 48816
rect 273438 48764 273444 48816
rect 273496 48804 273502 48816
rect 274542 48804 274548 48816
rect 273496 48776 274548 48804
rect 273496 48764 273502 48776
rect 274542 48764 274548 48776
rect 274600 48764 274606 48816
rect 274634 48764 274640 48816
rect 274692 48804 274698 48816
rect 275830 48804 275836 48816
rect 274692 48776 275836 48804
rect 274692 48764 274698 48776
rect 275830 48764 275836 48776
rect 275888 48764 275894 48816
rect 280614 48764 280620 48816
rect 280672 48804 280678 48816
rect 281442 48804 281448 48816
rect 280672 48776 281448 48804
rect 280672 48764 280678 48776
rect 281442 48764 281448 48776
rect 281500 48764 281506 48816
rect 281810 48764 281816 48816
rect 281868 48804 281874 48816
rect 282822 48804 282828 48816
rect 281868 48776 282828 48804
rect 281868 48764 281874 48776
rect 282822 48764 282828 48776
rect 282880 48764 282886 48816
rect 283006 48764 283012 48816
rect 283064 48804 283070 48816
rect 284202 48804 284208 48816
rect 283064 48776 284208 48804
rect 283064 48764 283070 48776
rect 284202 48764 284208 48776
rect 284260 48764 284266 48816
rect 290182 48764 290188 48816
rect 290240 48804 290246 48816
rect 291102 48804 291108 48816
rect 290240 48776 291108 48804
rect 290240 48764 290246 48776
rect 291102 48764 291108 48776
rect 291160 48764 291166 48816
rect 291378 48764 291384 48816
rect 291436 48804 291442 48816
rect 292482 48804 292488 48816
rect 291436 48776 292488 48804
rect 291436 48764 291442 48776
rect 292482 48764 292488 48776
rect 292540 48764 292546 48816
rect 292574 48764 292580 48816
rect 292632 48804 292638 48816
rect 293862 48804 293868 48816
rect 292632 48776 293868 48804
rect 292632 48764 292638 48776
rect 293862 48764 293868 48776
rect 293920 48764 293926 48816
rect 298462 48764 298468 48816
rect 298520 48804 298526 48816
rect 299382 48804 299388 48816
rect 298520 48776 299388 48804
rect 298520 48764 298526 48776
rect 299382 48764 299388 48776
rect 299440 48764 299446 48816
rect 299658 48764 299664 48816
rect 299716 48804 299722 48816
rect 300762 48804 300768 48816
rect 299716 48776 300768 48804
rect 299716 48764 299722 48776
rect 300762 48764 300768 48776
rect 300820 48764 300826 48816
rect 300854 48764 300860 48816
rect 300912 48804 300918 48816
rect 302142 48804 302148 48816
rect 300912 48776 302148 48804
rect 300912 48764 300918 48776
rect 302142 48764 302148 48776
rect 302200 48764 302206 48816
rect 306834 48764 306840 48816
rect 306892 48804 306898 48816
rect 307662 48804 307668 48816
rect 306892 48776 307668 48804
rect 306892 48764 306898 48776
rect 307662 48764 307668 48776
rect 307720 48764 307726 48816
rect 308030 48764 308036 48816
rect 308088 48804 308094 48816
rect 309042 48804 309048 48816
rect 308088 48776 309048 48804
rect 308088 48764 308094 48776
rect 309042 48764 309048 48776
rect 309100 48764 309106 48816
rect 309226 48764 309232 48816
rect 309284 48804 309290 48816
rect 310330 48804 310336 48816
rect 309284 48776 310336 48804
rect 309284 48764 309290 48776
rect 310330 48764 310336 48776
rect 310388 48764 310394 48816
rect 316402 48764 316408 48816
rect 316460 48804 316466 48816
rect 317322 48804 317328 48816
rect 316460 48776 317328 48804
rect 316460 48764 316466 48776
rect 317322 48764 317328 48776
rect 317380 48764 317386 48816
rect 323486 48764 323492 48816
rect 323544 48804 323550 48816
rect 324222 48804 324228 48816
rect 323544 48776 324228 48804
rect 323544 48764 323550 48776
rect 324222 48764 324228 48776
rect 324280 48764 324286 48816
rect 324682 48764 324688 48816
rect 324740 48804 324746 48816
rect 325602 48804 325608 48816
rect 324740 48776 325608 48804
rect 324740 48764 324746 48776
rect 325602 48764 325608 48776
rect 325660 48764 325666 48816
rect 325878 48764 325884 48816
rect 325936 48804 325942 48816
rect 326982 48804 326988 48816
rect 325936 48776 326988 48804
rect 325936 48764 325942 48776
rect 326982 48764 326988 48776
rect 327040 48764 327046 48816
rect 327074 48764 327080 48816
rect 327132 48804 327138 48816
rect 328270 48804 328276 48816
rect 327132 48776 328276 48804
rect 327132 48764 327138 48776
rect 328270 48764 328276 48776
rect 328328 48764 328334 48816
rect 329466 48764 329472 48816
rect 329524 48804 329530 48816
rect 330478 48804 330484 48816
rect 329524 48776 330484 48804
rect 329524 48764 329530 48776
rect 330478 48764 330484 48776
rect 330536 48764 330542 48816
rect 333054 48764 333060 48816
rect 333112 48804 333118 48816
rect 333882 48804 333888 48816
rect 333112 48776 333888 48804
rect 333112 48764 333118 48776
rect 333882 48764 333888 48776
rect 333940 48764 333946 48816
rect 334250 48764 334256 48816
rect 334308 48804 334314 48816
rect 335262 48804 335268 48816
rect 334308 48776 335268 48804
rect 334308 48764 334314 48776
rect 335262 48764 335268 48776
rect 335320 48764 335326 48816
rect 335446 48764 335452 48816
rect 335504 48804 335510 48816
rect 336642 48804 336648 48816
rect 335504 48776 336648 48804
rect 335504 48764 335510 48776
rect 336642 48764 336648 48776
rect 336700 48764 336706 48816
rect 342622 48764 342628 48816
rect 342680 48804 342686 48816
rect 343542 48804 343548 48816
rect 342680 48776 343548 48804
rect 342680 48764 342686 48776
rect 343542 48764 343548 48776
rect 343600 48764 343606 48816
rect 343726 48764 343732 48816
rect 343784 48804 343790 48816
rect 344830 48804 344836 48816
rect 343784 48776 344836 48804
rect 343784 48764 343790 48776
rect 344830 48764 344836 48776
rect 344888 48764 344894 48816
rect 350902 48764 350908 48816
rect 350960 48804 350966 48816
rect 351822 48804 351828 48816
rect 350960 48776 351828 48804
rect 350960 48764 350966 48776
rect 351822 48764 351828 48776
rect 351880 48764 351886 48816
rect 352098 48764 352104 48816
rect 352156 48804 352162 48816
rect 353202 48804 353208 48816
rect 352156 48776 353208 48804
rect 352156 48764 352162 48776
rect 353202 48764 353208 48776
rect 353260 48764 353266 48816
rect 353294 48764 353300 48816
rect 353352 48804 353358 48816
rect 354582 48804 354588 48816
rect 353352 48776 354588 48804
rect 353352 48764 353358 48776
rect 354582 48764 354588 48776
rect 354640 48764 354646 48816
rect 359274 48764 359280 48816
rect 359332 48804 359338 48816
rect 360102 48804 360108 48816
rect 359332 48776 360108 48804
rect 359332 48764 359338 48776
rect 360102 48764 360108 48776
rect 360160 48764 360166 48816
rect 360470 48764 360476 48816
rect 360528 48804 360534 48816
rect 361482 48804 361488 48816
rect 360528 48776 361488 48804
rect 360528 48764 360534 48776
rect 361482 48764 361488 48776
rect 361540 48764 361546 48816
rect 361666 48764 361672 48816
rect 361724 48804 361730 48816
rect 362862 48804 362868 48816
rect 361724 48776 362868 48804
rect 361724 48764 361730 48776
rect 362862 48764 362868 48776
rect 362920 48764 362926 48816
rect 369946 48764 369952 48816
rect 370004 48804 370010 48816
rect 371878 48804 371884 48816
rect 370004 48776 371884 48804
rect 370004 48764 370010 48776
rect 371878 48764 371884 48776
rect 371936 48764 371942 48816
rect 377122 48764 377128 48816
rect 377180 48804 377186 48816
rect 378042 48804 378048 48816
rect 377180 48776 378048 48804
rect 377180 48764 377186 48776
rect 378042 48764 378048 48776
rect 378100 48764 378106 48816
rect 378318 48764 378324 48816
rect 378376 48804 378382 48816
rect 379422 48804 379428 48816
rect 378376 48776 379428 48804
rect 378376 48764 378382 48776
rect 379422 48764 379428 48776
rect 379480 48764 379486 48816
rect 379514 48764 379520 48816
rect 379572 48804 379578 48816
rect 380802 48804 380808 48816
rect 379572 48776 380808 48804
rect 379572 48764 379578 48776
rect 380802 48764 380808 48776
rect 380860 48764 380866 48816
rect 386690 48764 386696 48816
rect 386748 48804 386754 48816
rect 387702 48804 387708 48816
rect 386748 48776 387708 48804
rect 386748 48764 386754 48776
rect 387702 48764 387708 48776
rect 387760 48764 387766 48816
rect 394970 48764 394976 48816
rect 395028 48804 395034 48816
rect 395982 48804 395988 48816
rect 395028 48776 395988 48804
rect 395028 48764 395034 48776
rect 395982 48764 395988 48776
rect 396040 48764 396046 48816
rect 405734 48764 405740 48816
rect 405792 48804 405798 48816
rect 406930 48804 406936 48816
rect 405792 48776 406936 48804
rect 405792 48764 405798 48776
rect 406930 48764 406936 48776
rect 406988 48764 406994 48816
rect 412910 48764 412916 48816
rect 412968 48804 412974 48816
rect 413922 48804 413928 48816
rect 412968 48776 413928 48804
rect 412968 48764 412974 48776
rect 413922 48764 413928 48776
rect 413980 48764 413986 48816
rect 414106 48764 414112 48816
rect 414164 48804 414170 48816
rect 415302 48804 415308 48816
rect 414164 48776 415308 48804
rect 414164 48764 414170 48776
rect 415302 48764 415308 48776
rect 415360 48764 415366 48816
rect 420086 48764 420092 48816
rect 420144 48804 420150 48816
rect 420822 48804 420828 48816
rect 420144 48776 420828 48804
rect 420144 48764 420150 48776
rect 420822 48764 420828 48776
rect 420880 48764 420886 48816
rect 421190 48764 421196 48816
rect 421248 48804 421254 48816
rect 422202 48804 422208 48816
rect 421248 48776 422208 48804
rect 421248 48764 421254 48776
rect 422202 48764 422208 48776
rect 422260 48764 422266 48816
rect 428366 48764 428372 48816
rect 428424 48804 428430 48816
rect 429102 48804 429108 48816
rect 428424 48776 429108 48804
rect 428424 48764 428430 48776
rect 429102 48764 429108 48776
rect 429160 48764 429166 48816
rect 429562 48764 429568 48816
rect 429620 48804 429626 48816
rect 430482 48804 430488 48816
rect 429620 48776 430488 48804
rect 429620 48764 429626 48776
rect 430482 48764 430488 48776
rect 430540 48764 430546 48816
rect 430758 48764 430764 48816
rect 430816 48804 430822 48816
rect 431862 48804 431868 48816
rect 430816 48776 431868 48804
rect 430816 48764 430822 48776
rect 431862 48764 431868 48776
rect 431920 48764 431926 48816
rect 431954 48764 431960 48816
rect 432012 48804 432018 48816
rect 433150 48804 433156 48816
rect 432012 48776 433156 48804
rect 432012 48764 432018 48776
rect 433150 48764 433156 48776
rect 433208 48764 433214 48816
rect 439130 48764 439136 48816
rect 439188 48804 439194 48816
rect 440142 48804 440148 48816
rect 439188 48776 440148 48804
rect 439188 48764 439194 48776
rect 440142 48764 440148 48776
rect 440200 48764 440206 48816
rect 440326 48764 440332 48816
rect 440384 48804 440390 48816
rect 441522 48804 441528 48816
rect 440384 48776 441528 48804
rect 440384 48764 440390 48776
rect 441522 48764 441528 48776
rect 441580 48764 441586 48816
rect 446214 48764 446220 48816
rect 446272 48804 446278 48816
rect 447042 48804 447048 48816
rect 446272 48776 447048 48804
rect 446272 48764 446278 48776
rect 447042 48764 447048 48776
rect 447100 48764 447106 48816
rect 447410 48764 447416 48816
rect 447468 48804 447474 48816
rect 448422 48804 448428 48816
rect 447468 48776 448428 48804
rect 447468 48764 447474 48776
rect 448422 48764 448428 48776
rect 448480 48764 448486 48816
rect 448606 48764 448612 48816
rect 448664 48804 448670 48816
rect 449710 48804 449716 48816
rect 448664 48776 449716 48804
rect 448664 48764 448670 48776
rect 449710 48764 449716 48776
rect 449768 48764 449774 48816
rect 455782 48764 455788 48816
rect 455840 48804 455846 48816
rect 456702 48804 456708 48816
rect 455840 48776 456708 48804
rect 455840 48764 455846 48776
rect 456702 48764 456708 48776
rect 456760 48764 456766 48816
rect 456978 48764 456984 48816
rect 457036 48804 457042 48816
rect 458082 48804 458088 48816
rect 457036 48776 458088 48804
rect 457036 48764 457042 48776
rect 458082 48764 458088 48776
rect 458140 48764 458146 48816
rect 458174 48764 458180 48816
rect 458232 48804 458238 48816
rect 459462 48804 459468 48816
rect 458232 48776 459468 48804
rect 458232 48764 458238 48776
rect 459462 48764 459468 48776
rect 459520 48764 459526 48816
rect 464154 48764 464160 48816
rect 464212 48804 464218 48816
rect 464982 48804 464988 48816
rect 464212 48776 464988 48804
rect 464212 48764 464218 48776
rect 464982 48764 464988 48776
rect 465040 48764 465046 48816
rect 465350 48764 465356 48816
rect 465408 48804 465414 48816
rect 466362 48804 466368 48816
rect 465408 48776 466368 48804
rect 465408 48764 465414 48776
rect 466362 48764 466368 48776
rect 466420 48764 466426 48816
rect 466546 48764 466552 48816
rect 466604 48804 466610 48816
rect 467742 48804 467748 48816
rect 466604 48776 467748 48804
rect 466604 48764 466610 48776
rect 467742 48764 467748 48776
rect 467800 48764 467806 48816
rect 473630 48764 473636 48816
rect 473688 48804 473694 48816
rect 474642 48804 474648 48816
rect 473688 48776 474648 48804
rect 473688 48764 473694 48776
rect 474642 48764 474648 48776
rect 474700 48764 474706 48816
rect 480806 48764 480812 48816
rect 480864 48804 480870 48816
rect 481542 48804 481548 48816
rect 480864 48776 481548 48804
rect 480864 48764 480870 48776
rect 481542 48764 481548 48776
rect 481600 48764 481606 48816
rect 483198 48764 483204 48816
rect 483256 48804 483262 48816
rect 484302 48804 484308 48816
rect 483256 48776 484308 48804
rect 483256 48764 483262 48776
rect 484302 48764 484308 48776
rect 484360 48764 484366 48816
rect 491570 48764 491576 48816
rect 491628 48804 491634 48816
rect 492582 48804 492588 48816
rect 491628 48776 492588 48804
rect 491628 48764 491634 48776
rect 492582 48764 492588 48776
rect 492640 48764 492646 48816
rect 492766 48764 492772 48816
rect 492824 48804 492830 48816
rect 493962 48804 493968 48816
rect 492824 48776 493968 48804
rect 492824 48764 492830 48776
rect 493962 48764 493968 48776
rect 494020 48764 494026 48816
rect 498654 48764 498660 48816
rect 498712 48804 498718 48816
rect 499482 48804 499488 48816
rect 498712 48776 499488 48804
rect 498712 48764 498718 48776
rect 499482 48764 499488 48776
rect 499540 48764 499546 48816
rect 499850 48764 499856 48816
rect 499908 48804 499914 48816
rect 500862 48804 500868 48816
rect 499908 48776 500868 48804
rect 499908 48764 499914 48776
rect 500862 48764 500868 48776
rect 500920 48764 500926 48816
rect 501046 48764 501052 48816
rect 501104 48804 501110 48816
rect 502242 48804 502248 48816
rect 501104 48776 502248 48804
rect 501104 48764 501110 48776
rect 502242 48764 502248 48776
rect 502300 48764 502306 48816
rect 508222 48764 508228 48816
rect 508280 48804 508286 48816
rect 509142 48804 509148 48816
rect 508280 48776 509148 48804
rect 508280 48764 508286 48776
rect 509142 48764 509148 48776
rect 509200 48764 509206 48816
rect 509418 48764 509424 48816
rect 509476 48804 509482 48816
rect 510522 48804 510528 48816
rect 509476 48776 510528 48804
rect 509476 48764 509482 48776
rect 510522 48764 510528 48776
rect 510580 48764 510586 48816
rect 516594 48764 516600 48816
rect 516652 48804 516658 48816
rect 517422 48804 517428 48816
rect 516652 48776 517428 48804
rect 516652 48764 516658 48776
rect 517422 48764 517428 48776
rect 517480 48764 517486 48816
rect 517790 48764 517796 48816
rect 517848 48804 517854 48816
rect 518802 48804 518808 48816
rect 517848 48776 518808 48804
rect 517848 48764 517854 48776
rect 518802 48764 518808 48776
rect 518860 48764 518866 48816
rect 518986 48764 518992 48816
rect 519044 48804 519050 48816
rect 520090 48804 520096 48816
rect 519044 48776 520096 48804
rect 519044 48764 519050 48776
rect 520090 48764 520096 48776
rect 520148 48764 520154 48816
rect 64874 48696 64880 48748
rect 64932 48736 64938 48748
rect 66162 48736 66168 48748
rect 64932 48708 66168 48736
rect 64932 48696 64938 48708
rect 66162 48696 66168 48708
rect 66220 48696 66226 48748
rect 238938 48696 238944 48748
rect 238996 48736 239002 48748
rect 240042 48736 240048 48748
rect 238996 48708 240048 48736
rect 238996 48696 239002 48708
rect 240042 48696 240048 48708
rect 240100 48696 240106 48748
rect 271046 48696 271052 48748
rect 271104 48736 271110 48748
rect 272518 48736 272524 48748
rect 271104 48708 272524 48736
rect 271104 48696 271110 48708
rect 272518 48696 272524 48708
rect 272576 48696 272582 48748
rect 315206 48696 315212 48748
rect 315264 48736 315270 48748
rect 315942 48736 315948 48748
rect 315264 48708 315948 48736
rect 315264 48696 315270 48708
rect 315942 48696 315948 48708
rect 316000 48696 316006 48748
rect 375926 48696 375932 48748
rect 375984 48736 375990 48748
rect 376662 48736 376668 48748
rect 375984 48708 376668 48736
rect 375984 48696 375990 48708
rect 376662 48696 376668 48708
rect 376720 48696 376726 48748
rect 472434 48696 472440 48748
rect 472492 48736 472498 48748
rect 473998 48736 474004 48748
rect 472492 48708 474004 48736
rect 472492 48696 472498 48708
rect 473998 48696 474004 48708
rect 474056 48696 474062 48748
rect 82814 48628 82820 48680
rect 82872 48668 82878 48680
rect 84010 48668 84016 48680
rect 82872 48640 84016 48668
rect 82872 48628 82878 48640
rect 84010 48628 84016 48640
rect 84068 48628 84074 48680
rect 125686 48628 125692 48680
rect 125744 48668 125750 48680
rect 126882 48668 126888 48680
rect 125744 48640 126888 48668
rect 125744 48628 125750 48640
rect 126882 48628 126888 48640
rect 126940 48628 126946 48680
rect 195974 48628 195980 48680
rect 196032 48668 196038 48680
rect 197262 48668 197268 48680
rect 196032 48640 197268 48668
rect 196032 48628 196038 48640
rect 197262 48628 197268 48640
rect 197320 48628 197326 48680
rect 230566 48628 230572 48680
rect 230624 48668 230630 48680
rect 231670 48668 231676 48680
rect 230624 48640 231676 48668
rect 230624 48628 230630 48640
rect 231670 48628 231676 48640
rect 231728 48628 231734 48680
rect 383102 48628 383108 48680
rect 383160 48668 383166 48680
rect 384298 48668 384304 48680
rect 383160 48640 384304 48668
rect 383160 48628 383166 48640
rect 384298 48628 384304 48640
rect 384356 48628 384362 48680
rect 387886 48628 387892 48680
rect 387944 48668 387950 48680
rect 389082 48668 389088 48680
rect 387944 48640 389088 48668
rect 387944 48628 387950 48640
rect 389082 48628 389088 48640
rect 389140 48628 389146 48680
rect 404538 48628 404544 48680
rect 404596 48668 404602 48680
rect 405642 48668 405648 48680
rect 404596 48640 405648 48668
rect 404596 48628 404602 48640
rect 405642 48628 405648 48640
rect 405700 48628 405706 48680
rect 135254 48492 135260 48544
rect 135312 48532 135318 48544
rect 136450 48532 136456 48544
rect 135312 48504 136456 48532
rect 135312 48492 135318 48504
rect 136450 48492 136456 48504
rect 136508 48492 136514 48544
rect 143534 48492 143540 48544
rect 143592 48532 143598 48544
rect 144822 48532 144828 48544
rect 143592 48504 144828 48532
rect 143592 48492 143598 48504
rect 144822 48492 144828 48504
rect 144880 48492 144886 48544
rect 166166 48492 166172 48544
rect 166224 48532 166230 48544
rect 167638 48532 167644 48544
rect 166224 48504 167644 48532
rect 166224 48492 166230 48504
rect 167638 48492 167644 48504
rect 167696 48492 167702 48544
rect 510614 48492 510620 48544
rect 510672 48532 510678 48544
rect 511902 48532 511908 48544
rect 510672 48504 511908 48532
rect 510672 48492 510678 48504
rect 511902 48492 511908 48504
rect 511960 48492 511966 48544
rect 411714 48424 411720 48476
rect 411772 48464 411778 48476
rect 412542 48464 412548 48476
rect 411772 48436 412548 48464
rect 411772 48424 411778 48436
rect 412542 48424 412548 48436
rect 412600 48424 412606 48476
rect 437934 48424 437940 48476
rect 437992 48464 437998 48476
rect 438762 48464 438768 48476
rect 437992 48436 438768 48464
rect 437992 48424 437998 48436
rect 438762 48424 438768 48436
rect 438820 48424 438826 48476
rect 385494 48356 385500 48408
rect 385552 48396 385558 48408
rect 386322 48396 386328 48408
rect 385552 48368 386328 48396
rect 385552 48356 385558 48368
rect 386322 48356 386328 48368
rect 386380 48356 386386 48408
rect 240134 48288 240140 48340
rect 240192 48328 240198 48340
rect 241422 48328 241428 48340
rect 240192 48300 241428 48328
rect 240192 48288 240198 48300
rect 241422 48288 241428 48300
rect 241480 48288 241486 48340
rect 262766 48288 262772 48340
rect 262824 48328 262830 48340
rect 263502 48328 263508 48340
rect 262824 48300 263508 48328
rect 262824 48288 262830 48300
rect 263502 48288 263508 48300
rect 263560 48288 263566 48340
rect 317598 48288 317604 48340
rect 317656 48328 317662 48340
rect 318702 48328 318708 48340
rect 317656 48300 318708 48328
rect 317656 48288 317662 48300
rect 318702 48288 318708 48300
rect 318760 48288 318766 48340
rect 368842 48288 368848 48340
rect 368900 48328 368906 48340
rect 369762 48328 369768 48340
rect 368900 48300 369768 48328
rect 368900 48288 368906 48300
rect 369762 48288 369768 48300
rect 369820 48288 369826 48340
rect 422386 48288 422392 48340
rect 422444 48328 422450 48340
rect 423582 48328 423588 48340
rect 422444 48300 423588 48328
rect 422444 48288 422450 48300
rect 423582 48288 423588 48300
rect 423640 48288 423646 48340
rect 427906 48328 427912 48340
rect 427867 48300 427912 48328
rect 427906 48288 427912 48300
rect 427964 48288 427970 48340
rect 434806 48328 434812 48340
rect 434767 48300 434812 48328
rect 434806 48288 434812 48300
rect 434864 48288 434870 48340
rect 484394 48288 484400 48340
rect 484452 48328 484458 48340
rect 485590 48328 485596 48340
rect 484452 48300 485596 48328
rect 484452 48288 484458 48300
rect 485590 48288 485596 48300
rect 485648 48288 485654 48340
rect 76834 47608 76840 47660
rect 76892 47648 76898 47660
rect 138014 47648 138020 47660
rect 76892 47620 138020 47648
rect 76892 47608 76898 47620
rect 138014 47608 138020 47620
rect 138072 47608 138078 47660
rect 194778 47608 194784 47660
rect 194836 47648 194842 47660
rect 255314 47648 255320 47660
rect 194836 47620 255320 47648
rect 194836 47608 194842 47620
rect 255314 47608 255320 47620
rect 255372 47608 255378 47660
rect 490374 47608 490380 47660
rect 490432 47648 490438 47660
rect 550634 47648 550640 47660
rect 490432 47620 550640 47648
rect 490432 47608 490438 47620
rect 550634 47608 550640 47620
rect 550692 47608 550698 47660
rect 136542 47540 136548 47592
rect 136600 47580 136606 47592
rect 197354 47580 197360 47592
rect 136600 47552 197360 47580
rect 136600 47540 136606 47552
rect 197354 47540 197360 47552
rect 197412 47540 197418 47592
rect 275922 47540 275928 47592
rect 275980 47580 275986 47592
rect 336734 47580 336740 47592
rect 275980 47552 336740 47580
rect 275980 47540 275986 47552
rect 336734 47540 336740 47552
rect 336792 47540 336798 47592
rect 347314 47540 347320 47592
rect 347372 47580 347378 47592
rect 408494 47580 408500 47592
rect 347372 47552 408500 47580
rect 347372 47540 347378 47552
rect 408494 47540 408500 47552
rect 408552 47540 408558 47592
rect 433242 47540 433248 47592
rect 433300 47580 433306 47592
rect 494054 47580 494060 47592
rect 433300 47552 494060 47580
rect 433300 47540 433306 47552
rect 494054 47540 494060 47552
rect 494112 47540 494118 47592
rect 219802 46316 219808 46368
rect 219860 46356 219866 46368
rect 280154 46356 280160 46368
rect 219860 46328 280160 46356
rect 219860 46316 219866 46328
rect 280154 46316 280160 46328
rect 280212 46316 280218 46368
rect 112622 46248 112628 46300
rect 112680 46288 112686 46300
rect 173894 46288 173900 46300
rect 112680 46260 173900 46288
rect 112680 46248 112686 46260
rect 173894 46248 173900 46260
rect 173952 46248 173958 46300
rect 278222 46248 278228 46300
rect 278280 46288 278286 46300
rect 339494 46288 339500 46300
rect 278280 46260 339500 46288
rect 278280 46248 278286 46260
rect 339494 46248 339500 46260
rect 339552 46248 339558 46300
rect 162670 46180 162676 46232
rect 162728 46220 162734 46232
rect 223574 46220 223580 46232
rect 162728 46192 223580 46220
rect 162728 46180 162734 46192
rect 223574 46180 223580 46192
rect 223632 46180 223638 46232
rect 293678 46180 293684 46232
rect 293736 46220 293742 46232
rect 354674 46220 354680 46232
rect 293736 46192 354680 46220
rect 293736 46180 293742 46192
rect 354674 46180 354680 46192
rect 354732 46180 354738 46232
rect 365254 46180 365260 46232
rect 365312 46220 365318 46232
rect 425054 46220 425060 46232
rect 365312 46192 425060 46220
rect 365312 46180 365318 46192
rect 425054 46180 425060 46192
rect 425112 46180 425118 46232
rect 436738 46180 436744 46232
rect 436796 46220 436802 46232
rect 496814 46220 496820 46232
rect 436796 46192 496820 46220
rect 436796 46180 436802 46192
rect 496814 46180 496820 46192
rect 496872 46180 496878 46232
rect 497458 46180 497464 46232
rect 497516 46220 497522 46232
rect 557534 46220 557540 46232
rect 497516 46192 557540 46220
rect 497516 46180 497522 46192
rect 557534 46180 557540 46192
rect 557592 46180 557598 46232
rect 184842 44956 184848 45008
rect 184900 44996 184906 45008
rect 244274 44996 244280 45008
rect 184900 44968 244280 44996
rect 184900 44956 184906 44968
rect 244274 44956 244280 44968
rect 244332 44956 244338 45008
rect 238662 44888 238668 44940
rect 238720 44928 238726 44940
rect 298094 44928 298100 44940
rect 238720 44900 298100 44928
rect 238720 44888 238726 44900
rect 298094 44888 298100 44900
rect 298152 44888 298158 44940
rect 338022 44888 338028 44940
rect 338080 44928 338086 44940
rect 398834 44928 398840 44940
rect 338080 44900 398840 44928
rect 338080 44888 338086 44900
rect 398834 44888 398840 44900
rect 398892 44888 398898 44940
rect 509142 44888 509148 44940
rect 509200 44928 509206 44940
rect 568574 44928 568580 44940
rect 509200 44900 568580 44928
rect 509200 44888 509206 44900
rect 568574 44888 568580 44900
rect 568632 44888 568638 44940
rect 131022 44820 131028 44872
rect 131080 44860 131086 44872
rect 191834 44860 191840 44872
rect 131080 44832 191840 44860
rect 131080 44820 131086 44832
rect 191834 44820 191840 44832
rect 191892 44820 191898 44872
rect 284110 44820 284116 44872
rect 284168 44860 284174 44872
rect 345014 44860 345020 44872
rect 284168 44832 345020 44860
rect 284168 44820 284174 44832
rect 345014 44820 345020 44832
rect 345072 44820 345078 44872
rect 384942 44820 384948 44872
rect 385000 44860 385006 44872
rect 444374 44860 444380 44872
rect 385000 44832 444380 44860
rect 385000 44820 385006 44832
rect 444374 44820 444380 44832
rect 444432 44820 444438 44872
rect 451182 44820 451188 44872
rect 451240 44860 451246 44872
rect 511994 44860 512000 44872
rect 451240 44832 512000 44860
rect 451240 44820 451246 44832
rect 511994 44820 512000 44832
rect 512052 44820 512058 44872
rect 263502 43460 263508 43512
rect 263560 43500 263566 43512
rect 323026 43500 323032 43512
rect 263560 43472 323032 43500
rect 263560 43460 263566 43472
rect 323026 43460 323032 43472
rect 323084 43460 323090 43512
rect 148962 43392 148968 43444
rect 149020 43432 149026 43444
rect 209866 43432 209872 43444
rect 149020 43404 209872 43432
rect 149020 43392 149026 43404
rect 209866 43392 209872 43404
rect 209924 43392 209930 43444
rect 213822 43392 213828 43444
rect 213880 43432 213886 43444
rect 273254 43432 273260 43444
rect 213880 43404 273260 43432
rect 213880 43392 213886 43404
rect 273254 43392 273260 43404
rect 273312 43392 273318 43444
rect 313182 43392 313188 43444
rect 313240 43432 313246 43444
rect 374086 43432 374092 43444
rect 313240 43404 374092 43432
rect 313240 43392 313246 43404
rect 374086 43392 374092 43404
rect 374144 43392 374150 43444
rect 401502 43392 401508 43444
rect 401560 43432 401566 43444
rect 460934 43432 460940 43444
rect 401560 43404 460940 43432
rect 401560 43392 401566 43404
rect 460934 43392 460940 43404
rect 460992 43392 460998 43444
rect 473998 43392 474004 43444
rect 474056 43432 474062 43444
rect 532694 43432 532700 43444
rect 474056 43404 532700 43432
rect 474056 43392 474062 43404
rect 532694 43392 532700 43404
rect 532752 43392 532758 43444
rect 256602 42168 256608 42220
rect 256660 42208 256666 42220
rect 316034 42208 316040 42220
rect 256660 42180 316040 42208
rect 256660 42168 256666 42180
rect 316034 42168 316040 42180
rect 316092 42168 316098 42220
rect 202782 42100 202788 42152
rect 202840 42140 202846 42152
rect 262214 42140 262220 42152
rect 202840 42112 262220 42140
rect 202840 42100 202846 42112
rect 262214 42100 262220 42112
rect 262272 42100 262278 42152
rect 81342 42032 81348 42084
rect 81400 42072 81406 42084
rect 140774 42072 140780 42084
rect 81400 42044 140780 42072
rect 81400 42032 81406 42044
rect 140774 42032 140780 42044
rect 140832 42032 140838 42084
rect 144730 42032 144736 42084
rect 144788 42072 144794 42084
rect 205634 42072 205640 42084
rect 144788 42044 205640 42072
rect 144788 42032 144794 42044
rect 205634 42032 205640 42044
rect 205692 42032 205698 42084
rect 310330 42032 310336 42084
rect 310388 42072 310394 42084
rect 369854 42072 369860 42084
rect 310388 42044 369860 42072
rect 310388 42032 310394 42044
rect 369854 42032 369860 42044
rect 369912 42032 369918 42084
rect 415210 42032 415216 42084
rect 415268 42072 415274 42084
rect 476114 42072 476120 42084
rect 415268 42044 476120 42072
rect 415268 42032 415274 42044
rect 476114 42032 476120 42044
rect 476172 42032 476178 42084
rect 493870 42032 493876 42084
rect 493928 42072 493934 42084
rect 554774 42072 554780 42084
rect 493928 42044 554780 42072
rect 493928 42032 493934 42044
rect 554774 42032 554780 42044
rect 554832 42032 554838 42084
rect 523678 41352 523684 41404
rect 523736 41392 523742 41404
rect 580166 41392 580172 41404
rect 523736 41364 580172 41392
rect 523736 41352 523742 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 299382 40808 299388 40860
rect 299440 40848 299446 40860
rect 358814 40848 358820 40860
rect 299440 40820 358820 40848
rect 299440 40808 299446 40820
rect 358814 40808 358820 40820
rect 358872 40808 358878 40860
rect 142062 40740 142068 40792
rect 142120 40780 142126 40792
rect 201494 40780 201500 40792
rect 142120 40752 201500 40780
rect 142120 40740 142126 40752
rect 201494 40740 201500 40752
rect 201552 40740 201558 40792
rect 249610 40740 249616 40792
rect 249668 40780 249674 40792
rect 309134 40780 309140 40792
rect 249668 40752 309140 40780
rect 249668 40740 249674 40752
rect 309134 40740 309140 40752
rect 309192 40740 309198 40792
rect 74442 40672 74448 40724
rect 74500 40712 74506 40724
rect 133874 40712 133880 40724
rect 74500 40684 133880 40712
rect 74500 40672 74506 40684
rect 133874 40672 133880 40684
rect 133932 40672 133938 40724
rect 198642 40672 198648 40724
rect 198700 40712 198706 40724
rect 259454 40712 259460 40724
rect 198700 40684 259460 40712
rect 198700 40672 198706 40684
rect 259454 40672 259460 40684
rect 259512 40672 259518 40724
rect 355962 40672 355968 40724
rect 356020 40712 356026 40724
rect 416866 40712 416872 40724
rect 356020 40684 416872 40712
rect 356020 40672 356026 40684
rect 416866 40672 416872 40684
rect 416924 40672 416930 40724
rect 419442 40672 419448 40724
rect 419500 40712 419506 40724
rect 478874 40712 478880 40724
rect 419500 40684 478880 40712
rect 419500 40672 419506 40684
rect 478874 40672 478880 40684
rect 478932 40672 478938 40724
rect 331122 39448 331128 39500
rect 331180 39488 331186 39500
rect 390554 39488 390560 39500
rect 331180 39460 390560 39488
rect 331180 39448 331186 39460
rect 390554 39448 390560 39460
rect 390612 39448 390618 39500
rect 180702 39380 180708 39432
rect 180760 39420 180766 39432
rect 241514 39420 241520 39432
rect 180760 39392 241520 39420
rect 180760 39380 180766 39392
rect 241514 39380 241520 39392
rect 241572 39380 241578 39432
rect 281442 39380 281448 39432
rect 281500 39420 281506 39432
rect 340874 39420 340880 39432
rect 281500 39392 340880 39420
rect 281500 39380 281506 39392
rect 340874 39380 340880 39392
rect 340932 39380 340938 39432
rect 420822 39380 420828 39432
rect 420880 39420 420886 39432
rect 480254 39420 480260 39432
rect 420880 39392 480260 39420
rect 420880 39380 420886 39392
rect 480254 39380 480260 39392
rect 480312 39380 480318 39432
rect 126790 39312 126796 39364
rect 126848 39352 126854 39364
rect 187694 39352 187700 39364
rect 126848 39324 187700 39352
rect 126848 39312 126854 39324
rect 187694 39312 187700 39324
rect 187752 39312 187758 39364
rect 234522 39312 234528 39364
rect 234580 39352 234586 39364
rect 295334 39352 295340 39364
rect 234580 39324 295340 39352
rect 234580 39312 234586 39324
rect 295334 39312 295340 39324
rect 295392 39312 295398 39364
rect 380710 39312 380716 39364
rect 380768 39352 380774 39364
rect 441614 39352 441620 39364
rect 380768 39324 441620 39352
rect 380768 39312 380774 39324
rect 441614 39312 441620 39324
rect 441672 39312 441678 39364
rect 511810 39312 511816 39364
rect 511868 39352 511874 39364
rect 571426 39352 571432 39364
rect 511868 39324 571432 39352
rect 511868 39312 511874 39324
rect 571426 39312 571432 39324
rect 571484 39312 571490 39364
rect 369854 38564 369860 38616
rect 369912 38604 369918 38616
rect 369946 38604 369952 38616
rect 369912 38576 369952 38604
rect 369912 38564 369918 38576
rect 369946 38564 369952 38576
rect 370004 38564 370010 38616
rect 427906 38604 427912 38616
rect 427867 38576 427912 38604
rect 427906 38564 427912 38576
rect 427964 38564 427970 38616
rect 434806 38604 434812 38616
rect 434767 38576 434812 38604
rect 434806 38564 434812 38576
rect 434864 38564 434870 38616
rect 188982 37952 188988 38004
rect 189040 37992 189046 38004
rect 248414 37992 248420 38004
rect 189040 37964 248420 37992
rect 189040 37952 189046 37964
rect 248414 37952 248420 37964
rect 248472 37952 248478 38004
rect 288342 37952 288348 38004
rect 288400 37992 288406 38004
rect 347774 37992 347780 38004
rect 288400 37964 347780 37992
rect 288400 37952 288406 37964
rect 347774 37952 347780 37964
rect 347832 37952 347838 38004
rect 389082 37952 389088 38004
rect 389140 37992 389146 38004
rect 448514 37992 448520 38004
rect 389140 37964 448520 37992
rect 389140 37952 389146 37964
rect 448514 37952 448520 37964
rect 448572 37952 448578 38004
rect 70302 37884 70308 37936
rect 70360 37924 70366 37936
rect 131114 37924 131120 37936
rect 70360 37896 131120 37924
rect 70360 37884 70366 37896
rect 131114 37884 131120 37896
rect 131172 37884 131178 37936
rect 135162 37884 135168 37936
rect 135220 37924 135226 37936
rect 194594 37924 194600 37936
rect 135220 37896 194600 37924
rect 135220 37884 135226 37896
rect 194594 37884 194600 37896
rect 194652 37884 194658 37936
rect 241330 37884 241336 37936
rect 241388 37924 241394 37936
rect 302234 37924 302240 37936
rect 241388 37896 302240 37924
rect 241388 37884 241394 37896
rect 302234 37884 302240 37896
rect 302292 37884 302298 37936
rect 342162 37884 342168 37936
rect 342220 37924 342226 37936
rect 401594 37924 401600 37936
rect 342220 37896 401600 37924
rect 342220 37884 342226 37896
rect 401594 37884 401600 37896
rect 401652 37884 401658 37936
rect 424962 37884 424968 37936
rect 425020 37924 425026 37936
rect 485774 37924 485780 37936
rect 425020 37896 485780 37924
rect 425020 37884 425026 37896
rect 485774 37884 485780 37896
rect 485832 37884 485838 37936
rect 520090 37884 520096 37936
rect 520148 37924 520154 37936
rect 578878 37924 578884 37936
rect 520148 37896 578884 37924
rect 520148 37884 520154 37896
rect 578878 37884 578884 37896
rect 578936 37884 578942 37936
rect 177942 36660 177948 36712
rect 178000 36700 178006 36712
rect 237374 36700 237380 36712
rect 178000 36672 237380 36700
rect 178000 36660 178006 36672
rect 237374 36660 237380 36672
rect 237432 36660 237438 36712
rect 231670 36592 231676 36644
rect 231728 36632 231734 36644
rect 291194 36632 291200 36644
rect 231728 36604 291200 36632
rect 231728 36592 231734 36604
rect 291194 36592 291200 36604
rect 291252 36592 291258 36644
rect 328270 36592 328276 36644
rect 328328 36632 328334 36644
rect 387794 36632 387800 36644
rect 328328 36604 387800 36632
rect 328328 36592 328334 36604
rect 387794 36592 387800 36604
rect 387852 36592 387858 36644
rect 409782 36592 409788 36644
rect 409840 36632 409846 36644
rect 469214 36632 469220 36644
rect 409840 36604 469220 36632
rect 409840 36592 409846 36604
rect 469214 36592 469220 36604
rect 469272 36592 469278 36644
rect 124122 36524 124128 36576
rect 124180 36564 124186 36576
rect 183554 36564 183560 36576
rect 124180 36536 183560 36564
rect 124180 36524 124186 36536
rect 183554 36524 183560 36536
rect 183612 36524 183618 36576
rect 277302 36524 277308 36576
rect 277360 36564 277366 36576
rect 338114 36564 338120 36576
rect 277360 36536 338120 36564
rect 277360 36524 277366 36536
rect 338114 36524 338120 36536
rect 338172 36524 338178 36576
rect 378042 36524 378048 36576
rect 378100 36564 378106 36576
rect 437474 36564 437480 36576
rect 378100 36536 437480 36564
rect 378100 36524 378106 36536
rect 437474 36524 437480 36536
rect 437532 36524 437538 36576
rect 470502 36524 470508 36576
rect 470560 36564 470566 36576
rect 529934 36564 529940 36576
rect 470560 36536 529940 36564
rect 470560 36524 470566 36536
rect 529934 36524 529940 36536
rect 529992 36524 529998 36576
rect 3326 35844 3332 35896
rect 3384 35884 3390 35896
rect 59998 35884 60004 35896
rect 3384 35856 60004 35884
rect 3384 35844 3390 35856
rect 59998 35844 60004 35856
rect 60056 35844 60062 35896
rect 227622 35300 227628 35352
rect 227680 35340 227686 35352
rect 287054 35340 287060 35352
rect 227680 35312 287060 35340
rect 227680 35300 227686 35312
rect 287054 35300 287060 35312
rect 287112 35300 287118 35352
rect 324222 35300 324228 35352
rect 324280 35340 324286 35352
rect 383654 35340 383660 35352
rect 324280 35312 383660 35340
rect 324280 35300 324286 35312
rect 383654 35300 383660 35312
rect 383712 35300 383718 35352
rect 170950 35232 170956 35284
rect 171008 35272 171014 35284
rect 230474 35272 230480 35284
rect 171008 35244 230480 35272
rect 171008 35232 171014 35244
rect 230474 35232 230480 35244
rect 230532 35232 230538 35284
rect 373902 35232 373908 35284
rect 373960 35272 373966 35284
rect 433334 35272 433340 35284
rect 373960 35244 433340 35272
rect 373960 35232 373966 35244
rect 433334 35232 433340 35244
rect 433392 35232 433398 35284
rect 119982 35164 119988 35216
rect 120040 35204 120046 35216
rect 180794 35204 180800 35216
rect 120040 35176 180800 35204
rect 120040 35164 120046 35176
rect 180794 35164 180800 35176
rect 180852 35164 180858 35216
rect 274542 35164 274548 35216
rect 274600 35204 274606 35216
rect 333974 35204 333980 35216
rect 274600 35176 333980 35204
rect 274600 35164 274606 35176
rect 333974 35164 333980 35176
rect 334032 35164 334038 35216
rect 406930 35164 406936 35216
rect 406988 35204 406994 35216
rect 466454 35204 466460 35216
rect 406988 35176 466460 35204
rect 406988 35164 406994 35176
rect 466454 35164 466460 35176
rect 466512 35164 466518 35216
rect 467742 35164 467748 35216
rect 467800 35204 467806 35216
rect 527174 35204 527180 35216
rect 467800 35176 527180 35204
rect 467800 35164 467806 35176
rect 527174 35164 527180 35176
rect 527232 35164 527238 35216
rect 167638 33804 167644 33856
rect 167696 33844 167702 33856
rect 227806 33844 227812 33856
rect 167696 33816 227812 33844
rect 167696 33804 167702 33816
rect 227806 33804 227812 33816
rect 227864 33804 227870 33856
rect 270402 33804 270408 33856
rect 270460 33844 270466 33856
rect 331214 33844 331220 33856
rect 270460 33816 331220 33844
rect 270460 33804 270466 33816
rect 331214 33804 331220 33816
rect 331272 33804 331278 33856
rect 371878 33804 371884 33856
rect 371936 33844 371942 33856
rect 430574 33844 430580 33856
rect 371936 33816 430580 33844
rect 371936 33804 371942 33816
rect 430574 33804 430580 33816
rect 430632 33804 430638 33856
rect 117222 33736 117228 33788
rect 117280 33776 117286 33788
rect 176654 33776 176660 33788
rect 117280 33748 176660 33776
rect 117280 33736 117286 33748
rect 176654 33736 176660 33748
rect 176712 33736 176718 33788
rect 223390 33736 223396 33788
rect 223448 33776 223454 33788
rect 284294 33776 284300 33788
rect 223448 33748 284300 33776
rect 223448 33736 223454 33748
rect 284294 33736 284300 33748
rect 284352 33736 284358 33788
rect 320082 33736 320088 33788
rect 320140 33776 320146 33788
rect 380894 33776 380900 33788
rect 320140 33748 380900 33776
rect 320140 33736 320146 33748
rect 380894 33736 380900 33748
rect 380952 33736 380958 33788
rect 459370 33736 459376 33788
rect 459428 33776 459434 33788
rect 520366 33776 520372 33788
rect 459428 33748 520372 33776
rect 459428 33736 459434 33748
rect 520366 33736 520372 33748
rect 520424 33736 520430 33788
rect 317322 32512 317328 32564
rect 317380 32552 317386 32564
rect 376754 32552 376760 32564
rect 317380 32524 376760 32552
rect 317380 32512 317386 32524
rect 376754 32512 376760 32524
rect 376812 32512 376818 32564
rect 160002 32444 160008 32496
rect 160060 32484 160066 32496
rect 219434 32484 219440 32496
rect 160060 32456 219440 32484
rect 160060 32444 160066 32456
rect 219434 32444 219440 32456
rect 219492 32444 219498 32496
rect 267550 32444 267556 32496
rect 267608 32484 267614 32496
rect 327074 32484 327080 32496
rect 267608 32456 327080 32484
rect 267608 32444 267614 32456
rect 327074 32444 327080 32456
rect 327132 32444 327138 32496
rect 413922 32444 413928 32496
rect 413980 32484 413986 32496
rect 473354 32484 473360 32496
rect 413980 32456 473360 32484
rect 413980 32444 413986 32456
rect 473354 32444 473360 32456
rect 473412 32444 473418 32496
rect 110322 32376 110328 32428
rect 110380 32416 110386 32428
rect 169754 32416 169760 32428
rect 110380 32388 169760 32416
rect 110380 32376 110386 32388
rect 169754 32376 169760 32388
rect 169812 32376 169818 32428
rect 216582 32376 216588 32428
rect 216640 32416 216646 32428
rect 277394 32416 277400 32428
rect 216640 32388 277400 32416
rect 216640 32376 216646 32388
rect 277394 32376 277400 32388
rect 277452 32376 277458 32428
rect 367002 32376 367008 32428
rect 367060 32416 367066 32428
rect 426434 32416 426440 32428
rect 367060 32388 426440 32416
rect 367060 32376 367066 32388
rect 426434 32376 426440 32388
rect 426492 32376 426498 32428
rect 456702 32376 456708 32428
rect 456760 32416 456766 32428
rect 516134 32416 516140 32428
rect 456760 32388 516140 32416
rect 456760 32376 456766 32388
rect 516134 32376 516140 32388
rect 516192 32376 516198 32428
rect 306282 31152 306288 31204
rect 306340 31192 306346 31204
rect 365714 31192 365720 31204
rect 306340 31164 365720 31192
rect 306340 31152 306346 31164
rect 365714 31152 365720 31164
rect 365772 31152 365778 31204
rect 155862 31084 155868 31136
rect 155920 31124 155926 31136
rect 216674 31124 216680 31136
rect 155920 31096 216680 31124
rect 155920 31084 155926 31096
rect 216674 31084 216680 31096
rect 216732 31084 216738 31136
rect 259362 31084 259368 31136
rect 259420 31124 259426 31136
rect 320174 31124 320180 31136
rect 259420 31096 320180 31124
rect 259420 31084 259426 31096
rect 320174 31084 320180 31096
rect 320232 31084 320238 31136
rect 510522 31084 510528 31136
rect 510580 31124 510586 31136
rect 569954 31124 569960 31136
rect 510580 31096 569960 31124
rect 510580 31084 510586 31096
rect 569954 31084 569960 31096
rect 570012 31084 570018 31136
rect 106182 31016 106188 31068
rect 106240 31056 106246 31068
rect 167086 31056 167092 31068
rect 106240 31028 167092 31056
rect 106240 31016 106246 31028
rect 167086 31016 167092 31028
rect 167144 31016 167150 31068
rect 205450 31016 205456 31068
rect 205508 31056 205514 31068
rect 266354 31056 266360 31068
rect 205508 31028 266360 31056
rect 205508 31016 205514 31028
rect 266354 31016 266360 31028
rect 266412 31016 266418 31068
rect 362770 31016 362776 31068
rect 362828 31056 362834 31068
rect 423674 31056 423680 31068
rect 362828 31028 423680 31056
rect 362828 31016 362834 31028
rect 423674 31016 423680 31028
rect 423732 31016 423738 31068
rect 452562 31016 452568 31068
rect 452620 31056 452626 31068
rect 512086 31056 512092 31068
rect 452620 31028 512092 31056
rect 452620 31016 452626 31028
rect 512086 31016 512092 31028
rect 512144 31016 512150 31068
rect 523770 30268 523776 30320
rect 523828 30308 523834 30320
rect 580166 30308 580172 30320
rect 523828 30280 580172 30308
rect 523828 30268 523834 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 245562 29724 245568 29776
rect 245620 29764 245626 29776
rect 304994 29764 305000 29776
rect 245620 29736 305000 29764
rect 245620 29724 245626 29736
rect 304994 29724 305000 29736
rect 305052 29724 305058 29776
rect 153010 29656 153016 29708
rect 153068 29696 153074 29708
rect 212534 29696 212540 29708
rect 153068 29668 212540 29696
rect 153068 29656 153074 29668
rect 212534 29656 212540 29668
rect 212592 29656 212598 29708
rect 292482 29656 292488 29708
rect 292540 29696 292546 29708
rect 351914 29696 351920 29708
rect 292540 29668 351920 29696
rect 292540 29656 292546 29668
rect 351914 29656 351920 29668
rect 351972 29656 351978 29708
rect 402882 29656 402888 29708
rect 402940 29696 402946 29708
rect 462314 29696 462320 29708
rect 402940 29668 462320 29696
rect 402940 29656 402946 29668
rect 462314 29656 462320 29668
rect 462372 29656 462378 29708
rect 102042 29588 102048 29640
rect 102100 29628 102106 29640
rect 162854 29628 162860 29640
rect 102100 29600 162860 29628
rect 102100 29588 102106 29600
rect 162854 29588 162860 29600
rect 162912 29588 162918 29640
rect 191742 29588 191748 29640
rect 191800 29628 191806 29640
rect 252646 29628 252652 29640
rect 191800 29600 252652 29628
rect 191800 29588 191806 29600
rect 252646 29588 252652 29600
rect 252704 29588 252710 29640
rect 349062 29588 349068 29640
rect 349120 29628 349126 29640
rect 408586 29628 408592 29640
rect 349120 29600 408592 29628
rect 349120 29588 349126 29600
rect 408586 29588 408592 29600
rect 408644 29588 408650 29640
rect 441430 29588 441436 29640
rect 441488 29628 441494 29640
rect 502426 29628 502432 29640
rect 441488 29600 502432 29628
rect 441488 29588 441494 29600
rect 502426 29588 502432 29600
rect 502484 29588 502490 29640
rect 427906 29016 427912 29028
rect 427867 28988 427912 29016
rect 427906 28976 427912 28988
rect 427964 28976 427970 29028
rect 434806 29016 434812 29028
rect 434767 28988 434812 29016
rect 434806 28976 434812 28988
rect 434864 28976 434870 29028
rect 252462 28296 252468 28348
rect 252520 28336 252526 28348
rect 313366 28336 313372 28348
rect 252520 28308 313372 28336
rect 252520 28296 252526 28308
rect 313366 28296 313372 28308
rect 313424 28296 313430 28348
rect 353202 28296 353208 28348
rect 353260 28336 353266 28348
rect 412634 28336 412640 28348
rect 353260 28308 412640 28336
rect 353260 28296 353266 28308
rect 412634 28296 412640 28308
rect 412692 28296 412698 28348
rect 449710 28296 449716 28348
rect 449768 28336 449774 28348
rect 509234 28336 509240 28348
rect 449768 28308 509240 28336
rect 449768 28296 449774 28308
rect 509234 28296 509240 28308
rect 509292 28296 509298 28348
rect 97902 28228 97908 28280
rect 97960 28268 97966 28280
rect 158806 28268 158812 28280
rect 97960 28240 158812 28268
rect 97960 28228 97966 28240
rect 158806 28228 158812 28240
rect 158864 28228 158870 28280
rect 201402 28228 201408 28280
rect 201460 28268 201466 28280
rect 262306 28268 262312 28280
rect 201460 28240 262312 28268
rect 201460 28228 201466 28240
rect 262306 28228 262312 28240
rect 262364 28228 262370 28280
rect 302050 28228 302056 28280
rect 302108 28268 302114 28280
rect 362954 28268 362960 28280
rect 302108 28240 362960 28268
rect 302108 28228 302114 28240
rect 362954 28228 362960 28240
rect 363012 28228 363018 28280
rect 398742 28228 398748 28280
rect 398800 28268 398806 28280
rect 459646 28268 459652 28280
rect 398800 28240 459652 28268
rect 398800 28228 398806 28240
rect 459646 28228 459652 28240
rect 459704 28228 459710 28280
rect 506382 28228 506388 28280
rect 506440 28268 506446 28280
rect 565814 28268 565820 28280
rect 506440 28240 565820 28268
rect 506440 28228 506446 28240
rect 565814 28228 565820 28240
rect 565872 28228 565878 28280
rect 369854 27548 369860 27600
rect 369912 27588 369918 27600
rect 370498 27588 370504 27600
rect 369912 27560 370504 27588
rect 369912 27548 369918 27560
rect 370498 27548 370504 27560
rect 370556 27548 370562 27600
rect 445662 27004 445668 27056
rect 445720 27044 445726 27056
rect 505094 27044 505100 27056
rect 445720 27016 505100 27044
rect 445720 27004 445726 27016
rect 505094 27004 505100 27016
rect 505152 27004 505158 27056
rect 272518 26936 272524 26988
rect 272576 26976 272582 26988
rect 331306 26976 331312 26988
rect 272576 26948 331312 26976
rect 272576 26936 272582 26948
rect 331306 26936 331312 26948
rect 331364 26936 331370 26988
rect 391842 26936 391848 26988
rect 391900 26976 391906 26988
rect 451274 26976 451280 26988
rect 391900 26948 451280 26976
rect 391900 26936 391906 26948
rect 451274 26936 451280 26948
rect 451332 26936 451338 26988
rect 93762 26868 93768 26920
rect 93820 26908 93826 26920
rect 154574 26908 154580 26920
rect 93820 26880 154580 26908
rect 93820 26868 93826 26880
rect 154574 26868 154580 26880
rect 154632 26868 154638 26920
rect 165522 26868 165528 26920
rect 165580 26908 165586 26920
rect 226334 26908 226340 26920
rect 165580 26880 226340 26908
rect 165580 26868 165586 26880
rect 226334 26868 226340 26880
rect 226392 26868 226398 26920
rect 244182 26868 244188 26920
rect 244240 26908 244246 26920
rect 305086 26908 305092 26920
rect 244240 26880 305092 26908
rect 244240 26868 244246 26880
rect 305086 26868 305092 26880
rect 305144 26868 305150 26920
rect 344830 26868 344836 26920
rect 344888 26908 344894 26920
rect 404354 26908 404360 26920
rect 344888 26880 404360 26908
rect 344888 26868 344894 26880
rect 404354 26868 404360 26880
rect 404412 26868 404418 26920
rect 502150 26868 502156 26920
rect 502208 26908 502214 26920
rect 563146 26908 563152 26920
rect 502208 26880 563152 26908
rect 502208 26868 502214 26880
rect 563146 26868 563152 26880
rect 563204 26868 563210 26920
rect 438762 25644 438768 25696
rect 438820 25684 438826 25696
rect 498194 25684 498200 25696
rect 438820 25656 498200 25684
rect 438820 25644 438826 25656
rect 498194 25644 498200 25656
rect 498252 25644 498258 25696
rect 237282 25576 237288 25628
rect 237340 25616 237346 25628
rect 296806 25616 296812 25628
rect 237340 25588 296812 25616
rect 237340 25576 237346 25588
rect 296806 25576 296812 25588
rect 296864 25576 296870 25628
rect 395982 25576 395988 25628
rect 396040 25616 396046 25628
rect 455414 25616 455420 25628
rect 396040 25588 455420 25616
rect 396040 25576 396046 25588
rect 455414 25576 455420 25588
rect 455472 25576 455478 25628
rect 91002 25508 91008 25560
rect 91060 25548 91066 25560
rect 150526 25548 150532 25560
rect 91060 25520 150532 25548
rect 91060 25508 91066 25520
rect 150526 25508 150532 25520
rect 150584 25508 150590 25560
rect 158622 25508 158628 25560
rect 158680 25548 158686 25560
rect 218146 25548 218152 25560
rect 158680 25520 218152 25548
rect 158680 25508 158686 25520
rect 218146 25508 218152 25520
rect 218204 25508 218210 25560
rect 267642 25508 267648 25560
rect 267700 25548 267706 25560
rect 328546 25548 328552 25560
rect 267700 25520 328552 25548
rect 267700 25508 267706 25520
rect 328546 25508 328552 25520
rect 328604 25508 328610 25560
rect 336550 25508 336556 25560
rect 336608 25548 336614 25560
rect 397546 25548 397552 25560
rect 336608 25520 397552 25548
rect 336608 25508 336614 25520
rect 397546 25508 397552 25520
rect 397604 25508 397610 25560
rect 495342 25508 495348 25560
rect 495400 25548 495406 25560
rect 554866 25548 554872 25560
rect 495400 25520 554872 25548
rect 495400 25508 495406 25520
rect 554866 25508 554872 25520
rect 554924 25508 554930 25560
rect 275830 24148 275836 24200
rect 275888 24188 275894 24200
rect 335354 24188 335360 24200
rect 275888 24160 335360 24188
rect 275888 24148 275894 24160
rect 335354 24148 335360 24160
rect 335412 24148 335418 24200
rect 360102 24148 360108 24200
rect 360160 24188 360166 24200
rect 419534 24188 419540 24200
rect 360160 24160 419540 24188
rect 360160 24148 360166 24160
rect 419534 24148 419540 24160
rect 419592 24148 419598 24200
rect 492582 24148 492588 24200
rect 492640 24188 492646 24200
rect 552014 24188 552020 24200
rect 492640 24160 552020 24188
rect 492640 24148 492646 24160
rect 552014 24148 552020 24160
rect 552072 24148 552078 24200
rect 86862 24080 86868 24132
rect 86920 24120 86926 24132
rect 147674 24120 147680 24132
rect 86920 24092 147680 24120
rect 86920 24080 86926 24092
rect 147674 24080 147680 24092
rect 147732 24080 147738 24132
rect 154482 24080 154488 24132
rect 154540 24120 154546 24132
rect 215294 24120 215300 24132
rect 154540 24092 215300 24120
rect 154540 24080 154546 24092
rect 215294 24080 215300 24092
rect 215352 24080 215358 24132
rect 226242 24080 226248 24132
rect 226300 24120 226306 24132
rect 287146 24120 287152 24132
rect 226300 24092 287152 24120
rect 226300 24080 226306 24092
rect 287146 24080 287152 24092
rect 287204 24080 287210 24132
rect 304902 24080 304908 24132
rect 304960 24120 304966 24132
rect 365806 24120 365812 24132
rect 304960 24092 365812 24120
rect 304960 24080 304966 24092
rect 365806 24080 365812 24092
rect 365864 24080 365870 24132
rect 434622 24080 434628 24132
rect 434680 24120 434686 24132
rect 494146 24120 494152 24132
rect 434680 24092 494152 24120
rect 434680 24080 434686 24092
rect 494146 24080 494152 24092
rect 494204 24080 494210 24132
rect 335262 22788 335268 22840
rect 335320 22828 335326 22840
rect 394786 22828 394792 22840
rect 335320 22800 394792 22828
rect 335320 22788 335326 22800
rect 394786 22788 394792 22800
rect 394844 22788 394850 22840
rect 431862 22788 431868 22840
rect 431920 22828 431926 22840
rect 491294 22828 491300 22840
rect 431920 22800 491300 22828
rect 431920 22788 431926 22800
rect 491294 22788 491300 22800
rect 491352 22788 491358 22840
rect 84010 22720 84016 22772
rect 84068 22760 84074 22772
rect 143534 22760 143540 22772
rect 84068 22732 143540 22760
rect 84068 22720 84074 22732
rect 143534 22720 143540 22732
rect 143592 22720 143598 22772
rect 151722 22720 151728 22772
rect 151780 22760 151786 22772
rect 211154 22760 211160 22772
rect 151780 22732 211160 22760
rect 151780 22720 151786 22732
rect 211154 22720 211160 22732
rect 211212 22720 211218 22772
rect 215110 22720 215116 22772
rect 215168 22760 215174 22772
rect 276014 22760 276020 22772
rect 215168 22732 276020 22760
rect 215168 22720 215174 22732
rect 276014 22720 276020 22732
rect 276072 22720 276078 22772
rect 286962 22720 286968 22772
rect 287020 22760 287026 22772
rect 347866 22760 347872 22772
rect 287020 22732 347872 22760
rect 287020 22720 287026 22732
rect 347866 22720 347872 22732
rect 347924 22720 347930 22772
rect 488442 22720 488448 22772
rect 488500 22760 488506 22772
rect 547874 22760 547880 22772
rect 488500 22732 547880 22760
rect 488500 22720 488506 22732
rect 547874 22720 547880 22732
rect 547932 22720 547938 22772
rect 427722 21428 427728 21480
rect 427780 21468 427786 21480
rect 487154 21468 487160 21480
rect 427780 21440 487160 21468
rect 427780 21428 427786 21440
rect 487154 21428 487160 21440
rect 487212 21428 487218 21480
rect 79962 21360 79968 21412
rect 80020 21400 80026 21412
rect 140866 21400 140872 21412
rect 80020 21372 140872 21400
rect 80020 21360 80026 21372
rect 140866 21360 140872 21372
rect 140924 21360 140930 21412
rect 147582 21360 147588 21412
rect 147640 21400 147646 21412
rect 208394 21400 208400 21412
rect 147640 21372 208400 21400
rect 147640 21360 147646 21372
rect 208394 21360 208400 21372
rect 208452 21360 208458 21412
rect 212442 21360 212448 21412
rect 212500 21400 212506 21412
rect 271874 21400 271880 21412
rect 212500 21372 271880 21400
rect 212500 21360 212506 21372
rect 271874 21360 271880 21372
rect 271932 21360 271938 21412
rect 273162 21360 273168 21412
rect 273220 21400 273226 21412
rect 332594 21400 332600 21412
rect 273220 21372 332600 21400
rect 273220 21360 273226 21372
rect 332594 21360 332600 21372
rect 332652 21360 332658 21412
rect 333882 21360 333888 21412
rect 333940 21400 333946 21412
rect 393314 21400 393320 21412
rect 333940 21372 393320 21400
rect 333940 21360 333946 21372
rect 393314 21360 393320 21372
rect 393372 21360 393378 21412
rect 485590 21360 485596 21412
rect 485648 21400 485654 21412
rect 545114 21400 545120 21412
rect 485648 21372 545120 21400
rect 485648 21360 485654 21372
rect 545114 21360 545120 21372
rect 545172 21360 545178 21412
rect 481542 20000 481548 20052
rect 481600 20040 481606 20052
rect 540974 20040 540980 20052
rect 481600 20012 540980 20040
rect 481600 20000 481606 20012
rect 540974 20000 540980 20012
rect 541032 20000 541038 20052
rect 75822 19932 75828 19984
rect 75880 19972 75886 19984
rect 136634 19972 136640 19984
rect 75880 19944 136640 19972
rect 75880 19932 75886 19944
rect 136634 19932 136640 19944
rect 136692 19932 136698 19984
rect 144822 19932 144828 19984
rect 144880 19972 144886 19984
rect 204254 19972 204260 19984
rect 144880 19944 204260 19972
rect 144880 19932 144886 19944
rect 204254 19932 204260 19944
rect 204312 19932 204318 19984
rect 205542 19932 205548 19984
rect 205600 19972 205606 19984
rect 264974 19972 264980 19984
rect 205600 19944 264980 19972
rect 205600 19932 205606 19944
rect 264974 19932 264980 19944
rect 265032 19932 265038 19984
rect 266262 19932 266268 19984
rect 266320 19972 266326 19984
rect 325694 19972 325700 19984
rect 266320 19944 325700 19972
rect 266320 19932 266326 19944
rect 325694 19932 325700 19944
rect 325752 19932 325758 19984
rect 326982 19932 326988 19984
rect 327040 19972 327046 19984
rect 386414 19972 386420 19984
rect 327040 19944 386420 19972
rect 327040 19932 327046 19944
rect 386414 19932 386420 19944
rect 386472 19932 386478 19984
rect 423490 19932 423496 19984
rect 423548 19972 423554 19984
rect 484394 19972 484400 19984
rect 423548 19944 484400 19972
rect 423548 19932 423554 19944
rect 484394 19932 484400 19944
rect 484452 19932 484458 19984
rect 328454 19252 328460 19304
rect 328512 19292 328518 19304
rect 394694 19292 394700 19304
rect 328512 19264 328557 19292
rect 394655 19264 394700 19292
rect 328512 19252 328518 19264
rect 394694 19252 394700 19264
rect 394752 19252 394758 19304
rect 397454 19292 397460 19304
rect 397415 19264 397460 19292
rect 397454 19252 397460 19264
rect 397512 19252 397518 19304
rect 427906 19292 427912 19304
rect 427867 19264 427912 19292
rect 427906 19252 427912 19264
rect 427964 19252 427970 19304
rect 434806 19292 434812 19304
rect 434767 19264 434812 19292
rect 434806 19252 434812 19264
rect 434864 19252 434870 19304
rect 269022 18640 269028 18692
rect 269080 18680 269086 18692
rect 330021 18683 330079 18689
rect 330021 18680 330033 18683
rect 269080 18652 330033 18680
rect 269080 18640 269086 18652
rect 330021 18649 330033 18652
rect 330067 18649 330079 18683
rect 330021 18643 330079 18649
rect 73062 18572 73068 18624
rect 73120 18612 73126 18624
rect 132586 18612 132592 18624
rect 73120 18584 132592 18612
rect 73120 18572 73126 18584
rect 132586 18572 132592 18584
rect 132644 18572 132650 18624
rect 140682 18572 140688 18624
rect 140740 18612 140746 18624
rect 201586 18612 201592 18624
rect 140740 18584 201592 18612
rect 140740 18572 140746 18584
rect 201586 18572 201592 18584
rect 201644 18572 201650 18624
rect 208302 18572 208308 18624
rect 208360 18612 208366 18624
rect 269114 18612 269120 18624
rect 208360 18584 269120 18612
rect 208360 18572 208366 18584
rect 269114 18572 269120 18584
rect 269172 18572 269178 18624
rect 330478 18572 330484 18624
rect 330536 18612 330542 18624
rect 390646 18612 390652 18624
rect 330536 18584 390652 18612
rect 330536 18572 330542 18584
rect 390646 18572 390652 18584
rect 390704 18572 390710 18624
rect 412542 18572 412548 18624
rect 412600 18612 412606 18624
rect 471974 18612 471980 18624
rect 412600 18584 471980 18612
rect 412600 18572 412606 18584
rect 471974 18572 471980 18584
rect 472032 18572 472038 18624
rect 474642 18572 474648 18624
rect 474700 18612 474706 18624
rect 534074 18612 534080 18624
rect 474700 18584 534080 18612
rect 474700 18572 474706 18584
rect 534074 18572 534080 18584
rect 534132 18572 534138 18624
rect 523862 17892 523868 17944
rect 523920 17932 523926 17944
rect 579798 17932 579804 17944
rect 523920 17904 579804 17932
rect 523920 17892 523926 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 129642 17212 129648 17264
rect 129700 17252 129706 17264
rect 190454 17252 190460 17264
rect 129700 17224 190460 17252
rect 129700 17212 129706 17224
rect 190454 17212 190460 17224
rect 190512 17212 190518 17264
rect 197170 17212 197176 17264
rect 197228 17252 197234 17264
rect 258074 17252 258080 17264
rect 197228 17224 258080 17252
rect 197228 17212 197234 17224
rect 258074 17212 258080 17224
rect 258132 17212 258138 17264
rect 262122 17212 262128 17264
rect 262180 17252 262186 17264
rect 321646 17252 321652 17264
rect 262180 17224 321652 17252
rect 262180 17212 262186 17224
rect 321646 17212 321652 17224
rect 321704 17212 321710 17264
rect 322842 17212 322848 17264
rect 322900 17252 322906 17264
rect 382366 17252 382372 17264
rect 322900 17224 382372 17252
rect 322900 17212 322906 17224
rect 382366 17212 382372 17224
rect 382424 17212 382430 17264
rect 408402 17212 408408 17264
rect 408460 17252 408466 17264
rect 467834 17252 467840 17264
rect 408460 17224 467840 17252
rect 408460 17212 408466 17224
rect 467834 17212 467840 17224
rect 467892 17212 467898 17264
rect 126882 15920 126888 15972
rect 126940 15960 126946 15972
rect 186314 15960 186320 15972
rect 126940 15932 186320 15960
rect 126940 15920 126946 15932
rect 186314 15920 186320 15932
rect 186372 15920 186378 15972
rect 318610 15920 318616 15972
rect 318668 15960 318674 15972
rect 379514 15960 379520 15972
rect 318668 15932 379520 15960
rect 318668 15920 318674 15932
rect 379514 15920 379520 15932
rect 379572 15920 379578 15972
rect 66898 15852 66904 15904
rect 66956 15892 66962 15904
rect 126974 15892 126980 15904
rect 66956 15864 126980 15892
rect 66956 15852 66962 15864
rect 126974 15852 126980 15864
rect 127032 15852 127038 15904
rect 194502 15852 194508 15904
rect 194560 15892 194566 15904
rect 253934 15892 253940 15904
rect 194560 15864 253940 15892
rect 194560 15852 194566 15864
rect 253934 15852 253940 15864
rect 253992 15852 253998 15904
rect 257890 15852 257896 15904
rect 257948 15892 257954 15904
rect 318794 15892 318800 15904
rect 257948 15864 318800 15892
rect 257948 15852 257954 15864
rect 318794 15852 318800 15864
rect 318852 15852 318858 15904
rect 405642 15852 405648 15904
rect 405700 15892 405706 15904
rect 465074 15892 465080 15904
rect 405700 15864 465080 15892
rect 405700 15852 405706 15864
rect 465074 15852 465080 15864
rect 465132 15852 465138 15904
rect 505002 15852 505008 15904
rect 505060 15892 505066 15904
rect 564434 15892 564440 15904
rect 505060 15864 564440 15892
rect 505060 15852 505066 15864
rect 564434 15852 564440 15864
rect 564492 15852 564498 15904
rect 122742 14424 122748 14476
rect 122800 14464 122806 14476
rect 183646 14464 183652 14476
rect 122800 14436 183652 14464
rect 122800 14424 122806 14436
rect 183646 14424 183652 14436
rect 183704 14424 183710 14476
rect 187602 14424 187608 14476
rect 187660 14464 187666 14476
rect 247034 14464 247040 14476
rect 187660 14436 247040 14464
rect 187660 14424 187666 14436
rect 247034 14424 247040 14436
rect 247092 14424 247098 14476
rect 248322 14424 248328 14476
rect 248380 14464 248386 14476
rect 307754 14464 307760 14476
rect 248380 14436 307760 14464
rect 248380 14424 248386 14436
rect 307754 14424 307760 14436
rect 307812 14424 307818 14476
rect 309042 14424 309048 14476
rect 309100 14464 309106 14476
rect 368474 14464 368480 14476
rect 309100 14436 368480 14464
rect 309100 14424 309106 14436
rect 368474 14424 368480 14436
rect 368532 14424 368538 14476
rect 397362 14424 397368 14476
rect 397420 14464 397426 14476
rect 458174 14464 458180 14476
rect 397420 14436 458180 14464
rect 397420 14424 397426 14436
rect 458174 14424 458180 14436
rect 458232 14424 458238 14476
rect 469122 14424 469128 14476
rect 469180 14464 469186 14476
rect 528646 14464 528652 14476
rect 469180 14436 528652 14464
rect 469180 14424 469186 14436
rect 528646 14424 528652 14436
rect 528704 14424 528710 14476
rect 118510 13064 118516 13116
rect 118568 13104 118574 13116
rect 179414 13104 179420 13116
rect 118568 13076 179420 13104
rect 118568 13064 118574 13076
rect 179414 13064 179420 13076
rect 179472 13064 179478 13116
rect 183462 13064 183468 13116
rect 183520 13104 183526 13116
rect 244366 13104 244372 13116
rect 183520 13076 244372 13104
rect 183520 13064 183526 13076
rect 244366 13064 244372 13076
rect 244424 13064 244430 13116
rect 251082 13064 251088 13116
rect 251140 13104 251146 13116
rect 311894 13104 311900 13116
rect 251140 13076 311900 13104
rect 251140 13064 251146 13076
rect 311894 13064 311900 13076
rect 311952 13064 311958 13116
rect 315942 13064 315948 13116
rect 316000 13104 316006 13116
rect 375374 13104 375380 13116
rect 316000 13076 375380 13104
rect 316000 13064 316006 13076
rect 375374 13064 375380 13076
rect 375432 13064 375438 13116
rect 384298 13064 384304 13116
rect 384356 13104 384362 13116
rect 443086 13104 443092 13116
rect 384356 13076 443092 13104
rect 384356 13064 384362 13076
rect 443086 13064 443092 13076
rect 443144 13064 443150 13116
rect 448422 13064 448428 13116
rect 448480 13104 448486 13116
rect 507854 13104 507860 13116
rect 448480 13076 507860 13104
rect 448480 13064 448486 13076
rect 507854 13064 507860 13076
rect 507912 13064 507918 13116
rect 322934 12452 322940 12504
rect 322992 12452 322998 12504
rect 325694 12452 325700 12504
rect 325752 12452 325758 12504
rect 327074 12452 327080 12504
rect 327132 12452 327138 12504
rect 322952 12424 322980 12452
rect 324038 12424 324044 12436
rect 322952 12396 324044 12424
rect 324038 12384 324044 12396
rect 324096 12384 324102 12436
rect 325712 12424 325740 12452
rect 326430 12424 326436 12436
rect 325712 12396 326436 12424
rect 326430 12384 326436 12396
rect 326488 12384 326494 12436
rect 327092 12356 327120 12452
rect 375374 12384 375380 12436
rect 375432 12424 375438 12436
rect 376386 12424 376392 12436
rect 375432 12396 376392 12424
rect 375432 12384 375438 12396
rect 376386 12384 376392 12396
rect 376444 12384 376450 12436
rect 376754 12384 376760 12436
rect 376812 12424 376818 12436
rect 377582 12424 377588 12436
rect 376812 12396 377588 12424
rect 376812 12384 376818 12396
rect 377582 12384 377588 12396
rect 377640 12384 377646 12436
rect 393314 12384 393320 12436
rect 393372 12424 393378 12436
rect 394234 12424 394240 12436
rect 393372 12396 394240 12424
rect 393372 12384 393378 12396
rect 394234 12384 394240 12396
rect 394292 12384 394298 12436
rect 408586 12384 408592 12436
rect 408644 12424 408650 12436
rect 409690 12424 409696 12436
rect 408644 12396 409696 12424
rect 408644 12384 408650 12396
rect 409690 12384 409696 12396
rect 409748 12384 409754 12436
rect 412634 12384 412640 12436
rect 412692 12424 412698 12436
rect 413278 12424 413284 12436
rect 412692 12396 413284 12424
rect 412692 12384 412698 12396
rect 413278 12384 413284 12396
rect 413336 12384 413342 12436
rect 327626 12356 327632 12368
rect 327092 12328 327632 12356
rect 327626 12316 327632 12328
rect 327684 12316 327690 12368
rect 302142 11772 302148 11824
rect 302200 11812 302206 11824
rect 361574 11812 361580 11824
rect 302200 11784 361580 11812
rect 302200 11772 302206 11784
rect 361574 11772 361580 11784
rect 361632 11772 361638 11824
rect 115842 11704 115848 11756
rect 115900 11744 115906 11756
rect 175366 11744 175372 11756
rect 115900 11716 175372 11744
rect 115900 11704 115906 11716
rect 175366 11704 175372 11716
rect 175424 11704 175430 11756
rect 179230 11704 179236 11756
rect 179288 11744 179294 11756
rect 240134 11744 240140 11756
rect 179288 11716 240140 11744
rect 179288 11704 179294 11716
rect 240134 11704 240140 11716
rect 240192 11704 240198 11756
rect 241422 11704 241428 11756
rect 241480 11744 241486 11756
rect 300854 11744 300860 11756
rect 241480 11716 300860 11744
rect 241480 11704 241486 11716
rect 300854 11704 300860 11716
rect 300912 11704 300918 11756
rect 303522 11704 303528 11756
rect 303580 11744 303586 11756
rect 364334 11744 364340 11756
rect 303580 11716 364340 11744
rect 303580 11704 303586 11716
rect 364334 11704 364340 11716
rect 364392 11704 364398 11756
rect 376662 11704 376668 11756
rect 376720 11744 376726 11756
rect 437014 11744 437020 11756
rect 376720 11716 437020 11744
rect 376720 11704 376726 11716
rect 437014 11704 437020 11716
rect 437072 11704 437078 11756
rect 444282 11704 444288 11756
rect 444340 11744 444346 11756
rect 503714 11744 503720 11756
rect 444340 11716 503720 11744
rect 444340 11704 444346 11716
rect 503714 11704 503720 11716
rect 503772 11704 503778 11756
rect 176562 10344 176568 10396
rect 176620 10384 176626 10396
rect 236086 10384 236092 10396
rect 176620 10356 236092 10384
rect 176620 10344 176626 10356
rect 236086 10344 236092 10356
rect 236144 10344 236150 10396
rect 285582 10344 285588 10396
rect 285640 10384 285646 10396
rect 346394 10384 346400 10396
rect 285640 10356 346400 10384
rect 285640 10344 285646 10356
rect 346394 10344 346400 10356
rect 346452 10344 346458 10396
rect 441522 10344 441528 10396
rect 441580 10384 441586 10396
rect 500954 10384 500960 10396
rect 441580 10356 500960 10384
rect 441580 10344 441586 10356
rect 500954 10344 500960 10356
rect 501012 10344 501018 10396
rect 111702 10276 111708 10328
rect 111760 10316 111766 10328
rect 172514 10316 172520 10328
rect 111760 10288 172520 10316
rect 111760 10276 111766 10288
rect 172514 10276 172520 10288
rect 172572 10276 172578 10328
rect 233142 10276 233148 10328
rect 233200 10316 233206 10328
rect 293954 10316 293960 10328
rect 233200 10288 293960 10316
rect 233200 10276 233206 10288
rect 293954 10276 293960 10288
rect 294012 10276 294018 10328
rect 298002 10276 298008 10328
rect 298060 10316 298066 10328
rect 357434 10316 357440 10328
rect 298060 10288 357440 10316
rect 298060 10276 298066 10288
rect 357434 10276 357440 10288
rect 357492 10276 357498 10328
rect 367738 10276 367744 10328
rect 367796 10316 367802 10328
rect 415394 10316 415400 10328
rect 367796 10288 415400 10316
rect 367796 10276 367802 10288
rect 415394 10276 415400 10288
rect 415452 10276 415458 10328
rect 416682 10276 416688 10328
rect 416740 10316 416746 10328
rect 477586 10316 477592 10328
rect 416740 10288 477592 10316
rect 416740 10276 416746 10288
rect 477586 10276 477592 10288
rect 477644 10276 477650 10328
rect 516042 10276 516048 10328
rect 516100 10316 516106 10328
rect 575474 10316 575480 10328
rect 516100 10288 575480 10316
rect 516100 10276 516106 10288
rect 575474 10276 575480 10288
rect 575532 10276 575538 10328
rect 434806 9772 434812 9784
rect 434767 9744 434812 9772
rect 434806 9732 434812 9744
rect 434864 9732 434870 9784
rect 328457 9707 328515 9713
rect 328457 9673 328469 9707
rect 328503 9704 328515 9707
rect 328822 9704 328828 9716
rect 328503 9676 328828 9704
rect 328503 9673 328515 9676
rect 328457 9667 328515 9673
rect 328822 9664 328828 9676
rect 328880 9664 328886 9716
rect 330018 9704 330024 9716
rect 329979 9676 330024 9704
rect 330018 9664 330024 9676
rect 330076 9664 330082 9716
rect 394697 9707 394755 9713
rect 394697 9673 394709 9707
rect 394743 9704 394755 9707
rect 395430 9704 395436 9716
rect 394743 9676 395436 9704
rect 394743 9673 394755 9676
rect 394697 9667 394755 9673
rect 395430 9664 395436 9676
rect 395488 9664 395494 9716
rect 397457 9707 397515 9713
rect 397457 9673 397469 9707
rect 397503 9704 397515 9707
rect 397822 9704 397828 9716
rect 397503 9676 397828 9704
rect 397503 9673 397515 9676
rect 397457 9667 397515 9673
rect 397822 9664 397828 9676
rect 397880 9664 397886 9716
rect 427906 9704 427912 9716
rect 427867 9676 427912 9704
rect 427906 9664 427912 9676
rect 427964 9664 427970 9716
rect 324038 9596 324044 9648
rect 324096 9596 324102 9648
rect 326430 9596 326436 9648
rect 326488 9596 326494 9648
rect 327626 9596 327632 9648
rect 327684 9596 327690 9648
rect 430574 9596 430580 9648
rect 430632 9636 430638 9648
rect 431129 9639 431187 9645
rect 431129 9636 431141 9639
rect 430632 9608 431141 9636
rect 430632 9596 430638 9608
rect 431129 9605 431141 9608
rect 431175 9605 431187 9639
rect 431129 9599 431187 9605
rect 434806 9596 434812 9648
rect 434864 9636 434870 9648
rect 435821 9639 435879 9645
rect 435821 9636 435833 9639
rect 434864 9608 435833 9636
rect 434864 9596 434870 9608
rect 435821 9605 435833 9608
rect 435867 9605 435879 9639
rect 435821 9599 435879 9605
rect 324056 9512 324084 9596
rect 326448 9512 326476 9596
rect 327644 9512 327672 9596
rect 324038 9460 324044 9512
rect 324096 9460 324102 9512
rect 326430 9460 326436 9512
rect 326488 9460 326494 9512
rect 327626 9460 327632 9512
rect 327684 9460 327690 9512
rect 230382 8984 230388 9036
rect 230440 9024 230446 9036
rect 290734 9024 290740 9036
rect 230440 8996 290740 9024
rect 230440 8984 230446 8996
rect 290734 8984 290740 8996
rect 290792 8984 290798 9036
rect 108942 8916 108948 8968
rect 109000 8956 109006 8968
rect 169386 8956 169392 8968
rect 109000 8928 169392 8956
rect 109000 8916 109006 8928
rect 169386 8916 169392 8928
rect 169444 8916 169450 8968
rect 172422 8916 172428 8968
rect 172480 8956 172486 8968
rect 233694 8956 233700 8968
rect 172480 8928 233700 8956
rect 172480 8916 172486 8928
rect 233694 8916 233700 8928
rect 233752 8916 233758 8968
rect 291102 8916 291108 8968
rect 291160 8956 291166 8968
rect 351362 8956 351368 8968
rect 291160 8928 351368 8956
rect 291160 8916 291166 8928
rect 351362 8916 351368 8928
rect 351420 8916 351426 8968
rect 351822 8916 351828 8968
rect 351880 8956 351886 8968
rect 412082 8956 412088 8968
rect 351880 8928 412088 8956
rect 351880 8916 351886 8928
rect 412082 8916 412088 8928
rect 412140 8916 412146 8968
rect 430482 8916 430488 8968
rect 430540 8956 430546 8968
rect 490558 8956 490564 8968
rect 430540 8928 490564 8956
rect 430540 8916 430546 8928
rect 490558 8916 490564 8928
rect 490616 8916 490622 8968
rect 499482 8916 499488 8968
rect 499540 8956 499546 8968
rect 559558 8956 559564 8968
rect 499540 8928 559564 8956
rect 499540 8916 499546 8928
rect 559558 8916 559564 8928
rect 559616 8916 559622 8968
rect 325234 7732 325240 7744
rect 321572 7704 325240 7732
rect 104802 7624 104808 7676
rect 104860 7664 104866 7676
rect 165890 7664 165896 7676
rect 104860 7636 165896 7664
rect 104860 7624 104866 7636
rect 165890 7624 165896 7636
rect 165948 7624 165954 7676
rect 169662 7624 169668 7676
rect 169720 7664 169726 7676
rect 230106 7664 230112 7676
rect 169720 7636 230112 7664
rect 169720 7624 169726 7636
rect 230106 7624 230112 7636
rect 230164 7624 230170 7676
rect 264882 7624 264888 7676
rect 264940 7664 264946 7676
rect 321572 7664 321600 7704
rect 325234 7692 325240 7704
rect 325292 7692 325298 7744
rect 264940 7636 321600 7664
rect 264940 7624 264946 7636
rect 321646 7624 321652 7676
rect 321704 7664 321710 7676
rect 322842 7664 322848 7676
rect 321704 7636 322848 7664
rect 321704 7624 321710 7636
rect 322842 7624 322848 7636
rect 322900 7624 322906 7676
rect 340782 7624 340788 7676
rect 340840 7664 340846 7676
rect 401318 7664 401324 7676
rect 340840 7636 401324 7664
rect 340840 7624 340846 7636
rect 401318 7624 401324 7636
rect 401376 7624 401382 7676
rect 433334 7624 433340 7676
rect 433392 7664 433398 7676
rect 434622 7664 434628 7676
rect 433392 7636 434628 7664
rect 433392 7624 433398 7636
rect 434622 7624 434628 7636
rect 434680 7624 434686 7676
rect 482278 7624 482284 7676
rect 482336 7664 482342 7676
rect 538122 7664 538128 7676
rect 482336 7636 538128 7664
rect 482336 7624 482342 7636
rect 538122 7624 538128 7636
rect 538180 7624 538186 7676
rect 137922 7556 137928 7608
rect 137980 7596 137986 7608
rect 199194 7596 199200 7608
rect 137980 7568 199200 7596
rect 137980 7556 137986 7568
rect 199194 7556 199200 7568
rect 199252 7556 199258 7608
rect 223482 7556 223488 7608
rect 223540 7596 223546 7608
rect 283650 7596 283656 7608
rect 223540 7568 283656 7596
rect 223540 7556 223546 7568
rect 283650 7556 283656 7568
rect 283708 7556 283714 7608
rect 284202 7556 284208 7608
rect 284260 7596 284266 7608
rect 344278 7596 344284 7608
rect 284260 7568 344284 7596
rect 284260 7556 284266 7568
rect 344278 7556 344284 7568
rect 344336 7556 344342 7608
rect 390554 7556 390560 7608
rect 390612 7596 390618 7608
rect 391842 7596 391848 7608
rect 390612 7568 391848 7596
rect 390612 7556 390618 7568
rect 391842 7556 391848 7568
rect 391900 7556 391906 7608
rect 423582 7556 423588 7608
rect 423640 7596 423646 7608
rect 483474 7596 483480 7608
rect 423640 7568 483480 7596
rect 423640 7556 423646 7568
rect 483474 7556 483480 7568
rect 483532 7556 483538 7608
rect 162762 6264 162768 6316
rect 162820 6304 162826 6316
rect 222930 6304 222936 6316
rect 162820 6276 222936 6304
rect 162820 6264 162826 6276
rect 222930 6264 222936 6276
rect 222988 6264 222994 6316
rect 219342 6196 219348 6248
rect 219400 6236 219406 6248
rect 279970 6236 279976 6248
rect 219400 6208 279976 6236
rect 219400 6196 219406 6208
rect 279970 6196 279976 6208
rect 280028 6196 280034 6248
rect 282822 6196 282828 6248
rect 282880 6236 282886 6248
rect 343082 6236 343088 6248
rect 282880 6208 343088 6236
rect 282880 6196 282886 6208
rect 343082 6196 343088 6208
rect 343140 6196 343146 6248
rect 345658 6196 345664 6248
rect 345716 6236 345722 6248
rect 372798 6236 372804 6248
rect 345716 6208 372804 6236
rect 345716 6196 345722 6208
rect 372798 6196 372804 6208
rect 372856 6196 372862 6248
rect 100570 6128 100576 6180
rect 100628 6168 100634 6180
rect 162302 6168 162308 6180
rect 100628 6140 162308 6168
rect 100628 6128 100634 6140
rect 162302 6128 162308 6140
rect 162360 6128 162366 6180
rect 209682 6128 209688 6180
rect 209740 6168 209746 6180
rect 270586 6168 270592 6180
rect 209740 6140 270592 6168
rect 209740 6128 209746 6140
rect 270586 6128 270592 6140
rect 270644 6128 270650 6180
rect 280062 6128 280068 6180
rect 280120 6168 280126 6180
rect 340690 6168 340696 6180
rect 280120 6140 340696 6168
rect 280120 6128 280126 6140
rect 340690 6128 340696 6140
rect 340748 6128 340754 6180
rect 344922 6128 344928 6180
rect 344980 6168 344986 6180
rect 406102 6168 406108 6180
rect 344980 6140 406108 6168
rect 344980 6128 344986 6140
rect 406102 6128 406108 6140
rect 406160 6128 406166 6180
rect 426342 6128 426348 6180
rect 426400 6168 426406 6180
rect 486970 6168 486976 6180
rect 426400 6140 486976 6168
rect 426400 6128 426406 6140
rect 486970 6128 486976 6140
rect 487028 6128 487034 6180
rect 502242 6128 502248 6180
rect 502300 6168 502306 6180
rect 561950 6168 561956 6180
rect 502300 6140 561956 6168
rect 502300 6128 502306 6140
rect 561950 6128 561956 6140
rect 562008 6128 562014 6180
rect 480162 5312 480168 5364
rect 480220 5352 480226 5364
rect 540514 5352 540520 5364
rect 480220 5324 540520 5352
rect 480220 5312 480226 5324
rect 540514 5312 540520 5324
rect 540572 5312 540578 5364
rect 362862 5244 362868 5296
rect 362920 5284 362926 5296
rect 422754 5284 422760 5296
rect 362920 5256 422760 5284
rect 362920 5244 362926 5256
rect 422754 5244 422760 5256
rect 422812 5244 422818 5296
rect 484302 5244 484308 5296
rect 484360 5284 484366 5296
rect 544102 5284 544108 5296
rect 484360 5256 544108 5284
rect 484360 5244 484366 5256
rect 544102 5244 544108 5256
rect 544160 5244 544166 5296
rect 369762 5176 369768 5228
rect 369820 5216 369826 5228
rect 429930 5216 429936 5228
rect 369820 5188 429936 5216
rect 369820 5176 369826 5188
rect 429930 5176 429936 5188
rect 429988 5176 429994 5228
rect 487062 5176 487068 5228
rect 487120 5216 487126 5228
rect 547690 5216 547696 5228
rect 487120 5188 547696 5216
rect 487120 5176 487126 5188
rect 547690 5176 547696 5188
rect 547748 5176 547754 5228
rect 394602 5108 394608 5160
rect 394660 5148 394666 5160
rect 454862 5148 454868 5160
rect 394660 5120 454868 5148
rect 394660 5108 394666 5120
rect 454862 5108 454868 5120
rect 454920 5108 454926 5160
rect 463602 5108 463608 5160
rect 463660 5148 463666 5160
rect 523862 5148 523868 5160
rect 463660 5120 523868 5148
rect 463660 5108 463666 5120
rect 523862 5108 523868 5120
rect 523920 5108 523926 5160
rect 380802 5040 380808 5092
rect 380860 5080 380866 5092
rect 440602 5080 440608 5092
rect 380860 5052 440608 5080
rect 380860 5040 380866 5052
rect 440602 5040 440608 5052
rect 440660 5040 440666 5092
rect 455322 5040 455328 5092
rect 455380 5080 455386 5092
rect 515582 5080 515588 5092
rect 455380 5052 515588 5080
rect 455380 5040 455386 5052
rect 515582 5040 515588 5052
rect 515640 5040 515646 5092
rect 358722 4972 358728 5024
rect 358780 5012 358786 5024
rect 419166 5012 419172 5024
rect 358780 4984 419172 5012
rect 358780 4972 358786 4984
rect 419166 4972 419172 4984
rect 419224 4972 419230 5024
rect 422297 5015 422355 5021
rect 422297 4981 422309 5015
rect 422343 5012 422355 5015
rect 428185 5015 428243 5021
rect 428185 5012 428197 5015
rect 422343 4984 428197 5012
rect 422343 4981 422355 4984
rect 422297 4975 422355 4981
rect 428185 4981 428197 4984
rect 428231 4981 428243 5015
rect 428185 4975 428243 4981
rect 466362 4972 466368 5024
rect 466420 5012 466426 5024
rect 526254 5012 526260 5024
rect 466420 4984 526260 5012
rect 466420 4972 466426 4984
rect 526254 4972 526260 4984
rect 526312 4972 526318 5024
rect 133782 4904 133788 4956
rect 133840 4944 133846 4956
rect 194410 4944 194416 4956
rect 133840 4916 194416 4944
rect 133840 4904 133846 4916
rect 194410 4904 194416 4916
rect 194468 4904 194474 4956
rect 376757 4947 376815 4953
rect 376757 4913 376769 4947
rect 376803 4944 376815 4947
rect 386325 4947 386383 4953
rect 386325 4944 386337 4947
rect 376803 4916 386337 4944
rect 376803 4913 376815 4916
rect 376757 4907 376815 4913
rect 386325 4913 386337 4916
rect 386371 4913 386383 4947
rect 386325 4907 386383 4913
rect 387702 4904 387708 4956
rect 387760 4944 387766 4956
rect 447778 4944 447784 4956
rect 387760 4916 447784 4944
rect 387760 4904 387766 4916
rect 447778 4904 447784 4916
rect 447836 4904 447842 4956
rect 462222 4904 462228 4956
rect 462280 4944 462286 4956
rect 522666 4944 522672 4956
rect 462280 4916 522672 4944
rect 462280 4904 462286 4916
rect 522666 4904 522672 4916
rect 522724 4904 522730 4956
rect 66162 4836 66168 4888
rect 66220 4876 66226 4888
rect 126606 4876 126612 4888
rect 66220 4848 126612 4876
rect 66220 4836 66226 4848
rect 126606 4836 126612 4848
rect 126664 4836 126670 4888
rect 173802 4836 173808 4888
rect 173860 4876 173866 4888
rect 234798 4876 234804 4888
rect 173860 4848 234804 4876
rect 173860 4836 173866 4848
rect 234798 4836 234804 4848
rect 234856 4836 234862 4888
rect 255222 4836 255228 4888
rect 255280 4876 255286 4888
rect 315758 4876 315764 4888
rect 255280 4848 315764 4876
rect 255280 4836 255286 4848
rect 315758 4836 315764 4848
rect 315816 4836 315822 4888
rect 390462 4836 390468 4888
rect 390520 4876 390526 4888
rect 402977 4879 403035 4885
rect 402977 4876 402989 4879
rect 390520 4848 402989 4876
rect 390520 4836 390526 4848
rect 402977 4845 402989 4848
rect 403023 4845 403035 4879
rect 402977 4839 403035 4845
rect 406381 4879 406439 4885
rect 406381 4845 406393 4879
rect 406427 4876 406439 4879
rect 422297 4879 422355 4885
rect 422297 4876 422309 4879
rect 406427 4848 422309 4876
rect 406427 4845 406439 4848
rect 406381 4839 406439 4845
rect 422297 4845 422309 4848
rect 422343 4845 422355 4879
rect 422297 4839 422355 4845
rect 428185 4879 428243 4885
rect 428185 4845 428197 4879
rect 428231 4876 428243 4879
rect 428231 4848 441660 4876
rect 428231 4845 428243 4848
rect 428185 4839 428243 4845
rect 68922 4768 68928 4820
rect 68980 4808 68986 4820
rect 130194 4808 130200 4820
rect 68980 4780 130200 4808
rect 68980 4768 68986 4780
rect 130194 4768 130200 4780
rect 130252 4768 130258 4820
rect 190362 4768 190368 4820
rect 190420 4808 190426 4820
rect 251450 4808 251456 4820
rect 190420 4780 251456 4808
rect 190420 4768 190426 4780
rect 251450 4768 251456 4780
rect 251508 4768 251514 4820
rect 295242 4768 295248 4820
rect 295300 4808 295306 4820
rect 356146 4808 356152 4820
rect 295300 4780 356152 4808
rect 295300 4768 295306 4780
rect 356146 4768 356152 4780
rect 356204 4768 356210 4820
rect 372522 4768 372528 4820
rect 372580 4808 372586 4820
rect 376757 4811 376815 4817
rect 376757 4808 376769 4811
rect 372580 4780 376769 4808
rect 372580 4768 372586 4780
rect 376757 4777 376769 4780
rect 376803 4777 376815 4811
rect 376757 4771 376815 4777
rect 386325 4743 386383 4749
rect 386325 4709 386337 4743
rect 386371 4740 386383 4743
rect 424965 4743 425023 4749
rect 386371 4712 386460 4740
rect 386371 4709 386383 4712
rect 386325 4703 386383 4709
rect 386432 4681 386460 4712
rect 402900 4712 408356 4740
rect 386417 4675 386475 4681
rect 386417 4641 386429 4675
rect 386463 4641 386475 4675
rect 386417 4635 386475 4641
rect 386601 4675 386659 4681
rect 386601 4641 386613 4675
rect 386647 4672 386659 4675
rect 402900 4672 402928 4712
rect 386647 4644 402928 4672
rect 402977 4675 403035 4681
rect 386647 4641 386659 4644
rect 386601 4635 386659 4641
rect 402977 4641 402989 4675
rect 403023 4672 403035 4675
rect 406381 4675 406439 4681
rect 406381 4672 406393 4675
rect 403023 4644 406393 4672
rect 403023 4641 403035 4644
rect 402977 4635 403035 4641
rect 406381 4641 406393 4644
rect 406427 4641 406439 4675
rect 408328 4672 408356 4712
rect 424965 4709 424977 4743
rect 425011 4740 425023 4743
rect 441632 4740 441660 4848
rect 459462 4836 459468 4888
rect 459520 4876 459526 4888
rect 519078 4876 519084 4888
rect 459520 4848 519084 4876
rect 459520 4836 459526 4848
rect 519078 4836 519084 4848
rect 519136 4836 519142 4888
rect 476022 4768 476028 4820
rect 476080 4808 476086 4820
rect 536926 4808 536932 4820
rect 476080 4780 536932 4808
rect 476080 4768 476086 4780
rect 536926 4768 536932 4780
rect 536984 4768 536990 4820
rect 451366 4740 451372 4752
rect 425011 4712 425100 4740
rect 441632 4712 451372 4740
rect 425011 4709 425023 4712
rect 424965 4703 425023 4709
rect 425072 4681 425100 4712
rect 451366 4700 451372 4712
rect 451424 4700 451430 4752
rect 415397 4675 415455 4681
rect 415397 4672 415409 4675
rect 408328 4644 415409 4672
rect 406381 4635 406439 4641
rect 415397 4641 415409 4644
rect 415443 4641 415455 4675
rect 415397 4635 415455 4641
rect 425057 4675 425115 4681
rect 425057 4641 425069 4675
rect 425103 4641 425115 4675
rect 425057 4635 425115 4641
rect 415397 4539 415455 4545
rect 415397 4505 415409 4539
rect 415443 4536 415455 4539
rect 424965 4539 425023 4545
rect 424965 4536 424977 4539
rect 415443 4508 424977 4536
rect 415443 4505 415455 4508
rect 415397 4499 415455 4505
rect 424965 4505 424977 4508
rect 425011 4505 425023 4539
rect 424965 4499 425023 4505
rect 143442 4088 143448 4140
rect 143500 4128 143506 4140
rect 203886 4128 203892 4140
rect 143500 4100 203892 4128
rect 143500 4088 143506 4100
rect 203886 4088 203892 4100
rect 203944 4088 203950 4140
rect 240042 4088 240048 4140
rect 240100 4128 240106 4140
rect 300302 4128 300308 4140
rect 240100 4100 300308 4128
rect 240100 4088 240106 4100
rect 300302 4088 300308 4100
rect 300360 4088 300366 4140
rect 347501 4131 347559 4137
rect 347501 4097 347513 4131
rect 347547 4128 347559 4131
rect 353754 4128 353760 4140
rect 347547 4100 353760 4128
rect 347547 4097 347559 4100
rect 347501 4091 347559 4097
rect 353754 4088 353760 4100
rect 353812 4088 353818 4140
rect 361482 4088 361488 4140
rect 361540 4128 361546 4140
rect 421558 4128 421564 4140
rect 361540 4100 421564 4128
rect 361540 4088 361546 4100
rect 421558 4088 421564 4100
rect 421616 4088 421622 4140
rect 443086 4088 443092 4140
rect 443144 4128 443150 4140
rect 444190 4128 444196 4140
rect 443144 4100 444196 4128
rect 443144 4088 443150 4100
rect 444190 4088 444196 4100
rect 444248 4088 444254 4140
rect 447042 4088 447048 4140
rect 447100 4128 447106 4140
rect 507210 4128 507216 4140
rect 447100 4100 507216 4128
rect 447100 4088 447106 4100
rect 507210 4088 507216 4100
rect 507268 4088 507274 4140
rect 507762 4088 507768 4140
rect 507820 4128 507826 4140
rect 567838 4128 567844 4140
rect 507820 4100 567844 4128
rect 507820 4088 507826 4100
rect 567838 4088 567844 4100
rect 567896 4088 567902 4140
rect 132586 4020 132592 4072
rect 132644 4060 132650 4072
rect 133782 4060 133788 4072
rect 132644 4032 133788 4060
rect 132644 4020 132650 4032
rect 133782 4020 133788 4032
rect 133840 4020 133846 4072
rect 150342 4020 150348 4072
rect 150400 4060 150406 4072
rect 211062 4060 211068 4072
rect 150400 4032 211068 4060
rect 150400 4020 150406 4032
rect 211062 4020 211068 4032
rect 211120 4020 211126 4072
rect 257982 4020 257988 4072
rect 258040 4060 258046 4072
rect 318058 4060 318064 4072
rect 258040 4032 318064 4060
rect 258040 4020 258046 4032
rect 318058 4020 318064 4032
rect 318116 4020 318122 4072
rect 350442 4020 350448 4072
rect 350500 4060 350506 4072
rect 410886 4060 410892 4072
rect 350500 4032 410892 4060
rect 350500 4020 350506 4032
rect 410886 4020 410892 4032
rect 410944 4020 410950 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 471514 4060 471520 4072
rect 411220 4032 471520 4060
rect 411220 4020 411226 4032
rect 471514 4020 471520 4032
rect 471572 4020 471578 4072
rect 503622 4020 503628 4072
rect 503680 4060 503686 4072
rect 564342 4060 564348 4072
rect 503680 4032 564348 4060
rect 503680 4020 503686 4032
rect 564342 4020 564348 4032
rect 564400 4020 564406 4072
rect 92290 3952 92296 4004
rect 92348 3992 92354 4004
rect 152734 3992 152740 4004
rect 92348 3964 152740 3992
rect 92348 3952 92354 3964
rect 152734 3952 152740 3964
rect 152792 3952 152798 4004
rect 161382 3952 161388 4004
rect 161440 3992 161446 4004
rect 221734 3992 221740 4004
rect 161440 3964 221740 3992
rect 161440 3952 161446 3964
rect 221734 3952 221740 3964
rect 221792 3952 221798 4004
rect 246942 3952 246948 4004
rect 247000 3992 247006 4004
rect 307386 3992 307392 4004
rect 247000 3964 307392 3992
rect 247000 3952 247006 3964
rect 307386 3952 307392 3964
rect 307444 3952 307450 4004
rect 314562 3952 314568 4004
rect 314620 3992 314626 4004
rect 375190 3992 375196 4004
rect 314620 3964 375196 3992
rect 314620 3952 314626 3964
rect 375190 3952 375196 3964
rect 375248 3952 375254 4004
rect 400122 3952 400128 4004
rect 400180 3992 400186 4004
rect 460750 3992 460756 4004
rect 400180 3964 460756 3992
rect 400180 3952 400186 3964
rect 460750 3952 460756 3964
rect 460808 3952 460814 4004
rect 460842 3952 460848 4004
rect 460900 3992 460906 4004
rect 521470 3992 521476 4004
rect 460900 3964 521476 3992
rect 460900 3952 460906 3964
rect 521470 3952 521476 3964
rect 521528 3952 521534 4004
rect 521562 3952 521568 4004
rect 521620 3992 521626 4004
rect 582190 3992 582196 4004
rect 521620 3964 582196 3992
rect 521620 3952 521626 3964
rect 582190 3952 582196 3964
rect 582248 3952 582254 4004
rect 71682 3884 71688 3936
rect 71740 3924 71746 3936
rect 132494 3924 132500 3936
rect 71740 3896 132500 3924
rect 71740 3884 71746 3896
rect 132494 3884 132500 3896
rect 132552 3884 132558 3936
rect 132604 3896 133920 3924
rect 78582 3816 78588 3868
rect 78640 3856 78646 3868
rect 132604 3856 132632 3896
rect 78640 3828 132632 3856
rect 133892 3856 133920 3896
rect 136450 3884 136456 3936
rect 136508 3924 136514 3936
rect 196802 3924 196808 3936
rect 136508 3896 196808 3924
rect 136508 3884 136514 3896
rect 196802 3884 196808 3896
rect 196860 3884 196866 3936
rect 200022 3884 200028 3936
rect 200080 3924 200086 3936
rect 261018 3924 261024 3936
rect 200080 3896 261024 3924
rect 200080 3884 200086 3896
rect 261018 3884 261024 3896
rect 261076 3884 261082 3936
rect 262214 3884 262220 3936
rect 262272 3924 262278 3936
rect 263410 3924 263416 3936
rect 262272 3896 263416 3924
rect 262272 3884 262278 3896
rect 263410 3884 263416 3896
rect 263468 3884 263474 3936
rect 307662 3884 307668 3936
rect 307720 3924 307726 3936
rect 368014 3924 368020 3936
rect 307720 3896 368020 3924
rect 307720 3884 307726 3896
rect 368014 3884 368020 3896
rect 368072 3884 368078 3936
rect 393222 3884 393228 3936
rect 393280 3924 393286 3936
rect 453666 3924 453672 3936
rect 393280 3896 453672 3924
rect 393280 3884 393286 3896
rect 453666 3884 453672 3896
rect 453724 3884 453730 3936
rect 464982 3884 464988 3936
rect 465040 3924 465046 3936
rect 525058 3924 525064 3936
rect 465040 3896 525064 3924
rect 465040 3884 465046 3896
rect 525058 3884 525064 3896
rect 525116 3884 525122 3936
rect 139670 3856 139676 3868
rect 133892 3828 139676 3856
rect 78640 3816 78646 3828
rect 139670 3816 139676 3828
rect 139728 3816 139734 3868
rect 140774 3816 140780 3868
rect 140832 3856 140838 3868
rect 142062 3856 142068 3868
rect 140832 3828 142068 3856
rect 140832 3816 140838 3828
rect 142062 3816 142068 3828
rect 142120 3816 142126 3868
rect 157242 3816 157248 3868
rect 157300 3856 157306 3868
rect 218054 3856 218060 3868
rect 157300 3828 218060 3856
rect 157300 3816 157306 3828
rect 218054 3816 218060 3828
rect 218112 3816 218118 3868
rect 229002 3816 229008 3868
rect 229060 3856 229066 3868
rect 289538 3856 289544 3868
rect 229060 3828 289544 3856
rect 229060 3816 229066 3828
rect 289538 3816 289544 3828
rect 289596 3816 289602 3868
rect 293862 3816 293868 3868
rect 293920 3856 293926 3868
rect 347501 3859 347559 3865
rect 347501 3856 347513 3859
rect 293920 3828 347513 3856
rect 293920 3816 293926 3828
rect 347501 3825 347513 3828
rect 347547 3825 347559 3859
rect 350258 3856 350264 3868
rect 347501 3819 347559 3825
rect 347608 3828 350264 3856
rect 84102 3748 84108 3800
rect 84160 3788 84166 3800
rect 145650 3788 145656 3800
rect 84160 3760 145656 3788
rect 84160 3748 84166 3760
rect 145650 3748 145656 3760
rect 145708 3748 145714 3800
rect 150526 3748 150532 3800
rect 150584 3788 150590 3800
rect 151538 3788 151544 3800
rect 150584 3760 151544 3788
rect 150584 3748 150590 3760
rect 151538 3748 151544 3760
rect 151596 3748 151602 3800
rect 153102 3748 153108 3800
rect 153160 3788 153166 3800
rect 214650 3788 214656 3800
rect 153160 3760 214656 3788
rect 153160 3748 153166 3760
rect 214650 3748 214656 3760
rect 214708 3748 214714 3800
rect 222102 3748 222108 3800
rect 222160 3788 222166 3800
rect 282454 3788 282460 3800
rect 222160 3760 282460 3788
rect 222160 3748 222166 3760
rect 282454 3748 282460 3760
rect 282512 3748 282518 3800
rect 289722 3748 289728 3800
rect 289780 3788 289786 3800
rect 347608 3788 347636 3828
rect 350258 3816 350264 3828
rect 350316 3816 350322 3868
rect 354582 3816 354588 3868
rect 354640 3856 354646 3868
rect 414474 3856 414480 3868
rect 354640 3828 414480 3856
rect 354640 3816 354646 3828
rect 414474 3816 414480 3828
rect 414532 3816 414538 3868
rect 415302 3816 415308 3868
rect 415360 3856 415366 3868
rect 475102 3856 475108 3868
rect 415360 3828 475108 3856
rect 415360 3816 415366 3828
rect 475102 3816 475108 3828
rect 475160 3816 475166 3868
rect 500862 3816 500868 3868
rect 500920 3856 500926 3868
rect 560754 3856 560760 3868
rect 500920 3828 560760 3856
rect 500920 3816 500926 3828
rect 560754 3816 560760 3828
rect 560812 3816 560818 3868
rect 289780 3760 347636 3788
rect 289780 3748 289786 3760
rect 347774 3748 347780 3800
rect 347832 3788 347838 3800
rect 349062 3788 349068 3800
rect 347832 3760 349068 3788
rect 347832 3748 347838 3760
rect 349062 3748 349068 3760
rect 349120 3748 349126 3800
rect 379422 3748 379428 3800
rect 379480 3788 379486 3800
rect 439406 3788 439412 3800
rect 379480 3760 439412 3788
rect 379480 3748 379486 3760
rect 439406 3748 439412 3760
rect 439464 3748 439470 3800
rect 446582 3788 446588 3800
rect 443104 3760 446588 3788
rect 114462 3680 114468 3732
rect 114520 3720 114526 3732
rect 175274 3720 175280 3732
rect 114520 3692 175280 3720
rect 114520 3680 114526 3692
rect 175274 3680 175280 3692
rect 175332 3680 175338 3732
rect 206922 3680 206928 3732
rect 206980 3720 206986 3732
rect 268102 3720 268108 3732
rect 206980 3692 268108 3720
rect 206980 3680 206986 3692
rect 268102 3680 268108 3692
rect 268160 3680 268166 3732
rect 296622 3680 296628 3732
rect 296680 3720 296686 3732
rect 357342 3720 357348 3732
rect 296680 3692 357348 3720
rect 296680 3680 296686 3692
rect 357342 3680 357348 3692
rect 357400 3680 357406 3732
rect 357434 3680 357440 3732
rect 357492 3720 357498 3732
rect 417970 3720 417976 3732
rect 357492 3692 417976 3720
rect 357492 3680 357498 3692
rect 417970 3680 417976 3692
rect 418028 3680 418034 3732
rect 418062 3680 418068 3732
rect 418120 3720 418126 3732
rect 442905 3723 442963 3729
rect 442905 3720 442917 3723
rect 418120 3692 442917 3720
rect 418120 3680 418126 3692
rect 442905 3689 442917 3692
rect 442951 3689 442963 3723
rect 442905 3683 442963 3689
rect 121362 3612 121368 3664
rect 121420 3652 121426 3664
rect 182542 3652 182548 3664
rect 121420 3624 182548 3652
rect 121420 3612 121426 3624
rect 182542 3612 182548 3624
rect 182600 3612 182606 3664
rect 189626 3652 189632 3664
rect 183480 3624 189632 3652
rect 128262 3544 128268 3596
rect 128320 3584 128326 3596
rect 183480 3584 183508 3624
rect 189626 3612 189632 3624
rect 189684 3612 189690 3664
rect 231762 3612 231768 3664
rect 231820 3652 231826 3664
rect 293126 3652 293132 3664
rect 231820 3624 293132 3652
rect 231820 3612 231826 3624
rect 293126 3612 293132 3624
rect 293184 3612 293190 3664
rect 382274 3652 382280 3664
rect 326356 3624 382280 3652
rect 128320 3556 183508 3584
rect 128320 3544 128326 3556
rect 183554 3544 183560 3596
rect 183612 3584 183618 3596
rect 184842 3584 184848 3596
rect 183612 3556 184848 3584
rect 183612 3544 183618 3556
rect 184842 3544 184848 3556
rect 184900 3544 184906 3596
rect 201494 3544 201500 3596
rect 201552 3584 201558 3596
rect 202690 3584 202696 3596
rect 201552 3556 202696 3584
rect 201552 3544 201558 3556
rect 202690 3544 202696 3556
rect 202748 3544 202754 3596
rect 218146 3544 218152 3596
rect 218204 3584 218210 3596
rect 219342 3584 219348 3596
rect 218204 3556 219348 3584
rect 218204 3544 218210 3556
rect 219342 3544 219348 3556
rect 219400 3544 219406 3596
rect 236086 3544 236092 3596
rect 236144 3584 236150 3596
rect 237190 3584 237196 3596
rect 236144 3556 237196 3584
rect 236144 3544 236150 3556
rect 237190 3544 237196 3556
rect 237248 3544 237254 3596
rect 242802 3544 242808 3596
rect 242860 3584 242866 3596
rect 303798 3584 303804 3596
rect 242860 3556 303804 3584
rect 242860 3544 242866 3556
rect 303798 3544 303804 3556
rect 303856 3544 303862 3596
rect 304994 3544 305000 3596
rect 305052 3584 305058 3596
rect 306190 3584 306196 3596
rect 305052 3556 306196 3584
rect 305052 3544 305058 3556
rect 306190 3544 306196 3556
rect 306248 3544 306254 3596
rect 310422 3544 310428 3596
rect 310480 3584 310486 3596
rect 326249 3587 326307 3593
rect 326249 3584 326261 3587
rect 310480 3556 326261 3584
rect 310480 3544 310486 3556
rect 326249 3553 326261 3556
rect 326295 3553 326307 3587
rect 326249 3547 326307 3553
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 63494 3516 63500 3528
rect 1728 3488 63500 3516
rect 1728 3476 1734 3488
rect 63494 3476 63500 3488
rect 63552 3476 63558 3528
rect 88242 3476 88248 3528
rect 88300 3516 88306 3528
rect 149238 3516 149244 3528
rect 88300 3488 149244 3516
rect 88300 3476 88306 3488
rect 149238 3476 149244 3488
rect 149296 3476 149302 3528
rect 171042 3476 171048 3528
rect 171100 3516 171106 3528
rect 232498 3516 232504 3528
rect 171100 3488 232504 3516
rect 171100 3476 171106 3488
rect 232498 3476 232504 3488
rect 232556 3476 232562 3528
rect 244274 3476 244280 3528
rect 244332 3516 244338 3528
rect 245562 3516 245568 3528
rect 244332 3488 245568 3516
rect 244332 3476 244338 3488
rect 245562 3476 245568 3488
rect 245620 3476 245626 3528
rect 249702 3476 249708 3528
rect 249760 3516 249766 3528
rect 310974 3516 310980 3528
rect 249760 3488 310980 3516
rect 249760 3476 249766 3488
rect 310974 3476 310980 3488
rect 311032 3476 311038 3528
rect 321462 3476 321468 3528
rect 321520 3516 321526 3528
rect 326356 3516 326384 3624
rect 382274 3612 382280 3624
rect 382332 3612 382338 3664
rect 386322 3612 386328 3664
rect 386380 3652 386386 3664
rect 443104 3652 443132 3760
rect 446582 3748 446588 3760
rect 446640 3748 446646 3800
rect 471882 3748 471888 3800
rect 471940 3788 471946 3800
rect 528557 3791 528615 3797
rect 528557 3788 528569 3791
rect 471940 3760 528569 3788
rect 471940 3748 471946 3760
rect 528557 3757 528569 3760
rect 528603 3757 528615 3791
rect 528557 3751 528615 3757
rect 528646 3748 528652 3800
rect 528704 3788 528710 3800
rect 529842 3788 529848 3800
rect 528704 3760 529848 3788
rect 528704 3748 528710 3760
rect 529842 3748 529848 3760
rect 529900 3748 529906 3800
rect 443181 3723 443239 3729
rect 443181 3689 443193 3723
rect 443227 3720 443239 3723
rect 478690 3720 478696 3732
rect 443227 3692 478696 3720
rect 443227 3689 443239 3692
rect 443181 3683 443239 3689
rect 478690 3680 478696 3692
rect 478748 3680 478754 3732
rect 513282 3680 513288 3732
rect 513340 3720 513346 3732
rect 573818 3720 573824 3732
rect 513340 3692 573824 3720
rect 513340 3680 513346 3692
rect 573818 3680 573824 3692
rect 573876 3680 573882 3732
rect 386380 3624 443132 3652
rect 386380 3612 386386 3624
rect 451274 3612 451280 3664
rect 451332 3652 451338 3664
rect 452470 3652 452476 3664
rect 451332 3624 452476 3652
rect 451332 3612 451338 3624
rect 452470 3612 452476 3624
rect 452528 3612 452534 3664
rect 467834 3612 467840 3664
rect 467892 3652 467898 3664
rect 469122 3652 469128 3664
rect 467892 3624 469128 3652
rect 467892 3612 467898 3624
rect 469122 3612 469128 3624
rect 469180 3612 469186 3664
rect 478782 3612 478788 3664
rect 478840 3652 478846 3664
rect 539318 3652 539324 3664
rect 478840 3624 539324 3652
rect 478840 3612 478846 3624
rect 539318 3612 539324 3624
rect 539376 3612 539382 3664
rect 326433 3587 326491 3593
rect 326433 3553 326445 3587
rect 326479 3584 326491 3587
rect 371602 3584 371608 3596
rect 326479 3556 371608 3584
rect 326479 3553 326491 3556
rect 326433 3547 326491 3553
rect 371602 3544 371608 3556
rect 371660 3544 371666 3596
rect 382366 3544 382372 3596
rect 382424 3584 382430 3596
rect 383562 3584 383568 3596
rect 382424 3556 383568 3584
rect 382424 3544 382430 3556
rect 383562 3544 383568 3556
rect 383620 3544 383626 3596
rect 422202 3544 422208 3596
rect 422260 3584 422266 3596
rect 482278 3584 482284 3596
rect 422260 3556 482284 3584
rect 422260 3544 422266 3556
rect 482278 3544 482284 3556
rect 482336 3544 482342 3596
rect 494146 3544 494152 3596
rect 494204 3584 494210 3596
rect 495342 3584 495348 3596
rect 494204 3556 495348 3584
rect 494204 3544 494210 3556
rect 495342 3544 495348 3556
rect 495400 3544 495406 3596
rect 496722 3544 496728 3596
rect 496780 3584 496786 3596
rect 557166 3584 557172 3596
rect 496780 3556 557172 3584
rect 496780 3544 496786 3556
rect 557166 3544 557172 3556
rect 557224 3544 557230 3596
rect 321520 3488 326384 3516
rect 321520 3476 321526 3488
rect 328362 3476 328368 3528
rect 328420 3516 328426 3528
rect 389450 3516 389456 3528
rect 328420 3488 389456 3516
rect 328420 3476 328426 3488
rect 389450 3476 389456 3488
rect 389508 3476 389514 3528
rect 425054 3476 425060 3528
rect 425112 3516 425118 3528
rect 426342 3516 426348 3528
rect 425112 3488 426348 3516
rect 425112 3476 425118 3488
rect 426342 3476 426348 3488
rect 426400 3476 426406 3528
rect 429102 3476 429108 3528
rect 429160 3516 429166 3528
rect 489362 3516 489368 3528
rect 429160 3488 489368 3516
rect 429160 3476 429166 3488
rect 489362 3476 489368 3488
rect 489420 3476 489426 3528
rect 493962 3476 493968 3528
rect 494020 3516 494026 3528
rect 553578 3516 553584 3528
rect 494020 3488 553584 3516
rect 494020 3476 494026 3488
rect 553578 3476 553584 3488
rect 553636 3476 553642 3528
rect 571426 3476 571432 3528
rect 571484 3516 571490 3528
rect 572622 3516 572628 3528
rect 571484 3488 572628 3516
rect 571484 3476 571490 3488
rect 572622 3476 572628 3488
rect 572680 3476 572686 3528
rect 578878 3476 578884 3528
rect 578936 3516 578942 3528
rect 579798 3516 579804 3528
rect 578936 3488 579804 3516
rect 578936 3476 578942 3488
rect 579798 3476 579804 3488
rect 579856 3476 579862 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 62114 3448 62120 3460
rect 624 3420 62120 3448
rect 624 3408 630 3420
rect 62114 3408 62120 3420
rect 62172 3408 62178 3460
rect 95142 3408 95148 3460
rect 95200 3448 95206 3460
rect 156322 3448 156328 3460
rect 95200 3420 156328 3448
rect 95200 3408 95206 3420
rect 156322 3408 156328 3420
rect 156380 3408 156386 3460
rect 164142 3408 164148 3460
rect 164200 3448 164206 3460
rect 225322 3448 225328 3460
rect 164200 3420 225328 3448
rect 164200 3408 164206 3420
rect 225322 3408 225328 3420
rect 225380 3408 225386 3460
rect 235902 3408 235908 3460
rect 235960 3448 235966 3460
rect 296714 3448 296720 3460
rect 235960 3420 296720 3448
rect 235960 3408 235966 3420
rect 296714 3408 296720 3420
rect 296772 3408 296778 3460
rect 300762 3408 300768 3460
rect 300820 3448 300826 3460
rect 360930 3448 360936 3460
rect 300820 3420 360936 3448
rect 300820 3408 300826 3420
rect 360930 3408 360936 3420
rect 360988 3408 360994 3460
rect 365714 3408 365720 3460
rect 365772 3448 365778 3460
rect 366910 3448 366916 3460
rect 365772 3420 366916 3448
rect 365772 3408 365778 3420
rect 366910 3408 366916 3420
rect 366968 3408 366974 3460
rect 371142 3408 371148 3460
rect 371200 3448 371206 3460
rect 432322 3448 432328 3460
rect 371200 3420 432328 3448
rect 371200 3408 371206 3420
rect 432322 3408 432328 3420
rect 432380 3408 432386 3460
rect 440142 3408 440148 3460
rect 440200 3448 440206 3460
rect 500126 3448 500132 3460
rect 440200 3420 500132 3448
rect 440200 3408 440206 3420
rect 500126 3408 500132 3420
rect 500184 3408 500190 3460
rect 517422 3408 517428 3460
rect 517480 3448 517486 3460
rect 577406 3448 577412 3460
rect 517480 3420 577412 3448
rect 517480 3408 517486 3420
rect 577406 3408 577412 3420
rect 577464 3408 577470 3460
rect 125502 3340 125508 3392
rect 125560 3380 125566 3392
rect 186038 3380 186044 3392
rect 125560 3352 186044 3380
rect 125560 3340 125566 3352
rect 186038 3340 186044 3352
rect 186096 3340 186102 3392
rect 215202 3340 215208 3392
rect 215260 3380 215266 3392
rect 215260 3352 267780 3380
rect 215260 3340 215266 3352
rect 118602 3272 118608 3324
rect 118660 3312 118666 3324
rect 118660 3284 173020 3312
rect 118660 3272 118666 3284
rect 107562 3204 107568 3256
rect 107620 3244 107626 3256
rect 168190 3244 168196 3256
rect 107620 3216 168196 3244
rect 107620 3204 107626 3216
rect 168190 3204 168196 3216
rect 168248 3204 168254 3256
rect 172992 3244 173020 3284
rect 175366 3272 175372 3324
rect 175424 3312 175430 3324
rect 176562 3312 176568 3324
rect 175424 3284 176568 3312
rect 175424 3272 175430 3284
rect 176562 3272 176568 3284
rect 176620 3272 176626 3324
rect 204162 3272 204168 3324
rect 204220 3312 204226 3324
rect 264606 3312 264612 3324
rect 204220 3284 264612 3312
rect 204220 3272 204226 3284
rect 264606 3272 264612 3284
rect 264664 3272 264670 3324
rect 178954 3244 178960 3256
rect 172992 3216 178960 3244
rect 178954 3204 178960 3216
rect 179012 3204 179018 3256
rect 197262 3204 197268 3256
rect 197320 3244 197326 3256
rect 257430 3244 257436 3256
rect 197320 3216 257436 3244
rect 197320 3204 197326 3216
rect 257430 3204 257436 3216
rect 257488 3204 257494 3256
rect 267752 3244 267780 3352
rect 270494 3340 270500 3392
rect 270552 3380 270558 3392
rect 271690 3380 271696 3392
rect 270552 3352 271696 3380
rect 270552 3340 270558 3352
rect 271690 3340 271696 3352
rect 271748 3340 271754 3392
rect 287054 3340 287060 3392
rect 287112 3380 287118 3392
rect 288342 3380 288348 3392
rect 287112 3352 288348 3380
rect 287112 3340 287118 3352
rect 288342 3340 288348 3352
rect 288400 3340 288406 3392
rect 336642 3340 336648 3392
rect 336700 3380 336706 3392
rect 396626 3380 396632 3392
rect 336700 3352 396632 3380
rect 336700 3340 336706 3352
rect 396626 3340 396632 3352
rect 396684 3340 396690 3392
rect 436002 3340 436008 3392
rect 436060 3380 436066 3392
rect 496538 3380 496544 3392
rect 436060 3352 496544 3380
rect 436060 3340 436066 3352
rect 496538 3340 496544 3352
rect 496596 3340 496602 3392
rect 511902 3340 511908 3392
rect 511960 3380 511966 3392
rect 571426 3380 571432 3392
rect 511960 3352 571432 3380
rect 511960 3340 511966 3352
rect 571426 3340 571432 3352
rect 571484 3340 571490 3392
rect 318702 3272 318708 3324
rect 318760 3312 318766 3324
rect 378778 3312 378784 3324
rect 318760 3284 378784 3312
rect 318760 3272 318766 3284
rect 378778 3272 378784 3284
rect 378836 3272 378842 3324
rect 453942 3272 453948 3324
rect 454000 3312 454006 3324
rect 514386 3312 514392 3324
rect 454000 3284 514392 3312
rect 454000 3272 454006 3284
rect 514386 3272 514392 3284
rect 514444 3272 514450 3324
rect 514662 3272 514668 3324
rect 514720 3312 514726 3324
rect 575014 3312 575020 3324
rect 514720 3284 575020 3312
rect 514720 3272 514726 3284
rect 575014 3272 575020 3284
rect 575072 3272 575078 3324
rect 275278 3244 275284 3256
rect 267752 3216 275284 3244
rect 275278 3204 275284 3216
rect 275336 3204 275342 3256
rect 325602 3204 325608 3256
rect 325660 3244 325666 3256
rect 385862 3244 385868 3256
rect 325660 3216 385868 3244
rect 325660 3204 325666 3216
rect 385862 3204 385868 3216
rect 385920 3204 385926 3256
rect 458082 3204 458088 3256
rect 458140 3244 458146 3256
rect 517882 3244 517888 3256
rect 458140 3216 517888 3244
rect 458140 3204 458146 3216
rect 517882 3204 517888 3216
rect 517940 3204 517946 3256
rect 518802 3204 518808 3256
rect 518860 3244 518866 3256
rect 578602 3244 578608 3256
rect 518860 3216 578608 3244
rect 518860 3204 518866 3216
rect 578602 3204 578608 3216
rect 578660 3204 578666 3256
rect 100662 3136 100668 3188
rect 100720 3176 100726 3188
rect 161106 3176 161112 3188
rect 100720 3148 161112 3176
rect 100720 3136 100726 3148
rect 161106 3136 161112 3148
rect 161164 3136 161170 3188
rect 193122 3136 193128 3188
rect 193180 3176 193186 3188
rect 253842 3176 253848 3188
rect 193180 3148 253848 3176
rect 193180 3136 193186 3148
rect 253842 3136 253848 3148
rect 253900 3136 253906 3188
rect 332502 3136 332508 3188
rect 332560 3176 332566 3188
rect 393038 3176 393044 3188
rect 332560 3148 393044 3176
rect 332560 3136 332566 3148
rect 393038 3136 393044 3148
rect 393096 3136 393102 3188
rect 442902 3136 442908 3188
rect 442960 3176 442966 3188
rect 503622 3176 503628 3188
rect 442960 3148 503628 3176
rect 442960 3136 442966 3148
rect 503622 3136 503628 3148
rect 503680 3136 503686 3188
rect 528557 3179 528615 3185
rect 528557 3145 528569 3179
rect 528603 3176 528615 3179
rect 532234 3176 532240 3188
rect 528603 3148 532240 3176
rect 528603 3145 528615 3148
rect 528557 3139 528615 3145
rect 532234 3136 532240 3148
rect 532292 3136 532298 3188
rect 99282 3068 99288 3120
rect 99340 3108 99346 3120
rect 159910 3108 159916 3120
rect 99340 3080 159916 3108
rect 99340 3068 99346 3080
rect 159910 3068 159916 3080
rect 159968 3068 159974 3120
rect 179322 3068 179328 3120
rect 179380 3108 179386 3120
rect 239582 3108 239588 3120
rect 179380 3080 239588 3108
rect 179380 3068 179386 3080
rect 239582 3068 239588 3080
rect 239640 3068 239646 3120
rect 343542 3068 343548 3120
rect 343600 3108 343606 3120
rect 403710 3108 403716 3120
rect 343600 3080 403716 3108
rect 343600 3068 343606 3080
rect 403710 3068 403716 3080
rect 403768 3068 403774 3120
rect 433150 3068 433156 3120
rect 433208 3108 433214 3120
rect 492950 3108 492956 3120
rect 433208 3080 492956 3108
rect 433208 3068 433214 3080
rect 492950 3068 492956 3080
rect 493008 3068 493014 3120
rect 186222 3000 186228 3052
rect 186280 3040 186286 3052
rect 246758 3040 246764 3052
rect 186280 3012 246764 3040
rect 186280 3000 186286 3012
rect 246758 3000 246764 3012
rect 246816 3000 246822 3052
rect 374086 2836 374092 2848
rect 374012 2808 374092 2836
rect 374012 2780 374040 2808
rect 374086 2796 374092 2808
rect 374144 2796 374150 2848
rect 427906 2796 427912 2848
rect 427964 2836 427970 2848
rect 427964 2808 428780 2836
rect 427964 2796 427970 2808
rect 428752 2780 428780 2808
rect 373994 2728 374000 2780
rect 374052 2728 374058 2780
rect 428734 2728 428740 2780
rect 428792 2728 428798 2780
rect 425057 2363 425115 2369
rect 425057 2329 425069 2363
rect 425103 2360 425115 2363
rect 433518 2360 433524 2372
rect 425103 2332 433524 2360
rect 425103 2329 425115 2332
rect 425057 2323 425115 2329
rect 433518 2320 433524 2332
rect 433576 2320 433582 2372
rect 328822 552 328828 604
rect 328880 592 328886 604
rect 328914 592 328920 604
rect 328880 564 328920 592
rect 328880 552 328886 564
rect 328914 552 328920 564
rect 328972 552 328978 604
rect 354674 552 354680 604
rect 354732 592 354738 604
rect 354950 592 354956 604
rect 354732 564 354956 592
rect 354732 552 354738 564
rect 354950 552 354956 564
rect 355008 552 355014 604
rect 357526 552 357532 604
rect 357584 592 357590 604
rect 358538 592 358544 604
rect 357584 564 358544 592
rect 357584 552 357590 564
rect 358538 552 358544 564
rect 358596 552 358602 604
rect 358814 552 358820 604
rect 358872 592 358878 604
rect 359734 592 359740 604
rect 358872 564 359740 592
rect 358872 552 358878 564
rect 359734 552 359740 564
rect 359792 552 359798 604
rect 361574 552 361580 604
rect 361632 592 361638 604
rect 362126 592 362132 604
rect 361632 564 362132 592
rect 361632 552 361638 564
rect 362126 552 362132 564
rect 362184 552 362190 604
rect 383654 552 383660 604
rect 383712 592 383718 604
rect 384666 592 384672 604
rect 383712 564 384672 592
rect 383712 552 383718 564
rect 384666 552 384672 564
rect 384724 552 384730 604
rect 386414 552 386420 604
rect 386472 592 386478 604
rect 387058 592 387064 604
rect 386472 564 387064 592
rect 386472 552 386478 564
rect 387058 552 387064 564
rect 387116 552 387122 604
rect 387794 552 387800 604
rect 387852 592 387858 604
rect 388254 592 388260 604
rect 387852 564 388260 592
rect 387852 552 387858 564
rect 388254 552 388260 564
rect 388312 552 388318 604
rect 431126 592 431132 604
rect 431087 564 431132 592
rect 431126 552 431132 564
rect 431184 552 431190 604
rect 435818 592 435824 604
rect 435779 564 435824 592
rect 435818 552 435824 564
rect 435876 552 435882 604
rect 455414 552 455420 604
rect 455472 592 455478 604
rect 456058 592 456064 604
rect 455472 564 456064 592
rect 455472 552 455478 564
rect 456058 552 456064 564
rect 456116 552 456122 604
rect 456886 552 456892 604
rect 456944 592 456950 604
rect 457254 592 457260 604
rect 456944 564 457260 592
rect 456944 552 456950 564
rect 457254 552 457260 564
rect 457312 552 457318 604
rect 471974 552 471980 604
rect 472032 592 472038 604
rect 472710 592 472716 604
rect 472032 564 472716 592
rect 472032 552 472038 564
rect 472710 552 472716 564
rect 472768 552 472774 604
rect 473354 552 473360 604
rect 473412 592 473418 604
rect 473906 592 473912 604
rect 473412 564 473912 592
rect 473412 552 473418 564
rect 473906 552 473912 564
rect 473964 552 473970 604
rect 478874 552 478880 604
rect 478932 592 478938 604
rect 479886 592 479892 604
rect 478932 564 479892 592
rect 478932 552 478938 564
rect 479886 552 479892 564
rect 479944 552 479950 604
rect 557534 552 557540 604
rect 557592 592 557598 604
rect 558362 592 558368 604
rect 557592 564 558368 592
rect 557592 552 557598 564
rect 558362 552 558368 564
rect 558420 552 558426 604
rect 564434 552 564440 604
rect 564492 592 564498 604
rect 565538 592 565544 604
rect 564492 564 565544 592
rect 564492 552 564498 564
rect 565538 552 565544 564
rect 565596 552 565602 604
rect 565814 552 565820 604
rect 565872 592 565878 604
rect 566734 592 566740 604
rect 565872 564 566740 592
rect 565872 552 565878 564
rect 566734 552 566740 564
rect 566792 552 566798 604
<< via1 >>
rect 411168 700408 411220 700460
rect 429844 700408 429896 700460
rect 463608 700408 463660 700460
rect 494796 700408 494848 700460
rect 514668 700408 514720 700460
rect 559656 700408 559708 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 394608 700340 394660 700392
rect 413652 700340 413704 700392
rect 445668 700340 445720 700392
rect 478512 700340 478564 700392
rect 496728 700340 496780 700392
rect 543464 700340 543516 700392
rect 343548 700272 343600 700324
rect 348792 700272 348844 700324
rect 378048 700272 378100 700324
rect 397460 700272 397512 700324
rect 429108 700272 429160 700324
rect 462320 700272 462372 700324
rect 480168 700272 480220 700324
rect 527180 700272 527232 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 326988 699660 327040 699712
rect 332508 699660 332560 699712
rect 360108 699660 360160 699712
rect 364984 699660 365036 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 523776 696940 523828 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 692724 72752 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 523684 685856 523736 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 683247 72568 683256
rect 72516 683213 72525 683247
rect 72525 683213 72559 683247
rect 72559 683213 72568 683247
rect 72516 683204 72568 683213
rect 72516 683068 72568 683120
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 219072 678988 219124 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 218980 678920 219032 678972
rect 72700 678895 72752 678904
rect 72700 678861 72709 678895
rect 72709 678861 72743 678895
rect 72743 678861 72752 678895
rect 72700 678852 72752 678861
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 72700 669264 72752 669316
rect 72884 669264 72936 669316
rect 218980 669264 219032 669316
rect 219164 669264 219216 669316
rect 72884 666476 72936 666528
rect 219164 666476 219216 666528
rect 72792 656931 72844 656940
rect 72792 656897 72801 656931
rect 72801 656897 72835 656931
rect 72835 656897 72844 656931
rect 72792 656888 72844 656897
rect 219072 656931 219124 656940
rect 219072 656897 219081 656931
rect 219081 656897 219115 656931
rect 219115 656897 219124 656931
rect 219072 656888 219124 656897
rect 377128 655460 377180 655512
rect 378048 655460 378100 655512
rect 428188 655460 428240 655512
rect 429108 655460 429160 655512
rect 462320 655460 462372 655512
rect 463608 655460 463660 655512
rect 479340 655460 479392 655512
rect 480168 655460 480220 655512
rect 513380 655256 513432 655308
rect 514668 655256 514720 655308
rect 325976 655120 326028 655172
rect 326988 655120 327040 655172
rect 8024 654916 8076 654968
rect 70492 654916 70544 654968
rect 72792 654916 72844 654968
rect 121552 654916 121604 654968
rect 137744 654916 137796 654968
rect 172704 654916 172756 654968
rect 41328 654848 41380 654900
rect 104532 654848 104584 654900
rect 106188 654848 106240 654900
rect 155592 654848 155644 654900
rect 171048 654848 171100 654900
rect 206744 654848 206796 654900
rect 219072 654848 219124 654900
rect 240784 654848 240836 654900
rect 24768 654780 24820 654832
rect 87512 654780 87564 654832
rect 89628 654780 89680 654832
rect 138572 654780 138624 654832
rect 154304 654780 154356 654832
rect 189724 654780 189776 654832
rect 202788 654780 202840 654832
rect 223764 654780 223816 654832
rect 235908 654780 235960 654832
rect 257896 654780 257948 654832
rect 267648 654780 267700 654832
rect 274916 654780 274968 654832
rect 284024 654780 284076 654832
rect 291936 654780 291988 654832
rect 300768 654100 300820 654152
rect 308956 654100 309008 654152
rect 3608 645804 3660 645856
rect 59360 645804 59412 645856
rect 523776 638936 523828 638988
rect 580172 638936 580224 638988
rect 3424 630572 3476 630624
rect 59360 630572 59412 630624
rect 524328 619556 524380 619608
rect 580264 619556 580316 619608
rect 3516 616768 3568 616820
rect 59360 616768 59412 616820
rect 523132 605752 523184 605804
rect 580448 605752 580500 605804
rect 3608 603032 3660 603084
rect 59360 603032 59412 603084
rect 523684 592016 523736 592068
rect 579804 592016 579856 592068
rect 3424 587800 3476 587852
rect 59360 587800 59412 587852
rect 524328 579572 524380 579624
rect 580356 579572 580408 579624
rect 3516 573996 3568 574048
rect 59360 573996 59412 574048
rect 523132 565768 523184 565820
rect 580448 565768 580500 565820
rect 3424 560192 3476 560244
rect 59360 560192 59412 560244
rect 523776 556180 523828 556232
rect 580172 556180 580224 556232
rect 523500 545096 523552 545148
rect 580172 545096 580224 545148
rect 3424 545028 3476 545080
rect 59360 545028 59412 545080
rect 523684 539520 523736 539572
rect 580264 539520 580316 539572
rect 3424 531224 3476 531276
rect 59360 531224 59412 531276
rect 3424 516128 3476 516180
rect 59360 516128 59412 516180
rect 523776 509260 523828 509312
rect 580172 509260 580224 509312
rect 3332 500964 3384 501016
rect 59360 500964 59412 501016
rect 523684 499468 523736 499520
rect 580264 499468 580316 499520
rect 523684 498176 523736 498228
rect 580172 498176 580224 498228
rect 3424 487160 3476 487212
rect 59360 487160 59412 487212
rect 3424 473356 3476 473408
rect 59360 473356 59412 473408
rect 523684 462340 523736 462392
rect 580172 462340 580224 462392
rect 524328 459484 524380 459536
rect 580264 459484 580316 459536
rect 3516 458192 3568 458244
rect 59360 458192 59412 458244
rect 523776 451256 523828 451308
rect 580172 451256 580224 451308
rect 3424 444388 3476 444440
rect 59360 444388 59412 444440
rect 523684 438880 523736 438932
rect 580172 438880 580224 438932
rect 3516 429156 3568 429208
rect 59360 429156 59412 429208
rect 3424 415420 3476 415472
rect 59360 415420 59412 415472
rect 523684 415420 523736 415472
rect 580172 415420 580224 415472
rect 523776 404336 523828 404388
rect 580172 404336 580224 404388
rect 3608 401616 3660 401668
rect 59360 401616 59412 401668
rect 523684 391960 523736 392012
rect 580172 391960 580224 392012
rect 3516 372580 3568 372632
rect 59360 372580 59412 372632
rect 524236 368500 524288 368552
rect 580172 368500 580224 368552
rect 3424 358776 3476 358828
rect 59360 358776 59412 358828
rect 523684 357416 523736 357468
rect 580172 357416 580224 357468
rect 523776 345040 523828 345092
rect 580172 345040 580224 345092
rect 3608 338036 3660 338088
rect 60004 338036 60056 338088
rect 3608 329808 3660 329860
rect 59360 329808 59412 329860
rect 524328 322872 524380 322924
rect 580172 322872 580224 322924
rect 3700 316004 3752 316056
rect 59360 316004 59412 316056
rect 524328 311788 524380 311840
rect 580172 311788 580224 311840
rect 524328 298732 524380 298784
rect 580172 298732 580224 298784
rect 3056 295264 3108 295316
rect 60188 295264 60240 295316
rect 3516 287036 3568 287088
rect 59360 287036 59412 287088
rect 523684 275952 523736 276004
rect 580172 275952 580224 276004
rect 3608 273232 3660 273284
rect 59360 273232 59412 273284
rect 523684 264868 523736 264920
rect 580172 264868 580224 264920
rect 3148 252492 3200 252544
rect 60096 252492 60148 252544
rect 523684 252492 523736 252544
rect 579804 252492 579856 252544
rect 3424 244264 3476 244316
rect 59360 244264 59412 244316
rect 3700 229100 3752 229152
rect 59360 229100 59412 229152
rect 523684 229032 523736 229084
rect 580172 229032 580224 229084
rect 523776 217948 523828 218000
rect 580172 217948 580224 218000
rect 3148 208292 3200 208344
rect 60004 208292 60056 208344
rect 523868 205572 523920 205624
rect 579804 205572 579856 205624
rect 3516 201492 3568 201544
rect 59360 201492 59412 201544
rect 3608 186328 3660 186380
rect 59360 186328 59412 186380
rect 523684 182112 523736 182164
rect 580172 182112 580224 182164
rect 523776 171028 523828 171080
rect 580172 171028 580224 171080
rect 3424 165520 3476 165572
rect 60096 165520 60148 165572
rect 3424 158720 3476 158772
rect 59360 158720 59412 158772
rect 523868 158652 523920 158704
rect 579804 158652 579856 158704
rect 3700 143556 3752 143608
rect 59360 143556 59412 143608
rect 523684 135192 523736 135244
rect 580172 135192 580224 135244
rect 523776 124108 523828 124160
rect 580172 124108 580224 124160
rect 2964 122748 3016 122800
rect 60004 122748 60056 122800
rect 3516 115948 3568 116000
rect 59360 115948 59412 116000
rect 523868 111732 523920 111784
rect 579804 111732 579856 111784
rect 3608 100716 3660 100768
rect 59360 100716 59412 100768
rect 523684 88272 523736 88324
rect 580172 88272 580224 88324
rect 3056 79976 3108 80028
rect 60096 79976 60148 80028
rect 523776 77188 523828 77240
rect 580172 77188 580224 77240
rect 3424 73176 3476 73228
rect 59360 73176 59412 73228
rect 523868 64812 523920 64864
rect 579804 64812 579856 64864
rect 3516 57944 3568 57996
rect 59360 57944 59412 57996
rect 477224 49648 477276 49700
rect 482284 49648 482336 49700
rect 167368 49444 167420 49496
rect 227904 49444 227956 49496
rect 110236 49376 110288 49428
rect 171232 49376 171284 49428
rect 396172 49376 396224 49428
rect 456892 49376 456944 49428
rect 88708 49308 88760 49360
rect 150624 49308 150676 49360
rect 188896 49308 188948 49360
rect 249892 49308 249944 49360
rect 403348 49308 403400 49360
rect 463792 49308 463844 49360
rect 103060 49240 103112 49292
rect 164332 49240 164384 49292
rect 174544 49240 174596 49292
rect 236184 49240 236236 49292
rect 253204 49240 253256 49292
rect 313464 49240 313516 49292
rect 374736 49240 374788 49292
rect 81624 49172 81676 49224
rect 142252 49172 142304 49224
rect 145932 49172 145984 49224
rect 207112 49172 207164 49224
rect 210332 49172 210384 49224
rect 270500 49172 270552 49224
rect 367652 49172 367704 49224
rect 474832 49172 474884 49224
rect 535460 49172 535512 49224
rect 74448 49104 74500 49156
rect 135444 49104 135496 49156
rect 138848 49104 138900 49156
rect 200212 49104 200264 49156
rect 224592 49104 224644 49156
rect 285772 49104 285824 49156
rect 311624 49104 311676 49156
rect 345664 49104 345716 49156
rect 389088 49104 389140 49156
rect 449992 49104 450044 49156
rect 482008 49104 482060 49156
rect 542360 49104 542412 49156
rect 67272 49036 67324 49088
rect 128452 49036 128504 49088
rect 131672 49036 131724 49088
rect 193404 49036 193456 49088
rect 217416 49036 217468 49088
rect 278964 49036 279016 49088
rect 346124 49036 346176 49088
rect 407212 49036 407264 49088
rect 489184 49036 489236 49088
rect 549260 49036 549312 49088
rect 95884 48968 95936 49020
rect 157432 48968 157484 49020
rect 181720 48968 181772 49020
rect 242992 48968 243044 49020
rect 260380 48968 260432 49020
rect 321744 48968 321796 49020
rect 354496 48968 354548 49020
rect 367744 48968 367796 49020
rect 381912 48968 381964 49020
rect 443184 48968 443236 49020
rect 467748 48968 467800 49020
rect 528560 48968 528612 49020
rect 66076 48764 66128 48816
rect 66904 48764 66956 48816
rect 70860 48764 70912 48816
rect 71688 48764 71740 48816
rect 72056 48764 72108 48816
rect 73068 48764 73120 48816
rect 73252 48764 73304 48816
rect 74448 48764 74500 48816
rect 80428 48764 80480 48816
rect 81348 48764 81400 48816
rect 89904 48764 89956 48816
rect 91008 48764 91060 48816
rect 91100 48764 91152 48816
rect 92296 48764 92348 48816
rect 97080 48764 97132 48816
rect 97908 48764 97960 48816
rect 98276 48764 98328 48816
rect 99288 48764 99340 48816
rect 99472 48764 99524 48816
rect 100668 48764 100720 48816
rect 105452 48764 105504 48816
rect 106188 48764 106240 48816
rect 106648 48764 106700 48816
rect 107568 48764 107620 48816
rect 107844 48764 107896 48816
rect 108948 48764 109000 48816
rect 109040 48764 109092 48816
rect 110328 48764 110380 48816
rect 113732 48764 113784 48816
rect 114468 48764 114520 48816
rect 114928 48764 114980 48816
rect 115848 48764 115900 48816
rect 116124 48764 116176 48816
rect 117228 48764 117280 48816
rect 117320 48764 117372 48816
rect 118608 48764 118660 48816
rect 123300 48764 123352 48816
rect 124128 48764 124180 48816
rect 124496 48764 124548 48816
rect 125508 48764 125560 48816
rect 132868 48764 132920 48816
rect 133788 48764 133840 48816
rect 134064 48764 134116 48816
rect 135168 48764 135220 48816
rect 141148 48764 141200 48816
rect 142068 48764 142120 48816
rect 142344 48764 142396 48816
rect 143448 48764 143500 48816
rect 149520 48764 149572 48816
rect 150348 48764 150400 48816
rect 150716 48764 150768 48816
rect 151728 48764 151780 48816
rect 151912 48764 151964 48816
rect 153016 48764 153068 48816
rect 157892 48764 157944 48816
rect 158628 48764 158680 48816
rect 159088 48764 159140 48816
rect 160008 48764 160060 48816
rect 160284 48764 160336 48816
rect 161388 48764 161440 48816
rect 161480 48764 161532 48816
rect 162768 48764 162820 48816
rect 168564 48764 168616 48816
rect 169668 48764 169720 48816
rect 169760 48764 169812 48816
rect 170956 48764 171008 48816
rect 175740 48764 175792 48816
rect 176568 48764 176620 48816
rect 176936 48764 176988 48816
rect 177948 48764 178000 48816
rect 178132 48764 178184 48816
rect 179328 48764 179380 48816
rect 185308 48764 185360 48816
rect 186228 48764 186280 48816
rect 186504 48764 186556 48816
rect 187608 48764 187660 48816
rect 187700 48764 187752 48816
rect 188988 48764 189040 48816
rect 193588 48764 193640 48816
rect 194508 48764 194560 48816
rect 201960 48764 202012 48816
rect 202788 48764 202840 48816
rect 203156 48764 203208 48816
rect 204168 48764 204220 48816
rect 204352 48764 204404 48816
rect 205548 48764 205600 48816
rect 211528 48764 211580 48816
rect 212448 48764 212500 48816
rect 212724 48764 212776 48816
rect 213828 48764 213880 48816
rect 213920 48764 213972 48816
rect 215208 48764 215260 48816
rect 218612 48764 218664 48816
rect 219348 48764 219400 48816
rect 221004 48764 221056 48816
rect 222108 48764 222160 48816
rect 222200 48764 222252 48816
rect 223488 48764 223540 48816
rect 228180 48764 228232 48816
rect 229008 48764 229060 48816
rect 229376 48764 229428 48816
rect 230388 48764 230440 48816
rect 237748 48764 237800 48816
rect 238668 48764 238720 48816
rect 246028 48764 246080 48816
rect 246948 48764 247000 48816
rect 247224 48764 247276 48816
rect 248328 48764 248380 48816
rect 248420 48764 248472 48816
rect 249616 48764 249668 48816
rect 254400 48764 254452 48816
rect 255228 48764 255280 48816
rect 255596 48764 255648 48816
rect 256608 48764 256660 48816
rect 256792 48764 256844 48816
rect 257988 48764 258040 48816
rect 263968 48764 264020 48816
rect 264888 48764 264940 48816
rect 265164 48764 265216 48816
rect 266268 48764 266320 48816
rect 266360 48764 266412 48816
rect 267556 48764 267608 48816
rect 272248 48764 272300 48816
rect 273168 48764 273220 48816
rect 273444 48764 273496 48816
rect 274548 48764 274600 48816
rect 274640 48764 274692 48816
rect 275836 48764 275888 48816
rect 280620 48764 280672 48816
rect 281448 48764 281500 48816
rect 281816 48764 281868 48816
rect 282828 48764 282880 48816
rect 283012 48764 283064 48816
rect 284208 48764 284260 48816
rect 290188 48764 290240 48816
rect 291108 48764 291160 48816
rect 291384 48764 291436 48816
rect 292488 48764 292540 48816
rect 292580 48764 292632 48816
rect 293868 48764 293920 48816
rect 298468 48764 298520 48816
rect 299388 48764 299440 48816
rect 299664 48764 299716 48816
rect 300768 48764 300820 48816
rect 300860 48764 300912 48816
rect 302148 48764 302200 48816
rect 306840 48764 306892 48816
rect 307668 48764 307720 48816
rect 308036 48764 308088 48816
rect 309048 48764 309100 48816
rect 309232 48764 309284 48816
rect 310336 48764 310388 48816
rect 316408 48764 316460 48816
rect 317328 48764 317380 48816
rect 323492 48764 323544 48816
rect 324228 48764 324280 48816
rect 324688 48764 324740 48816
rect 325608 48764 325660 48816
rect 325884 48764 325936 48816
rect 326988 48764 327040 48816
rect 327080 48764 327132 48816
rect 328276 48764 328328 48816
rect 329472 48764 329524 48816
rect 330484 48764 330536 48816
rect 333060 48764 333112 48816
rect 333888 48764 333940 48816
rect 334256 48764 334308 48816
rect 335268 48764 335320 48816
rect 335452 48764 335504 48816
rect 336648 48764 336700 48816
rect 342628 48764 342680 48816
rect 343548 48764 343600 48816
rect 343732 48764 343784 48816
rect 344836 48764 344888 48816
rect 350908 48764 350960 48816
rect 351828 48764 351880 48816
rect 352104 48764 352156 48816
rect 353208 48764 353260 48816
rect 353300 48764 353352 48816
rect 354588 48764 354640 48816
rect 359280 48764 359332 48816
rect 360108 48764 360160 48816
rect 360476 48764 360528 48816
rect 361488 48764 361540 48816
rect 361672 48764 361724 48816
rect 362868 48764 362920 48816
rect 369952 48764 370004 48816
rect 371884 48764 371936 48816
rect 377128 48764 377180 48816
rect 378048 48764 378100 48816
rect 378324 48764 378376 48816
rect 379428 48764 379480 48816
rect 379520 48764 379572 48816
rect 380808 48764 380860 48816
rect 386696 48764 386748 48816
rect 387708 48764 387760 48816
rect 394976 48764 395028 48816
rect 395988 48764 396040 48816
rect 405740 48764 405792 48816
rect 406936 48764 406988 48816
rect 412916 48764 412968 48816
rect 413928 48764 413980 48816
rect 414112 48764 414164 48816
rect 415308 48764 415360 48816
rect 420092 48764 420144 48816
rect 420828 48764 420880 48816
rect 421196 48764 421248 48816
rect 422208 48764 422260 48816
rect 428372 48764 428424 48816
rect 429108 48764 429160 48816
rect 429568 48764 429620 48816
rect 430488 48764 430540 48816
rect 430764 48764 430816 48816
rect 431868 48764 431920 48816
rect 431960 48764 432012 48816
rect 433156 48764 433208 48816
rect 439136 48764 439188 48816
rect 440148 48764 440200 48816
rect 440332 48764 440384 48816
rect 441528 48764 441580 48816
rect 446220 48764 446272 48816
rect 447048 48764 447100 48816
rect 447416 48764 447468 48816
rect 448428 48764 448480 48816
rect 448612 48764 448664 48816
rect 449716 48764 449768 48816
rect 455788 48764 455840 48816
rect 456708 48764 456760 48816
rect 456984 48764 457036 48816
rect 458088 48764 458140 48816
rect 458180 48764 458232 48816
rect 459468 48764 459520 48816
rect 464160 48764 464212 48816
rect 464988 48764 465040 48816
rect 465356 48764 465408 48816
rect 466368 48764 466420 48816
rect 466552 48764 466604 48816
rect 467748 48764 467800 48816
rect 473636 48764 473688 48816
rect 474648 48764 474700 48816
rect 480812 48764 480864 48816
rect 481548 48764 481600 48816
rect 483204 48764 483256 48816
rect 484308 48764 484360 48816
rect 491576 48764 491628 48816
rect 492588 48764 492640 48816
rect 492772 48764 492824 48816
rect 493968 48764 494020 48816
rect 498660 48764 498712 48816
rect 499488 48764 499540 48816
rect 499856 48764 499908 48816
rect 500868 48764 500920 48816
rect 501052 48764 501104 48816
rect 502248 48764 502300 48816
rect 508228 48764 508280 48816
rect 509148 48764 509200 48816
rect 509424 48764 509476 48816
rect 510528 48764 510580 48816
rect 516600 48764 516652 48816
rect 517428 48764 517480 48816
rect 517796 48764 517848 48816
rect 518808 48764 518860 48816
rect 518992 48764 519044 48816
rect 520096 48764 520148 48816
rect 64880 48696 64932 48748
rect 66168 48696 66220 48748
rect 238944 48696 238996 48748
rect 240048 48696 240100 48748
rect 271052 48696 271104 48748
rect 272524 48696 272576 48748
rect 315212 48696 315264 48748
rect 315948 48696 316000 48748
rect 375932 48696 375984 48748
rect 376668 48696 376720 48748
rect 472440 48696 472492 48748
rect 474004 48696 474056 48748
rect 82820 48628 82872 48680
rect 84016 48628 84068 48680
rect 125692 48628 125744 48680
rect 126888 48628 126940 48680
rect 195980 48628 196032 48680
rect 197268 48628 197320 48680
rect 230572 48628 230624 48680
rect 231676 48628 231728 48680
rect 383108 48628 383160 48680
rect 384304 48628 384356 48680
rect 387892 48628 387944 48680
rect 389088 48628 389140 48680
rect 404544 48628 404596 48680
rect 405648 48628 405700 48680
rect 135260 48492 135312 48544
rect 136456 48492 136508 48544
rect 143540 48492 143592 48544
rect 144828 48492 144880 48544
rect 166172 48492 166224 48544
rect 167644 48492 167696 48544
rect 510620 48492 510672 48544
rect 511908 48492 511960 48544
rect 411720 48424 411772 48476
rect 412548 48424 412600 48476
rect 437940 48424 437992 48476
rect 438768 48424 438820 48476
rect 385500 48356 385552 48408
rect 386328 48356 386380 48408
rect 240140 48288 240192 48340
rect 241428 48288 241480 48340
rect 262772 48288 262824 48340
rect 263508 48288 263560 48340
rect 317604 48288 317656 48340
rect 318708 48288 318760 48340
rect 368848 48288 368900 48340
rect 369768 48288 369820 48340
rect 422392 48288 422444 48340
rect 423588 48288 423640 48340
rect 427912 48331 427964 48340
rect 427912 48297 427921 48331
rect 427921 48297 427955 48331
rect 427955 48297 427964 48331
rect 427912 48288 427964 48297
rect 434812 48331 434864 48340
rect 434812 48297 434821 48331
rect 434821 48297 434855 48331
rect 434855 48297 434864 48331
rect 434812 48288 434864 48297
rect 484400 48288 484452 48340
rect 485596 48288 485648 48340
rect 76840 47608 76892 47660
rect 138020 47608 138072 47660
rect 194784 47608 194836 47660
rect 255320 47608 255372 47660
rect 490380 47608 490432 47660
rect 550640 47608 550692 47660
rect 136548 47540 136600 47592
rect 197360 47540 197412 47592
rect 275928 47540 275980 47592
rect 336740 47540 336792 47592
rect 347320 47540 347372 47592
rect 408500 47540 408552 47592
rect 433248 47540 433300 47592
rect 494060 47540 494112 47592
rect 219808 46316 219860 46368
rect 280160 46316 280212 46368
rect 112628 46248 112680 46300
rect 173900 46248 173952 46300
rect 278228 46248 278280 46300
rect 339500 46248 339552 46300
rect 162676 46180 162728 46232
rect 223580 46180 223632 46232
rect 293684 46180 293736 46232
rect 354680 46180 354732 46232
rect 365260 46180 365312 46232
rect 425060 46180 425112 46232
rect 436744 46180 436796 46232
rect 496820 46180 496872 46232
rect 497464 46180 497516 46232
rect 557540 46180 557592 46232
rect 184848 44956 184900 45008
rect 244280 44956 244332 45008
rect 238668 44888 238720 44940
rect 298100 44888 298152 44940
rect 338028 44888 338080 44940
rect 398840 44888 398892 44940
rect 509148 44888 509200 44940
rect 568580 44888 568632 44940
rect 131028 44820 131080 44872
rect 191840 44820 191892 44872
rect 284116 44820 284168 44872
rect 345020 44820 345072 44872
rect 384948 44820 385000 44872
rect 444380 44820 444432 44872
rect 451188 44820 451240 44872
rect 512000 44820 512052 44872
rect 263508 43460 263560 43512
rect 323032 43460 323084 43512
rect 148968 43392 149020 43444
rect 209872 43392 209924 43444
rect 213828 43392 213880 43444
rect 273260 43392 273312 43444
rect 313188 43392 313240 43444
rect 374092 43392 374144 43444
rect 401508 43392 401560 43444
rect 460940 43392 460992 43444
rect 474004 43392 474056 43444
rect 532700 43392 532752 43444
rect 256608 42168 256660 42220
rect 316040 42168 316092 42220
rect 202788 42100 202840 42152
rect 262220 42100 262272 42152
rect 81348 42032 81400 42084
rect 140780 42032 140832 42084
rect 144736 42032 144788 42084
rect 205640 42032 205692 42084
rect 310336 42032 310388 42084
rect 369860 42032 369912 42084
rect 415216 42032 415268 42084
rect 476120 42032 476172 42084
rect 493876 42032 493928 42084
rect 554780 42032 554832 42084
rect 523684 41352 523736 41404
rect 580172 41352 580224 41404
rect 299388 40808 299440 40860
rect 358820 40808 358872 40860
rect 142068 40740 142120 40792
rect 201500 40740 201552 40792
rect 249616 40740 249668 40792
rect 309140 40740 309192 40792
rect 74448 40672 74500 40724
rect 133880 40672 133932 40724
rect 198648 40672 198700 40724
rect 259460 40672 259512 40724
rect 355968 40672 356020 40724
rect 416872 40672 416924 40724
rect 419448 40672 419500 40724
rect 478880 40672 478932 40724
rect 331128 39448 331180 39500
rect 390560 39448 390612 39500
rect 180708 39380 180760 39432
rect 241520 39380 241572 39432
rect 281448 39380 281500 39432
rect 340880 39380 340932 39432
rect 420828 39380 420880 39432
rect 480260 39380 480312 39432
rect 126796 39312 126848 39364
rect 187700 39312 187752 39364
rect 234528 39312 234580 39364
rect 295340 39312 295392 39364
rect 380716 39312 380768 39364
rect 441620 39312 441672 39364
rect 511816 39312 511868 39364
rect 571432 39312 571484 39364
rect 369860 38564 369912 38616
rect 369952 38564 370004 38616
rect 427912 38607 427964 38616
rect 427912 38573 427921 38607
rect 427921 38573 427955 38607
rect 427955 38573 427964 38607
rect 427912 38564 427964 38573
rect 434812 38607 434864 38616
rect 434812 38573 434821 38607
rect 434821 38573 434855 38607
rect 434855 38573 434864 38607
rect 434812 38564 434864 38573
rect 188988 37952 189040 38004
rect 248420 37952 248472 38004
rect 288348 37952 288400 38004
rect 347780 37952 347832 38004
rect 389088 37952 389140 38004
rect 448520 37952 448572 38004
rect 70308 37884 70360 37936
rect 131120 37884 131172 37936
rect 135168 37884 135220 37936
rect 194600 37884 194652 37936
rect 241336 37884 241388 37936
rect 302240 37884 302292 37936
rect 342168 37884 342220 37936
rect 401600 37884 401652 37936
rect 424968 37884 425020 37936
rect 485780 37884 485832 37936
rect 520096 37884 520148 37936
rect 578884 37884 578936 37936
rect 177948 36660 178000 36712
rect 237380 36660 237432 36712
rect 231676 36592 231728 36644
rect 291200 36592 291252 36644
rect 328276 36592 328328 36644
rect 387800 36592 387852 36644
rect 409788 36592 409840 36644
rect 469220 36592 469272 36644
rect 124128 36524 124180 36576
rect 183560 36524 183612 36576
rect 277308 36524 277360 36576
rect 338120 36524 338172 36576
rect 378048 36524 378100 36576
rect 437480 36524 437532 36576
rect 470508 36524 470560 36576
rect 529940 36524 529992 36576
rect 3332 35844 3384 35896
rect 60004 35844 60056 35896
rect 227628 35300 227680 35352
rect 287060 35300 287112 35352
rect 324228 35300 324280 35352
rect 383660 35300 383712 35352
rect 170956 35232 171008 35284
rect 230480 35232 230532 35284
rect 373908 35232 373960 35284
rect 433340 35232 433392 35284
rect 119988 35164 120040 35216
rect 180800 35164 180852 35216
rect 274548 35164 274600 35216
rect 333980 35164 334032 35216
rect 406936 35164 406988 35216
rect 466460 35164 466512 35216
rect 467748 35164 467800 35216
rect 527180 35164 527232 35216
rect 167644 33804 167696 33856
rect 227812 33804 227864 33856
rect 270408 33804 270460 33856
rect 331220 33804 331272 33856
rect 371884 33804 371936 33856
rect 430580 33804 430632 33856
rect 117228 33736 117280 33788
rect 176660 33736 176712 33788
rect 223396 33736 223448 33788
rect 284300 33736 284352 33788
rect 320088 33736 320140 33788
rect 380900 33736 380952 33788
rect 459376 33736 459428 33788
rect 520372 33736 520424 33788
rect 317328 32512 317380 32564
rect 376760 32512 376812 32564
rect 160008 32444 160060 32496
rect 219440 32444 219492 32496
rect 267556 32444 267608 32496
rect 327080 32444 327132 32496
rect 413928 32444 413980 32496
rect 473360 32444 473412 32496
rect 110328 32376 110380 32428
rect 169760 32376 169812 32428
rect 216588 32376 216640 32428
rect 277400 32376 277452 32428
rect 367008 32376 367060 32428
rect 426440 32376 426492 32428
rect 456708 32376 456760 32428
rect 516140 32376 516192 32428
rect 306288 31152 306340 31204
rect 365720 31152 365772 31204
rect 155868 31084 155920 31136
rect 216680 31084 216732 31136
rect 259368 31084 259420 31136
rect 320180 31084 320232 31136
rect 510528 31084 510580 31136
rect 569960 31084 570012 31136
rect 106188 31016 106240 31068
rect 167092 31016 167144 31068
rect 205456 31016 205508 31068
rect 266360 31016 266412 31068
rect 362776 31016 362828 31068
rect 423680 31016 423732 31068
rect 452568 31016 452620 31068
rect 512092 31016 512144 31068
rect 523776 30268 523828 30320
rect 580172 30268 580224 30320
rect 245568 29724 245620 29776
rect 305000 29724 305052 29776
rect 153016 29656 153068 29708
rect 212540 29656 212592 29708
rect 292488 29656 292540 29708
rect 351920 29656 351972 29708
rect 402888 29656 402940 29708
rect 462320 29656 462372 29708
rect 102048 29588 102100 29640
rect 162860 29588 162912 29640
rect 191748 29588 191800 29640
rect 252652 29588 252704 29640
rect 349068 29588 349120 29640
rect 408592 29588 408644 29640
rect 441436 29588 441488 29640
rect 502432 29588 502484 29640
rect 427912 29019 427964 29028
rect 427912 28985 427921 29019
rect 427921 28985 427955 29019
rect 427955 28985 427964 29019
rect 427912 28976 427964 28985
rect 434812 29019 434864 29028
rect 434812 28985 434821 29019
rect 434821 28985 434855 29019
rect 434855 28985 434864 29019
rect 434812 28976 434864 28985
rect 252468 28296 252520 28348
rect 313372 28296 313424 28348
rect 353208 28296 353260 28348
rect 412640 28296 412692 28348
rect 449716 28296 449768 28348
rect 509240 28296 509292 28348
rect 97908 28228 97960 28280
rect 158812 28228 158864 28280
rect 201408 28228 201460 28280
rect 262312 28228 262364 28280
rect 302056 28228 302108 28280
rect 362960 28228 363012 28280
rect 398748 28228 398800 28280
rect 459652 28228 459704 28280
rect 506388 28228 506440 28280
rect 565820 28228 565872 28280
rect 369860 27548 369912 27600
rect 370504 27548 370556 27600
rect 445668 27004 445720 27056
rect 505100 27004 505152 27056
rect 272524 26936 272576 26988
rect 331312 26936 331364 26988
rect 391848 26936 391900 26988
rect 451280 26936 451332 26988
rect 93768 26868 93820 26920
rect 154580 26868 154632 26920
rect 165528 26868 165580 26920
rect 226340 26868 226392 26920
rect 244188 26868 244240 26920
rect 305092 26868 305144 26920
rect 344836 26868 344888 26920
rect 404360 26868 404412 26920
rect 502156 26868 502208 26920
rect 563152 26868 563204 26920
rect 438768 25644 438820 25696
rect 498200 25644 498252 25696
rect 237288 25576 237340 25628
rect 296812 25576 296864 25628
rect 395988 25576 396040 25628
rect 455420 25576 455472 25628
rect 91008 25508 91060 25560
rect 150532 25508 150584 25560
rect 158628 25508 158680 25560
rect 218152 25508 218204 25560
rect 267648 25508 267700 25560
rect 328552 25508 328604 25560
rect 336556 25508 336608 25560
rect 397552 25508 397604 25560
rect 495348 25508 495400 25560
rect 554872 25508 554924 25560
rect 275836 24148 275888 24200
rect 335360 24148 335412 24200
rect 360108 24148 360160 24200
rect 419540 24148 419592 24200
rect 492588 24148 492640 24200
rect 552020 24148 552072 24200
rect 86868 24080 86920 24132
rect 147680 24080 147732 24132
rect 154488 24080 154540 24132
rect 215300 24080 215352 24132
rect 226248 24080 226300 24132
rect 287152 24080 287204 24132
rect 304908 24080 304960 24132
rect 365812 24080 365864 24132
rect 434628 24080 434680 24132
rect 494152 24080 494204 24132
rect 335268 22788 335320 22840
rect 394792 22788 394844 22840
rect 431868 22788 431920 22840
rect 491300 22788 491352 22840
rect 84016 22720 84068 22772
rect 143540 22720 143592 22772
rect 151728 22720 151780 22772
rect 211160 22720 211212 22772
rect 215116 22720 215168 22772
rect 276020 22720 276072 22772
rect 286968 22720 287020 22772
rect 347872 22720 347924 22772
rect 488448 22720 488500 22772
rect 547880 22720 547932 22772
rect 427728 21428 427780 21480
rect 487160 21428 487212 21480
rect 79968 21360 80020 21412
rect 140872 21360 140924 21412
rect 147588 21360 147640 21412
rect 208400 21360 208452 21412
rect 212448 21360 212500 21412
rect 271880 21360 271932 21412
rect 273168 21360 273220 21412
rect 332600 21360 332652 21412
rect 333888 21360 333940 21412
rect 393320 21360 393372 21412
rect 485596 21360 485648 21412
rect 545120 21360 545172 21412
rect 481548 20000 481600 20052
rect 540980 20000 541032 20052
rect 75828 19932 75880 19984
rect 136640 19932 136692 19984
rect 144828 19932 144880 19984
rect 204260 19932 204312 19984
rect 205548 19932 205600 19984
rect 264980 19932 265032 19984
rect 266268 19932 266320 19984
rect 325700 19932 325752 19984
rect 326988 19932 327040 19984
rect 386420 19932 386472 19984
rect 423496 19932 423548 19984
rect 484400 19932 484452 19984
rect 328460 19295 328512 19304
rect 328460 19261 328469 19295
rect 328469 19261 328503 19295
rect 328503 19261 328512 19295
rect 394700 19295 394752 19304
rect 328460 19252 328512 19261
rect 394700 19261 394709 19295
rect 394709 19261 394743 19295
rect 394743 19261 394752 19295
rect 394700 19252 394752 19261
rect 397460 19295 397512 19304
rect 397460 19261 397469 19295
rect 397469 19261 397503 19295
rect 397503 19261 397512 19295
rect 397460 19252 397512 19261
rect 427912 19295 427964 19304
rect 427912 19261 427921 19295
rect 427921 19261 427955 19295
rect 427955 19261 427964 19295
rect 427912 19252 427964 19261
rect 434812 19295 434864 19304
rect 434812 19261 434821 19295
rect 434821 19261 434855 19295
rect 434855 19261 434864 19295
rect 434812 19252 434864 19261
rect 269028 18640 269080 18692
rect 73068 18572 73120 18624
rect 132592 18572 132644 18624
rect 140688 18572 140740 18624
rect 201592 18572 201644 18624
rect 208308 18572 208360 18624
rect 269120 18572 269172 18624
rect 330484 18572 330536 18624
rect 390652 18572 390704 18624
rect 412548 18572 412600 18624
rect 471980 18572 472032 18624
rect 474648 18572 474700 18624
rect 534080 18572 534132 18624
rect 523868 17892 523920 17944
rect 579804 17892 579856 17944
rect 129648 17212 129700 17264
rect 190460 17212 190512 17264
rect 197176 17212 197228 17264
rect 258080 17212 258132 17264
rect 262128 17212 262180 17264
rect 321652 17212 321704 17264
rect 322848 17212 322900 17264
rect 382372 17212 382424 17264
rect 408408 17212 408460 17264
rect 467840 17212 467892 17264
rect 126888 15920 126940 15972
rect 186320 15920 186372 15972
rect 318616 15920 318668 15972
rect 379520 15920 379572 15972
rect 66904 15852 66956 15904
rect 126980 15852 127032 15904
rect 194508 15852 194560 15904
rect 253940 15852 253992 15904
rect 257896 15852 257948 15904
rect 318800 15852 318852 15904
rect 405648 15852 405700 15904
rect 465080 15852 465132 15904
rect 505008 15852 505060 15904
rect 564440 15852 564492 15904
rect 122748 14424 122800 14476
rect 183652 14424 183704 14476
rect 187608 14424 187660 14476
rect 247040 14424 247092 14476
rect 248328 14424 248380 14476
rect 307760 14424 307812 14476
rect 309048 14424 309100 14476
rect 368480 14424 368532 14476
rect 397368 14424 397420 14476
rect 458180 14424 458232 14476
rect 469128 14424 469180 14476
rect 528652 14424 528704 14476
rect 118516 13064 118568 13116
rect 179420 13064 179472 13116
rect 183468 13064 183520 13116
rect 244372 13064 244424 13116
rect 251088 13064 251140 13116
rect 311900 13064 311952 13116
rect 315948 13064 316000 13116
rect 375380 13064 375432 13116
rect 384304 13064 384356 13116
rect 443092 13064 443144 13116
rect 448428 13064 448480 13116
rect 507860 13064 507912 13116
rect 322940 12452 322992 12504
rect 325700 12452 325752 12504
rect 327080 12452 327132 12504
rect 324044 12384 324096 12436
rect 326436 12384 326488 12436
rect 375380 12384 375432 12436
rect 376392 12384 376444 12436
rect 376760 12384 376812 12436
rect 377588 12384 377640 12436
rect 393320 12384 393372 12436
rect 394240 12384 394292 12436
rect 408592 12384 408644 12436
rect 409696 12384 409748 12436
rect 412640 12384 412692 12436
rect 413284 12384 413336 12436
rect 327632 12316 327684 12368
rect 302148 11772 302200 11824
rect 361580 11772 361632 11824
rect 115848 11704 115900 11756
rect 175372 11704 175424 11756
rect 179236 11704 179288 11756
rect 240140 11704 240192 11756
rect 241428 11704 241480 11756
rect 300860 11704 300912 11756
rect 303528 11704 303580 11756
rect 364340 11704 364392 11756
rect 376668 11704 376720 11756
rect 437020 11704 437072 11756
rect 444288 11704 444340 11756
rect 503720 11704 503772 11756
rect 176568 10344 176620 10396
rect 236092 10344 236144 10396
rect 285588 10344 285640 10396
rect 346400 10344 346452 10396
rect 441528 10344 441580 10396
rect 500960 10344 501012 10396
rect 111708 10276 111760 10328
rect 172520 10276 172572 10328
rect 233148 10276 233200 10328
rect 293960 10276 294012 10328
rect 298008 10276 298060 10328
rect 357440 10276 357492 10328
rect 367744 10276 367796 10328
rect 415400 10276 415452 10328
rect 416688 10276 416740 10328
rect 477592 10276 477644 10328
rect 516048 10276 516100 10328
rect 575480 10276 575532 10328
rect 434812 9775 434864 9784
rect 434812 9741 434821 9775
rect 434821 9741 434855 9775
rect 434855 9741 434864 9775
rect 434812 9732 434864 9741
rect 328828 9664 328880 9716
rect 330024 9707 330076 9716
rect 330024 9673 330033 9707
rect 330033 9673 330067 9707
rect 330067 9673 330076 9707
rect 330024 9664 330076 9673
rect 395436 9664 395488 9716
rect 397828 9664 397880 9716
rect 427912 9707 427964 9716
rect 427912 9673 427921 9707
rect 427921 9673 427955 9707
rect 427955 9673 427964 9707
rect 427912 9664 427964 9673
rect 324044 9596 324096 9648
rect 326436 9596 326488 9648
rect 327632 9596 327684 9648
rect 430580 9596 430632 9648
rect 434812 9596 434864 9648
rect 324044 9460 324096 9512
rect 326436 9460 326488 9512
rect 327632 9460 327684 9512
rect 230388 8984 230440 9036
rect 290740 8984 290792 9036
rect 108948 8916 109000 8968
rect 169392 8916 169444 8968
rect 172428 8916 172480 8968
rect 233700 8916 233752 8968
rect 291108 8916 291160 8968
rect 351368 8916 351420 8968
rect 351828 8916 351880 8968
rect 412088 8916 412140 8968
rect 430488 8916 430540 8968
rect 490564 8916 490616 8968
rect 499488 8916 499540 8968
rect 559564 8916 559616 8968
rect 104808 7624 104860 7676
rect 165896 7624 165948 7676
rect 169668 7624 169720 7676
rect 230112 7624 230164 7676
rect 264888 7624 264940 7676
rect 325240 7692 325292 7744
rect 321652 7624 321704 7676
rect 322848 7624 322900 7676
rect 340788 7624 340840 7676
rect 401324 7624 401376 7676
rect 433340 7624 433392 7676
rect 434628 7624 434680 7676
rect 482284 7624 482336 7676
rect 538128 7624 538180 7676
rect 137928 7556 137980 7608
rect 199200 7556 199252 7608
rect 223488 7556 223540 7608
rect 283656 7556 283708 7608
rect 284208 7556 284260 7608
rect 344284 7556 344336 7608
rect 390560 7556 390612 7608
rect 391848 7556 391900 7608
rect 423588 7556 423640 7608
rect 483480 7556 483532 7608
rect 162768 6264 162820 6316
rect 222936 6264 222988 6316
rect 219348 6196 219400 6248
rect 279976 6196 280028 6248
rect 282828 6196 282880 6248
rect 343088 6196 343140 6248
rect 345664 6196 345716 6248
rect 372804 6196 372856 6248
rect 100576 6128 100628 6180
rect 162308 6128 162360 6180
rect 209688 6128 209740 6180
rect 270592 6128 270644 6180
rect 280068 6128 280120 6180
rect 340696 6128 340748 6180
rect 344928 6128 344980 6180
rect 406108 6128 406160 6180
rect 426348 6128 426400 6180
rect 486976 6128 487028 6180
rect 502248 6128 502300 6180
rect 561956 6128 562008 6180
rect 480168 5312 480220 5364
rect 540520 5312 540572 5364
rect 362868 5244 362920 5296
rect 422760 5244 422812 5296
rect 484308 5244 484360 5296
rect 544108 5244 544160 5296
rect 369768 5176 369820 5228
rect 429936 5176 429988 5228
rect 487068 5176 487120 5228
rect 547696 5176 547748 5228
rect 394608 5108 394660 5160
rect 454868 5108 454920 5160
rect 463608 5108 463660 5160
rect 523868 5108 523920 5160
rect 380808 5040 380860 5092
rect 440608 5040 440660 5092
rect 455328 5040 455380 5092
rect 515588 5040 515640 5092
rect 358728 4972 358780 5024
rect 419172 4972 419224 5024
rect 466368 4972 466420 5024
rect 526260 4972 526312 5024
rect 133788 4904 133840 4956
rect 194416 4904 194468 4956
rect 387708 4904 387760 4956
rect 447784 4904 447836 4956
rect 462228 4904 462280 4956
rect 522672 4904 522724 4956
rect 66168 4836 66220 4888
rect 126612 4836 126664 4888
rect 173808 4836 173860 4888
rect 234804 4836 234856 4888
rect 255228 4836 255280 4888
rect 315764 4836 315816 4888
rect 390468 4836 390520 4888
rect 68928 4768 68980 4820
rect 130200 4768 130252 4820
rect 190368 4768 190420 4820
rect 251456 4768 251508 4820
rect 295248 4768 295300 4820
rect 356152 4768 356204 4820
rect 372528 4768 372580 4820
rect 459468 4836 459520 4888
rect 519084 4836 519136 4888
rect 476028 4768 476080 4820
rect 536932 4768 536984 4820
rect 451372 4700 451424 4752
rect 143448 4088 143500 4140
rect 203892 4088 203944 4140
rect 240048 4088 240100 4140
rect 300308 4088 300360 4140
rect 353760 4088 353812 4140
rect 361488 4088 361540 4140
rect 421564 4088 421616 4140
rect 443092 4088 443144 4140
rect 444196 4088 444248 4140
rect 447048 4088 447100 4140
rect 507216 4088 507268 4140
rect 507768 4088 507820 4140
rect 567844 4088 567896 4140
rect 132592 4020 132644 4072
rect 133788 4020 133840 4072
rect 150348 4020 150400 4072
rect 211068 4020 211120 4072
rect 257988 4020 258040 4072
rect 318064 4020 318116 4072
rect 350448 4020 350500 4072
rect 410892 4020 410944 4072
rect 411168 4020 411220 4072
rect 471520 4020 471572 4072
rect 503628 4020 503680 4072
rect 564348 4020 564400 4072
rect 92296 3952 92348 4004
rect 152740 3952 152792 4004
rect 161388 3952 161440 4004
rect 221740 3952 221792 4004
rect 246948 3952 247000 4004
rect 307392 3952 307444 4004
rect 314568 3952 314620 4004
rect 375196 3952 375248 4004
rect 400128 3952 400180 4004
rect 460756 3952 460808 4004
rect 460848 3952 460900 4004
rect 521476 3952 521528 4004
rect 521568 3952 521620 4004
rect 582196 3952 582248 4004
rect 71688 3884 71740 3936
rect 132500 3884 132552 3936
rect 78588 3816 78640 3868
rect 136456 3884 136508 3936
rect 196808 3884 196860 3936
rect 200028 3884 200080 3936
rect 261024 3884 261076 3936
rect 262220 3884 262272 3936
rect 263416 3884 263468 3936
rect 307668 3884 307720 3936
rect 368020 3884 368072 3936
rect 393228 3884 393280 3936
rect 453672 3884 453724 3936
rect 464988 3884 465040 3936
rect 525064 3884 525116 3936
rect 139676 3816 139728 3868
rect 140780 3816 140832 3868
rect 142068 3816 142120 3868
rect 157248 3816 157300 3868
rect 218060 3816 218112 3868
rect 229008 3816 229060 3868
rect 289544 3816 289596 3868
rect 293868 3816 293920 3868
rect 84108 3748 84160 3800
rect 145656 3748 145708 3800
rect 150532 3748 150584 3800
rect 151544 3748 151596 3800
rect 153108 3748 153160 3800
rect 214656 3748 214708 3800
rect 222108 3748 222160 3800
rect 282460 3748 282512 3800
rect 289728 3748 289780 3800
rect 350264 3816 350316 3868
rect 354588 3816 354640 3868
rect 414480 3816 414532 3868
rect 415308 3816 415360 3868
rect 475108 3816 475160 3868
rect 500868 3816 500920 3868
rect 560760 3816 560812 3868
rect 347780 3748 347832 3800
rect 349068 3748 349120 3800
rect 379428 3748 379480 3800
rect 439412 3748 439464 3800
rect 114468 3680 114520 3732
rect 175280 3680 175332 3732
rect 206928 3680 206980 3732
rect 268108 3680 268160 3732
rect 296628 3680 296680 3732
rect 357348 3680 357400 3732
rect 357440 3680 357492 3732
rect 417976 3680 418028 3732
rect 418068 3680 418120 3732
rect 121368 3612 121420 3664
rect 182548 3612 182600 3664
rect 128268 3544 128320 3596
rect 189632 3612 189684 3664
rect 231768 3612 231820 3664
rect 293132 3612 293184 3664
rect 183560 3544 183612 3596
rect 184848 3544 184900 3596
rect 201500 3544 201552 3596
rect 202696 3544 202748 3596
rect 218152 3544 218204 3596
rect 219348 3544 219400 3596
rect 236092 3544 236144 3596
rect 237196 3544 237248 3596
rect 242808 3544 242860 3596
rect 303804 3544 303856 3596
rect 305000 3544 305052 3596
rect 306196 3544 306248 3596
rect 310428 3544 310480 3596
rect 1676 3476 1728 3528
rect 63500 3476 63552 3528
rect 88248 3476 88300 3528
rect 149244 3476 149296 3528
rect 171048 3476 171100 3528
rect 232504 3476 232556 3528
rect 244280 3476 244332 3528
rect 245568 3476 245620 3528
rect 249708 3476 249760 3528
rect 310980 3476 311032 3528
rect 321468 3476 321520 3528
rect 382280 3612 382332 3664
rect 386328 3612 386380 3664
rect 446588 3748 446640 3800
rect 471888 3748 471940 3800
rect 528652 3748 528704 3800
rect 529848 3748 529900 3800
rect 478696 3680 478748 3732
rect 513288 3680 513340 3732
rect 573824 3680 573876 3732
rect 451280 3612 451332 3664
rect 452476 3612 452528 3664
rect 467840 3612 467892 3664
rect 469128 3612 469180 3664
rect 478788 3612 478840 3664
rect 539324 3612 539376 3664
rect 371608 3544 371660 3596
rect 382372 3544 382424 3596
rect 383568 3544 383620 3596
rect 422208 3544 422260 3596
rect 482284 3544 482336 3596
rect 494152 3544 494204 3596
rect 495348 3544 495400 3596
rect 496728 3544 496780 3596
rect 557172 3544 557224 3596
rect 328368 3476 328420 3528
rect 389456 3476 389508 3528
rect 425060 3476 425112 3528
rect 426348 3476 426400 3528
rect 429108 3476 429160 3528
rect 489368 3476 489420 3528
rect 493968 3476 494020 3528
rect 553584 3476 553636 3528
rect 571432 3476 571484 3528
rect 572628 3476 572680 3528
rect 578884 3476 578936 3528
rect 579804 3476 579856 3528
rect 572 3408 624 3460
rect 62120 3408 62172 3460
rect 95148 3408 95200 3460
rect 156328 3408 156380 3460
rect 164148 3408 164200 3460
rect 225328 3408 225380 3460
rect 235908 3408 235960 3460
rect 296720 3408 296772 3460
rect 300768 3408 300820 3460
rect 360936 3408 360988 3460
rect 365720 3408 365772 3460
rect 366916 3408 366968 3460
rect 371148 3408 371200 3460
rect 432328 3408 432380 3460
rect 440148 3408 440200 3460
rect 500132 3408 500184 3460
rect 517428 3408 517480 3460
rect 577412 3408 577464 3460
rect 125508 3340 125560 3392
rect 186044 3340 186096 3392
rect 215208 3340 215260 3392
rect 118608 3272 118660 3324
rect 107568 3204 107620 3256
rect 168196 3204 168248 3256
rect 175372 3272 175424 3324
rect 176568 3272 176620 3324
rect 204168 3272 204220 3324
rect 264612 3272 264664 3324
rect 178960 3204 179012 3256
rect 197268 3204 197320 3256
rect 257436 3204 257488 3256
rect 270500 3340 270552 3392
rect 271696 3340 271748 3392
rect 287060 3340 287112 3392
rect 288348 3340 288400 3392
rect 336648 3340 336700 3392
rect 396632 3340 396684 3392
rect 436008 3340 436060 3392
rect 496544 3340 496596 3392
rect 511908 3340 511960 3392
rect 571432 3340 571484 3392
rect 318708 3272 318760 3324
rect 378784 3272 378836 3324
rect 453948 3272 454000 3324
rect 514392 3272 514444 3324
rect 514668 3272 514720 3324
rect 575020 3272 575072 3324
rect 275284 3204 275336 3256
rect 325608 3204 325660 3256
rect 385868 3204 385920 3256
rect 458088 3204 458140 3256
rect 517888 3204 517940 3256
rect 518808 3204 518860 3256
rect 578608 3204 578660 3256
rect 100668 3136 100720 3188
rect 161112 3136 161164 3188
rect 193128 3136 193180 3188
rect 253848 3136 253900 3188
rect 332508 3136 332560 3188
rect 393044 3136 393096 3188
rect 442908 3136 442960 3188
rect 503628 3136 503680 3188
rect 532240 3136 532292 3188
rect 99288 3068 99340 3120
rect 159916 3068 159968 3120
rect 179328 3068 179380 3120
rect 239588 3068 239640 3120
rect 343548 3068 343600 3120
rect 403716 3068 403768 3120
rect 433156 3068 433208 3120
rect 492956 3068 493008 3120
rect 186228 3000 186280 3052
rect 246764 3000 246816 3052
rect 374092 2796 374144 2848
rect 427912 2796 427964 2848
rect 374000 2728 374052 2780
rect 428740 2728 428792 2780
rect 433524 2320 433576 2372
rect 328828 552 328880 604
rect 328920 552 328972 604
rect 354680 552 354732 604
rect 354956 552 355008 604
rect 357532 552 357584 604
rect 358544 552 358596 604
rect 358820 552 358872 604
rect 359740 552 359792 604
rect 361580 552 361632 604
rect 362132 552 362184 604
rect 383660 552 383712 604
rect 384672 552 384724 604
rect 386420 552 386472 604
rect 387064 552 387116 604
rect 387800 552 387852 604
rect 388260 552 388312 604
rect 431132 595 431184 604
rect 431132 561 431141 595
rect 431141 561 431175 595
rect 431175 561 431184 595
rect 431132 552 431184 561
rect 435824 595 435876 604
rect 435824 561 435833 595
rect 435833 561 435867 595
rect 435867 561 435876 595
rect 435824 552 435876 561
rect 455420 552 455472 604
rect 456064 552 456116 604
rect 456892 552 456944 604
rect 457260 552 457312 604
rect 471980 552 472032 604
rect 472716 552 472768 604
rect 473360 552 473412 604
rect 473912 552 473964 604
rect 478880 552 478932 604
rect 479892 552 479944 604
rect 557540 552 557592 604
rect 558368 552 558420 604
rect 564440 552 564492 604
rect 565544 552 565596 604
rect 565820 552 565872 604
rect 566740 552 566792 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3606 682272 3662 682281
rect 3606 682207 3662 682216
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3436 630630 3464 667927
rect 3514 653576 3570 653585
rect 3514 653511 3570 653520
rect 3424 630624 3476 630630
rect 3424 630566 3476 630572
rect 3528 616826 3556 653511
rect 3620 645862 3648 682207
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654974 8064 663734
rect 8024 654968 8076 654974
rect 8024 654910 8076 654916
rect 24780 654838 24808 699654
rect 41340 654906 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 692782 72740 698278
rect 72700 692776 72752 692782
rect 72700 692718 72752 692724
rect 72516 683256 72568 683262
rect 72516 683198 72568 683204
rect 72528 683126 72556 683198
rect 72516 683120 72568 683126
rect 72516 683062 72568 683068
rect 72700 678904 72752 678910
rect 72700 678846 72752 678852
rect 72712 669322 72740 678846
rect 72700 669316 72752 669322
rect 72700 669258 72752 669264
rect 72884 669316 72936 669322
rect 72884 669258 72936 669264
rect 72896 666534 72924 669258
rect 72884 666528 72936 666534
rect 72884 666470 72936 666476
rect 72792 656940 72844 656946
rect 72792 656882 72844 656888
rect 72804 654974 72832 656882
rect 70492 654968 70544 654974
rect 70492 654910 70544 654916
rect 72792 654968 72844 654974
rect 72792 654910 72844 654916
rect 41328 654900 41380 654906
rect 41328 654842 41380 654848
rect 24768 654832 24820 654838
rect 24768 654774 24820 654780
rect 70504 651916 70532 654910
rect 89640 654838 89668 699654
rect 106200 654906 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654974 137784 663734
rect 121552 654968 121604 654974
rect 121552 654910 121604 654916
rect 137744 654968 137796 654974
rect 137744 654910 137796 654916
rect 104532 654900 104584 654906
rect 104532 654842 104584 654848
rect 106188 654900 106240 654906
rect 106188 654842 106240 654848
rect 87512 654832 87564 654838
rect 87512 654774 87564 654780
rect 89628 654832 89680 654838
rect 89628 654774 89680 654780
rect 87524 651916 87552 654774
rect 104544 651916 104572 654842
rect 121564 651916 121592 654910
rect 154316 654838 154344 663734
rect 171060 654906 171088 700198
rect 172704 654968 172756 654974
rect 172704 654910 172756 654916
rect 155592 654900 155644 654906
rect 155592 654842 155644 654848
rect 171048 654900 171100 654906
rect 171048 654842 171100 654848
rect 138572 654832 138624 654838
rect 138572 654774 138624 654780
rect 154304 654832 154356 654838
rect 154304 654774 154356 654780
rect 138584 651916 138612 654774
rect 155604 651916 155632 654842
rect 172716 651916 172744 654910
rect 202800 654838 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 679046 219112 685850
rect 219072 679040 219124 679046
rect 219072 678982 219124 678988
rect 218980 678972 219032 678978
rect 218980 678914 219032 678920
rect 218992 669322 219020 678914
rect 218980 669316 219032 669322
rect 218980 669258 219032 669264
rect 219164 669316 219216 669322
rect 219164 669258 219216 669264
rect 219176 666534 219204 669258
rect 219164 666528 219216 666534
rect 219164 666470 219216 666476
rect 219072 656940 219124 656946
rect 219072 656882 219124 656888
rect 219084 654906 219112 656882
rect 206744 654900 206796 654906
rect 206744 654842 206796 654848
rect 219072 654900 219124 654906
rect 219072 654842 219124 654848
rect 189724 654832 189776 654838
rect 189724 654774 189776 654780
rect 202788 654832 202840 654838
rect 202788 654774 202840 654780
rect 189736 651916 189764 654774
rect 206756 651916 206784 654842
rect 235920 654838 235948 699654
rect 240784 654900 240836 654906
rect 240784 654842 240836 654848
rect 223764 654832 223816 654838
rect 223764 654774 223816 654780
rect 235908 654832 235960 654838
rect 235908 654774 235960 654780
rect 223776 651916 223804 654774
rect 240796 651916 240824 654842
rect 267660 654838 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 343548 700324 343600 700330
rect 343548 700266 343600 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 326988 699712 327040 699718
rect 326988 699654 327040 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654838 284064 663734
rect 257896 654832 257948 654838
rect 257896 654774 257948 654780
rect 267648 654832 267700 654838
rect 267648 654774 267700 654780
rect 274916 654832 274968 654838
rect 274916 654774 274968 654780
rect 284024 654832 284076 654838
rect 284024 654774 284076 654780
rect 291936 654832 291988 654838
rect 291936 654774 291988 654780
rect 257908 651916 257936 654774
rect 274928 651916 274956 654774
rect 291948 651916 291976 654774
rect 300780 654158 300808 699654
rect 327000 655178 327028 699654
rect 325976 655172 326028 655178
rect 325976 655114 326028 655120
rect 326988 655172 327040 655178
rect 326988 655114 327040 655120
rect 300768 654152 300820 654158
rect 300768 654094 300820 654100
rect 308956 654152 309008 654158
rect 308956 654094 309008 654100
rect 308968 651916 308996 654094
rect 325988 651916 326016 655114
rect 343560 651794 343588 700266
rect 364996 699718 365024 703520
rect 394608 700392 394660 700398
rect 394608 700334 394660 700340
rect 378048 700324 378100 700330
rect 378048 700266 378100 700272
rect 360108 699712 360160 699718
rect 360108 699654 360160 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 360120 651916 360148 699654
rect 378060 655518 378088 700266
rect 377128 655512 377180 655518
rect 377128 655454 377180 655460
rect 378048 655512 378100 655518
rect 378048 655454 378100 655460
rect 377140 651916 377168 655454
rect 394620 651794 394648 700334
rect 397472 700330 397500 703520
rect 411168 700460 411220 700466
rect 411168 700402 411220 700408
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 411180 651916 411208 700402
rect 413664 700398 413692 703520
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 445668 700392 445720 700398
rect 445668 700334 445720 700340
rect 429108 700324 429160 700330
rect 429108 700266 429160 700272
rect 429120 655518 429148 700266
rect 428188 655512 428240 655518
rect 428188 655454 428240 655460
rect 429108 655512 429160 655518
rect 429108 655454 429160 655460
rect 428200 651916 428228 655454
rect 445680 651930 445708 700334
rect 462332 700330 462360 703520
rect 463608 700460 463660 700466
rect 463608 700402 463660 700408
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 463620 655518 463648 700402
rect 478524 700398 478552 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 514668 700460 514720 700466
rect 514668 700402 514720 700408
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 496728 700392 496780 700398
rect 496728 700334 496780 700340
rect 480168 700324 480220 700330
rect 480168 700266 480220 700272
rect 480180 655518 480208 700266
rect 462320 655512 462372 655518
rect 462320 655454 462372 655460
rect 463608 655512 463660 655518
rect 463608 655454 463660 655460
rect 479340 655512 479392 655518
rect 479340 655454 479392 655460
rect 480168 655512 480220 655518
rect 480168 655454 480220 655460
rect 445326 651902 445708 651930
rect 462332 651916 462360 655454
rect 479352 651916 479380 655454
rect 496740 651930 496768 700334
rect 514680 655314 514708 700402
rect 527192 700330 527220 703520
rect 543476 700398 543504 703520
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 523776 696992 523828 696998
rect 523776 696934 523828 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 523684 685908 523736 685914
rect 523684 685850 523736 685856
rect 513380 655308 513432 655314
rect 513380 655250 513432 655256
rect 514668 655308 514720 655314
rect 514668 655250 514720 655256
rect 496386 651902 496768 651930
rect 513392 651916 513420 655250
rect 343022 651766 343588 651794
rect 394174 651766 394648 651794
rect 3608 645856 3660 645862
rect 3608 645798 3660 645804
rect 59360 645856 59412 645862
rect 59360 645798 59412 645804
rect 59372 644745 59400 645798
rect 59358 644736 59414 644745
rect 59358 644671 59414 644680
rect 523696 631961 523724 685850
rect 523788 645289 523816 696934
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 523774 645280 523830 645289
rect 523774 645215 523830 645224
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 523776 638988 523828 638994
rect 523776 638930 523828 638936
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 523682 631952 523738 631961
rect 523682 631887 523738 631896
rect 59360 630624 59412 630630
rect 59360 630566 59412 630572
rect 59372 630465 59400 630566
rect 59358 630456 59414 630465
rect 59358 630391 59414 630400
rect 3606 624880 3662 624889
rect 3606 624815 3662 624824
rect 3516 616820 3568 616826
rect 3516 616762 3568 616768
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 587858 3464 610399
rect 3620 603090 3648 624815
rect 59360 616820 59412 616826
rect 59360 616762 59412 616768
rect 59372 616185 59400 616762
rect 59358 616176 59414 616185
rect 59358 616111 59414 616120
rect 523132 605804 523184 605810
rect 523132 605746 523184 605752
rect 523144 605305 523172 605746
rect 523130 605296 523186 605305
rect 523130 605231 523186 605240
rect 3608 603084 3660 603090
rect 3608 603026 3660 603032
rect 59360 603084 59412 603090
rect 59360 603026 59412 603032
rect 59372 601905 59400 603026
rect 59358 601896 59414 601905
rect 59358 601831 59414 601840
rect 3514 596048 3570 596057
rect 3514 595983 3570 595992
rect 3424 587852 3476 587858
rect 3424 587794 3476 587800
rect 3528 574054 3556 595983
rect 523684 592068 523736 592074
rect 523684 592010 523736 592016
rect 59360 587852 59412 587858
rect 59360 587794 59412 587800
rect 59372 587625 59400 587794
rect 59358 587616 59414 587625
rect 59358 587551 59414 587560
rect 3516 574048 3568 574054
rect 3516 573990 3568 573996
rect 59360 574048 59412 574054
rect 59360 573990 59412 573996
rect 59372 573345 59400 573990
rect 59358 573336 59414 573345
rect 59358 573271 59414 573280
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 560250 3464 567287
rect 523132 565820 523184 565826
rect 523132 565762 523184 565768
rect 523144 565321 523172 565762
rect 523130 565312 523186 565321
rect 523130 565247 523186 565256
rect 3424 560244 3476 560250
rect 3424 560186 3476 560192
rect 59360 560244 59412 560250
rect 59360 560186 59412 560192
rect 59372 559065 59400 560186
rect 59358 559056 59414 559065
rect 59358 558991 59414 559000
rect 3422 553072 3478 553081
rect 3422 553007 3478 553016
rect 3436 545086 3464 553007
rect 523696 551993 523724 592010
rect 523788 591977 523816 638930
rect 580276 619614 580304 674591
rect 580446 651128 580502 651137
rect 580446 651063 580502 651072
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 524328 619608 524380 619614
rect 524328 619550 524380 619556
rect 580264 619608 580316 619614
rect 580264 619550 580316 619556
rect 524340 618633 524368 619550
rect 524326 618624 524382 618633
rect 524326 618559 524382 618568
rect 579802 592512 579858 592521
rect 579802 592447 579858 592456
rect 579816 592074 579844 592447
rect 579804 592068 579856 592074
rect 579804 592010 579856 592016
rect 523774 591968 523830 591977
rect 523774 591903 523830 591912
rect 580262 580816 580318 580825
rect 580262 580751 580318 580760
rect 524328 579624 524380 579630
rect 524328 579566 524380 579572
rect 524340 578649 524368 579566
rect 524326 578640 524382 578649
rect 524326 578575 524382 578584
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 523776 556232 523828 556238
rect 523776 556174 523828 556180
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 523682 551984 523738 551993
rect 523682 551919 523738 551928
rect 523500 545148 523552 545154
rect 523500 545090 523552 545096
rect 3424 545080 3476 545086
rect 3424 545022 3476 545028
rect 59360 545080 59412 545086
rect 59360 545022 59412 545028
rect 59372 544785 59400 545022
rect 59358 544776 59414 544785
rect 59358 544711 59414 544720
rect 3422 538656 3478 538665
rect 3422 538591 3478 538600
rect 3436 531282 3464 538591
rect 523512 538234 523540 545090
rect 523684 539572 523736 539578
rect 523684 539514 523736 539520
rect 523696 538665 523724 539514
rect 523682 538656 523738 538665
rect 523682 538591 523738 538600
rect 523512 538206 523724 538234
rect 3424 531276 3476 531282
rect 3424 531218 3476 531224
rect 59360 531276 59412 531282
rect 59360 531218 59412 531224
rect 59372 530505 59400 531218
rect 59358 530496 59414 530505
rect 59358 530431 59414 530440
rect 59358 516216 59414 516225
rect 3424 516180 3476 516186
rect 59358 516151 59360 516160
rect 3424 516122 3476 516128
rect 59412 516151 59414 516160
rect 59360 516122 59412 516128
rect 3436 509969 3464 516122
rect 523696 512009 523724 538206
rect 523788 525337 523816 556174
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580276 539578 580304 580751
rect 580368 579630 580396 627671
rect 580460 605810 580488 651063
rect 580448 605804 580500 605810
rect 580448 605746 580500 605752
rect 580446 604208 580502 604217
rect 580446 604143 580502 604152
rect 580356 579624 580408 579630
rect 580356 579566 580408 579572
rect 580460 565826 580488 604143
rect 580448 565820 580500 565826
rect 580448 565762 580500 565768
rect 580264 539572 580316 539578
rect 580264 539514 580316 539520
rect 580262 533896 580318 533905
rect 580262 533831 580318 533840
rect 523774 525328 523830 525337
rect 523774 525263 523830 525272
rect 523682 512000 523738 512009
rect 523682 511935 523738 511944
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 3422 509960 3478 509969
rect 3422 509895 3478 509904
rect 580184 509318 580212 510303
rect 523776 509312 523828 509318
rect 523776 509254 523828 509260
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 59358 501936 59414 501945
rect 59358 501871 59414 501880
rect 59372 501022 59400 501871
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 59360 501016 59412 501022
rect 59360 500958 59412 500964
rect 3344 495553 3372 500958
rect 523684 499520 523736 499526
rect 523684 499462 523736 499468
rect 523696 498681 523724 499462
rect 523682 498672 523738 498681
rect 523682 498607 523738 498616
rect 523684 498228 523736 498234
rect 523684 498170 523736 498176
rect 3330 495544 3386 495553
rect 3330 495479 3386 495488
rect 59358 487656 59414 487665
rect 59358 487591 59414 487600
rect 59372 487218 59400 487591
rect 3424 487212 3476 487218
rect 3424 487154 3476 487160
rect 59360 487212 59412 487218
rect 59360 487154 59412 487160
rect 3436 481137 3464 487154
rect 3422 481128 3478 481137
rect 3422 481063 3478 481072
rect 3424 473408 3476 473414
rect 59360 473408 59412 473414
rect 3424 473350 3476 473356
rect 59358 473376 59360 473385
rect 59412 473376 59414 473385
rect 3436 452441 3464 473350
rect 59358 473311 59414 473320
rect 523696 472025 523724 498170
rect 523788 485353 523816 509254
rect 580276 499526 580304 533831
rect 580264 499520 580316 499526
rect 580264 499462 580316 499468
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580262 486840 580318 486849
rect 580262 486775 580318 486784
rect 523774 485344 523830 485353
rect 523774 485279 523830 485288
rect 523682 472016 523738 472025
rect 523682 471951 523738 471960
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 523684 462392 523736 462398
rect 523684 462334 523736 462340
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 59358 459096 59414 459105
rect 59358 459031 59414 459040
rect 59372 458250 59400 459031
rect 3516 458244 3568 458250
rect 3516 458186 3568 458192
rect 59360 458244 59412 458250
rect 59360 458186 59412 458192
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 3424 444440 3476 444446
rect 3424 444382 3476 444388
rect 3436 423745 3464 444382
rect 3528 438025 3556 458186
rect 523696 445369 523724 462334
rect 580276 459542 580304 486775
rect 524328 459536 524380 459542
rect 524328 459478 524380 459484
rect 580264 459536 580316 459542
rect 580264 459478 580316 459484
rect 524340 458697 524368 459478
rect 524326 458688 524382 458697
rect 524326 458623 524382 458632
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 523776 451308 523828 451314
rect 523776 451250 523828 451256
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 523682 445360 523738 445369
rect 523682 445295 523738 445304
rect 59358 444816 59414 444825
rect 59358 444751 59414 444760
rect 59372 444446 59400 444751
rect 59360 444440 59412 444446
rect 59360 444382 59412 444388
rect 523684 438932 523736 438938
rect 523684 438874 523736 438880
rect 3514 438016 3570 438025
rect 3514 437951 3570 437960
rect 59358 430536 59414 430545
rect 59358 430471 59414 430480
rect 59372 429214 59400 430471
rect 3516 429208 3568 429214
rect 3516 429150 3568 429156
rect 59360 429208 59412 429214
rect 59360 429150 59412 429156
rect 3422 423736 3478 423745
rect 3422 423671 3478 423680
rect 3424 415472 3476 415478
rect 3424 415414 3476 415420
rect 3436 380633 3464 415414
rect 3528 395049 3556 429150
rect 523696 418713 523724 438874
rect 523788 432041 523816 451250
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 523774 432032 523830 432041
rect 523774 431967 523830 431976
rect 523682 418704 523738 418713
rect 523682 418639 523738 418648
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 59358 416256 59414 416265
rect 59358 416191 59414 416200
rect 59372 415478 59400 416191
rect 580184 415478 580212 416463
rect 59360 415472 59412 415478
rect 59360 415414 59412 415420
rect 523684 415472 523736 415478
rect 523684 415414 523736 415420
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 523696 405385 523724 415414
rect 523682 405376 523738 405385
rect 523682 405311 523738 405320
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 523776 404388 523828 404394
rect 523776 404330 523828 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 59358 401976 59414 401985
rect 59358 401911 59414 401920
rect 59372 401674 59400 401911
rect 3608 401668 3660 401674
rect 3608 401610 3660 401616
rect 59360 401668 59412 401674
rect 59360 401610 59412 401616
rect 3514 395040 3570 395049
rect 3514 394975 3570 394984
rect 3422 380624 3478 380633
rect 3422 380559 3478 380568
rect 3516 372632 3568 372638
rect 3516 372574 3568 372580
rect 3424 358828 3476 358834
rect 3424 358770 3476 358776
rect 3436 308825 3464 358770
rect 3528 323105 3556 372574
rect 3620 366217 3648 401610
rect 523788 392057 523816 404330
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 523774 392048 523830 392057
rect 523684 392012 523736 392018
rect 580184 392018 580212 392935
rect 523774 391983 523830 391992
rect 580172 392012 580224 392018
rect 523684 391954 523736 391960
rect 580172 391954 580224 391960
rect 60002 387696 60058 387705
rect 60002 387631 60058 387640
rect 59358 373416 59414 373425
rect 59358 373351 59414 373360
rect 59372 372638 59400 373351
rect 59360 372632 59412 372638
rect 59360 372574 59412 372580
rect 3606 366208 3662 366217
rect 3606 366143 3662 366152
rect 59358 359136 59414 359145
rect 59358 359071 59414 359080
rect 59372 358834 59400 359071
rect 59360 358828 59412 358834
rect 59360 358770 59412 358776
rect 60016 338094 60044 387631
rect 523696 378729 523724 391954
rect 523682 378720 523738 378729
rect 523682 378655 523738 378664
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 524236 368552 524288 368558
rect 524236 368494 524288 368500
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 524248 365401 524276 368494
rect 524234 365392 524290 365401
rect 524234 365327 524290 365336
rect 580170 357912 580226 357921
rect 580170 357847 580226 357856
rect 580184 357474 580212 357847
rect 523684 357468 523736 357474
rect 523684 357410 523736 357416
rect 580172 357468 580224 357474
rect 580172 357410 580224 357416
rect 523696 351937 523724 357410
rect 523682 351928 523738 351937
rect 523682 351863 523738 351872
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345098 580212 346015
rect 523776 345092 523828 345098
rect 523776 345034 523828 345040
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 60186 344720 60242 344729
rect 60186 344655 60242 344664
rect 3608 338088 3660 338094
rect 3608 338030 3660 338036
rect 60004 338088 60056 338094
rect 60004 338030 60056 338036
rect 3620 337521 3648 338030
rect 3606 337512 3662 337521
rect 3606 337447 3662 337456
rect 59358 330440 59414 330449
rect 59358 330375 59414 330384
rect 59372 329866 59400 330375
rect 3608 329860 3660 329866
rect 3608 329802 3660 329808
rect 59360 329860 59412 329866
rect 59360 329802 59412 329808
rect 3514 323096 3570 323105
rect 3514 323031 3570 323040
rect 3422 308816 3478 308825
rect 3422 308751 3478 308760
rect 3056 295316 3108 295322
rect 3056 295258 3108 295264
rect 3068 294409 3096 295258
rect 3054 294400 3110 294409
rect 3054 294335 3110 294344
rect 3516 287088 3568 287094
rect 3516 287030 3568 287036
rect 3148 252544 3200 252550
rect 3148 252486 3200 252492
rect 3160 251297 3188 252486
rect 3146 251288 3202 251297
rect 3146 251223 3202 251232
rect 3424 244316 3476 244322
rect 3424 244258 3476 244264
rect 3148 208344 3200 208350
rect 3148 208286 3200 208292
rect 3160 208185 3188 208286
rect 3146 208176 3202 208185
rect 3146 208111 3202 208120
rect 3436 193905 3464 244258
rect 3528 237017 3556 287030
rect 3620 280129 3648 329802
rect 59358 316160 59414 316169
rect 59358 316095 59414 316104
rect 59372 316062 59400 316095
rect 3700 316056 3752 316062
rect 3700 315998 3752 316004
rect 59360 316056 59412 316062
rect 59360 315998 59412 316004
rect 3606 280120 3662 280129
rect 3606 280055 3662 280064
rect 3608 273284 3660 273290
rect 3608 273226 3660 273232
rect 3514 237008 3570 237017
rect 3514 236943 3570 236952
rect 3620 222601 3648 273226
rect 3712 265713 3740 315998
rect 60094 301880 60150 301889
rect 60094 301815 60150 301824
rect 59358 287600 59414 287609
rect 59358 287535 59414 287544
rect 59372 287094 59400 287535
rect 59360 287088 59412 287094
rect 59360 287030 59412 287036
rect 59358 273320 59414 273329
rect 59358 273255 59360 273264
rect 59412 273255 59414 273264
rect 59360 273226 59412 273232
rect 3698 265704 3754 265713
rect 3698 265639 3754 265648
rect 60002 259040 60058 259049
rect 60002 258975 60058 258984
rect 59358 244760 59414 244769
rect 59358 244695 59414 244704
rect 59372 244322 59400 244695
rect 59360 244316 59412 244322
rect 59360 244258 59412 244264
rect 59358 230480 59414 230489
rect 59358 230415 59414 230424
rect 59372 229158 59400 230415
rect 3700 229152 3752 229158
rect 3700 229094 3752 229100
rect 59360 229152 59412 229158
rect 59360 229094 59412 229100
rect 3606 222592 3662 222601
rect 3606 222527 3662 222536
rect 3516 201544 3568 201550
rect 3516 201486 3568 201492
rect 3422 193896 3478 193905
rect 3422 193831 3478 193840
rect 3424 165572 3476 165578
rect 3424 165514 3476 165520
rect 3436 165073 3464 165514
rect 3422 165064 3478 165073
rect 3422 164999 3478 165008
rect 3424 158772 3476 158778
rect 3424 158714 3476 158720
rect 2964 122800 3016 122806
rect 2964 122742 3016 122748
rect 2976 122097 3004 122742
rect 2962 122088 3018 122097
rect 2962 122023 3018 122032
rect 3436 107681 3464 158714
rect 3528 150793 3556 201486
rect 3608 186380 3660 186386
rect 3608 186322 3660 186328
rect 3514 150784 3570 150793
rect 3514 150719 3570 150728
rect 3620 136377 3648 186322
rect 3712 179489 3740 229094
rect 60016 208350 60044 258975
rect 60108 252550 60136 301815
rect 60200 295322 60228 344655
rect 523788 338609 523816 345034
rect 523774 338600 523830 338609
rect 523774 338535 523830 338544
rect 524326 325272 524382 325281
rect 524326 325207 524382 325216
rect 524340 322930 524368 325207
rect 524328 322924 524380 322930
rect 524328 322866 524380 322872
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 524326 311944 524382 311953
rect 524326 311879 524382 311888
rect 524340 311846 524368 311879
rect 524328 311840 524380 311846
rect 524328 311782 524380 311788
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580184 298790 580212 299095
rect 524328 298784 524380 298790
rect 524328 298726 524380 298732
rect 580172 298784 580224 298790
rect 580172 298726 580224 298732
rect 524340 298625 524368 298726
rect 524326 298616 524382 298625
rect 524326 298551 524382 298560
rect 60188 295316 60240 295322
rect 60188 295258 60240 295264
rect 523682 285288 523738 285297
rect 523682 285223 523738 285232
rect 523696 276010 523724 285223
rect 523684 276004 523736 276010
rect 523684 275946 523736 275952
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 523682 271960 523738 271969
rect 523682 271895 523738 271904
rect 523696 264926 523724 271895
rect 523684 264920 523736 264926
rect 523684 264862 523736 264868
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 523682 258632 523738 258641
rect 523682 258567 523738 258576
rect 523696 252550 523724 258567
rect 60096 252544 60148 252550
rect 60096 252486 60148 252492
rect 523684 252544 523736 252550
rect 523684 252486 523736 252492
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 523682 245304 523738 245313
rect 523682 245239 523738 245248
rect 523696 229090 523724 245239
rect 523774 231976 523830 231985
rect 523774 231911 523830 231920
rect 523684 229084 523736 229090
rect 523684 229026 523736 229032
rect 523788 218006 523816 231911
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 523866 218648 523922 218657
rect 523866 218583 523922 218592
rect 523776 218000 523828 218006
rect 523776 217942 523828 217948
rect 60094 216200 60150 216209
rect 60094 216135 60150 216144
rect 60004 208344 60056 208350
rect 60004 208286 60056 208292
rect 59358 201920 59414 201929
rect 59358 201855 59414 201864
rect 59372 201550 59400 201855
rect 59360 201544 59412 201550
rect 59360 201486 59412 201492
rect 59358 187640 59414 187649
rect 59358 187575 59414 187584
rect 59372 186386 59400 187575
rect 59360 186380 59412 186386
rect 59360 186322 59412 186328
rect 3698 179480 3754 179489
rect 3698 179415 3754 179424
rect 60002 173360 60058 173369
rect 60002 173295 60058 173304
rect 59358 159080 59414 159089
rect 59358 159015 59414 159024
rect 59372 158778 59400 159015
rect 59360 158772 59412 158778
rect 59360 158714 59412 158720
rect 59358 144800 59414 144809
rect 59358 144735 59414 144744
rect 59372 143614 59400 144735
rect 3700 143608 3752 143614
rect 3700 143550 3752 143556
rect 59360 143608 59412 143614
rect 59360 143550 59412 143556
rect 3606 136368 3662 136377
rect 3606 136303 3662 136312
rect 3516 116000 3568 116006
rect 3516 115942 3568 115948
rect 3422 107672 3478 107681
rect 3422 107607 3478 107616
rect 3056 80028 3108 80034
rect 3056 79970 3108 79976
rect 3068 78985 3096 79970
rect 3054 78976 3110 78985
rect 3054 78911 3110 78920
rect 3424 73228 3476 73234
rect 3424 73170 3476 73176
rect 3332 35896 3384 35902
rect 3330 35864 3332 35873
rect 3384 35864 3386 35873
rect 3330 35799 3386 35808
rect 3436 21457 3464 73170
rect 3528 64569 3556 115942
rect 3608 100768 3660 100774
rect 3608 100710 3660 100716
rect 3514 64560 3570 64569
rect 3514 64495 3570 64504
rect 3516 57996 3568 58002
rect 3516 57938 3568 57944
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3528 7177 3556 57938
rect 3620 50153 3648 100710
rect 3712 93265 3740 143550
rect 60016 122806 60044 173295
rect 60108 165578 60136 216135
rect 523880 205630 523908 218583
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 523868 205624 523920 205630
rect 523868 205566 523920 205572
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 523682 205320 523738 205329
rect 523682 205255 523738 205264
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 523696 182170 523724 205255
rect 523774 191992 523830 192001
rect 523774 191927 523830 191936
rect 523684 182164 523736 182170
rect 523684 182106 523736 182112
rect 523788 171086 523816 191927
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 523866 178664 523922 178673
rect 523866 178599 523922 178608
rect 523776 171080 523828 171086
rect 523776 171022 523828 171028
rect 60096 165572 60148 165578
rect 60096 165514 60148 165520
rect 523682 165336 523738 165345
rect 523682 165271 523738 165280
rect 523696 135250 523724 165271
rect 523880 158710 523908 178599
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 523868 158704 523920 158710
rect 523868 158646 523920 158652
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 523774 152008 523830 152017
rect 523774 151943 523830 151952
rect 523684 135244 523736 135250
rect 523684 135186 523736 135192
rect 60094 130520 60150 130529
rect 60094 130455 60150 130464
rect 60004 122800 60056 122806
rect 60004 122742 60056 122748
rect 59358 116240 59414 116249
rect 59358 116175 59414 116184
rect 59372 116006 59400 116175
rect 59360 116000 59412 116006
rect 59360 115942 59412 115948
rect 59358 101960 59414 101969
rect 59358 101895 59414 101904
rect 59372 100774 59400 101895
rect 59360 100768 59412 100774
rect 59360 100710 59412 100716
rect 3698 93256 3754 93265
rect 3698 93191 3754 93200
rect 60002 87680 60058 87689
rect 60002 87615 60058 87624
rect 59358 73400 59414 73409
rect 59358 73335 59414 73344
rect 59372 73234 59400 73335
rect 59360 73228 59412 73234
rect 59360 73170 59412 73176
rect 59358 59120 59414 59129
rect 59358 59055 59414 59064
rect 59372 58002 59400 59055
rect 59360 57996 59412 58002
rect 59360 57938 59412 57944
rect 3606 50144 3662 50153
rect 3606 50079 3662 50088
rect 60016 35902 60044 87615
rect 60108 80034 60136 130455
rect 523682 125352 523738 125361
rect 523682 125287 523738 125296
rect 523696 88330 523724 125287
rect 523788 124166 523816 151943
rect 523866 138680 523922 138689
rect 523866 138615 523922 138624
rect 523776 124160 523828 124166
rect 523776 124102 523828 124108
rect 523774 112024 523830 112033
rect 523774 111959 523830 111968
rect 523684 88324 523736 88330
rect 523684 88266 523736 88272
rect 523682 85368 523738 85377
rect 523682 85303 523738 85312
rect 60096 80028 60148 80034
rect 60096 79970 60148 79976
rect 62132 52006 62606 52034
rect 63512 52006 63710 52034
rect 60004 35896 60056 35902
rect 60004 35838 60056 35844
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 62132 3466 62160 52006
rect 63512 3534 63540 52006
rect 64892 48754 64920 52020
rect 66088 48822 66116 52020
rect 67284 49094 67312 52020
rect 68494 52006 68968 52034
rect 69690 52006 70348 52034
rect 67272 49088 67324 49094
rect 67272 49030 67324 49036
rect 66076 48816 66128 48822
rect 66076 48758 66128 48764
rect 66904 48816 66956 48822
rect 66904 48758 66956 48764
rect 64880 48748 64932 48754
rect 64880 48690 64932 48696
rect 66168 48748 66220 48754
rect 66168 48690 66220 48696
rect 66180 4894 66208 48690
rect 66916 15910 66944 48758
rect 66904 15904 66956 15910
rect 66904 15846 66956 15852
rect 66168 4888 66220 4894
rect 66168 4830 66220 4836
rect 68940 4826 68968 52006
rect 70320 37942 70348 52006
rect 70872 48822 70900 52020
rect 72068 48822 72096 52020
rect 73264 48822 73292 52020
rect 74460 49162 74488 52020
rect 75670 52006 75868 52034
rect 74448 49156 74500 49162
rect 74448 49098 74500 49104
rect 70860 48816 70912 48822
rect 70860 48758 70912 48764
rect 71688 48816 71740 48822
rect 71688 48758 71740 48764
rect 72056 48816 72108 48822
rect 72056 48758 72108 48764
rect 73068 48816 73120 48822
rect 73068 48758 73120 48764
rect 73252 48816 73304 48822
rect 73252 48758 73304 48764
rect 74448 48816 74500 48822
rect 74448 48758 74500 48764
rect 70308 37936 70360 37942
rect 70308 37878 70360 37884
rect 68928 4820 68980 4826
rect 68928 4762 68980 4768
rect 71700 3942 71728 48758
rect 73080 18630 73108 48758
rect 74460 40730 74488 48758
rect 74448 40724 74500 40730
rect 74448 40666 74500 40672
rect 75840 19990 75868 52006
rect 76852 47666 76880 52020
rect 78062 52006 78628 52034
rect 79258 52006 80008 52034
rect 76840 47660 76892 47666
rect 76840 47602 76892 47608
rect 75828 19984 75880 19990
rect 75828 19926 75880 19932
rect 73068 18624 73120 18630
rect 73068 18566 73120 18572
rect 71688 3936 71740 3942
rect 71688 3878 71740 3884
rect 78600 3874 78628 52006
rect 79980 21418 80008 52006
rect 80440 48822 80468 52020
rect 81636 49230 81664 52020
rect 81624 49224 81676 49230
rect 81624 49166 81676 49172
rect 80428 48816 80480 48822
rect 80428 48758 80480 48764
rect 81348 48816 81400 48822
rect 81348 48758 81400 48764
rect 81360 42090 81388 48758
rect 82832 48686 82860 52020
rect 84042 52006 84148 52034
rect 85238 52006 85528 52034
rect 86434 52006 86908 52034
rect 87630 52006 88288 52034
rect 82820 48680 82872 48686
rect 82820 48622 82872 48628
rect 84016 48680 84068 48686
rect 84016 48622 84068 48628
rect 81348 42084 81400 42090
rect 81348 42026 81400 42032
rect 84028 22778 84056 48622
rect 84016 22772 84068 22778
rect 84016 22714 84068 22720
rect 79968 21412 80020 21418
rect 79968 21354 80020 21360
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 84120 3806 84148 52006
rect 84108 3800 84160 3806
rect 84108 3742 84160 3748
rect 63500 3528 63552 3534
rect 85500 3505 85528 52006
rect 86880 24138 86908 52006
rect 86868 24132 86920 24138
rect 86868 24074 86920 24080
rect 88260 3534 88288 52006
rect 88720 49366 88748 52020
rect 88708 49360 88760 49366
rect 88708 49302 88760 49308
rect 89916 48822 89944 52020
rect 91112 48822 91140 52020
rect 92322 52006 92428 52034
rect 93518 52006 93808 52034
rect 94714 52006 95188 52034
rect 89904 48816 89956 48822
rect 89904 48758 89956 48764
rect 91008 48816 91060 48822
rect 91008 48758 91060 48764
rect 91100 48816 91152 48822
rect 91100 48758 91152 48764
rect 92296 48816 92348 48822
rect 92296 48758 92348 48764
rect 91020 25566 91048 48758
rect 91008 25560 91060 25566
rect 91008 25502 91060 25508
rect 92308 4010 92336 48758
rect 92296 4004 92348 4010
rect 92296 3946 92348 3952
rect 88248 3528 88300 3534
rect 63500 3470 63552 3476
rect 85486 3496 85542 3505
rect 62120 3460 62172 3466
rect 88248 3470 88300 3476
rect 85486 3431 85542 3440
rect 62120 3402 62172 3408
rect 92400 3369 92428 52006
rect 93780 26926 93808 52006
rect 93768 26920 93820 26926
rect 93768 26862 93820 26868
rect 95160 3466 95188 52006
rect 95896 49026 95924 52020
rect 95884 49020 95936 49026
rect 95884 48962 95936 48968
rect 97092 48822 97120 52020
rect 98288 48822 98316 52020
rect 99484 48822 99512 52020
rect 100588 52006 100694 52034
rect 101890 52006 102088 52034
rect 97080 48816 97132 48822
rect 97080 48758 97132 48764
rect 97908 48816 97960 48822
rect 97908 48758 97960 48764
rect 98276 48816 98328 48822
rect 98276 48758 98328 48764
rect 99288 48816 99340 48822
rect 99288 48758 99340 48764
rect 99472 48816 99524 48822
rect 99472 48758 99524 48764
rect 97920 28286 97948 48758
rect 97908 28280 97960 28286
rect 97908 28222 97960 28228
rect 95148 3460 95200 3466
rect 95148 3402 95200 3408
rect 92386 3360 92442 3369
rect 92386 3295 92442 3304
rect 99300 3126 99328 48758
rect 100588 6186 100616 52006
rect 100668 48816 100720 48822
rect 100668 48758 100720 48764
rect 100576 6180 100628 6186
rect 100576 6122 100628 6128
rect 100680 3194 100708 48758
rect 102060 29646 102088 52006
rect 103072 49298 103100 52020
rect 104282 52006 104848 52034
rect 103060 49292 103112 49298
rect 103060 49234 103112 49240
rect 102048 29640 102100 29646
rect 102048 29582 102100 29588
rect 104820 7682 104848 52006
rect 105464 48822 105492 52020
rect 106660 48822 106688 52020
rect 107856 48822 107884 52020
rect 109052 48822 109080 52020
rect 110248 49434 110276 52020
rect 111458 52006 111748 52034
rect 110236 49428 110288 49434
rect 110236 49370 110288 49376
rect 105452 48816 105504 48822
rect 105452 48758 105504 48764
rect 106188 48816 106240 48822
rect 106188 48758 106240 48764
rect 106648 48816 106700 48822
rect 106648 48758 106700 48764
rect 107568 48816 107620 48822
rect 107568 48758 107620 48764
rect 107844 48816 107896 48822
rect 107844 48758 107896 48764
rect 108948 48816 109000 48822
rect 108948 48758 109000 48764
rect 109040 48816 109092 48822
rect 109040 48758 109092 48764
rect 110328 48816 110380 48822
rect 110328 48758 110380 48764
rect 106200 31074 106228 48758
rect 106188 31068 106240 31074
rect 106188 31010 106240 31016
rect 104808 7676 104860 7682
rect 104808 7618 104860 7624
rect 107580 3262 107608 48758
rect 108960 8974 108988 48758
rect 110340 32434 110368 48758
rect 110328 32428 110380 32434
rect 110328 32370 110380 32376
rect 111720 10334 111748 52006
rect 112640 46306 112668 52020
rect 113744 48822 113772 52020
rect 114940 48822 114968 52020
rect 116136 48822 116164 52020
rect 117332 48822 117360 52020
rect 113732 48816 113784 48822
rect 113732 48758 113784 48764
rect 114468 48816 114520 48822
rect 114468 48758 114520 48764
rect 114928 48816 114980 48822
rect 114928 48758 114980 48764
rect 115848 48816 115900 48822
rect 115848 48758 115900 48764
rect 116124 48816 116176 48822
rect 116124 48758 116176 48764
rect 117228 48816 117280 48822
rect 117228 48758 117280 48764
rect 117320 48816 117372 48822
rect 117320 48758 117372 48764
rect 112628 46300 112680 46306
rect 112628 46242 112680 46248
rect 111708 10328 111760 10334
rect 111708 10270 111760 10276
rect 108948 8968 109000 8974
rect 108948 8910 109000 8916
rect 114480 3738 114508 48758
rect 115860 11762 115888 48758
rect 117240 33794 117268 48758
rect 117228 33788 117280 33794
rect 117228 33730 117280 33736
rect 118528 13122 118556 52020
rect 119738 52006 120028 52034
rect 120934 52006 121408 52034
rect 122130 52006 122788 52034
rect 118608 48816 118660 48822
rect 118608 48758 118660 48764
rect 118516 13116 118568 13122
rect 118516 13058 118568 13064
rect 115848 11756 115900 11762
rect 115848 11698 115900 11704
rect 114468 3732 114520 3738
rect 114468 3674 114520 3680
rect 118620 3330 118648 48758
rect 120000 35222 120028 52006
rect 119988 35216 120040 35222
rect 119988 35158 120040 35164
rect 121380 3670 121408 52006
rect 122760 14482 122788 52006
rect 123312 48822 123340 52020
rect 124508 48822 124536 52020
rect 123300 48816 123352 48822
rect 123300 48758 123352 48764
rect 124128 48816 124180 48822
rect 124128 48758 124180 48764
rect 124496 48816 124548 48822
rect 124496 48758 124548 48764
rect 125508 48816 125560 48822
rect 125508 48758 125560 48764
rect 124140 36582 124168 48758
rect 124128 36576 124180 36582
rect 124128 36518 124180 36524
rect 122748 14476 122800 14482
rect 122748 14418 122800 14424
rect 121368 3664 121420 3670
rect 121368 3606 121420 3612
rect 125520 3398 125548 48758
rect 125704 48686 125732 52020
rect 126808 52006 126914 52034
rect 128110 52006 128308 52034
rect 129306 52006 129688 52034
rect 130502 52006 131068 52034
rect 125692 48680 125744 48686
rect 125692 48622 125744 48628
rect 126808 39370 126836 52006
rect 126888 48680 126940 48686
rect 126888 48622 126940 48628
rect 126796 39364 126848 39370
rect 126796 39306 126848 39312
rect 126900 15978 126928 48622
rect 126888 15972 126940 15978
rect 126888 15914 126940 15920
rect 126980 15904 127032 15910
rect 126980 15846 127032 15852
rect 126612 4888 126664 4894
rect 126612 4830 126664 4836
rect 125508 3392 125560 3398
rect 125508 3334 125560 3340
rect 118608 3324 118660 3330
rect 118608 3266 118660 3272
rect 107568 3256 107620 3262
rect 107568 3198 107620 3204
rect 100668 3188 100720 3194
rect 100668 3130 100720 3136
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 126624 480 126652 4830
rect 126992 3482 127020 15846
rect 128280 3602 128308 52006
rect 128452 49088 128504 49094
rect 128452 49030 128504 49036
rect 128268 3596 128320 3602
rect 128268 3538 128320 3544
rect 128464 3482 128492 49030
rect 129660 17270 129688 52006
rect 131040 44878 131068 52006
rect 131684 49094 131712 52020
rect 131672 49088 131724 49094
rect 131672 49030 131724 49036
rect 132880 48822 132908 52020
rect 134076 48822 134104 52020
rect 132868 48816 132920 48822
rect 132868 48758 132920 48764
rect 133788 48816 133840 48822
rect 133788 48758 133840 48764
rect 134064 48816 134116 48822
rect 134064 48758 134116 48764
rect 135168 48816 135220 48822
rect 135168 48758 135220 48764
rect 131028 44872 131080 44878
rect 131028 44814 131080 44820
rect 131120 37936 131172 37942
rect 131120 37878 131172 37884
rect 129648 17264 129700 17270
rect 129648 17206 129700 17212
rect 130200 4820 130252 4826
rect 130200 4762 130252 4768
rect 126992 3454 127848 3482
rect 128464 3454 129044 3482
rect 127820 480 127848 3454
rect 129016 480 129044 3454
rect 130212 480 130240 4762
rect 131132 3482 131160 37878
rect 132592 18624 132644 18630
rect 132592 18566 132644 18572
rect 132604 4078 132632 18566
rect 133800 4962 133828 48758
rect 133880 40724 133932 40730
rect 133880 40666 133932 40672
rect 133788 4956 133840 4962
rect 133788 4898 133840 4904
rect 132592 4072 132644 4078
rect 132592 4014 132644 4020
rect 133788 4072 133840 4078
rect 133788 4014 133840 4020
rect 132500 3936 132552 3942
rect 132500 3878 132552 3884
rect 132512 3754 132540 3878
rect 132512 3726 132632 3754
rect 131132 3454 131436 3482
rect 131408 480 131436 3454
rect 132604 480 132632 3726
rect 133800 480 133828 4014
rect 133892 3346 133920 40666
rect 135180 37942 135208 48758
rect 135272 48550 135300 52020
rect 136482 52006 136588 52034
rect 137678 52006 137968 52034
rect 135444 49156 135496 49162
rect 135444 49098 135496 49104
rect 135260 48544 135312 48550
rect 135260 48486 135312 48492
rect 135168 37936 135220 37942
rect 135168 37878 135220 37884
rect 135456 3346 135484 49098
rect 136456 48544 136508 48550
rect 136456 48486 136508 48492
rect 136468 3942 136496 48486
rect 136560 47598 136588 52006
rect 136548 47592 136600 47598
rect 136548 47534 136600 47540
rect 136640 19984 136692 19990
rect 136640 19926 136692 19932
rect 136456 3936 136508 3942
rect 136456 3878 136508 3884
rect 136652 3346 136680 19926
rect 137940 7614 137968 52006
rect 138860 49162 138888 52020
rect 139978 52006 140728 52034
rect 138848 49156 138900 49162
rect 138848 49098 138900 49104
rect 138020 47660 138072 47666
rect 138020 47602 138072 47608
rect 137928 7608 137980 7614
rect 137928 7550 137980 7556
rect 138032 3346 138060 47602
rect 140700 18630 140728 52006
rect 141160 48822 141188 52020
rect 142252 49224 142304 49230
rect 142252 49166 142304 49172
rect 141148 48816 141200 48822
rect 141148 48758 141200 48764
rect 142068 48816 142120 48822
rect 142068 48758 142120 48764
rect 140780 42084 140832 42090
rect 140780 42026 140832 42032
rect 140688 18624 140740 18630
rect 140688 18566 140740 18572
rect 140792 3874 140820 42026
rect 142080 40798 142108 48758
rect 142068 40792 142120 40798
rect 142068 40734 142120 40740
rect 140872 21412 140924 21418
rect 140872 21354 140924 21360
rect 139676 3868 139728 3874
rect 139676 3810 139728 3816
rect 140780 3868 140832 3874
rect 140780 3810 140832 3816
rect 133892 3318 134932 3346
rect 135456 3318 136128 3346
rect 136652 3318 137324 3346
rect 138032 3318 138520 3346
rect 134904 480 134932 3318
rect 136100 480 136128 3318
rect 137296 480 137324 3318
rect 138492 480 138520 3318
rect 139688 480 139716 3810
rect 140884 480 140912 21354
rect 142068 3868 142120 3874
rect 142068 3810 142120 3816
rect 142080 480 142108 3810
rect 142264 3346 142292 49166
rect 142356 48822 142384 52020
rect 142344 48816 142396 48822
rect 142344 48758 142396 48764
rect 143448 48816 143500 48822
rect 143448 48758 143500 48764
rect 143460 4146 143488 48758
rect 143552 48550 143580 52020
rect 143540 48544 143592 48550
rect 143540 48486 143592 48492
rect 144748 42090 144776 52020
rect 145944 49230 145972 52020
rect 147154 52006 147628 52034
rect 148350 52006 149008 52034
rect 145932 49224 145984 49230
rect 145932 49166 145984 49172
rect 144828 48544 144880 48550
rect 144828 48486 144880 48492
rect 144736 42084 144788 42090
rect 144736 42026 144788 42032
rect 143540 22772 143592 22778
rect 143540 22714 143592 22720
rect 143448 4140 143500 4146
rect 143448 4082 143500 4088
rect 143552 3346 143580 22714
rect 144840 19990 144868 48486
rect 147600 21418 147628 52006
rect 148980 43450 149008 52006
rect 149532 48822 149560 52020
rect 150624 49360 150676 49366
rect 150624 49302 150676 49308
rect 149520 48816 149572 48822
rect 149520 48758 149572 48764
rect 150348 48816 150400 48822
rect 150348 48758 150400 48764
rect 148968 43444 149020 43450
rect 148968 43386 149020 43392
rect 147680 24132 147732 24138
rect 147680 24074 147732 24080
rect 147588 21412 147640 21418
rect 147588 21354 147640 21360
rect 144828 19984 144880 19990
rect 144828 19926 144880 19932
rect 145656 3800 145708 3806
rect 145656 3742 145708 3748
rect 142264 3318 143304 3346
rect 143552 3318 144500 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3742
rect 146850 3496 146906 3505
rect 146850 3431 146906 3440
rect 146864 480 146892 3431
rect 147692 3346 147720 24074
rect 150360 4078 150388 48758
rect 150532 25560 150584 25566
rect 150532 25502 150584 25508
rect 150348 4072 150400 4078
rect 150348 4014 150400 4020
rect 150544 3806 150572 25502
rect 150532 3800 150584 3806
rect 150532 3742 150584 3748
rect 149244 3528 149296 3534
rect 150636 3482 150664 49302
rect 150728 48822 150756 52020
rect 151924 48822 151952 52020
rect 150716 48816 150768 48822
rect 150716 48758 150768 48764
rect 151728 48816 151780 48822
rect 151728 48758 151780 48764
rect 151912 48816 151964 48822
rect 151912 48758 151964 48764
rect 153016 48816 153068 48822
rect 153016 48758 153068 48764
rect 151740 22778 151768 48758
rect 153028 29714 153056 48758
rect 153016 29708 153068 29714
rect 153016 29650 153068 29656
rect 151728 22772 151780 22778
rect 151728 22714 151780 22720
rect 152740 4004 152792 4010
rect 152740 3946 152792 3952
rect 151544 3800 151596 3806
rect 151544 3742 151596 3748
rect 149244 3470 149296 3476
rect 147692 3318 148088 3346
rect 148060 480 148088 3318
rect 149256 480 149284 3470
rect 150452 3454 150664 3482
rect 150452 480 150480 3454
rect 151556 480 151584 3742
rect 152752 480 152780 3946
rect 153120 3806 153148 52020
rect 154330 52006 154528 52034
rect 155526 52006 155908 52034
rect 156722 52006 157288 52034
rect 154500 24138 154528 52006
rect 155880 31142 155908 52006
rect 155868 31136 155920 31142
rect 155868 31078 155920 31084
rect 154580 26920 154632 26926
rect 154580 26862 154632 26868
rect 154488 24132 154540 24138
rect 154488 24074 154540 24080
rect 153108 3800 153160 3806
rect 153108 3742 153160 3748
rect 153934 3360 153990 3369
rect 154592 3346 154620 26862
rect 157260 3874 157288 52006
rect 157432 49020 157484 49026
rect 157432 48962 157484 48968
rect 157248 3868 157300 3874
rect 157248 3810 157300 3816
rect 156328 3460 156380 3466
rect 156328 3402 156380 3408
rect 154592 3318 155172 3346
rect 153934 3295 153990 3304
rect 153948 480 153976 3295
rect 155144 480 155172 3318
rect 156340 480 156368 3402
rect 157444 1578 157472 48962
rect 157904 48822 157932 52020
rect 159100 48822 159128 52020
rect 160296 48822 160324 52020
rect 161492 48822 161520 52020
rect 157892 48816 157944 48822
rect 157892 48758 157944 48764
rect 158628 48816 158680 48822
rect 158628 48758 158680 48764
rect 159088 48816 159140 48822
rect 159088 48758 159140 48764
rect 160008 48816 160060 48822
rect 160008 48758 160060 48764
rect 160284 48816 160336 48822
rect 160284 48758 160336 48764
rect 161388 48816 161440 48822
rect 161388 48758 161440 48764
rect 161480 48816 161532 48822
rect 161480 48758 161532 48764
rect 158640 25566 158668 48758
rect 160020 32502 160048 48758
rect 160008 32496 160060 32502
rect 160008 32438 160060 32444
rect 158812 28280 158864 28286
rect 158812 28222 158864 28228
rect 158628 25560 158680 25566
rect 158628 25502 158680 25508
rect 158824 1578 158852 28222
rect 161400 4010 161428 48758
rect 162688 46238 162716 52020
rect 163898 52006 164188 52034
rect 165002 52006 165568 52034
rect 162768 48816 162820 48822
rect 162768 48758 162820 48764
rect 162676 46232 162728 46238
rect 162676 46174 162728 46180
rect 162780 6322 162808 48758
rect 162860 29640 162912 29646
rect 162860 29582 162912 29588
rect 162768 6316 162820 6322
rect 162768 6258 162820 6264
rect 162308 6180 162360 6186
rect 162308 6122 162360 6128
rect 161388 4004 161440 4010
rect 161388 3946 161440 3952
rect 161112 3188 161164 3194
rect 161112 3130 161164 3136
rect 159916 3120 159968 3126
rect 159916 3062 159968 3068
rect 157444 1550 157564 1578
rect 157536 480 157564 1550
rect 158732 1550 158852 1578
rect 158732 480 158760 1550
rect 159928 480 159956 3062
rect 161124 480 161152 3130
rect 162320 480 162348 6122
rect 162872 3482 162900 29582
rect 162872 3454 163544 3482
rect 164160 3466 164188 52006
rect 164332 49292 164384 49298
rect 164332 49234 164384 49240
rect 164344 3482 164372 49234
rect 165540 26926 165568 52006
rect 166184 48550 166212 52020
rect 167380 49502 167408 52020
rect 167368 49496 167420 49502
rect 167368 49438 167420 49444
rect 168576 48822 168604 52020
rect 169772 48822 169800 52020
rect 170982 52006 171088 52034
rect 172178 52006 172468 52034
rect 173374 52006 173848 52034
rect 168564 48816 168616 48822
rect 168564 48758 168616 48764
rect 169668 48816 169720 48822
rect 169668 48758 169720 48764
rect 169760 48816 169812 48822
rect 169760 48758 169812 48764
rect 170956 48816 171008 48822
rect 170956 48758 171008 48764
rect 166172 48544 166224 48550
rect 166172 48486 166224 48492
rect 167644 48544 167696 48550
rect 167644 48486 167696 48492
rect 167656 33862 167684 48486
rect 167644 33856 167696 33862
rect 167644 33798 167696 33804
rect 167092 31068 167144 31074
rect 167092 31010 167144 31016
rect 165528 26920 165580 26926
rect 165528 26862 165580 26868
rect 165896 7676 165948 7682
rect 165896 7618 165948 7624
rect 163516 480 163544 3454
rect 164148 3460 164200 3466
rect 164344 3454 164740 3482
rect 164148 3402 164200 3408
rect 164712 480 164740 3454
rect 165908 480 165936 7618
rect 167104 480 167132 31010
rect 169392 8968 169444 8974
rect 169392 8910 169444 8916
rect 168196 3256 168248 3262
rect 168196 3198 168248 3204
rect 168208 480 168236 3198
rect 169404 480 169432 8910
rect 169680 7682 169708 48758
rect 170968 35290 170996 48758
rect 170956 35284 171008 35290
rect 170956 35226 171008 35232
rect 169760 32428 169812 32434
rect 169760 32370 169812 32376
rect 169668 7676 169720 7682
rect 169668 7618 169720 7624
rect 169772 3482 169800 32370
rect 171060 3534 171088 52006
rect 171232 49428 171284 49434
rect 171232 49370 171284 49376
rect 171048 3528 171100 3534
rect 169772 3454 170628 3482
rect 171048 3470 171100 3476
rect 170600 480 170628 3454
rect 171244 3346 171272 49370
rect 172440 8974 172468 52006
rect 172520 10328 172572 10334
rect 172520 10270 172572 10276
rect 172428 8968 172480 8974
rect 172428 8910 172480 8916
rect 172532 3346 172560 10270
rect 173820 4894 173848 52006
rect 174556 49298 174584 52020
rect 174544 49292 174596 49298
rect 174544 49234 174596 49240
rect 175752 48822 175780 52020
rect 176948 48822 176976 52020
rect 178144 48822 178172 52020
rect 179248 52006 179354 52034
rect 180550 52006 180748 52034
rect 175740 48816 175792 48822
rect 175740 48758 175792 48764
rect 176568 48816 176620 48822
rect 176568 48758 176620 48764
rect 176936 48816 176988 48822
rect 176936 48758 176988 48764
rect 177948 48816 178000 48822
rect 177948 48758 178000 48764
rect 178132 48816 178184 48822
rect 178132 48758 178184 48764
rect 173900 46300 173952 46306
rect 173900 46242 173952 46248
rect 173808 4888 173860 4894
rect 173808 4830 173860 4836
rect 173912 3346 173940 46242
rect 175372 11756 175424 11762
rect 175372 11698 175424 11704
rect 175280 3732 175332 3738
rect 175280 3674 175332 3680
rect 171244 3318 171824 3346
rect 172532 3318 173020 3346
rect 173912 3318 174216 3346
rect 171796 480 171824 3318
rect 172992 480 173020 3318
rect 174188 480 174216 3318
rect 175292 3210 175320 3674
rect 175384 3330 175412 11698
rect 176580 10402 176608 48758
rect 177960 36718 177988 48758
rect 177948 36712 178000 36718
rect 177948 36654 178000 36660
rect 176660 33788 176712 33794
rect 176660 33730 176712 33736
rect 176568 10396 176620 10402
rect 176568 10338 176620 10344
rect 176672 3346 176700 33730
rect 179248 11762 179276 52006
rect 179328 48816 179380 48822
rect 179328 48758 179380 48764
rect 179236 11756 179288 11762
rect 179236 11698 179288 11704
rect 175372 3324 175424 3330
rect 175372 3266 175424 3272
rect 176568 3324 176620 3330
rect 176672 3318 177804 3346
rect 176568 3266 176620 3272
rect 175292 3182 175412 3210
rect 175384 480 175412 3182
rect 176580 480 176608 3266
rect 177776 480 177804 3318
rect 178960 3256 179012 3262
rect 178960 3198 179012 3204
rect 178972 480 179000 3198
rect 179340 3126 179368 48758
rect 180720 39438 180748 52006
rect 181732 49026 181760 52020
rect 182942 52006 183508 52034
rect 184138 52006 184888 52034
rect 181720 49020 181772 49026
rect 181720 48962 181772 48968
rect 180708 39432 180760 39438
rect 180708 39374 180760 39380
rect 180800 35216 180852 35222
rect 180800 35158 180852 35164
rect 179420 13116 179472 13122
rect 179420 13058 179472 13064
rect 179432 3346 179460 13058
rect 180812 3346 180840 35158
rect 183480 13122 183508 52006
rect 184860 45014 184888 52006
rect 185320 48822 185348 52020
rect 186516 48822 186544 52020
rect 187712 48822 187740 52020
rect 188908 49366 188936 52020
rect 190118 52006 190408 52034
rect 191222 52006 191788 52034
rect 192418 52006 193168 52034
rect 188896 49360 188948 49366
rect 188896 49302 188948 49308
rect 185308 48816 185360 48822
rect 185308 48758 185360 48764
rect 186228 48816 186280 48822
rect 186228 48758 186280 48764
rect 186504 48816 186556 48822
rect 186504 48758 186556 48764
rect 187608 48816 187660 48822
rect 187608 48758 187660 48764
rect 187700 48816 187752 48822
rect 187700 48758 187752 48764
rect 188988 48816 189040 48822
rect 188988 48758 189040 48764
rect 184848 45008 184900 45014
rect 184848 44950 184900 44956
rect 183560 36576 183612 36582
rect 183560 36518 183612 36524
rect 183468 13116 183520 13122
rect 183468 13058 183520 13064
rect 182548 3664 182600 3670
rect 182548 3606 182600 3612
rect 179432 3318 180196 3346
rect 180812 3318 181392 3346
rect 179328 3120 179380 3126
rect 179328 3062 179380 3068
rect 180168 480 180196 3318
rect 181364 480 181392 3318
rect 182560 480 182588 3606
rect 183572 3602 183600 36518
rect 183652 14476 183704 14482
rect 183652 14418 183704 14424
rect 183560 3596 183612 3602
rect 183560 3538 183612 3544
rect 183664 3482 183692 14418
rect 184848 3596 184900 3602
rect 184848 3538 184900 3544
rect 183664 3454 183784 3482
rect 183756 480 183784 3454
rect 184860 480 184888 3538
rect 186044 3392 186096 3398
rect 186044 3334 186096 3340
rect 186056 480 186084 3334
rect 186240 3058 186268 48758
rect 186320 15972 186372 15978
rect 186320 15914 186372 15920
rect 186332 3346 186360 15914
rect 187620 14482 187648 48758
rect 187700 39364 187752 39370
rect 187700 39306 187752 39312
rect 187608 14476 187660 14482
rect 187608 14418 187660 14424
rect 187712 3346 187740 39306
rect 189000 38010 189028 48758
rect 188988 38004 189040 38010
rect 188988 37946 189040 37952
rect 190380 4826 190408 52006
rect 191760 29646 191788 52006
rect 191840 44872 191892 44878
rect 191840 44814 191892 44820
rect 191748 29640 191800 29646
rect 191748 29582 191800 29588
rect 190460 17264 190512 17270
rect 190460 17206 190512 17212
rect 190368 4820 190420 4826
rect 190368 4762 190420 4768
rect 189632 3664 189684 3670
rect 189632 3606 189684 3612
rect 186332 3318 187280 3346
rect 187712 3318 188476 3346
rect 186228 3052 186280 3058
rect 186228 2994 186280 3000
rect 187252 480 187280 3318
rect 188448 480 188476 3318
rect 189644 480 189672 3606
rect 190472 3346 190500 17206
rect 191852 3346 191880 44814
rect 190472 3318 190868 3346
rect 191852 3318 192064 3346
rect 190840 480 190868 3318
rect 192036 480 192064 3318
rect 193140 3194 193168 52006
rect 193404 49088 193456 49094
rect 193404 49030 193456 49036
rect 193416 3346 193444 49030
rect 193600 48822 193628 52020
rect 193588 48816 193640 48822
rect 193588 48758 193640 48764
rect 194508 48816 194560 48822
rect 194508 48758 194560 48764
rect 194520 15910 194548 48758
rect 194796 47666 194824 52020
rect 195992 48686 196020 52020
rect 195980 48680 196032 48686
rect 195980 48622 196032 48628
rect 194784 47660 194836 47666
rect 194784 47602 194836 47608
rect 194600 37936 194652 37942
rect 194600 37878 194652 37884
rect 194508 15904 194560 15910
rect 194508 15846 194560 15852
rect 194416 4956 194468 4962
rect 194416 4898 194468 4904
rect 193232 3318 193444 3346
rect 193128 3188 193180 3194
rect 193128 3130 193180 3136
rect 193232 480 193260 3318
rect 194428 480 194456 4898
rect 194612 3346 194640 37878
rect 197188 17270 197216 52020
rect 198398 52006 198688 52034
rect 199594 52006 200068 52034
rect 200790 52006 201448 52034
rect 197268 48680 197320 48686
rect 197268 48622 197320 48628
rect 197176 17264 197228 17270
rect 197176 17206 197228 17212
rect 196808 3936 196860 3942
rect 196808 3878 196860 3884
rect 194612 3318 195652 3346
rect 195624 480 195652 3318
rect 196820 480 196848 3878
rect 197280 3262 197308 48622
rect 197360 47592 197412 47598
rect 197360 47534 197412 47540
rect 197372 3346 197400 47534
rect 198660 40730 198688 52006
rect 198648 40724 198700 40730
rect 198648 40666 198700 40672
rect 199200 7608 199252 7614
rect 199200 7550 199252 7556
rect 197372 3318 198044 3346
rect 197268 3256 197320 3262
rect 197268 3198 197320 3204
rect 198016 480 198044 3318
rect 199212 480 199240 7550
rect 200040 3942 200068 52006
rect 200212 49156 200264 49162
rect 200212 49098 200264 49104
rect 200028 3936 200080 3942
rect 200028 3878 200080 3884
rect 200224 3346 200252 49098
rect 201420 28286 201448 52006
rect 201972 48822 202000 52020
rect 203168 48822 203196 52020
rect 204364 48822 204392 52020
rect 205468 52006 205574 52034
rect 206770 52006 206968 52034
rect 207966 52006 208348 52034
rect 209162 52006 209728 52034
rect 201960 48816 202012 48822
rect 201960 48758 202012 48764
rect 202788 48816 202840 48822
rect 202788 48758 202840 48764
rect 203156 48816 203208 48822
rect 203156 48758 203208 48764
rect 204168 48816 204220 48822
rect 204168 48758 204220 48764
rect 204352 48816 204404 48822
rect 204352 48758 204404 48764
rect 202800 42158 202828 48758
rect 202788 42152 202840 42158
rect 202788 42094 202840 42100
rect 201500 40792 201552 40798
rect 201500 40734 201552 40740
rect 201408 28280 201460 28286
rect 201408 28222 201460 28228
rect 201512 3602 201540 40734
rect 201592 18624 201644 18630
rect 201592 18566 201644 18572
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 201604 3482 201632 18566
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 202696 3596 202748 3602
rect 202696 3538 202748 3544
rect 201512 3454 201632 3482
rect 200224 3318 200436 3346
rect 200408 480 200436 3318
rect 201512 480 201540 3454
rect 202708 480 202736 3538
rect 203904 480 203932 4082
rect 204180 3330 204208 48758
rect 205468 31074 205496 52006
rect 205548 48816 205600 48822
rect 205548 48758 205600 48764
rect 205456 31068 205508 31074
rect 205456 31010 205508 31016
rect 205560 19990 205588 48758
rect 205640 42084 205692 42090
rect 205640 42026 205692 42032
rect 204260 19984 204312 19990
rect 204260 19926 204312 19932
rect 205548 19984 205600 19990
rect 205548 19926 205600 19932
rect 204272 3346 204300 19926
rect 205652 3346 205680 42026
rect 206940 3738 206968 52006
rect 207112 49224 207164 49230
rect 207112 49166 207164 49172
rect 206928 3732 206980 3738
rect 206928 3674 206980 3680
rect 207124 3346 207152 49166
rect 208320 18630 208348 52006
rect 208400 21412 208452 21418
rect 208400 21354 208452 21360
rect 208308 18624 208360 18630
rect 208308 18566 208360 18572
rect 208412 3346 208440 21354
rect 209700 6186 209728 52006
rect 210344 49230 210372 52020
rect 210332 49224 210384 49230
rect 210332 49166 210384 49172
rect 211540 48822 211568 52020
rect 212736 48822 212764 52020
rect 213932 48822 213960 52020
rect 211528 48816 211580 48822
rect 211528 48758 211580 48764
rect 212448 48816 212500 48822
rect 212448 48758 212500 48764
rect 212724 48816 212776 48822
rect 212724 48758 212776 48764
rect 213828 48816 213880 48822
rect 213828 48758 213880 48764
rect 213920 48816 213972 48822
rect 213920 48758 213972 48764
rect 209872 43444 209924 43450
rect 209872 43386 209924 43392
rect 209688 6180 209740 6186
rect 209688 6122 209740 6128
rect 204168 3324 204220 3330
rect 204272 3318 205128 3346
rect 205652 3318 206324 3346
rect 207124 3318 207520 3346
rect 208412 3318 208716 3346
rect 204168 3266 204220 3272
rect 205100 480 205128 3318
rect 206296 480 206324 3318
rect 207492 480 207520 3318
rect 208688 480 208716 3318
rect 209884 480 209912 43386
rect 211160 22772 211212 22778
rect 211160 22714 211212 22720
rect 211068 4072 211120 4078
rect 211068 4014 211120 4020
rect 211080 480 211108 4014
rect 211172 3346 211200 22714
rect 212460 21418 212488 48758
rect 213840 43450 213868 48758
rect 213828 43444 213880 43450
rect 213828 43386 213880 43392
rect 212540 29708 212592 29714
rect 212540 29650 212592 29656
rect 212448 21412 212500 21418
rect 212448 21354 212500 21360
rect 212552 3346 212580 29650
rect 215128 22778 215156 52020
rect 216246 52006 216628 52034
rect 215208 48816 215260 48822
rect 215208 48758 215260 48764
rect 215116 22772 215168 22778
rect 215116 22714 215168 22720
rect 214656 3800 214708 3806
rect 214656 3742 214708 3748
rect 211172 3318 212304 3346
rect 212552 3318 213500 3346
rect 212276 480 212304 3318
rect 213472 480 213500 3318
rect 214668 480 214696 3742
rect 215220 3398 215248 48758
rect 216600 32434 216628 52006
rect 217428 49094 217456 52020
rect 217416 49088 217468 49094
rect 217416 49030 217468 49036
rect 218624 48822 218652 52020
rect 218612 48816 218664 48822
rect 218612 48758 218664 48764
rect 219348 48816 219400 48822
rect 219348 48758 219400 48764
rect 216588 32428 216640 32434
rect 216588 32370 216640 32376
rect 216680 31136 216732 31142
rect 216680 31078 216732 31084
rect 215300 24132 215352 24138
rect 215300 24074 215352 24080
rect 215208 3392 215260 3398
rect 215208 3334 215260 3340
rect 215312 3346 215340 24074
rect 216692 3346 216720 31078
rect 218152 25560 218204 25566
rect 218152 25502 218204 25508
rect 218060 3868 218112 3874
rect 218060 3810 218112 3816
rect 218072 3482 218100 3810
rect 218164 3602 218192 25502
rect 219360 6254 219388 48758
rect 219820 46374 219848 52020
rect 221016 48822 221044 52020
rect 222212 48822 222240 52020
rect 221004 48816 221056 48822
rect 221004 48758 221056 48764
rect 222108 48816 222160 48822
rect 222108 48758 222160 48764
rect 222200 48816 222252 48822
rect 222200 48758 222252 48764
rect 219808 46368 219860 46374
rect 219808 46310 219860 46316
rect 219440 32496 219492 32502
rect 219440 32438 219492 32444
rect 219348 6248 219400 6254
rect 219348 6190 219400 6196
rect 218152 3596 218204 3602
rect 218152 3538 218204 3544
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 218072 3454 218192 3482
rect 215312 3318 215892 3346
rect 216692 3318 217088 3346
rect 215864 480 215892 3318
rect 217060 480 217088 3318
rect 218164 480 218192 3454
rect 219360 480 219388 3538
rect 219452 3346 219480 32438
rect 221740 4004 221792 4010
rect 221740 3946 221792 3952
rect 219452 3318 220584 3346
rect 220556 480 220584 3318
rect 221752 480 221780 3946
rect 222120 3806 222148 48758
rect 223408 33794 223436 52020
rect 224604 49162 224632 52020
rect 225814 52006 226288 52034
rect 227010 52006 227668 52034
rect 224592 49156 224644 49162
rect 224592 49098 224644 49104
rect 223488 48816 223540 48822
rect 223488 48758 223540 48764
rect 223396 33788 223448 33794
rect 223396 33730 223448 33736
rect 223500 7614 223528 48758
rect 223580 46232 223632 46238
rect 223580 46174 223632 46180
rect 223488 7608 223540 7614
rect 223488 7550 223540 7556
rect 222936 6316 222988 6322
rect 222936 6258 222988 6264
rect 222108 3800 222160 3806
rect 222108 3742 222160 3748
rect 222948 480 222976 6258
rect 223592 3346 223620 46174
rect 226260 24138 226288 52006
rect 227640 35358 227668 52006
rect 227904 49496 227956 49502
rect 227904 49438 227956 49444
rect 227628 35352 227680 35358
rect 227628 35294 227680 35300
rect 227812 33856 227864 33862
rect 227812 33798 227864 33804
rect 226340 26920 226392 26926
rect 226340 26862 226392 26868
rect 226248 24132 226300 24138
rect 226248 24074 226300 24080
rect 225328 3460 225380 3466
rect 225328 3402 225380 3408
rect 223592 3318 224172 3346
rect 224144 480 224172 3318
rect 225340 480 225368 3402
rect 226352 3346 226380 26862
rect 227824 3482 227852 33798
rect 227732 3454 227852 3482
rect 226352 3318 226564 3346
rect 226536 480 226564 3318
rect 227732 480 227760 3454
rect 227916 3346 227944 49438
rect 228192 48822 228220 52020
rect 229388 48822 229416 52020
rect 228180 48816 228232 48822
rect 228180 48758 228232 48764
rect 229008 48816 229060 48822
rect 229008 48758 229060 48764
rect 229376 48816 229428 48822
rect 229376 48758 229428 48764
rect 230388 48816 230440 48822
rect 230388 48758 230440 48764
rect 229020 3874 229048 48758
rect 230400 9042 230428 48758
rect 230584 48686 230612 52020
rect 230572 48680 230624 48686
rect 230572 48622 230624 48628
rect 231676 48680 231728 48686
rect 231676 48622 231728 48628
rect 231688 36650 231716 48622
rect 231676 36644 231728 36650
rect 231676 36586 231728 36592
rect 230480 35284 230532 35290
rect 230480 35226 230532 35232
rect 230388 9036 230440 9042
rect 230388 8978 230440 8984
rect 230112 7676 230164 7682
rect 230112 7618 230164 7624
rect 229008 3868 229060 3874
rect 229008 3810 229060 3816
rect 227916 3318 228956 3346
rect 228928 480 228956 3318
rect 230124 480 230152 7618
rect 230492 3482 230520 35226
rect 231780 3670 231808 52020
rect 232990 52006 233188 52034
rect 234186 52006 234568 52034
rect 235382 52006 235948 52034
rect 236578 52006 237328 52034
rect 233160 10334 233188 52006
rect 234540 39370 234568 52006
rect 234528 39364 234580 39370
rect 234528 39306 234580 39312
rect 233148 10328 233200 10334
rect 233148 10270 233200 10276
rect 233700 8968 233752 8974
rect 233700 8910 233752 8916
rect 231768 3664 231820 3670
rect 231768 3606 231820 3612
rect 232504 3528 232556 3534
rect 230492 3454 231348 3482
rect 232504 3470 232556 3476
rect 231320 480 231348 3454
rect 232516 480 232544 3470
rect 233712 480 233740 8910
rect 234804 4888 234856 4894
rect 234804 4830 234856 4836
rect 234816 480 234844 4830
rect 235920 3466 235948 52006
rect 236184 49292 236236 49298
rect 236184 49234 236236 49240
rect 236092 10396 236144 10402
rect 236092 10338 236144 10344
rect 236104 3602 236132 10338
rect 236092 3596 236144 3602
rect 236092 3538 236144 3544
rect 236196 3482 236224 49234
rect 237300 25634 237328 52006
rect 237760 48822 237788 52020
rect 237748 48816 237800 48822
rect 237748 48758 237800 48764
rect 238668 48816 238720 48822
rect 238668 48758 238720 48764
rect 238680 44946 238708 48758
rect 238956 48754 238984 52020
rect 238944 48748 238996 48754
rect 238944 48690 238996 48696
rect 240048 48748 240100 48754
rect 240048 48690 240100 48696
rect 238668 44940 238720 44946
rect 238668 44882 238720 44888
rect 237380 36712 237432 36718
rect 237380 36654 237432 36660
rect 237288 25628 237340 25634
rect 237288 25570 237340 25576
rect 237196 3596 237248 3602
rect 237196 3538 237248 3544
rect 235908 3460 235960 3466
rect 235908 3402 235960 3408
rect 236012 3454 236224 3482
rect 236012 480 236040 3454
rect 237208 480 237236 3538
rect 237392 3482 237420 36654
rect 240060 4146 240088 48690
rect 240152 48346 240180 52020
rect 240140 48340 240192 48346
rect 240140 48282 240192 48288
rect 241348 37942 241376 52020
rect 242466 52006 242848 52034
rect 243662 52006 244228 52034
rect 244858 52006 245608 52034
rect 241428 48340 241480 48346
rect 241428 48282 241480 48288
rect 241336 37936 241388 37942
rect 241336 37878 241388 37884
rect 241440 11762 241468 48282
rect 241520 39432 241572 39438
rect 241520 39374 241572 39380
rect 240140 11756 240192 11762
rect 240140 11698 240192 11704
rect 241428 11756 241480 11762
rect 241428 11698 241480 11704
rect 240048 4140 240100 4146
rect 240048 4082 240100 4088
rect 237392 3454 238432 3482
rect 238404 480 238432 3454
rect 240152 3346 240180 11698
rect 241532 3346 241560 39374
rect 242820 3602 242848 52006
rect 242992 49020 243044 49026
rect 242992 48962 243044 48968
rect 242808 3596 242860 3602
rect 242808 3538 242860 3544
rect 243004 3346 243032 48962
rect 244200 26926 244228 52006
rect 244280 45008 244332 45014
rect 244280 44950 244332 44956
rect 244188 26920 244240 26926
rect 244188 26862 244240 26868
rect 244292 3534 244320 44950
rect 245580 29782 245608 52006
rect 246040 48822 246068 52020
rect 247236 48822 247264 52020
rect 248432 48822 248460 52020
rect 249642 52006 249748 52034
rect 250838 52006 251128 52034
rect 252034 52006 252508 52034
rect 246028 48816 246080 48822
rect 246028 48758 246080 48764
rect 246948 48816 247000 48822
rect 246948 48758 247000 48764
rect 247224 48816 247276 48822
rect 247224 48758 247276 48764
rect 248328 48816 248380 48822
rect 248328 48758 248380 48764
rect 248420 48816 248472 48822
rect 248420 48758 248472 48764
rect 249616 48816 249668 48822
rect 249616 48758 249668 48764
rect 245568 29776 245620 29782
rect 245568 29718 245620 29724
rect 244372 13116 244424 13122
rect 244372 13058 244424 13064
rect 244280 3528 244332 3534
rect 244280 3470 244332 3476
rect 240152 3318 240824 3346
rect 241532 3318 242020 3346
rect 243004 3318 243216 3346
rect 239588 3120 239640 3126
rect 239588 3062 239640 3068
rect 239600 480 239628 3062
rect 240796 480 240824 3318
rect 241992 480 242020 3318
rect 243188 480 243216 3318
rect 244384 480 244412 13058
rect 246960 4010 246988 48758
rect 248340 14482 248368 48758
rect 249628 40798 249656 48758
rect 249616 40792 249668 40798
rect 249616 40734 249668 40740
rect 248420 38004 248472 38010
rect 248420 37946 248472 37952
rect 247040 14476 247092 14482
rect 247040 14418 247092 14424
rect 248328 14476 248380 14482
rect 248328 14418 248380 14424
rect 246948 4004 247000 4010
rect 246948 3946 247000 3952
rect 245568 3528 245620 3534
rect 245568 3470 245620 3476
rect 245580 480 245608 3470
rect 247052 3346 247080 14418
rect 248432 3346 248460 37946
rect 249720 3534 249748 52006
rect 249892 49360 249944 49366
rect 249892 49302 249944 49308
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 249904 3346 249932 49302
rect 251100 13122 251128 52006
rect 252480 28354 252508 52006
rect 253216 49298 253244 52020
rect 253204 49292 253256 49298
rect 253204 49234 253256 49240
rect 254412 48822 254440 52020
rect 255608 48822 255636 52020
rect 256804 48822 256832 52020
rect 257908 52006 258014 52034
rect 259210 52006 259408 52034
rect 254400 48816 254452 48822
rect 254400 48758 254452 48764
rect 255228 48816 255280 48822
rect 255228 48758 255280 48764
rect 255596 48816 255648 48822
rect 255596 48758 255648 48764
rect 256608 48816 256660 48822
rect 256608 48758 256660 48764
rect 256792 48816 256844 48822
rect 256792 48758 256844 48764
rect 252652 29640 252704 29646
rect 252652 29582 252704 29588
rect 252468 28348 252520 28354
rect 252468 28290 252520 28296
rect 251088 13116 251140 13122
rect 251088 13058 251140 13064
rect 251456 4820 251508 4826
rect 251456 4762 251508 4768
rect 247052 3318 248000 3346
rect 248432 3318 249196 3346
rect 249904 3318 250392 3346
rect 246764 3052 246816 3058
rect 246764 2994 246816 3000
rect 246776 480 246804 2994
rect 247972 480 248000 3318
rect 249168 480 249196 3318
rect 250364 480 250392 3318
rect 251468 480 251496 4762
rect 252664 480 252692 29582
rect 253940 15904 253992 15910
rect 253940 15846 253992 15852
rect 253952 3346 253980 15846
rect 255240 4894 255268 48758
rect 255320 47660 255372 47666
rect 255320 47602 255372 47608
rect 255228 4888 255280 4894
rect 255228 4830 255280 4836
rect 255332 3346 255360 47602
rect 256620 42226 256648 48758
rect 256608 42220 256660 42226
rect 256608 42162 256660 42168
rect 257908 15910 257936 52006
rect 257988 48816 258040 48822
rect 257988 48758 258040 48764
rect 257896 15904 257948 15910
rect 257896 15846 257948 15852
rect 258000 4078 258028 48758
rect 259380 31142 259408 52006
rect 260392 49026 260420 52020
rect 261602 52006 262168 52034
rect 260380 49020 260432 49026
rect 260380 48962 260432 48968
rect 259460 40724 259512 40730
rect 259460 40666 259512 40672
rect 259368 31136 259420 31142
rect 259368 31078 259420 31084
rect 258080 17264 258132 17270
rect 258080 17206 258132 17212
rect 257988 4072 258040 4078
rect 257988 4014 258040 4020
rect 258092 3482 258120 17206
rect 259472 3482 259500 40666
rect 262140 17270 262168 52006
rect 262784 48346 262812 52020
rect 263980 48822 264008 52020
rect 265176 48822 265204 52020
rect 266372 48822 266400 52020
rect 267490 52006 267688 52034
rect 268686 52006 269068 52034
rect 269882 52006 270448 52034
rect 263968 48816 264020 48822
rect 263968 48758 264020 48764
rect 264888 48816 264940 48822
rect 264888 48758 264940 48764
rect 265164 48816 265216 48822
rect 265164 48758 265216 48764
rect 266268 48816 266320 48822
rect 266268 48758 266320 48764
rect 266360 48816 266412 48822
rect 266360 48758 266412 48764
rect 267556 48816 267608 48822
rect 267556 48758 267608 48764
rect 262772 48340 262824 48346
rect 262772 48282 262824 48288
rect 263508 48340 263560 48346
rect 263508 48282 263560 48288
rect 263520 43518 263548 48282
rect 263508 43512 263560 43518
rect 263508 43454 263560 43460
rect 262220 42152 262272 42158
rect 262220 42094 262272 42100
rect 262128 17264 262180 17270
rect 262128 17206 262180 17212
rect 262232 3942 262260 42094
rect 262312 28280 262364 28286
rect 262312 28222 262364 28228
rect 261024 3936 261076 3942
rect 261024 3878 261076 3884
rect 262220 3936 262272 3942
rect 262220 3878 262272 3884
rect 258092 3454 258672 3482
rect 259472 3454 259868 3482
rect 253952 3318 255084 3346
rect 255332 3318 256280 3346
rect 253848 3188 253900 3194
rect 253848 3130 253900 3136
rect 253860 480 253888 3130
rect 255056 480 255084 3318
rect 256252 480 256280 3318
rect 257436 3256 257488 3262
rect 257436 3198 257488 3204
rect 257448 480 257476 3198
rect 258644 480 258672 3454
rect 259840 480 259868 3454
rect 261036 480 261064 3878
rect 262324 3482 262352 28222
rect 264900 7682 264928 48758
rect 266280 19990 266308 48758
rect 267568 32502 267596 48758
rect 267556 32496 267608 32502
rect 267556 32438 267608 32444
rect 266360 31068 266412 31074
rect 266360 31010 266412 31016
rect 264980 19984 265032 19990
rect 264980 19926 265032 19932
rect 266268 19984 266320 19990
rect 266268 19926 266320 19932
rect 264888 7676 264940 7682
rect 264888 7618 264940 7624
rect 263416 3936 263468 3942
rect 263416 3878 263468 3884
rect 262232 3454 262352 3482
rect 262232 480 262260 3454
rect 263428 480 263456 3878
rect 264992 3482 265020 19926
rect 266372 3482 266400 31010
rect 267660 25566 267688 52006
rect 267648 25560 267700 25566
rect 267648 25502 267700 25508
rect 269040 18698 269068 52006
rect 270420 33862 270448 52006
rect 270500 49224 270552 49230
rect 270500 49166 270552 49172
rect 270408 33856 270460 33862
rect 270408 33798 270460 33804
rect 269028 18692 269080 18698
rect 269028 18634 269080 18640
rect 269120 18624 269172 18630
rect 269120 18566 269172 18572
rect 268108 3732 268160 3738
rect 268108 3674 268160 3680
rect 264992 3454 265848 3482
rect 266372 3454 267044 3482
rect 264612 3324 264664 3330
rect 264612 3266 264664 3272
rect 264624 480 264652 3266
rect 265820 480 265848 3454
rect 267016 480 267044 3454
rect 268120 480 268148 3674
rect 269132 3482 269160 18566
rect 269132 3454 269344 3482
rect 269316 480 269344 3454
rect 270512 3398 270540 49166
rect 271064 48754 271092 52020
rect 272260 48822 272288 52020
rect 273456 48822 273484 52020
rect 274652 48822 274680 52020
rect 275862 52006 275968 52034
rect 277058 52006 277348 52034
rect 272248 48816 272300 48822
rect 272248 48758 272300 48764
rect 273168 48816 273220 48822
rect 273168 48758 273220 48764
rect 273444 48816 273496 48822
rect 273444 48758 273496 48764
rect 274548 48816 274600 48822
rect 274548 48758 274600 48764
rect 274640 48816 274692 48822
rect 274640 48758 274692 48764
rect 275836 48816 275888 48822
rect 275836 48758 275888 48764
rect 271052 48748 271104 48754
rect 271052 48690 271104 48696
rect 272524 48748 272576 48754
rect 272524 48690 272576 48696
rect 272536 26994 272564 48690
rect 272524 26988 272576 26994
rect 272524 26930 272576 26936
rect 273180 21418 273208 48758
rect 273260 43444 273312 43450
rect 273260 43386 273312 43392
rect 271880 21412 271932 21418
rect 271880 21354 271932 21360
rect 273168 21412 273220 21418
rect 273168 21354 273220 21360
rect 270592 6180 270644 6186
rect 270592 6122 270644 6128
rect 270500 3392 270552 3398
rect 270500 3334 270552 3340
rect 270604 3210 270632 6122
rect 271892 3482 271920 21354
rect 273272 3482 273300 43386
rect 274560 35222 274588 48758
rect 274548 35216 274600 35222
rect 274548 35158 274600 35164
rect 275848 24206 275876 48758
rect 275940 47598 275968 52006
rect 275928 47592 275980 47598
rect 275928 47534 275980 47540
rect 277320 36582 277348 52006
rect 278240 46306 278268 52020
rect 279450 52006 280108 52034
rect 278964 49088 279016 49094
rect 278964 49030 279016 49036
rect 278228 46300 278280 46306
rect 278228 46242 278280 46248
rect 277308 36576 277360 36582
rect 277308 36518 277360 36524
rect 277400 32428 277452 32434
rect 277400 32370 277452 32376
rect 275836 24200 275888 24206
rect 275836 24142 275888 24148
rect 276020 22772 276072 22778
rect 276020 22714 276072 22720
rect 276032 3482 276060 22714
rect 271892 3454 272932 3482
rect 273272 3454 274128 3482
rect 276032 3454 276520 3482
rect 271696 3392 271748 3398
rect 271696 3334 271748 3340
rect 270512 3182 270632 3210
rect 270512 480 270540 3182
rect 271708 480 271736 3334
rect 272904 480 272932 3454
rect 274100 480 274128 3454
rect 275284 3256 275336 3262
rect 275284 3198 275336 3204
rect 275296 480 275324 3198
rect 276492 480 276520 3454
rect 277412 3380 277440 32370
rect 278976 3482 279004 49030
rect 279976 6248 280028 6254
rect 279976 6190 280028 6196
rect 279988 6066 280016 6190
rect 280080 6186 280108 52006
rect 280632 48822 280660 52020
rect 281828 48822 281856 52020
rect 283024 48822 283052 52020
rect 284128 52006 284234 52034
rect 285430 52006 285628 52034
rect 286626 52006 287008 52034
rect 287822 52006 288388 52034
rect 289018 52006 289768 52034
rect 280620 48816 280672 48822
rect 280620 48758 280672 48764
rect 281448 48816 281500 48822
rect 281448 48758 281500 48764
rect 281816 48816 281868 48822
rect 281816 48758 281868 48764
rect 282828 48816 282880 48822
rect 282828 48758 282880 48764
rect 283012 48816 283064 48822
rect 283012 48758 283064 48764
rect 280160 46368 280212 46374
rect 280160 46310 280212 46316
rect 280068 6180 280120 6186
rect 280068 6122 280120 6128
rect 279988 6038 280108 6066
rect 278884 3454 279004 3482
rect 277412 3352 277716 3380
rect 277688 480 277716 3352
rect 278884 480 278912 3454
rect 280080 480 280108 6038
rect 280172 3380 280200 46310
rect 281460 39438 281488 48758
rect 281448 39432 281500 39438
rect 281448 39374 281500 39380
rect 282840 6254 282868 48758
rect 284128 44878 284156 52006
rect 284208 48816 284260 48822
rect 284208 48758 284260 48764
rect 284116 44872 284168 44878
rect 284116 44814 284168 44820
rect 284220 7614 284248 48758
rect 284300 33788 284352 33794
rect 284300 33730 284352 33736
rect 283656 7608 283708 7614
rect 283656 7550 283708 7556
rect 284208 7608 284260 7614
rect 284208 7550 284260 7556
rect 282828 6248 282880 6254
rect 282828 6190 282880 6196
rect 282460 3800 282512 3806
rect 282460 3742 282512 3748
rect 280172 3352 281304 3380
rect 281276 480 281304 3352
rect 282472 480 282500 3742
rect 283668 480 283696 7550
rect 284312 3380 284340 33730
rect 285600 10402 285628 52006
rect 285772 49156 285824 49162
rect 285772 49098 285824 49104
rect 285588 10396 285640 10402
rect 285588 10338 285640 10344
rect 285784 3380 285812 49098
rect 286980 22778 287008 52006
rect 288360 38010 288388 52006
rect 288348 38004 288400 38010
rect 288348 37946 288400 37952
rect 287060 35352 287112 35358
rect 287060 35294 287112 35300
rect 286968 22772 287020 22778
rect 286968 22714 287020 22720
rect 287072 3398 287100 35294
rect 287152 24132 287204 24138
rect 287152 24074 287204 24080
rect 287060 3392 287112 3398
rect 284312 3352 284800 3380
rect 285784 3352 285996 3380
rect 284772 480 284800 3352
rect 285968 480 285996 3352
rect 287060 3334 287112 3340
rect 287164 480 287192 24074
rect 289544 3868 289596 3874
rect 289544 3810 289596 3816
rect 288348 3392 288400 3398
rect 288348 3334 288400 3340
rect 288360 480 288388 3334
rect 289556 480 289584 3810
rect 289740 3806 289768 52006
rect 290200 48822 290228 52020
rect 291396 48822 291424 52020
rect 292592 48822 292620 52020
rect 290188 48816 290240 48822
rect 290188 48758 290240 48764
rect 291108 48816 291160 48822
rect 291108 48758 291160 48764
rect 291384 48816 291436 48822
rect 291384 48758 291436 48764
rect 292488 48816 292540 48822
rect 292488 48758 292540 48764
rect 292580 48816 292632 48822
rect 292580 48758 292632 48764
rect 290740 9036 290792 9042
rect 290740 8978 290792 8984
rect 289728 3800 289780 3806
rect 289728 3742 289780 3748
rect 290752 480 290780 8978
rect 291120 8974 291148 48758
rect 291200 36644 291252 36650
rect 291200 36586 291252 36592
rect 291108 8968 291160 8974
rect 291108 8910 291160 8916
rect 291212 3346 291240 36586
rect 292500 29714 292528 48758
rect 293696 46238 293724 52020
rect 294906 52006 295288 52034
rect 296102 52006 296668 52034
rect 297298 52006 298048 52034
rect 293868 48816 293920 48822
rect 293868 48758 293920 48764
rect 293684 46232 293736 46238
rect 293684 46174 293736 46180
rect 292488 29708 292540 29714
rect 292488 29650 292540 29656
rect 293880 3874 293908 48758
rect 293960 10328 294012 10334
rect 293960 10270 294012 10276
rect 293868 3868 293920 3874
rect 293868 3810 293920 3816
rect 293132 3664 293184 3670
rect 293132 3606 293184 3612
rect 291212 3318 291976 3346
rect 291948 480 291976 3318
rect 293144 480 293172 3606
rect 293972 3346 294000 10270
rect 295260 4826 295288 52006
rect 295340 39364 295392 39370
rect 295340 39306 295392 39312
rect 295248 4820 295300 4826
rect 295248 4762 295300 4768
rect 295352 3448 295380 39306
rect 296640 3738 296668 52006
rect 296812 25628 296864 25634
rect 296812 25570 296864 25576
rect 296628 3732 296680 3738
rect 296628 3674 296680 3680
rect 296824 3482 296852 25570
rect 298020 10334 298048 52006
rect 298480 48822 298508 52020
rect 299676 48822 299704 52020
rect 300872 48822 300900 52020
rect 298468 48816 298520 48822
rect 298468 48758 298520 48764
rect 299388 48816 299440 48822
rect 299388 48758 299440 48764
rect 299664 48816 299716 48822
rect 299664 48758 299716 48764
rect 300768 48816 300820 48822
rect 300768 48758 300820 48764
rect 300860 48816 300912 48822
rect 300860 48758 300912 48764
rect 298100 44940 298152 44946
rect 298100 44882 298152 44888
rect 298008 10328 298060 10334
rect 298008 10270 298060 10276
rect 298112 3482 298140 44882
rect 299400 40866 299428 48758
rect 299388 40860 299440 40866
rect 299388 40802 299440 40808
rect 300308 4140 300360 4146
rect 300308 4082 300360 4088
rect 296720 3460 296772 3466
rect 295352 3420 295564 3448
rect 293972 3318 294368 3346
rect 294340 480 294368 3318
rect 295536 480 295564 3420
rect 296824 3454 297956 3482
rect 298112 3454 299152 3482
rect 296720 3402 296772 3408
rect 296732 480 296760 3402
rect 297928 480 297956 3454
rect 299124 480 299152 3454
rect 300320 480 300348 4082
rect 300780 3466 300808 48758
rect 302068 28286 302096 52020
rect 303278 52006 303568 52034
rect 304474 52006 304948 52034
rect 305670 52006 306328 52034
rect 302148 48816 302200 48822
rect 302148 48758 302200 48764
rect 302056 28280 302108 28286
rect 302056 28222 302108 28228
rect 302160 11830 302188 48758
rect 302240 37936 302292 37942
rect 302240 37878 302292 37884
rect 302148 11824 302200 11830
rect 302148 11766 302200 11772
rect 300860 11756 300912 11762
rect 300860 11698 300912 11704
rect 300872 3482 300900 11698
rect 302252 3482 302280 37878
rect 303540 11762 303568 52006
rect 304920 24138 304948 52006
rect 306300 31210 306328 52006
rect 306852 48822 306880 52020
rect 308048 48822 308076 52020
rect 309244 48822 309272 52020
rect 306840 48816 306892 48822
rect 306840 48758 306892 48764
rect 307668 48816 307720 48822
rect 307668 48758 307720 48764
rect 308036 48816 308088 48822
rect 308036 48758 308088 48764
rect 309048 48816 309100 48822
rect 309048 48758 309100 48764
rect 309232 48816 309284 48822
rect 309232 48758 309284 48764
rect 310336 48816 310388 48822
rect 310336 48758 310388 48764
rect 306288 31204 306340 31210
rect 306288 31146 306340 31152
rect 305000 29776 305052 29782
rect 305000 29718 305052 29724
rect 304908 24132 304960 24138
rect 304908 24074 304960 24080
rect 303528 11756 303580 11762
rect 303528 11698 303580 11704
rect 305012 3602 305040 29718
rect 305092 26920 305144 26926
rect 305092 26862 305144 26868
rect 303804 3596 303856 3602
rect 303804 3538 303856 3544
rect 305000 3596 305052 3602
rect 305000 3538 305052 3544
rect 300768 3460 300820 3466
rect 300872 3454 301452 3482
rect 302252 3454 302648 3482
rect 300768 3402 300820 3408
rect 301424 480 301452 3454
rect 302620 480 302648 3454
rect 303816 480 303844 3538
rect 305104 3482 305132 26862
rect 307392 4004 307444 4010
rect 307392 3946 307444 3952
rect 306196 3596 306248 3602
rect 306196 3538 306248 3544
rect 305012 3454 305132 3482
rect 305012 480 305040 3454
rect 306208 480 306236 3538
rect 307404 480 307432 3946
rect 307680 3942 307708 48758
rect 309060 14482 309088 48758
rect 310348 42090 310376 48758
rect 310336 42084 310388 42090
rect 310336 42026 310388 42032
rect 309140 40792 309192 40798
rect 309140 40734 309192 40740
rect 307760 14476 307812 14482
rect 307760 14418 307812 14424
rect 309048 14476 309100 14482
rect 309048 14418 309100 14424
rect 307668 3936 307720 3942
rect 307668 3878 307720 3884
rect 307772 3346 307800 14418
rect 309152 3346 309180 40734
rect 310440 3602 310468 52020
rect 311636 49162 311664 52020
rect 312846 52006 313228 52034
rect 314042 52006 314608 52034
rect 311624 49156 311676 49162
rect 311624 49098 311676 49104
rect 313200 43450 313228 52006
rect 313464 49292 313516 49298
rect 313464 49234 313516 49240
rect 313188 43444 313240 43450
rect 313188 43386 313240 43392
rect 313372 28348 313424 28354
rect 313372 28290 313424 28296
rect 311900 13116 311952 13122
rect 311900 13058 311952 13064
rect 310428 3596 310480 3602
rect 310428 3538 310480 3544
rect 310980 3528 311032 3534
rect 310980 3470 311032 3476
rect 307772 3318 308628 3346
rect 309152 3318 309824 3346
rect 308600 480 308628 3318
rect 309796 480 309824 3318
rect 310992 480 311020 3470
rect 311912 3346 311940 13058
rect 311912 3318 312216 3346
rect 312188 480 312216 3318
rect 313384 480 313412 28290
rect 313476 3346 313504 49234
rect 314580 4010 314608 52006
rect 315224 48754 315252 52020
rect 316420 48822 316448 52020
rect 316408 48816 316460 48822
rect 316408 48758 316460 48764
rect 317328 48816 317380 48822
rect 317328 48758 317380 48764
rect 315212 48748 315264 48754
rect 315212 48690 315264 48696
rect 315948 48748 316000 48754
rect 315948 48690 316000 48696
rect 315960 13122 315988 48690
rect 316040 42220 316092 42226
rect 316040 42162 316092 42168
rect 315948 13116 316000 13122
rect 315948 13058 316000 13064
rect 315764 4888 315816 4894
rect 315764 4830 315816 4836
rect 314568 4004 314620 4010
rect 314568 3946 314620 3952
rect 313476 3318 314608 3346
rect 314580 480 314608 3318
rect 315776 480 315804 4830
rect 316052 3346 316080 42162
rect 317340 32570 317368 48758
rect 317616 48346 317644 52020
rect 318628 52006 318734 52034
rect 319930 52006 320128 52034
rect 321126 52006 321508 52034
rect 322322 52006 322888 52034
rect 317604 48340 317656 48346
rect 317604 48282 317656 48288
rect 317328 32564 317380 32570
rect 317328 32506 317380 32512
rect 318628 15978 318656 52006
rect 318708 48340 318760 48346
rect 318708 48282 318760 48288
rect 318616 15972 318668 15978
rect 318616 15914 318668 15920
rect 318064 4072 318116 4078
rect 318064 4014 318116 4020
rect 316052 3318 317000 3346
rect 316972 480 317000 3318
rect 318076 480 318104 4014
rect 318720 3330 318748 48282
rect 320100 33794 320128 52006
rect 320088 33788 320140 33794
rect 320088 33730 320140 33736
rect 320180 31136 320232 31142
rect 320180 31078 320232 31084
rect 318800 15904 318852 15910
rect 318800 15846 318852 15852
rect 318812 3346 318840 15846
rect 320192 3346 320220 31078
rect 321480 3534 321508 52006
rect 321744 49020 321796 49026
rect 321744 48962 321796 48968
rect 321652 17264 321704 17270
rect 321652 17206 321704 17212
rect 321664 7682 321692 17206
rect 321652 7676 321704 7682
rect 321652 7618 321704 7624
rect 321756 7562 321784 48962
rect 322860 17270 322888 52006
rect 323504 48822 323532 52020
rect 324700 48822 324728 52020
rect 325896 48822 325924 52020
rect 327092 48822 327120 52020
rect 328302 52006 328408 52034
rect 323492 48816 323544 48822
rect 323492 48758 323544 48764
rect 324228 48816 324280 48822
rect 324228 48758 324280 48764
rect 324688 48816 324740 48822
rect 324688 48758 324740 48764
rect 325608 48816 325660 48822
rect 325608 48758 325660 48764
rect 325884 48816 325936 48822
rect 325884 48758 325936 48764
rect 326988 48816 327040 48822
rect 326988 48758 327040 48764
rect 327080 48816 327132 48822
rect 327080 48758 327132 48764
rect 328276 48816 328328 48822
rect 328276 48758 328328 48764
rect 323032 43512 323084 43518
rect 323032 43454 323084 43460
rect 323044 38706 323072 43454
rect 322952 38678 323072 38706
rect 322848 17264 322900 17270
rect 322848 17206 322900 17212
rect 322952 12510 322980 38678
rect 324240 35358 324268 48758
rect 324228 35352 324280 35358
rect 324228 35294 324280 35300
rect 322940 12504 322992 12510
rect 322940 12446 322992 12452
rect 324044 12436 324096 12442
rect 324044 12378 324096 12384
rect 324056 9654 324084 12378
rect 324044 9648 324096 9654
rect 324044 9590 324096 9596
rect 324044 9512 324096 9518
rect 324044 9454 324096 9460
rect 322848 7676 322900 7682
rect 322848 7618 322900 7624
rect 321664 7534 321784 7562
rect 321468 3528 321520 3534
rect 321468 3470 321520 3476
rect 318708 3324 318760 3330
rect 318812 3318 319300 3346
rect 320192 3318 320496 3346
rect 318708 3266 318760 3272
rect 319272 480 319300 3318
rect 320468 480 320496 3318
rect 321664 480 321692 7534
rect 322860 480 322888 7618
rect 324056 480 324084 9454
rect 325240 7744 325292 7750
rect 325240 7686 325292 7692
rect 325252 480 325280 7686
rect 325620 3262 325648 48758
rect 327000 19990 327028 48758
rect 328288 36650 328316 48758
rect 328276 36644 328328 36650
rect 328276 36586 328328 36592
rect 327080 32496 327132 32502
rect 327080 32438 327132 32444
rect 325700 19984 325752 19990
rect 325700 19926 325752 19932
rect 326988 19984 327040 19990
rect 326988 19926 327040 19932
rect 325712 12510 325740 19926
rect 327092 12510 327120 32438
rect 325700 12504 325752 12510
rect 325700 12446 325752 12452
rect 327080 12504 327132 12510
rect 327080 12446 327132 12452
rect 326436 12436 326488 12442
rect 326436 12378 326488 12384
rect 326448 9654 326476 12378
rect 327632 12368 327684 12374
rect 327632 12310 327684 12316
rect 327644 9654 327672 12310
rect 326436 9648 326488 9654
rect 326436 9590 326488 9596
rect 327632 9648 327684 9654
rect 327632 9590 327684 9596
rect 326436 9512 326488 9518
rect 326436 9454 326488 9460
rect 327632 9512 327684 9518
rect 327632 9454 327684 9460
rect 325608 3256 325660 3262
rect 325608 3198 325660 3204
rect 326448 480 326476 9454
rect 327644 480 327672 9454
rect 328380 3534 328408 52006
rect 329484 48822 329512 52020
rect 330694 52006 331168 52034
rect 331890 52006 332548 52034
rect 329472 48816 329524 48822
rect 329472 48758 329524 48764
rect 330484 48816 330536 48822
rect 330484 48758 330536 48764
rect 328552 25560 328604 25566
rect 328552 25502 328604 25508
rect 328564 19394 328592 25502
rect 328472 19366 328592 19394
rect 328472 19310 328500 19366
rect 328460 19304 328512 19310
rect 328460 19246 328512 19252
rect 330496 18630 330524 48758
rect 331140 39506 331168 52006
rect 331128 39500 331180 39506
rect 331128 39442 331180 39448
rect 331220 33856 331272 33862
rect 331220 33798 331272 33804
rect 330484 18624 330536 18630
rect 330484 18566 330536 18572
rect 328828 9716 328880 9722
rect 328828 9658 328880 9664
rect 330024 9716 330076 9722
rect 330024 9658 330076 9664
rect 328840 9602 328868 9658
rect 328840 9574 328960 9602
rect 328368 3528 328420 3534
rect 328368 3470 328420 3476
rect 328932 610 328960 9574
rect 328828 604 328880 610
rect 328828 546 328880 552
rect 328920 604 328972 610
rect 328920 546 328972 552
rect 328840 480 328868 546
rect 330036 480 330064 9658
rect 331232 480 331260 33798
rect 331312 26988 331364 26994
rect 331312 26930 331364 26936
rect 331324 3346 331352 26930
rect 331324 3318 332456 3346
rect 332428 480 332456 3318
rect 332520 3194 332548 52006
rect 333072 48822 333100 52020
rect 334268 48822 334296 52020
rect 335464 48822 335492 52020
rect 336568 52006 336674 52034
rect 337870 52006 338068 52034
rect 339066 52006 339448 52034
rect 340262 52006 340828 52034
rect 341458 52006 342208 52034
rect 333060 48816 333112 48822
rect 333060 48758 333112 48764
rect 333888 48816 333940 48822
rect 333888 48758 333940 48764
rect 334256 48816 334308 48822
rect 334256 48758 334308 48764
rect 335268 48816 335320 48822
rect 335268 48758 335320 48764
rect 335452 48816 335504 48822
rect 335452 48758 335504 48764
rect 333900 21418 333928 48758
rect 333980 35216 334032 35222
rect 333980 35158 334032 35164
rect 332600 21412 332652 21418
rect 332600 21354 332652 21360
rect 333888 21412 333940 21418
rect 333888 21354 333940 21360
rect 332612 3346 332640 21354
rect 333992 3346 334020 35158
rect 335280 22846 335308 48758
rect 336568 25566 336596 52006
rect 336648 48816 336700 48822
rect 336648 48758 336700 48764
rect 336556 25560 336608 25566
rect 336556 25502 336608 25508
rect 335360 24200 335412 24206
rect 335360 24142 335412 24148
rect 335268 22840 335320 22846
rect 335268 22782 335320 22788
rect 335372 3482 335400 24142
rect 335372 3454 335952 3482
rect 332612 3318 333652 3346
rect 333992 3318 334756 3346
rect 332508 3188 332560 3194
rect 332508 3130 332560 3136
rect 333624 480 333652 3318
rect 334728 480 334756 3318
rect 335924 480 335952 3454
rect 336660 3398 336688 48758
rect 336740 47592 336792 47598
rect 336740 47534 336792 47540
rect 336752 3482 336780 47534
rect 338040 44946 338068 52006
rect 338028 44940 338080 44946
rect 338028 44882 338080 44888
rect 338120 36576 338172 36582
rect 338120 36518 338172 36524
rect 338132 3482 338160 36518
rect 336752 3454 337148 3482
rect 338132 3454 338344 3482
rect 336648 3392 336700 3398
rect 336648 3334 336700 3340
rect 337120 480 337148 3454
rect 338316 480 338344 3454
rect 339420 3369 339448 52006
rect 339500 46300 339552 46306
rect 339500 46242 339552 46248
rect 339406 3360 339462 3369
rect 339406 3295 339462 3304
rect 339512 480 339540 46242
rect 340800 7682 340828 52006
rect 340880 39432 340932 39438
rect 340880 39374 340932 39380
rect 340788 7676 340840 7682
rect 340788 7618 340840 7624
rect 340696 6180 340748 6186
rect 340696 6122 340748 6128
rect 340708 480 340736 6122
rect 340892 3482 340920 39374
rect 342180 37942 342208 52006
rect 342640 48822 342668 52020
rect 343744 48822 343772 52020
rect 342628 48816 342680 48822
rect 342628 48758 342680 48764
rect 343548 48816 343600 48822
rect 343548 48758 343600 48764
rect 343732 48816 343784 48822
rect 343732 48758 343784 48764
rect 344836 48816 344888 48822
rect 344836 48758 344888 48764
rect 342168 37936 342220 37942
rect 342168 37878 342220 37884
rect 343088 6248 343140 6254
rect 343088 6190 343140 6196
rect 340892 3454 341932 3482
rect 341904 480 341932 3454
rect 343100 480 343128 6190
rect 343560 3126 343588 48758
rect 344848 26926 344876 48758
rect 344836 26920 344888 26926
rect 344836 26862 344888 26868
rect 344284 7608 344336 7614
rect 344284 7550 344336 7556
rect 343548 3120 343600 3126
rect 343548 3062 343600 3068
rect 344296 480 344324 7550
rect 344940 6186 344968 52020
rect 345664 49156 345716 49162
rect 345664 49098 345716 49104
rect 345020 44872 345072 44878
rect 345020 44814 345072 44820
rect 344928 6180 344980 6186
rect 344928 6122 344980 6128
rect 345032 3482 345060 44814
rect 345676 6254 345704 49098
rect 346136 49094 346164 52020
rect 346124 49088 346176 49094
rect 346124 49030 346176 49036
rect 347332 47598 347360 52020
rect 348542 52006 349108 52034
rect 349738 52006 350488 52034
rect 347320 47592 347372 47598
rect 347320 47534 347372 47540
rect 347780 38004 347832 38010
rect 347780 37946 347832 37952
rect 346400 10396 346452 10402
rect 346400 10338 346452 10344
rect 345664 6248 345716 6254
rect 345664 6190 345716 6196
rect 346412 3482 346440 10338
rect 347792 3806 347820 37946
rect 349080 29646 349108 52006
rect 349068 29640 349120 29646
rect 349068 29582 349120 29588
rect 347872 22772 347924 22778
rect 347872 22714 347924 22720
rect 347780 3800 347832 3806
rect 347780 3742 347832 3748
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347884 480 347912 22714
rect 350460 4078 350488 52006
rect 350920 48822 350948 52020
rect 352116 48822 352144 52020
rect 353312 48822 353340 52020
rect 354508 49026 354536 52020
rect 355718 52006 356008 52034
rect 356914 52006 357388 52034
rect 358110 52006 358768 52034
rect 354496 49020 354548 49026
rect 354496 48962 354548 48968
rect 350908 48816 350960 48822
rect 350908 48758 350960 48764
rect 351828 48816 351880 48822
rect 351828 48758 351880 48764
rect 352104 48816 352156 48822
rect 352104 48758 352156 48764
rect 353208 48816 353260 48822
rect 353208 48758 353260 48764
rect 353300 48816 353352 48822
rect 353300 48758 353352 48764
rect 354588 48816 354640 48822
rect 354588 48758 354640 48764
rect 351840 8974 351868 48758
rect 351920 29708 351972 29714
rect 351920 29650 351972 29656
rect 351368 8968 351420 8974
rect 351368 8910 351420 8916
rect 351828 8968 351880 8974
rect 351828 8910 351880 8916
rect 350448 4072 350500 4078
rect 350448 4014 350500 4020
rect 350264 3868 350316 3874
rect 350264 3810 350316 3816
rect 349068 3800 349120 3806
rect 349068 3742 349120 3748
rect 349080 480 349108 3742
rect 350276 480 350304 3810
rect 351380 480 351408 8910
rect 351932 3482 351960 29650
rect 353220 28354 353248 48758
rect 353208 28348 353260 28354
rect 353208 28290 353260 28296
rect 353760 4140 353812 4146
rect 353760 4082 353812 4088
rect 351932 3454 352604 3482
rect 352576 480 352604 3454
rect 353772 480 353800 4082
rect 354600 3874 354628 48758
rect 354680 46232 354732 46238
rect 354680 46174 354732 46180
rect 354588 3868 354640 3874
rect 354588 3810 354640 3816
rect 354692 610 354720 46174
rect 355980 40730 356008 52006
rect 355968 40724 356020 40730
rect 355968 40666 356020 40672
rect 356152 4820 356204 4826
rect 356152 4762 356204 4768
rect 354680 604 354732 610
rect 354680 546 354732 552
rect 354956 604 355008 610
rect 354956 546 355008 552
rect 354968 480 354996 546
rect 356164 480 356192 4762
rect 357360 3856 357388 52006
rect 357440 10328 357492 10334
rect 357440 10270 357492 10276
rect 357452 4026 357480 10270
rect 358740 5030 358768 52006
rect 359292 48822 359320 52020
rect 360488 48822 360516 52020
rect 361684 48822 361712 52020
rect 362788 52006 362894 52034
rect 364090 52006 364288 52034
rect 359280 48816 359332 48822
rect 359280 48758 359332 48764
rect 360108 48816 360160 48822
rect 360108 48758 360160 48764
rect 360476 48816 360528 48822
rect 360476 48758 360528 48764
rect 361488 48816 361540 48822
rect 361488 48758 361540 48764
rect 361672 48816 361724 48822
rect 361672 48758 361724 48764
rect 358820 40860 358872 40866
rect 358820 40802 358872 40808
rect 358728 5024 358780 5030
rect 358728 4966 358780 4972
rect 357452 3998 357572 4026
rect 357360 3828 357480 3856
rect 357452 3738 357480 3828
rect 357348 3732 357400 3738
rect 357348 3674 357400 3680
rect 357440 3732 357492 3738
rect 357440 3674 357492 3680
rect 357360 480 357388 3674
rect 357544 610 357572 3998
rect 358832 610 358860 40802
rect 360120 24206 360148 48758
rect 360108 24200 360160 24206
rect 360108 24142 360160 24148
rect 361500 4146 361528 48758
rect 362788 31074 362816 52006
rect 362868 48816 362920 48822
rect 362868 48758 362920 48764
rect 362776 31068 362828 31074
rect 362776 31010 362828 31016
rect 361580 11824 361632 11830
rect 361580 11766 361632 11772
rect 361488 4140 361540 4146
rect 361488 4082 361540 4088
rect 360936 3460 360988 3466
rect 360936 3402 360988 3408
rect 357532 604 357584 610
rect 357532 546 357584 552
rect 358544 604 358596 610
rect 358544 546 358596 552
rect 358820 604 358872 610
rect 358820 546 358872 552
rect 359740 604 359792 610
rect 359740 546 359792 552
rect 358556 480 358584 546
rect 359752 480 359780 546
rect 360948 480 360976 3402
rect 361592 610 361620 11766
rect 362880 5302 362908 48758
rect 362960 28280 363012 28286
rect 362960 28222 363012 28228
rect 362868 5296 362920 5302
rect 362868 5238 362920 5244
rect 362972 626 363000 28222
rect 364260 3505 364288 52006
rect 365272 46238 365300 52020
rect 366482 52006 367048 52034
rect 365260 46232 365312 46238
rect 365260 46174 365312 46180
rect 367020 32434 367048 52006
rect 367664 49230 367692 52020
rect 367652 49224 367704 49230
rect 367652 49166 367704 49172
rect 367744 49020 367796 49026
rect 367744 48962 367796 48968
rect 367008 32428 367060 32434
rect 367008 32370 367060 32376
rect 365720 31204 365772 31210
rect 365720 31146 365772 31152
rect 364340 11756 364392 11762
rect 364340 11698 364392 11704
rect 364246 3496 364302 3505
rect 364246 3431 364302 3440
rect 364352 3346 364380 11698
rect 365732 3466 365760 31146
rect 365812 24132 365864 24138
rect 365812 24074 365864 24080
rect 365720 3460 365772 3466
rect 365720 3402 365772 3408
rect 364352 3318 364564 3346
rect 361580 604 361632 610
rect 361580 546 361632 552
rect 362132 604 362184 610
rect 362972 598 363368 626
rect 362132 546 362184 552
rect 362144 480 362172 546
rect 363340 480 363368 598
rect 364536 480 364564 3318
rect 365824 1442 365852 24074
rect 367756 10334 367784 48962
rect 368860 48346 368888 52020
rect 369964 48822 369992 52020
rect 369952 48816 370004 48822
rect 369952 48758 370004 48764
rect 368848 48340 368900 48346
rect 368848 48282 368900 48288
rect 369768 48340 369820 48346
rect 369768 48282 369820 48288
rect 368480 14476 368532 14482
rect 368480 14418 368532 14424
rect 367744 10328 367796 10334
rect 367744 10270 367796 10276
rect 368020 3936 368072 3942
rect 368020 3878 368072 3884
rect 366916 3460 366968 3466
rect 366916 3402 366968 3408
rect 365732 1414 365852 1442
rect 365732 480 365760 1414
rect 366928 480 366956 3402
rect 368032 480 368060 3878
rect 368492 3346 368520 14418
rect 369780 5234 369808 48282
rect 369860 42084 369912 42090
rect 369860 42026 369912 42032
rect 369872 38622 369900 42026
rect 369860 38616 369912 38622
rect 369860 38558 369912 38564
rect 369952 38616 370004 38622
rect 369952 38558 370004 38564
rect 369964 29050 369992 38558
rect 369872 29022 369992 29050
rect 369872 27606 369900 29022
rect 369860 27600 369912 27606
rect 369860 27542 369912 27548
rect 370504 27600 370556 27606
rect 370504 27542 370556 27548
rect 369768 5228 369820 5234
rect 369768 5170 369820 5176
rect 370516 3448 370544 27542
rect 371160 3466 371188 52020
rect 372370 52006 372568 52034
rect 373566 52006 373948 52034
rect 371884 48816 371936 48822
rect 371884 48758 371936 48764
rect 371896 33862 371924 48758
rect 371884 33856 371936 33862
rect 371884 33798 371936 33804
rect 372540 4826 372568 52006
rect 373920 35290 373948 52006
rect 374748 49298 374776 52020
rect 374736 49292 374788 49298
rect 374736 49234 374788 49240
rect 375944 48754 375972 52020
rect 377140 48822 377168 52020
rect 378336 48822 378364 52020
rect 379532 48822 379560 52020
rect 377128 48816 377180 48822
rect 377128 48758 377180 48764
rect 378048 48816 378100 48822
rect 378048 48758 378100 48764
rect 378324 48816 378376 48822
rect 378324 48758 378376 48764
rect 379428 48816 379480 48822
rect 379428 48758 379480 48764
rect 379520 48816 379572 48822
rect 379520 48758 379572 48764
rect 375932 48748 375984 48754
rect 375932 48690 375984 48696
rect 376668 48748 376720 48754
rect 376668 48690 376720 48696
rect 374092 43444 374144 43450
rect 374092 43386 374144 43392
rect 373908 35284 373960 35290
rect 373908 35226 373960 35232
rect 372804 6248 372856 6254
rect 372804 6190 372856 6196
rect 372528 4820 372580 4826
rect 372528 4762 372580 4768
rect 371608 3596 371660 3602
rect 371608 3538 371660 3544
rect 370424 3420 370544 3448
rect 371148 3460 371200 3466
rect 368492 3318 369256 3346
rect 369228 480 369256 3318
rect 370424 480 370452 3420
rect 371148 3402 371200 3408
rect 371620 480 371648 3538
rect 372816 480 372844 6190
rect 374104 2854 374132 43386
rect 375380 13116 375432 13122
rect 375380 13058 375432 13064
rect 375392 12442 375420 13058
rect 375380 12436 375432 12442
rect 375380 12378 375432 12384
rect 376392 12436 376444 12442
rect 376392 12378 376444 12384
rect 375196 4004 375248 4010
rect 375196 3946 375248 3952
rect 374092 2848 374144 2854
rect 374092 2790 374144 2796
rect 374000 2780 374052 2786
rect 374000 2722 374052 2728
rect 374012 480 374040 2722
rect 375208 480 375236 3946
rect 376404 480 376432 12378
rect 376680 11762 376708 48690
rect 378060 36582 378088 48758
rect 378048 36576 378100 36582
rect 378048 36518 378100 36524
rect 376760 32564 376812 32570
rect 376760 32506 376812 32512
rect 376772 12442 376800 32506
rect 376760 12436 376812 12442
rect 376760 12378 376812 12384
rect 377588 12436 377640 12442
rect 377588 12378 377640 12384
rect 376668 11756 376720 11762
rect 376668 11698 376720 11704
rect 377600 480 377628 12378
rect 379440 3806 379468 48758
rect 380728 39370 380756 52020
rect 381924 49026 381952 52020
rect 381912 49020 381964 49026
rect 381912 48962 381964 48968
rect 380808 48816 380860 48822
rect 380808 48758 380860 48764
rect 380716 39364 380768 39370
rect 380716 39306 380768 39312
rect 379520 15972 379572 15978
rect 379520 15914 379572 15920
rect 379428 3800 379480 3806
rect 379428 3742 379480 3748
rect 379532 3346 379560 15914
rect 380820 5098 380848 48758
rect 383120 48686 383148 52020
rect 384330 52006 384988 52034
rect 383108 48680 383160 48686
rect 383108 48622 383160 48628
rect 384304 48680 384356 48686
rect 384304 48622 384356 48628
rect 383660 35352 383712 35358
rect 383660 35294 383712 35300
rect 380900 33788 380952 33794
rect 380900 33730 380952 33736
rect 380808 5092 380860 5098
rect 380808 5034 380860 5040
rect 380912 3346 380940 33730
rect 382372 17264 382424 17270
rect 382372 17206 382424 17212
rect 382280 3664 382332 3670
rect 382280 3606 382332 3612
rect 382292 3482 382320 3606
rect 382384 3602 382412 17206
rect 382372 3596 382424 3602
rect 382372 3538 382424 3544
rect 383568 3596 383620 3602
rect 383568 3538 383620 3544
rect 382292 3454 382412 3482
rect 378784 3324 378836 3330
rect 379532 3318 380020 3346
rect 380912 3318 381216 3346
rect 378784 3266 378836 3272
rect 378796 480 378824 3266
rect 379992 480 380020 3318
rect 381188 480 381216 3318
rect 382384 480 382412 3454
rect 383580 480 383608 3538
rect 383672 610 383700 35294
rect 384316 13122 384344 48622
rect 384960 44878 384988 52006
rect 385512 48414 385540 52020
rect 386708 48822 386736 52020
rect 386696 48816 386748 48822
rect 386696 48758 386748 48764
rect 387708 48816 387760 48822
rect 387708 48758 387760 48764
rect 385500 48408 385552 48414
rect 385500 48350 385552 48356
rect 386328 48408 386380 48414
rect 386328 48350 386380 48356
rect 384948 44872 385000 44878
rect 384948 44814 385000 44820
rect 384304 13116 384356 13122
rect 384304 13058 384356 13064
rect 386340 3670 386368 48350
rect 386420 19984 386472 19990
rect 386420 19926 386472 19932
rect 386328 3664 386380 3670
rect 386328 3606 386380 3612
rect 385868 3256 385920 3262
rect 385868 3198 385920 3204
rect 383660 604 383712 610
rect 383660 546 383712 552
rect 384672 604 384724 610
rect 384672 546 384724 552
rect 384684 480 384712 546
rect 385880 480 385908 3198
rect 386432 610 386460 19926
rect 387720 4962 387748 48758
rect 387904 48686 387932 52020
rect 389100 49162 389128 52020
rect 390310 52006 390508 52034
rect 391506 52006 391888 52034
rect 392702 52006 393268 52034
rect 393898 52006 394648 52034
rect 389088 49156 389140 49162
rect 389088 49098 389140 49104
rect 387892 48680 387944 48686
rect 387892 48622 387944 48628
rect 389088 48680 389140 48686
rect 389088 48622 389140 48628
rect 389100 38010 389128 48622
rect 389088 38004 389140 38010
rect 389088 37946 389140 37952
rect 387800 36644 387852 36650
rect 387800 36586 387852 36592
rect 387708 4956 387760 4962
rect 387708 4898 387760 4904
rect 387812 610 387840 36586
rect 390480 4894 390508 52006
rect 390560 39500 390612 39506
rect 390560 39442 390612 39448
rect 390572 7614 390600 39442
rect 391860 26994 391888 52006
rect 391848 26988 391900 26994
rect 391848 26930 391900 26936
rect 390652 18624 390704 18630
rect 390652 18566 390704 18572
rect 390560 7608 390612 7614
rect 390560 7550 390612 7556
rect 390468 4888 390520 4894
rect 390468 4830 390520 4836
rect 389456 3528 389508 3534
rect 389456 3470 389508 3476
rect 386420 604 386472 610
rect 386420 546 386472 552
rect 387064 604 387116 610
rect 387064 546 387116 552
rect 387800 604 387852 610
rect 387800 546 387852 552
rect 388260 604 388312 610
rect 388260 546 388312 552
rect 387076 480 387104 546
rect 388272 480 388300 546
rect 389468 480 389496 3470
rect 390664 480 390692 18566
rect 391848 7608 391900 7614
rect 391848 7550 391900 7556
rect 391860 480 391888 7550
rect 393240 3942 393268 52006
rect 393320 21412 393372 21418
rect 393320 21354 393372 21360
rect 393332 12442 393360 21354
rect 393320 12436 393372 12442
rect 393320 12378 393372 12384
rect 394240 12436 394292 12442
rect 394240 12378 394292 12384
rect 393228 3936 393280 3942
rect 393228 3878 393280 3884
rect 393044 3188 393096 3194
rect 393044 3130 393096 3136
rect 393056 480 393084 3130
rect 394252 480 394280 12378
rect 394620 5166 394648 52006
rect 394988 48822 395016 52020
rect 396184 49434 396212 52020
rect 396172 49428 396224 49434
rect 396172 49370 396224 49376
rect 394976 48816 395028 48822
rect 394976 48758 395028 48764
rect 395988 48816 396040 48822
rect 395988 48758 396040 48764
rect 396000 25634 396028 48758
rect 395988 25628 396040 25634
rect 395988 25570 396040 25576
rect 394792 22840 394844 22846
rect 394792 22782 394844 22788
rect 394804 19394 394832 22782
rect 394712 19366 394832 19394
rect 394712 19310 394740 19366
rect 394700 19304 394752 19310
rect 394700 19246 394752 19252
rect 397380 14482 397408 52020
rect 398590 52006 398788 52034
rect 399786 52006 400168 52034
rect 400982 52006 401548 52034
rect 402178 52006 402928 52034
rect 398760 28286 398788 52006
rect 398840 44940 398892 44946
rect 398840 44882 398892 44888
rect 398748 28280 398800 28286
rect 398748 28222 398800 28228
rect 397552 25560 397604 25566
rect 397552 25502 397604 25508
rect 397564 19394 397592 25502
rect 397472 19366 397592 19394
rect 397472 19310 397500 19366
rect 397460 19304 397512 19310
rect 397460 19246 397512 19252
rect 397368 14476 397420 14482
rect 397368 14418 397420 14424
rect 395436 9716 395488 9722
rect 395436 9658 395488 9664
rect 397828 9716 397880 9722
rect 397828 9658 397880 9664
rect 394608 5160 394660 5166
rect 394608 5102 394660 5108
rect 395448 480 395476 9658
rect 396632 3392 396684 3398
rect 396632 3334 396684 3340
rect 396644 480 396672 3334
rect 397840 480 397868 9658
rect 398852 3346 398880 44882
rect 400140 4010 400168 52006
rect 401520 43450 401548 52006
rect 401508 43444 401560 43450
rect 401508 43386 401560 43392
rect 401600 37936 401652 37942
rect 401600 37878 401652 37884
rect 401324 7676 401376 7682
rect 401324 7618 401376 7624
rect 400128 4004 400180 4010
rect 400128 3946 400180 3952
rect 400218 3360 400274 3369
rect 398852 3318 399064 3346
rect 399036 480 399064 3318
rect 400218 3295 400274 3304
rect 400232 480 400260 3295
rect 401336 480 401364 7618
rect 401612 3346 401640 37878
rect 402900 29714 402928 52006
rect 403360 49366 403388 52020
rect 403348 49360 403400 49366
rect 403348 49302 403400 49308
rect 404556 48686 404584 52020
rect 405752 48822 405780 52020
rect 406962 52006 407068 52034
rect 408158 52006 408448 52034
rect 409354 52006 409828 52034
rect 410550 52006 411208 52034
rect 405740 48816 405792 48822
rect 405740 48758 405792 48764
rect 406936 48816 406988 48822
rect 406936 48758 406988 48764
rect 404544 48680 404596 48686
rect 404544 48622 404596 48628
rect 405648 48680 405700 48686
rect 405648 48622 405700 48628
rect 402888 29708 402940 29714
rect 402888 29650 402940 29656
rect 404360 26920 404412 26926
rect 404360 26862 404412 26868
rect 404372 3346 404400 26862
rect 405660 15910 405688 48622
rect 406948 35222 406976 48758
rect 406936 35216 406988 35222
rect 406936 35158 406988 35164
rect 405648 15904 405700 15910
rect 405648 15846 405700 15852
rect 406108 6180 406160 6186
rect 406108 6122 406160 6128
rect 401612 3318 402560 3346
rect 404372 3318 404952 3346
rect 402532 480 402560 3318
rect 403716 3120 403768 3126
rect 403716 3062 403768 3068
rect 403728 480 403756 3062
rect 404924 480 404952 3318
rect 406120 480 406148 6122
rect 407040 3369 407068 52006
rect 407212 49088 407264 49094
rect 407212 49030 407264 49036
rect 407224 3482 407252 49030
rect 408420 17270 408448 52006
rect 408500 47592 408552 47598
rect 408500 47534 408552 47540
rect 408408 17264 408460 17270
rect 408408 17206 408460 17212
rect 407224 3454 407344 3482
rect 407026 3360 407082 3369
rect 407026 3295 407082 3304
rect 407316 480 407344 3454
rect 408512 480 408540 47534
rect 409800 36650 409828 52006
rect 409788 36644 409840 36650
rect 409788 36586 409840 36592
rect 408592 29640 408644 29646
rect 408592 29582 408644 29588
rect 408604 12442 408632 29582
rect 408592 12436 408644 12442
rect 408592 12378 408644 12384
rect 409696 12436 409748 12442
rect 409696 12378 409748 12384
rect 409708 480 409736 12378
rect 411180 4078 411208 52006
rect 411732 48482 411760 52020
rect 412928 48822 412956 52020
rect 414124 48822 414152 52020
rect 415228 52006 415334 52034
rect 416530 52006 416728 52034
rect 417726 52006 418108 52034
rect 418922 52006 419488 52034
rect 412916 48816 412968 48822
rect 412916 48758 412968 48764
rect 413928 48816 413980 48822
rect 413928 48758 413980 48764
rect 414112 48816 414164 48822
rect 414112 48758 414164 48764
rect 411720 48476 411772 48482
rect 411720 48418 411772 48424
rect 412548 48476 412600 48482
rect 412548 48418 412600 48424
rect 412560 18630 412588 48418
rect 413940 32502 413968 48758
rect 415228 42090 415256 52006
rect 415308 48816 415360 48822
rect 415308 48758 415360 48764
rect 415216 42084 415268 42090
rect 415216 42026 415268 42032
rect 413928 32496 413980 32502
rect 413928 32438 413980 32444
rect 412640 28348 412692 28354
rect 412640 28290 412692 28296
rect 412548 18624 412600 18630
rect 412548 18566 412600 18572
rect 412652 12442 412680 28290
rect 412640 12436 412692 12442
rect 412640 12378 412692 12384
rect 413284 12436 413336 12442
rect 413284 12378 413336 12384
rect 412088 8968 412140 8974
rect 412088 8910 412140 8916
rect 410892 4072 410944 4078
rect 410892 4014 410944 4020
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 410904 480 410932 4014
rect 412100 480 412128 8910
rect 413296 480 413324 12378
rect 415320 3874 415348 48758
rect 416700 10334 416728 52006
rect 416872 40724 416924 40730
rect 416872 40666 416924 40672
rect 415400 10328 415452 10334
rect 415400 10270 415452 10276
rect 416688 10328 416740 10334
rect 416688 10270 416740 10276
rect 414480 3868 414532 3874
rect 414480 3810 414532 3816
rect 415308 3868 415360 3874
rect 415308 3810 415360 3816
rect 414492 480 414520 3810
rect 415412 898 415440 10270
rect 415412 870 415716 898
rect 415688 480 415716 870
rect 416884 480 416912 40666
rect 418080 3738 418108 52006
rect 419460 40730 419488 52006
rect 420104 48822 420132 52020
rect 421208 48822 421236 52020
rect 420092 48816 420144 48822
rect 420092 48758 420144 48764
rect 420828 48816 420880 48822
rect 420828 48758 420880 48764
rect 421196 48816 421248 48822
rect 421196 48758 421248 48764
rect 422208 48816 422260 48822
rect 422208 48758 422260 48764
rect 419448 40724 419500 40730
rect 419448 40666 419500 40672
rect 420840 39438 420868 48758
rect 420828 39432 420880 39438
rect 420828 39374 420880 39380
rect 419540 24200 419592 24206
rect 419540 24142 419592 24148
rect 419172 5024 419224 5030
rect 419172 4966 419224 4972
rect 417976 3732 418028 3738
rect 417976 3674 418028 3680
rect 418068 3732 418120 3738
rect 418068 3674 418120 3680
rect 417988 480 418016 3674
rect 419184 480 419212 4966
rect 419552 3346 419580 24142
rect 421564 4140 421616 4146
rect 421564 4082 421616 4088
rect 419552 3318 420408 3346
rect 420380 480 420408 3318
rect 421576 480 421604 4082
rect 422220 3602 422248 48758
rect 422404 48346 422432 52020
rect 423508 52006 423614 52034
rect 424810 52006 425008 52034
rect 426006 52006 426388 52034
rect 427202 52006 427768 52034
rect 422392 48340 422444 48346
rect 422392 48282 422444 48288
rect 423508 19990 423536 52006
rect 423588 48340 423640 48346
rect 423588 48282 423640 48288
rect 423496 19984 423548 19990
rect 423496 19926 423548 19932
rect 423600 7614 423628 48282
rect 424980 37942 425008 52006
rect 425060 46232 425112 46238
rect 425060 46174 425112 46180
rect 424968 37936 425020 37942
rect 424968 37878 425020 37884
rect 423680 31068 423732 31074
rect 423680 31010 423732 31016
rect 423588 7608 423640 7614
rect 423588 7550 423640 7556
rect 422760 5296 422812 5302
rect 422760 5238 422812 5244
rect 422208 3596 422260 3602
rect 422208 3538 422260 3544
rect 422772 480 422800 5238
rect 423692 3346 423720 31010
rect 425072 3534 425100 46174
rect 426360 6186 426388 52006
rect 426440 32428 426492 32434
rect 426440 32370 426492 32376
rect 426348 6180 426400 6186
rect 426348 6122 426400 6128
rect 425060 3528 425112 3534
rect 426348 3528 426400 3534
rect 425060 3470 425112 3476
rect 425150 3496 425206 3505
rect 426348 3470 426400 3476
rect 425150 3431 425206 3440
rect 423692 3318 423996 3346
rect 423968 480 423996 3318
rect 425164 480 425192 3431
rect 426360 480 426388 3470
rect 426452 3346 426480 32370
rect 427740 21486 427768 52006
rect 428384 48822 428412 52020
rect 429580 48822 429608 52020
rect 430776 48822 430804 52020
rect 431972 48822 432000 52020
rect 433182 52006 433288 52034
rect 434378 52006 434668 52034
rect 435574 52006 436048 52034
rect 428372 48816 428424 48822
rect 428372 48758 428424 48764
rect 429108 48816 429160 48822
rect 429108 48758 429160 48764
rect 429568 48816 429620 48822
rect 429568 48758 429620 48764
rect 430488 48816 430540 48822
rect 430488 48758 430540 48764
rect 430764 48816 430816 48822
rect 430764 48758 430816 48764
rect 431868 48816 431920 48822
rect 431868 48758 431920 48764
rect 431960 48816 432012 48822
rect 431960 48758 432012 48764
rect 433156 48816 433208 48822
rect 433156 48758 433208 48764
rect 427912 48340 427964 48346
rect 427912 48282 427964 48288
rect 427924 38622 427952 48282
rect 427912 38616 427964 38622
rect 427912 38558 427964 38564
rect 427912 29028 427964 29034
rect 427912 28970 427964 28976
rect 427728 21480 427780 21486
rect 427728 21422 427780 21428
rect 427924 19310 427952 28970
rect 427912 19304 427964 19310
rect 427912 19246 427964 19252
rect 427912 9716 427964 9722
rect 427912 9658 427964 9664
rect 426452 3318 427584 3346
rect 427556 480 427584 3318
rect 427924 2854 427952 9658
rect 429120 3534 429148 48758
rect 430500 8974 430528 48758
rect 430580 33856 430632 33862
rect 430580 33798 430632 33804
rect 430592 9654 430620 33798
rect 431880 22846 431908 48758
rect 431868 22840 431920 22846
rect 431868 22782 431920 22788
rect 430580 9648 430632 9654
rect 430580 9590 430632 9596
rect 430488 8968 430540 8974
rect 430488 8910 430540 8916
rect 429936 5228 429988 5234
rect 429936 5170 429988 5176
rect 429108 3528 429160 3534
rect 429108 3470 429160 3476
rect 427912 2848 427964 2854
rect 427912 2790 427964 2796
rect 428740 2780 428792 2786
rect 428740 2722 428792 2728
rect 428752 480 428780 2722
rect 429948 480 429976 5170
rect 432328 3460 432380 3466
rect 432328 3402 432380 3408
rect 431132 604 431184 610
rect 431132 546 431184 552
rect 431144 480 431172 546
rect 432340 480 432368 3402
rect 433168 3126 433196 48758
rect 433260 47598 433288 52006
rect 433248 47592 433300 47598
rect 433248 47534 433300 47540
rect 433340 35284 433392 35290
rect 433340 35226 433392 35232
rect 433352 7682 433380 35226
rect 434640 24138 434668 52006
rect 434812 48340 434864 48346
rect 434812 48282 434864 48288
rect 434824 38622 434852 48282
rect 434812 38616 434864 38622
rect 434812 38558 434864 38564
rect 434812 29028 434864 29034
rect 434812 28970 434864 28976
rect 434628 24132 434680 24138
rect 434628 24074 434680 24080
rect 434824 19310 434852 28970
rect 434812 19304 434864 19310
rect 434812 19246 434864 19252
rect 434812 9784 434864 9790
rect 434812 9726 434864 9732
rect 434824 9654 434852 9726
rect 434812 9648 434864 9654
rect 434812 9590 434864 9596
rect 433340 7676 433392 7682
rect 433340 7618 433392 7624
rect 434628 7676 434680 7682
rect 434628 7618 434680 7624
rect 433156 3120 433208 3126
rect 433156 3062 433208 3068
rect 433524 2372 433576 2378
rect 433524 2314 433576 2320
rect 433536 480 433564 2314
rect 434640 480 434668 7618
rect 436020 3398 436048 52006
rect 436756 46238 436784 52020
rect 437952 48482 437980 52020
rect 439148 48822 439176 52020
rect 440344 48822 440372 52020
rect 441448 52006 441554 52034
rect 442750 52006 442948 52034
rect 443946 52006 444328 52034
rect 445142 52006 445708 52034
rect 439136 48816 439188 48822
rect 439136 48758 439188 48764
rect 440148 48816 440200 48822
rect 440148 48758 440200 48764
rect 440332 48816 440384 48822
rect 440332 48758 440384 48764
rect 437940 48476 437992 48482
rect 437940 48418 437992 48424
rect 438768 48476 438820 48482
rect 438768 48418 438820 48424
rect 436744 46232 436796 46238
rect 436744 46174 436796 46180
rect 437480 36576 437532 36582
rect 437480 36518 437532 36524
rect 437020 11756 437072 11762
rect 437020 11698 437072 11704
rect 436008 3392 436060 3398
rect 436008 3334 436060 3340
rect 435824 604 435876 610
rect 435824 546 435876 552
rect 435836 480 435864 546
rect 437032 480 437060 11698
rect 437492 3346 437520 36518
rect 438780 25702 438808 48418
rect 438768 25696 438820 25702
rect 438768 25638 438820 25644
rect 439412 3800 439464 3806
rect 439412 3742 439464 3748
rect 437492 3318 438256 3346
rect 438228 480 438256 3318
rect 439424 480 439452 3742
rect 440160 3466 440188 48758
rect 441448 29646 441476 52006
rect 441528 48816 441580 48822
rect 441528 48758 441580 48764
rect 441436 29640 441488 29646
rect 441436 29582 441488 29588
rect 441540 10402 441568 48758
rect 441620 39364 441672 39370
rect 441620 39306 441672 39312
rect 441528 10396 441580 10402
rect 441528 10338 441580 10344
rect 440608 5092 440660 5098
rect 440608 5034 440660 5040
rect 440148 3460 440200 3466
rect 440148 3402 440200 3408
rect 440620 480 440648 5034
rect 441632 3346 441660 39306
rect 441632 3318 441844 3346
rect 441816 480 441844 3318
rect 442920 3194 442948 52006
rect 443184 49020 443236 49026
rect 443184 48962 443236 48968
rect 443092 13116 443144 13122
rect 443092 13058 443144 13064
rect 443104 4146 443132 13058
rect 443092 4140 443144 4146
rect 443092 4082 443144 4088
rect 443196 3482 443224 48962
rect 444300 11762 444328 52006
rect 444380 44872 444432 44878
rect 444380 44814 444432 44820
rect 444288 11756 444340 11762
rect 444288 11698 444340 11704
rect 444196 4140 444248 4146
rect 444196 4082 444248 4088
rect 443012 3454 443224 3482
rect 442908 3188 442960 3194
rect 442908 3130 442960 3136
rect 443012 480 443040 3454
rect 444208 480 444236 4082
rect 444392 3346 444420 44814
rect 445680 27062 445708 52006
rect 446232 48822 446260 52020
rect 447428 48822 447456 52020
rect 448624 48822 448652 52020
rect 446220 48816 446272 48822
rect 446220 48758 446272 48764
rect 447048 48816 447100 48822
rect 447048 48758 447100 48764
rect 447416 48816 447468 48822
rect 447416 48758 447468 48764
rect 448428 48816 448480 48822
rect 448428 48758 448480 48764
rect 448612 48816 448664 48822
rect 448612 48758 448664 48764
rect 449716 48816 449768 48822
rect 449716 48758 449768 48764
rect 445668 27056 445720 27062
rect 445668 26998 445720 27004
rect 447060 4146 447088 48758
rect 448440 13122 448468 48758
rect 448520 38004 448572 38010
rect 448520 37946 448572 37952
rect 448428 13116 448480 13122
rect 448428 13058 448480 13064
rect 447784 4956 447836 4962
rect 447784 4898 447836 4904
rect 447048 4140 447100 4146
rect 447048 4082 447100 4088
rect 446588 3800 446640 3806
rect 446588 3742 446640 3748
rect 444392 3318 445432 3346
rect 445404 480 445432 3318
rect 446600 480 446628 3742
rect 447796 480 447824 4898
rect 448532 3346 448560 37946
rect 449728 28354 449756 48758
rect 449716 28348 449768 28354
rect 449716 28290 449768 28296
rect 449820 3505 449848 52020
rect 451030 52006 451228 52034
rect 452226 52006 452608 52034
rect 453422 52006 453988 52034
rect 454618 52006 455368 52034
rect 449992 49156 450044 49162
rect 449992 49098 450044 49104
rect 449806 3496 449862 3505
rect 449806 3431 449862 3440
rect 450004 3346 450032 49098
rect 451200 44878 451228 52006
rect 451188 44872 451240 44878
rect 451188 44814 451240 44820
rect 452580 31074 452608 52006
rect 452568 31068 452620 31074
rect 452568 31010 452620 31016
rect 451280 26988 451332 26994
rect 451280 26930 451332 26936
rect 451292 3670 451320 26930
rect 451372 4752 451424 4758
rect 451372 4694 451424 4700
rect 451280 3664 451332 3670
rect 451280 3606 451332 3612
rect 448532 3318 449020 3346
rect 450004 3318 450216 3346
rect 448992 480 449020 3318
rect 450188 480 450216 3318
rect 451384 2530 451412 4694
rect 453672 3936 453724 3942
rect 453672 3878 453724 3884
rect 452476 3664 452528 3670
rect 452476 3606 452528 3612
rect 451292 2502 451412 2530
rect 451292 480 451320 2502
rect 452488 480 452516 3606
rect 453684 480 453712 3878
rect 453960 3330 453988 52006
rect 454868 5160 454920 5166
rect 454868 5102 454920 5108
rect 453948 3324 454000 3330
rect 453948 3266 454000 3272
rect 454880 480 454908 5102
rect 455340 5098 455368 52006
rect 455800 48822 455828 52020
rect 456892 49428 456944 49434
rect 456892 49370 456944 49376
rect 455788 48816 455840 48822
rect 455788 48758 455840 48764
rect 456708 48816 456760 48822
rect 456708 48758 456760 48764
rect 456720 32434 456748 48758
rect 456708 32428 456760 32434
rect 456708 32370 456760 32376
rect 455420 25628 455472 25634
rect 455420 25570 455472 25576
rect 455328 5092 455380 5098
rect 455328 5034 455380 5040
rect 455432 610 455460 25570
rect 456904 610 456932 49370
rect 456996 48822 457024 52020
rect 458192 48822 458220 52020
rect 456984 48816 457036 48822
rect 456984 48758 457036 48764
rect 458088 48816 458140 48822
rect 458088 48758 458140 48764
rect 458180 48816 458232 48822
rect 458180 48758 458232 48764
rect 458100 3262 458128 48758
rect 459388 33794 459416 52020
rect 460598 52006 460888 52034
rect 461794 52006 462268 52034
rect 462990 52006 463648 52034
rect 459468 48816 459520 48822
rect 459468 48758 459520 48764
rect 459376 33788 459428 33794
rect 459376 33730 459428 33736
rect 458180 14476 458232 14482
rect 458180 14418 458232 14424
rect 458088 3256 458140 3262
rect 458088 3198 458140 3204
rect 458192 626 458220 14418
rect 459480 4894 459508 48758
rect 459652 28280 459704 28286
rect 459652 28222 459704 28228
rect 459468 4888 459520 4894
rect 459468 4830 459520 4836
rect 455420 604 455472 610
rect 455420 546 455472 552
rect 456064 604 456116 610
rect 456064 546 456116 552
rect 456892 604 456944 610
rect 456892 546 456944 552
rect 457260 604 457312 610
rect 458192 598 458496 626
rect 457260 546 457312 552
rect 456076 480 456104 546
rect 457272 480 457300 546
rect 458468 480 458496 598
rect 459664 480 459692 28222
rect 460860 4010 460888 52006
rect 460940 43444 460992 43450
rect 460940 43386 460992 43392
rect 460756 4004 460808 4010
rect 460756 3946 460808 3952
rect 460848 4004 460900 4010
rect 460848 3946 460900 3952
rect 460768 3890 460796 3946
rect 460768 3862 460888 3890
rect 460860 480 460888 3862
rect 460952 3346 460980 43386
rect 462240 4962 462268 52006
rect 462320 29708 462372 29714
rect 462320 29650 462372 29656
rect 462228 4956 462280 4962
rect 462228 4898 462280 4904
rect 462332 3346 462360 29650
rect 463620 5166 463648 52006
rect 463792 49360 463844 49366
rect 463792 49302 463844 49308
rect 463608 5160 463660 5166
rect 463608 5102 463660 5108
rect 463804 3346 463832 49302
rect 464172 48822 464200 52020
rect 465368 48822 465396 52020
rect 466564 48822 466592 52020
rect 467760 49026 467788 52020
rect 468970 52006 469168 52034
rect 470166 52006 470548 52034
rect 471362 52006 471928 52034
rect 467748 49020 467800 49026
rect 467748 48962 467800 48968
rect 464160 48816 464212 48822
rect 464160 48758 464212 48764
rect 464988 48816 465040 48822
rect 464988 48758 465040 48764
rect 465356 48816 465408 48822
rect 465356 48758 465408 48764
rect 466368 48816 466420 48822
rect 466368 48758 466420 48764
rect 466552 48816 466604 48822
rect 466552 48758 466604 48764
rect 467748 48816 467800 48822
rect 467748 48758 467800 48764
rect 465000 3942 465028 48758
rect 465080 15904 465132 15910
rect 465080 15846 465132 15852
rect 464988 3936 465040 3942
rect 464988 3878 465040 3884
rect 460952 3318 462084 3346
rect 462332 3318 463280 3346
rect 463804 3318 464476 3346
rect 462056 480 462084 3318
rect 463252 480 463280 3318
rect 464448 480 464476 3318
rect 465092 1850 465120 15846
rect 466380 5030 466408 48758
rect 467760 35222 467788 48758
rect 466460 35216 466512 35222
rect 466460 35158 466512 35164
rect 467748 35216 467800 35222
rect 467748 35158 467800 35164
rect 466368 5024 466420 5030
rect 466368 4966 466420 4972
rect 466472 3346 466500 35158
rect 467840 17264 467892 17270
rect 467840 17206 467892 17212
rect 467852 3670 467880 17206
rect 469140 14482 469168 52006
rect 469220 36644 469272 36650
rect 469220 36586 469272 36592
rect 469128 14476 469180 14482
rect 469128 14418 469180 14424
rect 467840 3664 467892 3670
rect 467840 3606 467892 3612
rect 469128 3664 469180 3670
rect 469128 3606 469180 3612
rect 467930 3360 467986 3369
rect 466472 3318 466868 3346
rect 465092 1822 465672 1850
rect 465644 480 465672 1822
rect 466840 480 466868 3318
rect 467930 3295 467986 3304
rect 467944 480 467972 3295
rect 469140 480 469168 3606
rect 469232 3346 469260 36586
rect 470520 36582 470548 52006
rect 470508 36576 470560 36582
rect 470508 36518 470560 36524
rect 471520 4072 471572 4078
rect 471520 4014 471572 4020
rect 469232 3318 470364 3346
rect 470336 480 470364 3318
rect 471532 480 471560 4014
rect 471900 3806 471928 52006
rect 472452 48754 472480 52020
rect 473648 48822 473676 52020
rect 474844 49230 474872 52020
rect 474832 49224 474884 49230
rect 474832 49166 474884 49172
rect 473636 48816 473688 48822
rect 473636 48758 473688 48764
rect 474648 48816 474700 48822
rect 474648 48758 474700 48764
rect 472440 48748 472492 48754
rect 472440 48690 472492 48696
rect 474004 48748 474056 48754
rect 474004 48690 474056 48696
rect 474016 43450 474044 48690
rect 474004 43444 474056 43450
rect 474004 43386 474056 43392
rect 473360 32496 473412 32502
rect 473360 32438 473412 32444
rect 471980 18624 472032 18630
rect 471980 18566 472032 18572
rect 471888 3800 471940 3806
rect 471888 3742 471940 3748
rect 471992 610 472020 18566
rect 473372 610 473400 32438
rect 474660 18630 474688 48758
rect 474648 18624 474700 18630
rect 474648 18566 474700 18572
rect 476040 4826 476068 52020
rect 477236 49706 477264 52020
rect 478446 52006 478828 52034
rect 479642 52006 480208 52034
rect 477224 49700 477276 49706
rect 477224 49642 477276 49648
rect 476120 42084 476172 42090
rect 476120 42026 476172 42032
rect 476028 4820 476080 4826
rect 476028 4762 476080 4768
rect 475108 3868 475160 3874
rect 475108 3810 475160 3816
rect 471980 604 472032 610
rect 471980 546 472032 552
rect 472716 604 472768 610
rect 472716 546 472768 552
rect 473360 604 473412 610
rect 473360 546 473412 552
rect 473912 604 473964 610
rect 473912 546 473964 552
rect 472728 480 472756 546
rect 473924 480 473952 546
rect 475120 480 475148 3810
rect 476132 626 476160 42026
rect 477592 10328 477644 10334
rect 477592 10270 477644 10276
rect 477604 626 477632 10270
rect 478696 3732 478748 3738
rect 478696 3674 478748 3680
rect 476132 598 476344 626
rect 476316 480 476344 598
rect 477512 598 477632 626
rect 477512 480 477540 598
rect 478708 480 478736 3674
rect 478800 3670 478828 52006
rect 478880 40724 478932 40730
rect 478880 40666 478932 40672
rect 478788 3664 478840 3670
rect 478788 3606 478840 3612
rect 478892 610 478920 40666
rect 480180 5370 480208 52006
rect 480824 48822 480852 52020
rect 482020 49162 482048 52020
rect 482284 49700 482336 49706
rect 482284 49642 482336 49648
rect 482008 49156 482060 49162
rect 482008 49098 482060 49104
rect 480812 48816 480864 48822
rect 480812 48758 480864 48764
rect 481548 48816 481600 48822
rect 481548 48758 481600 48764
rect 480260 39432 480312 39438
rect 480260 39374 480312 39380
rect 480168 5364 480220 5370
rect 480168 5306 480220 5312
rect 480272 3482 480300 39374
rect 481560 20058 481588 48758
rect 481548 20052 481600 20058
rect 481548 19994 481600 20000
rect 482296 7682 482324 49642
rect 483216 48822 483244 52020
rect 483204 48816 483256 48822
rect 483204 48758 483256 48764
rect 484308 48816 484360 48822
rect 484308 48758 484360 48764
rect 482284 7676 482336 7682
rect 482284 7618 482336 7624
rect 483480 7608 483532 7614
rect 483480 7550 483532 7556
rect 482284 3596 482336 3602
rect 482284 3538 482336 3544
rect 480272 3454 481128 3482
rect 478880 604 478932 610
rect 478880 546 478932 552
rect 479892 604 479944 610
rect 479892 546 479944 552
rect 479904 480 479932 546
rect 481100 480 481128 3454
rect 482296 480 482324 3538
rect 483492 480 483520 7550
rect 484320 5302 484348 48758
rect 484412 48346 484440 52020
rect 485622 52006 485728 52034
rect 486818 52006 487108 52034
rect 488014 52006 488488 52034
rect 484400 48340 484452 48346
rect 484400 48282 484452 48288
rect 485596 48340 485648 48346
rect 485596 48282 485648 48288
rect 485608 21418 485636 48282
rect 485596 21412 485648 21418
rect 485596 21354 485648 21360
rect 484400 19984 484452 19990
rect 484400 19926 484452 19932
rect 484308 5296 484360 5302
rect 484308 5238 484360 5244
rect 484412 3482 484440 19926
rect 485700 3641 485728 52006
rect 485780 37936 485832 37942
rect 485780 37878 485832 37884
rect 485686 3632 485742 3641
rect 485686 3567 485742 3576
rect 484412 3454 484624 3482
rect 484596 480 484624 3454
rect 485792 480 485820 37878
rect 486976 6180 487028 6186
rect 486976 6122 487028 6128
rect 486988 480 487016 6122
rect 487080 5234 487108 52006
rect 488460 22778 488488 52006
rect 489196 49094 489224 52020
rect 489184 49088 489236 49094
rect 489184 49030 489236 49036
rect 490392 47666 490420 52020
rect 491588 48822 491616 52020
rect 492784 48822 492812 52020
rect 493888 52006 493994 52034
rect 495190 52006 495388 52034
rect 496386 52006 496768 52034
rect 491576 48816 491628 48822
rect 491576 48758 491628 48764
rect 492588 48816 492640 48822
rect 492588 48758 492640 48764
rect 492772 48816 492824 48822
rect 492772 48758 492824 48764
rect 490380 47660 490432 47666
rect 490380 47602 490432 47608
rect 492600 24206 492628 48758
rect 493888 42090 493916 52006
rect 493968 48816 494020 48822
rect 493968 48758 494020 48764
rect 493876 42084 493928 42090
rect 493876 42026 493928 42032
rect 492588 24200 492640 24206
rect 492588 24142 492640 24148
rect 491300 22840 491352 22846
rect 491300 22782 491352 22788
rect 488448 22772 488500 22778
rect 488448 22714 488500 22720
rect 487160 21480 487212 21486
rect 487160 21422 487212 21428
rect 487068 5228 487120 5234
rect 487068 5170 487120 5176
rect 487172 3482 487200 21422
rect 490564 8968 490616 8974
rect 490564 8910 490616 8916
rect 489368 3528 489420 3534
rect 487172 3454 488212 3482
rect 489368 3470 489420 3476
rect 488184 480 488212 3454
rect 489380 480 489408 3470
rect 490576 480 490604 8910
rect 491312 3482 491340 22782
rect 493980 3534 494008 48758
rect 494060 47592 494112 47598
rect 494060 47534 494112 47540
rect 493968 3528 494020 3534
rect 491312 3454 491800 3482
rect 493968 3470 494020 3476
rect 494072 3482 494100 47534
rect 495360 25566 495388 52006
rect 495348 25560 495400 25566
rect 495348 25502 495400 25508
rect 494152 24132 494204 24138
rect 494152 24074 494204 24080
rect 494164 3602 494192 24074
rect 496740 3602 496768 52006
rect 497476 46238 497504 52020
rect 498672 48822 498700 52020
rect 499868 48822 499896 52020
rect 501064 48822 501092 52020
rect 502168 52006 502274 52034
rect 503470 52006 503668 52034
rect 504666 52006 505048 52034
rect 505862 52006 506428 52034
rect 507058 52006 507808 52034
rect 498660 48816 498712 48822
rect 498660 48758 498712 48764
rect 499488 48816 499540 48822
rect 499488 48758 499540 48764
rect 499856 48816 499908 48822
rect 499856 48758 499908 48764
rect 500868 48816 500920 48822
rect 500868 48758 500920 48764
rect 501052 48816 501104 48822
rect 501052 48758 501104 48764
rect 496820 46232 496872 46238
rect 496820 46174 496872 46180
rect 497464 46232 497516 46238
rect 497464 46174 497516 46180
rect 494152 3596 494204 3602
rect 494152 3538 494204 3544
rect 495348 3596 495400 3602
rect 495348 3538 495400 3544
rect 496728 3596 496780 3602
rect 496728 3538 496780 3544
rect 494072 3454 494192 3482
rect 491772 480 491800 3454
rect 492956 3120 493008 3126
rect 492956 3062 493008 3068
rect 492968 480 492996 3062
rect 494164 480 494192 3454
rect 495360 480 495388 3538
rect 496832 3482 496860 46174
rect 498200 25696 498252 25702
rect 498200 25638 498252 25644
rect 498212 3482 498240 25638
rect 499500 8974 499528 48758
rect 499488 8968 499540 8974
rect 499488 8910 499540 8916
rect 500880 3874 500908 48758
rect 502168 26926 502196 52006
rect 502248 48816 502300 48822
rect 502248 48758 502300 48764
rect 502156 26920 502208 26926
rect 502156 26862 502208 26868
rect 500960 10396 501012 10402
rect 500960 10338 501012 10344
rect 500868 3868 500920 3874
rect 500868 3810 500920 3816
rect 496832 3454 497780 3482
rect 498212 3454 498976 3482
rect 496544 3392 496596 3398
rect 496544 3334 496596 3340
rect 496556 480 496584 3334
rect 497752 480 497780 3454
rect 498948 480 498976 3454
rect 500132 3460 500184 3466
rect 500132 3402 500184 3408
rect 500144 480 500172 3402
rect 500972 898 501000 10338
rect 502260 6186 502288 48758
rect 502432 29640 502484 29646
rect 502432 29582 502484 29588
rect 502248 6180 502300 6186
rect 502248 6122 502300 6128
rect 500972 870 501276 898
rect 501248 480 501276 870
rect 502444 480 502472 29582
rect 503640 4078 503668 52006
rect 505020 15910 505048 52006
rect 506400 28286 506428 52006
rect 506388 28280 506440 28286
rect 506388 28222 506440 28228
rect 505100 27056 505152 27062
rect 505100 26998 505152 27004
rect 505008 15904 505060 15910
rect 505008 15846 505060 15852
rect 503720 11756 503772 11762
rect 503720 11698 503772 11704
rect 503628 4072 503680 4078
rect 503628 4014 503680 4020
rect 503732 3346 503760 11698
rect 505112 3346 505140 26998
rect 507780 4146 507808 52006
rect 508240 48822 508268 52020
rect 509436 48822 509464 52020
rect 508228 48816 508280 48822
rect 508228 48758 508280 48764
rect 509148 48816 509200 48822
rect 509148 48758 509200 48764
rect 509424 48816 509476 48822
rect 509424 48758 509476 48764
rect 510528 48816 510580 48822
rect 510528 48758 510580 48764
rect 509160 44946 509188 48758
rect 509148 44940 509200 44946
rect 509148 44882 509200 44888
rect 510540 31142 510568 48758
rect 510632 48550 510660 52020
rect 510620 48544 510672 48550
rect 510620 48486 510672 48492
rect 511828 39370 511856 52020
rect 513038 52006 513328 52034
rect 514234 52006 514708 52034
rect 515430 52006 516088 52034
rect 511908 48544 511960 48550
rect 511908 48486 511960 48492
rect 511816 39364 511868 39370
rect 511816 39306 511868 39312
rect 510528 31136 510580 31142
rect 510528 31078 510580 31084
rect 509240 28348 509292 28354
rect 509240 28290 509292 28296
rect 507860 13116 507912 13122
rect 507860 13058 507912 13064
rect 507216 4140 507268 4146
rect 507216 4082 507268 4088
rect 507768 4140 507820 4146
rect 507768 4082 507820 4088
rect 503732 3318 504864 3346
rect 505112 3318 506060 3346
rect 503628 3188 503680 3194
rect 503628 3130 503680 3136
rect 503640 480 503668 3130
rect 504836 480 504864 3318
rect 506032 480 506060 3318
rect 507228 480 507256 4082
rect 507872 3346 507900 13058
rect 509252 3346 509280 28290
rect 510802 3496 510858 3505
rect 510802 3431 510858 3440
rect 507872 3318 508452 3346
rect 509252 3318 509648 3346
rect 508424 480 508452 3318
rect 509620 480 509648 3318
rect 510816 480 510844 3431
rect 511920 3398 511948 48486
rect 512000 44872 512052 44878
rect 512000 44814 512052 44820
rect 511908 3392 511960 3398
rect 511908 3334 511960 3340
rect 512012 480 512040 44814
rect 512092 31068 512144 31074
rect 512092 31010 512144 31016
rect 512104 3346 512132 31010
rect 513300 3738 513328 52006
rect 513288 3732 513340 3738
rect 513288 3674 513340 3680
rect 512104 3318 513236 3346
rect 514680 3330 514708 52006
rect 516060 10334 516088 52006
rect 516612 48822 516640 52020
rect 517808 48822 517836 52020
rect 519004 48822 519032 52020
rect 516600 48816 516652 48822
rect 516600 48758 516652 48764
rect 517428 48816 517480 48822
rect 517428 48758 517480 48764
rect 517796 48816 517848 48822
rect 517796 48758 517848 48764
rect 518808 48816 518860 48822
rect 518808 48758 518860 48764
rect 518992 48816 519044 48822
rect 518992 48758 519044 48764
rect 520096 48816 520148 48822
rect 520096 48758 520148 48764
rect 516140 32428 516192 32434
rect 516140 32370 516192 32376
rect 516048 10328 516100 10334
rect 516048 10270 516100 10276
rect 515588 5092 515640 5098
rect 515588 5034 515640 5040
rect 513208 480 513236 3318
rect 514392 3324 514444 3330
rect 514392 3266 514444 3272
rect 514668 3324 514720 3330
rect 514668 3266 514720 3272
rect 514404 480 514432 3266
rect 515600 480 515628 5034
rect 516152 3346 516180 32370
rect 517440 3466 517468 48758
rect 517428 3460 517480 3466
rect 517428 3402 517480 3408
rect 516152 3318 516824 3346
rect 516796 480 516824 3318
rect 518820 3262 518848 48758
rect 520108 37942 520136 48758
rect 520096 37936 520148 37942
rect 520096 37878 520148 37884
rect 519084 4888 519136 4894
rect 519084 4830 519136 4836
rect 517888 3256 517940 3262
rect 517888 3198 517940 3204
rect 518808 3256 518860 3262
rect 518808 3198 518860 3204
rect 517900 480 517928 3198
rect 519096 480 519124 4830
rect 520200 3369 520228 52020
rect 521410 52006 521608 52034
rect 520372 33788 520424 33794
rect 520372 33730 520424 33736
rect 520384 3482 520412 33730
rect 521580 4010 521608 52006
rect 523696 41410 523724 85303
rect 523788 77246 523816 111959
rect 523880 111790 523908 138615
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 523868 111784 523920 111790
rect 523868 111726 523920 111732
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 523866 98696 523922 98705
rect 523866 98631 523922 98640
rect 523776 77240 523828 77246
rect 523776 77182 523828 77188
rect 523774 72040 523830 72049
rect 523774 71975 523830 71984
rect 523684 41404 523736 41410
rect 523684 41346 523736 41352
rect 523788 30326 523816 71975
rect 523880 64870 523908 98631
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 523868 64864 523920 64870
rect 523868 64806 523920 64812
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 523866 58712 523922 58721
rect 523866 58647 523922 58656
rect 523776 30320 523828 30326
rect 523776 30262 523828 30268
rect 523880 17950 523908 58647
rect 535460 49224 535512 49230
rect 535460 49166 535512 49172
rect 528560 49020 528612 49026
rect 528560 48962 528612 48968
rect 527180 35216 527232 35222
rect 527180 35158 527232 35164
rect 523868 17944 523920 17950
rect 523868 17886 523920 17892
rect 523868 5160 523920 5166
rect 523868 5102 523920 5108
rect 522672 4956 522724 4962
rect 522672 4898 522724 4904
rect 521476 4004 521528 4010
rect 521476 3946 521528 3952
rect 521568 4004 521620 4010
rect 521568 3946 521620 3952
rect 520292 3454 520412 3482
rect 520186 3360 520242 3369
rect 520186 3295 520242 3304
rect 520292 480 520320 3454
rect 521488 480 521516 3946
rect 522684 480 522712 4898
rect 523880 480 523908 5102
rect 526260 5024 526312 5030
rect 526260 4966 526312 4972
rect 525064 3936 525116 3942
rect 525064 3878 525116 3884
rect 525076 480 525104 3878
rect 526272 480 526300 4966
rect 527192 3346 527220 35158
rect 528572 3482 528600 48962
rect 532700 43444 532752 43450
rect 532700 43386 532752 43392
rect 529940 36576 529992 36582
rect 529940 36518 529992 36524
rect 528652 14476 528704 14482
rect 528652 14418 528704 14424
rect 528664 3806 528692 14418
rect 528652 3800 528704 3806
rect 528652 3742 528704 3748
rect 529848 3800 529900 3806
rect 529848 3742 529900 3748
rect 528572 3454 528692 3482
rect 527192 3318 527496 3346
rect 527468 480 527496 3318
rect 528664 480 528692 3454
rect 529860 480 529888 3742
rect 529952 3482 529980 36518
rect 532712 3482 532740 43386
rect 534080 18624 534132 18630
rect 534080 18566 534132 18572
rect 534092 3482 534120 18566
rect 535472 3482 535500 49166
rect 542360 49156 542412 49162
rect 542360 49098 542412 49104
rect 540980 20052 541032 20058
rect 540980 19994 541032 20000
rect 538128 7676 538180 7682
rect 538128 7618 538180 7624
rect 536932 4820 536984 4826
rect 536932 4762 536984 4768
rect 529952 3454 531084 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 531056 480 531084 3454
rect 532240 3188 532292 3194
rect 532240 3130 532292 3136
rect 532252 480 532280 3130
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 4762
rect 538140 480 538168 7618
rect 540520 5364 540572 5370
rect 540520 5306 540572 5312
rect 539324 3664 539376 3670
rect 539324 3606 539376 3612
rect 539336 480 539364 3606
rect 540532 480 540560 5306
rect 540992 3482 541020 19994
rect 542372 3482 542400 49098
rect 549260 49088 549312 49094
rect 549260 49030 549312 49036
rect 547880 22772 547932 22778
rect 547880 22714 547932 22720
rect 545120 21412 545172 21418
rect 545120 21354 545172 21360
rect 544108 5296 544160 5302
rect 544108 5238 544160 5244
rect 540992 3454 541756 3482
rect 542372 3454 542952 3482
rect 541728 480 541756 3454
rect 542924 480 542952 3454
rect 544120 480 544148 5238
rect 545132 3482 545160 21354
rect 547696 5228 547748 5234
rect 547696 5170 547748 5176
rect 546498 3632 546554 3641
rect 546498 3567 546554 3576
rect 545132 3454 545344 3482
rect 545316 480 545344 3454
rect 546512 480 546540 3567
rect 547708 480 547736 5170
rect 547892 3482 547920 22714
rect 549272 3482 549300 49030
rect 550640 47660 550692 47666
rect 550640 47602 550692 47608
rect 550652 3482 550680 47602
rect 557540 46232 557592 46238
rect 557540 46174 557592 46180
rect 554780 42084 554832 42090
rect 554780 42026 554832 42032
rect 552020 24200 552072 24206
rect 552020 24142 552072 24148
rect 552032 3482 552060 24142
rect 553584 3528 553636 3534
rect 547892 3454 548932 3482
rect 549272 3454 550128 3482
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 553584 3470 553636 3476
rect 548904 480 548932 3454
rect 550100 480 550128 3454
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3470
rect 554792 480 554820 42026
rect 554872 25560 554924 25566
rect 554872 25502 554924 25508
rect 554884 3482 554912 25502
rect 557172 3596 557224 3602
rect 557172 3538 557224 3544
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3538
rect 557552 610 557580 46174
rect 568580 44940 568632 44946
rect 568580 44882 568632 44888
rect 565820 28280 565872 28286
rect 565820 28222 565872 28228
rect 563152 26920 563204 26926
rect 563152 26862 563204 26868
rect 559564 8968 559616 8974
rect 559564 8910 559616 8916
rect 557540 604 557592 610
rect 557540 546 557592 552
rect 558368 604 558420 610
rect 558368 546 558420 552
rect 558380 480 558408 546
rect 559576 480 559604 8910
rect 561956 6180 562008 6186
rect 561956 6122 562008 6128
rect 560760 3868 560812 3874
rect 560760 3810 560812 3816
rect 560772 480 560800 3810
rect 561968 480 561996 6122
rect 563164 480 563192 26862
rect 564440 15904 564492 15910
rect 564440 15846 564492 15852
rect 564348 4072 564400 4078
rect 564348 4014 564400 4020
rect 564360 480 564388 4014
rect 564452 610 564480 15846
rect 565832 610 565860 28222
rect 567844 4140 567896 4146
rect 567844 4082 567896 4088
rect 564440 604 564492 610
rect 564440 546 564492 552
rect 565544 604 565596 610
rect 565544 546 565596 552
rect 565820 604 565872 610
rect 565820 546 565872 552
rect 566740 604 566792 610
rect 566740 546 566792 552
rect 565556 480 565584 546
rect 566752 480 566780 546
rect 567856 480 567884 4082
rect 568592 1306 568620 44882
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 571432 39364 571484 39370
rect 571432 39306 571484 39312
rect 569960 31136 570012 31142
rect 569960 31078 570012 31084
rect 569972 3482 570000 31078
rect 571444 3534 571472 39306
rect 578884 37936 578936 37942
rect 578884 37878 578936 37884
rect 575480 10328 575532 10334
rect 575480 10270 575532 10276
rect 573824 3732 573876 3738
rect 573824 3674 573876 3680
rect 571432 3528 571484 3534
rect 569972 3454 570276 3482
rect 571432 3470 571484 3476
rect 572628 3528 572680 3534
rect 572628 3470 572680 3476
rect 568592 1278 569080 1306
rect 569052 480 569080 1278
rect 570248 480 570276 3454
rect 571432 3392 571484 3398
rect 571432 3334 571484 3340
rect 571444 480 571472 3334
rect 572640 480 572668 3470
rect 573836 480 573864 3674
rect 575492 3482 575520 10270
rect 578896 3534 578924 37878
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 582196 4004 582248 4010
rect 582196 3946 582248 3952
rect 578884 3528 578936 3534
rect 575492 3454 576256 3482
rect 578884 3470 578936 3476
rect 579804 3528 579856 3534
rect 579804 3470 579856 3476
rect 575020 3324 575072 3330
rect 575020 3266 575072 3272
rect 575032 480 575060 3266
rect 576228 480 576256 3454
rect 577412 3460 577464 3466
rect 577412 3402 577464 3408
rect 577424 480 577452 3402
rect 578608 3256 578660 3262
rect 578608 3198 578660 3204
rect 578620 480 578648 3198
rect 579816 480 579844 3470
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 3946
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3606 682216 3662 682272
rect 3422 667936 3478 667992
rect 3514 653520 3570 653576
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 580170 697992 580226 698048
rect 59358 644680 59414 644736
rect 580170 686296 580226 686352
rect 580262 674600 580318 674656
rect 523774 645224 523830 645280
rect 580170 639376 580226 639432
rect 523682 631896 523738 631952
rect 59358 630400 59414 630456
rect 3606 624824 3662 624880
rect 3422 610408 3478 610464
rect 59358 616120 59414 616176
rect 523130 605240 523186 605296
rect 59358 601840 59414 601896
rect 3514 595992 3570 596048
rect 59358 587560 59414 587616
rect 59358 573280 59414 573336
rect 3422 567296 3478 567352
rect 523130 565256 523186 565312
rect 59358 559000 59414 559056
rect 3422 553016 3478 553072
rect 580446 651072 580502 651128
rect 580354 627680 580410 627736
rect 524326 618568 524382 618624
rect 579802 592456 579858 592512
rect 523774 591912 523830 591968
rect 580262 580760 580318 580816
rect 524326 578584 524382 578640
rect 580170 557232 580226 557288
rect 523682 551928 523738 551984
rect 59358 544720 59414 544776
rect 3422 538600 3478 538656
rect 523682 538600 523738 538656
rect 59358 530440 59414 530496
rect 59358 516180 59414 516216
rect 59358 516160 59360 516180
rect 59360 516160 59412 516180
rect 59412 516160 59414 516180
rect 580170 545536 580226 545592
rect 580446 604152 580502 604208
rect 580262 533840 580318 533896
rect 523774 525272 523830 525328
rect 523682 511944 523738 512000
rect 580170 510312 580226 510368
rect 3422 509904 3478 509960
rect 59358 501880 59414 501936
rect 523682 498616 523738 498672
rect 3330 495488 3386 495544
rect 59358 487600 59414 487656
rect 3422 481072 3478 481128
rect 59358 473356 59360 473376
rect 59360 473356 59412 473376
rect 59412 473356 59414 473376
rect 59358 473320 59414 473356
rect 580170 498616 580226 498672
rect 580262 486784 580318 486840
rect 523774 485288 523830 485344
rect 523682 471960 523738 472016
rect 580170 463392 580226 463448
rect 59358 459040 59414 459096
rect 3422 452376 3478 452432
rect 524326 458632 524382 458688
rect 580170 451696 580226 451752
rect 523682 445304 523738 445360
rect 59358 444760 59414 444816
rect 3514 437960 3570 438016
rect 59358 430480 59414 430536
rect 3422 423680 3478 423736
rect 580170 439864 580226 439920
rect 523774 431976 523830 432032
rect 523682 418648 523738 418704
rect 580170 416472 580226 416528
rect 59358 416200 59414 416256
rect 523682 405320 523738 405376
rect 580170 404776 580226 404832
rect 59358 401920 59414 401976
rect 3514 394984 3570 395040
rect 3422 380568 3478 380624
rect 580170 392944 580226 393000
rect 523774 391992 523830 392048
rect 60002 387640 60058 387696
rect 59358 373360 59414 373416
rect 3606 366152 3662 366208
rect 59358 359080 59414 359136
rect 523682 378664 523738 378720
rect 580170 369552 580226 369608
rect 524234 365336 524290 365392
rect 580170 357856 580226 357912
rect 523682 351872 523738 351928
rect 580170 346024 580226 346080
rect 60186 344664 60242 344720
rect 3606 337456 3662 337512
rect 59358 330384 59414 330440
rect 3514 323040 3570 323096
rect 3422 308760 3478 308816
rect 3054 294344 3110 294400
rect 3146 251232 3202 251288
rect 3146 208120 3202 208176
rect 59358 316104 59414 316160
rect 3606 280064 3662 280120
rect 3514 236952 3570 237008
rect 60094 301824 60150 301880
rect 59358 287544 59414 287600
rect 59358 273284 59414 273320
rect 59358 273264 59360 273284
rect 59360 273264 59412 273284
rect 59412 273264 59414 273284
rect 3698 265648 3754 265704
rect 60002 258984 60058 259040
rect 59358 244704 59414 244760
rect 59358 230424 59414 230480
rect 3606 222536 3662 222592
rect 3422 193840 3478 193896
rect 3422 165008 3478 165064
rect 2962 122032 3018 122088
rect 3514 150728 3570 150784
rect 523774 338544 523830 338600
rect 524326 325216 524382 325272
rect 580170 322632 580226 322688
rect 524326 311888 524382 311944
rect 580170 310800 580226 310856
rect 580170 299104 580226 299160
rect 524326 298560 524382 298616
rect 523682 285232 523738 285288
rect 580170 275712 580226 275768
rect 523682 271904 523738 271960
rect 580170 263880 580226 263936
rect 523682 258576 523738 258632
rect 579802 252184 579858 252240
rect 523682 245248 523738 245304
rect 523774 231920 523830 231976
rect 580170 228792 580226 228848
rect 523866 218592 523922 218648
rect 60094 216144 60150 216200
rect 59358 201864 59414 201920
rect 59358 187584 59414 187640
rect 3698 179424 3754 179480
rect 60002 173304 60058 173360
rect 59358 159024 59414 159080
rect 59358 144744 59414 144800
rect 3606 136312 3662 136368
rect 3422 107616 3478 107672
rect 3054 78920 3110 78976
rect 3330 35844 3332 35864
rect 3332 35844 3384 35864
rect 3384 35844 3386 35864
rect 3330 35808 3386 35844
rect 3514 64504 3570 64560
rect 3422 21392 3478 21448
rect 580170 216960 580226 217016
rect 523682 205264 523738 205320
rect 579802 205264 579858 205320
rect 523774 191936 523830 191992
rect 580170 181872 580226 181928
rect 523866 178608 523922 178664
rect 523682 165280 523738 165336
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 523774 151952 523830 152008
rect 60094 130464 60150 130520
rect 59358 116184 59414 116240
rect 59358 101904 59414 101960
rect 3698 93200 3754 93256
rect 60002 87624 60058 87680
rect 59358 73344 59414 73400
rect 59358 59064 59414 59120
rect 3606 50088 3662 50144
rect 523682 125296 523738 125352
rect 523866 138624 523922 138680
rect 523774 111968 523830 112024
rect 523682 85312 523738 85368
rect 3514 7112 3570 7168
rect 85486 3440 85542 3496
rect 92386 3304 92442 3360
rect 146850 3440 146906 3496
rect 153934 3304 153990 3360
rect 339406 3304 339462 3360
rect 364246 3440 364302 3496
rect 400218 3304 400274 3360
rect 407026 3304 407082 3360
rect 425150 3440 425206 3496
rect 449806 3440 449862 3496
rect 467930 3304 467986 3360
rect 485686 3576 485742 3632
rect 510802 3440 510858 3496
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 523866 98640 523922 98696
rect 523774 71984 523830 72040
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 523866 58656 523922 58712
rect 520186 3304 520242 3360
rect 546498 3576 546554 3632
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
rect 580998 3304 581054 3360
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3601 682274 3667 682277
rect -960 682272 3667 682274
rect -960 682216 3606 682272
rect 3662 682216 3667 682272
rect -960 682214 3667 682216
rect -960 682124 480 682214
rect 3601 682211 3667 682214
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3509 653578 3575 653581
rect -960 653576 3575 653578
rect -960 653520 3514 653576
rect 3570 653520 3575 653576
rect -960 653518 3575 653520
rect -960 653428 480 653518
rect 3509 653515 3575 653518
rect 580441 651130 580507 651133
rect 583520 651130 584960 651220
rect 580441 651128 584960 651130
rect 580441 651072 580446 651128
rect 580502 651072 584960 651128
rect 580441 651070 584960 651072
rect 580441 651067 580507 651070
rect 583520 650980 584960 651070
rect 523769 645282 523835 645285
rect 521916 645280 523835 645282
rect 521916 645224 523774 645280
rect 523830 645224 523835 645280
rect 521916 645222 523835 645224
rect 523769 645219 523835 645222
rect 59353 644738 59419 644741
rect 59353 644736 62100 644738
rect 59353 644680 59358 644736
rect 59414 644680 62100 644736
rect 59353 644678 62100 644680
rect 59353 644675 59419 644678
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 523677 631954 523743 631957
rect 521916 631952 523743 631954
rect 521916 631896 523682 631952
rect 523738 631896 523743 631952
rect 521916 631894 523743 631896
rect 523677 631891 523743 631894
rect 59353 630458 59419 630461
rect 59353 630456 62100 630458
rect 59353 630400 59358 630456
rect 59414 630400 62100 630456
rect 59353 630398 62100 630400
rect 59353 630395 59419 630398
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3601 624882 3667 624885
rect -960 624880 3667 624882
rect -960 624824 3606 624880
rect 3662 624824 3667 624880
rect -960 624822 3667 624824
rect -960 624732 480 624822
rect 3601 624819 3667 624822
rect 524321 618626 524387 618629
rect 521916 618624 524387 618626
rect 521916 618568 524326 618624
rect 524382 618568 524387 618624
rect 521916 618566 524387 618568
rect 524321 618563 524387 618566
rect 59353 616178 59419 616181
rect 59353 616176 62100 616178
rect 59353 616120 59358 616176
rect 59414 616120 62100 616176
rect 59353 616118 62100 616120
rect 59353 616115 59419 616118
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 523125 605298 523191 605301
rect 521916 605296 523191 605298
rect 521916 605240 523130 605296
rect 523186 605240 523191 605296
rect 521916 605238 523191 605240
rect 523125 605235 523191 605238
rect 580441 604210 580507 604213
rect 583520 604210 584960 604300
rect 580441 604208 584960 604210
rect 580441 604152 580446 604208
rect 580502 604152 584960 604208
rect 580441 604150 584960 604152
rect 580441 604147 580507 604150
rect 583520 604060 584960 604150
rect 59353 601898 59419 601901
rect 59353 601896 62100 601898
rect 59353 601840 59358 601896
rect 59414 601840 62100 601896
rect 59353 601838 62100 601840
rect 59353 601835 59419 601838
rect -960 596050 480 596140
rect 3509 596050 3575 596053
rect -960 596048 3575 596050
rect -960 595992 3514 596048
rect 3570 595992 3575 596048
rect -960 595990 3575 595992
rect -960 595900 480 595990
rect 3509 595987 3575 595990
rect 579797 592514 579863 592517
rect 583520 592514 584960 592604
rect 579797 592512 584960 592514
rect 579797 592456 579802 592512
rect 579858 592456 584960 592512
rect 579797 592454 584960 592456
rect 579797 592451 579863 592454
rect 583520 592364 584960 592454
rect 523769 591970 523835 591973
rect 521916 591968 523835 591970
rect 521916 591912 523774 591968
rect 523830 591912 523835 591968
rect 521916 591910 523835 591912
rect 523769 591907 523835 591910
rect 59353 587618 59419 587621
rect 59353 587616 62100 587618
rect 59353 587560 59358 587616
rect 59414 587560 62100 587616
rect 59353 587558 62100 587560
rect 59353 587555 59419 587558
rect -960 581620 480 581860
rect 580257 580818 580323 580821
rect 583520 580818 584960 580908
rect 580257 580816 584960 580818
rect 580257 580760 580262 580816
rect 580318 580760 584960 580816
rect 580257 580758 584960 580760
rect 580257 580755 580323 580758
rect 583520 580668 584960 580758
rect 524321 578642 524387 578645
rect 521916 578640 524387 578642
rect 521916 578584 524326 578640
rect 524382 578584 524387 578640
rect 521916 578582 524387 578584
rect 524321 578579 524387 578582
rect 59353 573338 59419 573341
rect 59353 573336 62100 573338
rect 59353 573280 59358 573336
rect 59414 573280 62100 573336
rect 59353 573278 62100 573280
rect 59353 573275 59419 573278
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 523125 565314 523191 565317
rect 521916 565312 523191 565314
rect 521916 565256 523130 565312
rect 523186 565256 523191 565312
rect 521916 565254 523191 565256
rect 523125 565251 523191 565254
rect 59353 559058 59419 559061
rect 59353 559056 62100 559058
rect 59353 559000 59358 559056
rect 59414 559000 62100 559056
rect 59353 558998 62100 559000
rect 59353 558995 59419 558998
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3417 553074 3483 553077
rect -960 553072 3483 553074
rect -960 553016 3422 553072
rect 3478 553016 3483 553072
rect -960 553014 3483 553016
rect -960 552924 480 553014
rect 3417 553011 3483 553014
rect 523677 551986 523743 551989
rect 521916 551984 523743 551986
rect 521916 551928 523682 551984
rect 523738 551928 523743 551984
rect 521916 551926 523743 551928
rect 523677 551923 523743 551926
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 59353 544778 59419 544781
rect 59353 544776 62100 544778
rect 59353 544720 59358 544776
rect 59414 544720 62100 544776
rect 59353 544718 62100 544720
rect 59353 544715 59419 544718
rect -960 538658 480 538748
rect 3417 538658 3483 538661
rect 523677 538658 523743 538661
rect -960 538656 3483 538658
rect -960 538600 3422 538656
rect 3478 538600 3483 538656
rect -960 538598 3483 538600
rect 521916 538656 523743 538658
rect 521916 538600 523682 538656
rect 523738 538600 523743 538656
rect 521916 538598 523743 538600
rect -960 538508 480 538598
rect 3417 538595 3483 538598
rect 523677 538595 523743 538598
rect 580257 533898 580323 533901
rect 583520 533898 584960 533988
rect 580257 533896 584960 533898
rect 580257 533840 580262 533896
rect 580318 533840 584960 533896
rect 580257 533838 584960 533840
rect 580257 533835 580323 533838
rect 583520 533748 584960 533838
rect 59353 530498 59419 530501
rect 59353 530496 62100 530498
rect 59353 530440 59358 530496
rect 59414 530440 62100 530496
rect 59353 530438 62100 530440
rect 59353 530435 59419 530438
rect 523769 525330 523835 525333
rect 521916 525328 523835 525330
rect 521916 525272 523774 525328
rect 523830 525272 523835 525328
rect 521916 525270 523835 525272
rect 523769 525267 523835 525270
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 59353 516218 59419 516221
rect 59353 516216 62100 516218
rect 59353 516160 59358 516216
rect 59414 516160 62100 516216
rect 59353 516158 62100 516160
rect 59353 516155 59419 516158
rect 523677 512002 523743 512005
rect 521916 512000 523743 512002
rect 521916 511944 523682 512000
rect 523738 511944 523743 512000
rect 521916 511942 523743 511944
rect 523677 511939 523743 511942
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3417 509962 3483 509965
rect -960 509960 3483 509962
rect -960 509904 3422 509960
rect 3478 509904 3483 509960
rect -960 509902 3483 509904
rect -960 509812 480 509902
rect 3417 509899 3483 509902
rect 59353 501938 59419 501941
rect 59353 501936 62100 501938
rect 59353 501880 59358 501936
rect 59414 501880 62100 501936
rect 59353 501878 62100 501880
rect 59353 501875 59419 501878
rect 523677 498674 523743 498677
rect 521916 498672 523743 498674
rect 521916 498616 523682 498672
rect 523738 498616 523743 498672
rect 521916 498614 523743 498616
rect 523677 498611 523743 498614
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 59353 487658 59419 487661
rect 59353 487656 62100 487658
rect 59353 487600 59358 487656
rect 59414 487600 62100 487656
rect 59353 487598 62100 487600
rect 59353 487595 59419 487598
rect 580257 486842 580323 486845
rect 583520 486842 584960 486932
rect 580257 486840 584960 486842
rect 580257 486784 580262 486840
rect 580318 486784 584960 486840
rect 580257 486782 584960 486784
rect 580257 486779 580323 486782
rect 583520 486692 584960 486782
rect 523769 485346 523835 485349
rect 521916 485344 523835 485346
rect 521916 485288 523774 485344
rect 523830 485288 523835 485344
rect 521916 485286 523835 485288
rect 523769 485283 523835 485286
rect -960 481130 480 481220
rect 3417 481130 3483 481133
rect -960 481128 3483 481130
rect -960 481072 3422 481128
rect 3478 481072 3483 481128
rect -960 481070 3483 481072
rect -960 480980 480 481070
rect 3417 481067 3483 481070
rect 583520 474996 584960 475236
rect 59353 473378 59419 473381
rect 59353 473376 62100 473378
rect 59353 473320 59358 473376
rect 59414 473320 62100 473376
rect 59353 473318 62100 473320
rect 59353 473315 59419 473318
rect 523677 472018 523743 472021
rect 521916 472016 523743 472018
rect 521916 471960 523682 472016
rect 523738 471960 523743 472016
rect 521916 471958 523743 471960
rect 523677 471955 523743 471958
rect -960 466700 480 466940
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 59353 459098 59419 459101
rect 59353 459096 62100 459098
rect 59353 459040 59358 459096
rect 59414 459040 62100 459096
rect 59353 459038 62100 459040
rect 59353 459035 59419 459038
rect 524321 458690 524387 458693
rect 521916 458688 524387 458690
rect 521916 458632 524326 458688
rect 524382 458632 524387 458688
rect 521916 458630 524387 458632
rect 524321 458627 524387 458630
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 523677 445362 523743 445365
rect 521916 445360 523743 445362
rect 521916 445304 523682 445360
rect 523738 445304 523743 445360
rect 521916 445302 523743 445304
rect 523677 445299 523743 445302
rect 59353 444818 59419 444821
rect 59353 444816 62100 444818
rect 59353 444760 59358 444816
rect 59414 444760 62100 444816
rect 59353 444758 62100 444760
rect 59353 444755 59419 444758
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3509 438018 3575 438021
rect -960 438016 3575 438018
rect -960 437960 3514 438016
rect 3570 437960 3575 438016
rect -960 437958 3575 437960
rect -960 437868 480 437958
rect 3509 437955 3575 437958
rect 523769 432034 523835 432037
rect 521916 432032 523835 432034
rect 521916 431976 523774 432032
rect 523830 431976 523835 432032
rect 521916 431974 523835 431976
rect 523769 431971 523835 431974
rect 59353 430538 59419 430541
rect 59353 430536 62100 430538
rect 59353 430480 59358 430536
rect 59414 430480 62100 430536
rect 59353 430478 62100 430480
rect 59353 430475 59419 430478
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3417 423738 3483 423741
rect -960 423736 3483 423738
rect -960 423680 3422 423736
rect 3478 423680 3483 423736
rect -960 423678 3483 423680
rect -960 423588 480 423678
rect 3417 423675 3483 423678
rect 523677 418706 523743 418709
rect 521916 418704 523743 418706
rect 521916 418648 523682 418704
rect 523738 418648 523743 418704
rect 521916 418646 523743 418648
rect 523677 418643 523743 418646
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 59353 416258 59419 416261
rect 59353 416256 62100 416258
rect 59353 416200 59358 416256
rect 59414 416200 62100 416256
rect 59353 416198 62100 416200
rect 59353 416195 59419 416198
rect -960 409172 480 409412
rect 523677 405378 523743 405381
rect 521916 405376 523743 405378
rect 521916 405320 523682 405376
rect 523738 405320 523743 405376
rect 521916 405318 523743 405320
rect 523677 405315 523743 405318
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 59353 401978 59419 401981
rect 59353 401976 62100 401978
rect 59353 401920 59358 401976
rect 59414 401920 62100 401976
rect 59353 401918 62100 401920
rect 59353 401915 59419 401918
rect -960 395042 480 395132
rect 3509 395042 3575 395045
rect -960 395040 3575 395042
rect -960 394984 3514 395040
rect 3570 394984 3575 395040
rect -960 394982 3575 394984
rect -960 394892 480 394982
rect 3509 394979 3575 394982
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 523769 392050 523835 392053
rect 521916 392048 523835 392050
rect 521916 391992 523774 392048
rect 523830 391992 523835 392048
rect 521916 391990 523835 391992
rect 523769 391987 523835 391990
rect 59997 387698 60063 387701
rect 59997 387696 62100 387698
rect 59997 387640 60002 387696
rect 60058 387640 62100 387696
rect 59997 387638 62100 387640
rect 59997 387635 60063 387638
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3417 380626 3483 380629
rect -960 380624 3483 380626
rect -960 380568 3422 380624
rect 3478 380568 3483 380624
rect -960 380566 3483 380568
rect -960 380476 480 380566
rect 3417 380563 3483 380566
rect 523677 378722 523743 378725
rect 521916 378720 523743 378722
rect 521916 378664 523682 378720
rect 523738 378664 523743 378720
rect 521916 378662 523743 378664
rect 523677 378659 523743 378662
rect 59353 373418 59419 373421
rect 59353 373416 62100 373418
rect 59353 373360 59358 373416
rect 59414 373360 62100 373416
rect 59353 373358 62100 373360
rect 59353 373355 59419 373358
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3601 366210 3667 366213
rect -960 366208 3667 366210
rect -960 366152 3606 366208
rect 3662 366152 3667 366208
rect -960 366150 3667 366152
rect -960 366060 480 366150
rect 3601 366147 3667 366150
rect 524229 365394 524295 365397
rect 521916 365392 524295 365394
rect 521916 365336 524234 365392
rect 524290 365336 524295 365392
rect 521916 365334 524295 365336
rect 524229 365331 524295 365334
rect 59353 359138 59419 359141
rect 59353 359136 62100 359138
rect 59353 359080 59358 359136
rect 59414 359080 62100 359136
rect 59353 359078 62100 359080
rect 59353 359075 59419 359078
rect 580165 357914 580231 357917
rect 583520 357914 584960 358004
rect 580165 357912 584960 357914
rect 580165 357856 580170 357912
rect 580226 357856 584960 357912
rect 580165 357854 584960 357856
rect 580165 357851 580231 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 523677 351930 523743 351933
rect 521916 351928 523743 351930
rect 521916 351872 523682 351928
rect 523738 351872 523743 351928
rect 521916 351870 523743 351872
rect 523677 351867 523743 351870
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 60181 344722 60247 344725
rect 60181 344720 62100 344722
rect 60181 344664 60186 344720
rect 60242 344664 62100 344720
rect 60181 344662 62100 344664
rect 60181 344659 60247 344662
rect 523769 338602 523835 338605
rect 521916 338600 523835 338602
rect 521916 338544 523774 338600
rect 523830 338544 523835 338600
rect 521916 338542 523835 338544
rect 523769 338539 523835 338542
rect -960 337514 480 337604
rect 3601 337514 3667 337517
rect -960 337512 3667 337514
rect -960 337456 3606 337512
rect 3662 337456 3667 337512
rect -960 337454 3667 337456
rect -960 337364 480 337454
rect 3601 337451 3667 337454
rect 583520 334236 584960 334476
rect 59353 330442 59419 330445
rect 59353 330440 62100 330442
rect 59353 330384 59358 330440
rect 59414 330384 62100 330440
rect 59353 330382 62100 330384
rect 59353 330379 59419 330382
rect 524321 325274 524387 325277
rect 521916 325272 524387 325274
rect 521916 325216 524326 325272
rect 524382 325216 524387 325272
rect 521916 325214 524387 325216
rect 524321 325211 524387 325214
rect -960 323098 480 323188
rect 3509 323098 3575 323101
rect -960 323096 3575 323098
rect -960 323040 3514 323096
rect 3570 323040 3575 323096
rect -960 323038 3575 323040
rect -960 322948 480 323038
rect 3509 323035 3575 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 59353 316162 59419 316165
rect 59353 316160 62100 316162
rect 59353 316104 59358 316160
rect 59414 316104 62100 316160
rect 59353 316102 62100 316104
rect 59353 316099 59419 316102
rect 524321 311946 524387 311949
rect 521916 311944 524387 311946
rect 521916 311888 524326 311944
rect 524382 311888 524387 311944
rect 521916 311886 524387 311888
rect 524321 311883 524387 311886
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3417 308818 3483 308821
rect -960 308816 3483 308818
rect -960 308760 3422 308816
rect 3478 308760 3483 308816
rect -960 308758 3483 308760
rect -960 308668 480 308758
rect 3417 308755 3483 308758
rect 60089 301882 60155 301885
rect 60089 301880 62100 301882
rect 60089 301824 60094 301880
rect 60150 301824 62100 301880
rect 60089 301822 62100 301824
rect 60089 301819 60155 301822
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect 524321 298618 524387 298621
rect 521916 298616 524387 298618
rect 521916 298560 524326 298616
rect 524382 298560 524387 298616
rect 521916 298558 524387 298560
rect 524321 298555 524387 298558
rect -960 294402 480 294492
rect 3049 294402 3115 294405
rect -960 294400 3115 294402
rect -960 294344 3054 294400
rect 3110 294344 3115 294400
rect -960 294342 3115 294344
rect -960 294252 480 294342
rect 3049 294339 3115 294342
rect 59353 287602 59419 287605
rect 59353 287600 62100 287602
rect 59353 287544 59358 287600
rect 59414 287544 62100 287600
rect 59353 287542 62100 287544
rect 59353 287539 59419 287542
rect 583520 287316 584960 287556
rect 523677 285290 523743 285293
rect 521916 285288 523743 285290
rect 521916 285232 523682 285288
rect 523738 285232 523743 285288
rect 521916 285230 523743 285232
rect 523677 285227 523743 285230
rect -960 280122 480 280212
rect 3601 280122 3667 280125
rect -960 280120 3667 280122
rect -960 280064 3606 280120
rect 3662 280064 3667 280120
rect -960 280062 3667 280064
rect -960 279972 480 280062
rect 3601 280059 3667 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 59353 273322 59419 273325
rect 59353 273320 62100 273322
rect 59353 273264 59358 273320
rect 59414 273264 62100 273320
rect 59353 273262 62100 273264
rect 59353 273259 59419 273262
rect 523677 271962 523743 271965
rect 521916 271960 523743 271962
rect 521916 271904 523682 271960
rect 523738 271904 523743 271960
rect 521916 271902 523743 271904
rect 523677 271899 523743 271902
rect -960 265706 480 265796
rect 3693 265706 3759 265709
rect -960 265704 3759 265706
rect -960 265648 3698 265704
rect 3754 265648 3759 265704
rect -960 265646 3759 265648
rect -960 265556 480 265646
rect 3693 265643 3759 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 59997 259042 60063 259045
rect 59997 259040 62100 259042
rect 59997 258984 60002 259040
rect 60058 258984 62100 259040
rect 59997 258982 62100 258984
rect 59997 258979 60063 258982
rect 523677 258634 523743 258637
rect 521916 258632 523743 258634
rect 521916 258576 523682 258632
rect 523738 258576 523743 258632
rect 521916 258574 523743 258576
rect 523677 258571 523743 258574
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 523677 245306 523743 245309
rect 521916 245304 523743 245306
rect 521916 245248 523682 245304
rect 523738 245248 523743 245304
rect 521916 245246 523743 245248
rect 523677 245243 523743 245246
rect 59353 244762 59419 244765
rect 59353 244760 62100 244762
rect 59353 244704 59358 244760
rect 59414 244704 62100 244760
rect 59353 244702 62100 244704
rect 59353 244699 59419 244702
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3509 237010 3575 237013
rect -960 237008 3575 237010
rect -960 236952 3514 237008
rect 3570 236952 3575 237008
rect -960 236950 3575 236952
rect -960 236860 480 236950
rect 3509 236947 3575 236950
rect 523769 231978 523835 231981
rect 521916 231976 523835 231978
rect 521916 231920 523774 231976
rect 523830 231920 523835 231976
rect 521916 231918 523835 231920
rect 523769 231915 523835 231918
rect 59353 230482 59419 230485
rect 59353 230480 62100 230482
rect 59353 230424 59358 230480
rect 59414 230424 62100 230480
rect 59353 230422 62100 230424
rect 59353 230419 59419 230422
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3601 222594 3667 222597
rect -960 222592 3667 222594
rect -960 222536 3606 222592
rect 3662 222536 3667 222592
rect -960 222534 3667 222536
rect -960 222444 480 222534
rect 3601 222531 3667 222534
rect 523861 218650 523927 218653
rect 521916 218648 523927 218650
rect 521916 218592 523866 218648
rect 523922 218592 523927 218648
rect 521916 218590 523927 218592
rect 523861 218587 523927 218590
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 60089 216202 60155 216205
rect 60089 216200 62100 216202
rect 60089 216144 60094 216200
rect 60150 216144 62100 216200
rect 60089 216142 62100 216144
rect 60089 216139 60155 216142
rect -960 208178 480 208268
rect 3141 208178 3207 208181
rect -960 208176 3207 208178
rect -960 208120 3146 208176
rect 3202 208120 3207 208176
rect -960 208118 3207 208120
rect -960 208028 480 208118
rect 3141 208115 3207 208118
rect 523677 205322 523743 205325
rect 521916 205320 523743 205322
rect 521916 205264 523682 205320
rect 523738 205264 523743 205320
rect 521916 205262 523743 205264
rect 523677 205259 523743 205262
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 59353 201922 59419 201925
rect 59353 201920 62100 201922
rect 59353 201864 59358 201920
rect 59414 201864 62100 201920
rect 59353 201862 62100 201864
rect 59353 201859 59419 201862
rect -960 193898 480 193988
rect 3417 193898 3483 193901
rect -960 193896 3483 193898
rect -960 193840 3422 193896
rect 3478 193840 3483 193896
rect -960 193838 3483 193840
rect -960 193748 480 193838
rect 3417 193835 3483 193838
rect 583520 193476 584960 193716
rect 523769 191994 523835 191997
rect 521916 191992 523835 191994
rect 521916 191936 523774 191992
rect 523830 191936 523835 191992
rect 521916 191934 523835 191936
rect 523769 191931 523835 191934
rect 59353 187642 59419 187645
rect 59353 187640 62100 187642
rect 59353 187584 59358 187640
rect 59414 187584 62100 187640
rect 59353 187582 62100 187584
rect 59353 187579 59419 187582
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3693 179482 3759 179485
rect -960 179480 3759 179482
rect -960 179424 3698 179480
rect 3754 179424 3759 179480
rect -960 179422 3759 179424
rect -960 179332 480 179422
rect 3693 179419 3759 179422
rect 523861 178666 523927 178669
rect 521916 178664 523927 178666
rect 521916 178608 523866 178664
rect 523922 178608 523927 178664
rect 521916 178606 523927 178608
rect 523861 178603 523927 178606
rect 59997 173362 60063 173365
rect 59997 173360 62100 173362
rect 59997 173304 60002 173360
rect 60058 173304 62100 173360
rect 59997 173302 62100 173304
rect 59997 173299 60063 173302
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 523677 165338 523743 165341
rect 521916 165336 523743 165338
rect 521916 165280 523682 165336
rect 523738 165280 523743 165336
rect 521916 165278 523743 165280
rect 523677 165275 523743 165278
rect -960 165066 480 165156
rect 3417 165066 3483 165069
rect -960 165064 3483 165066
rect -960 165008 3422 165064
rect 3478 165008 3483 165064
rect -960 165006 3483 165008
rect -960 164916 480 165006
rect 3417 165003 3483 165006
rect 59353 159082 59419 159085
rect 59353 159080 62100 159082
rect 59353 159024 59358 159080
rect 59414 159024 62100 159080
rect 59353 159022 62100 159024
rect 59353 159019 59419 159022
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 523769 152010 523835 152013
rect 521916 152008 523835 152010
rect 521916 151952 523774 152008
rect 523830 151952 523835 152008
rect 521916 151950 523835 151952
rect 523769 151947 523835 151950
rect -960 150786 480 150876
rect 3509 150786 3575 150789
rect -960 150784 3575 150786
rect -960 150728 3514 150784
rect 3570 150728 3575 150784
rect -960 150726 3575 150728
rect -960 150636 480 150726
rect 3509 150723 3575 150726
rect 583520 146556 584960 146796
rect 59353 144802 59419 144805
rect 59353 144800 62100 144802
rect 59353 144744 59358 144800
rect 59414 144744 62100 144800
rect 59353 144742 62100 144744
rect 59353 144739 59419 144742
rect 523861 138682 523927 138685
rect 521916 138680 523927 138682
rect 521916 138624 523866 138680
rect 523922 138624 523927 138680
rect 521916 138622 523927 138624
rect 523861 138619 523927 138622
rect -960 136370 480 136460
rect 3601 136370 3667 136373
rect -960 136368 3667 136370
rect -960 136312 3606 136368
rect 3662 136312 3667 136368
rect -960 136310 3667 136312
rect -960 136220 480 136310
rect 3601 136307 3667 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 60089 130522 60155 130525
rect 60089 130520 62100 130522
rect 60089 130464 60094 130520
rect 60150 130464 62100 130520
rect 60089 130462 62100 130464
rect 60089 130459 60155 130462
rect 523677 125354 523743 125357
rect 521916 125352 523743 125354
rect 521916 125296 523682 125352
rect 523738 125296 523743 125352
rect 521916 125294 523743 125296
rect 523677 125291 523743 125294
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2957 122090 3023 122093
rect -960 122088 3023 122090
rect -960 122032 2962 122088
rect 3018 122032 3023 122088
rect -960 122030 3023 122032
rect -960 121940 480 122030
rect 2957 122027 3023 122030
rect 59353 116242 59419 116245
rect 59353 116240 62100 116242
rect 59353 116184 59358 116240
rect 59414 116184 62100 116240
rect 59353 116182 62100 116184
rect 59353 116179 59419 116182
rect 523769 112026 523835 112029
rect 521916 112024 523835 112026
rect 521916 111968 523774 112024
rect 523830 111968 523835 112024
rect 521916 111966 523835 111968
rect 523769 111963 523835 111966
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3417 107674 3483 107677
rect -960 107672 3483 107674
rect -960 107616 3422 107672
rect 3478 107616 3483 107672
rect -960 107614 3483 107616
rect -960 107524 480 107614
rect 3417 107611 3483 107614
rect 59353 101962 59419 101965
rect 59353 101960 62100 101962
rect 59353 101904 59358 101960
rect 59414 101904 62100 101960
rect 59353 101902 62100 101904
rect 59353 101899 59419 101902
rect 583520 99636 584960 99876
rect 523861 98698 523927 98701
rect 521916 98696 523927 98698
rect 521916 98640 523866 98696
rect 523922 98640 523927 98696
rect 521916 98638 523927 98640
rect 523861 98635 523927 98638
rect -960 93258 480 93348
rect 3693 93258 3759 93261
rect -960 93256 3759 93258
rect -960 93200 3698 93256
rect 3754 93200 3759 93256
rect -960 93198 3759 93200
rect -960 93108 480 93198
rect 3693 93195 3759 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 59997 87682 60063 87685
rect 59997 87680 62100 87682
rect 59997 87624 60002 87680
rect 60058 87624 62100 87680
rect 59997 87622 62100 87624
rect 59997 87619 60063 87622
rect 523677 85370 523743 85373
rect 521916 85368 523743 85370
rect 521916 85312 523682 85368
rect 523738 85312 523743 85368
rect 521916 85310 523743 85312
rect 523677 85307 523743 85310
rect -960 78978 480 79068
rect 3049 78978 3115 78981
rect -960 78976 3115 78978
rect -960 78920 3054 78976
rect 3110 78920 3115 78976
rect -960 78918 3115 78920
rect -960 78828 480 78918
rect 3049 78915 3115 78918
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 59353 73402 59419 73405
rect 59353 73400 62100 73402
rect 59353 73344 59358 73400
rect 59414 73344 62100 73400
rect 59353 73342 62100 73344
rect 59353 73339 59419 73342
rect 523769 72042 523835 72045
rect 521916 72040 523835 72042
rect 521916 71984 523774 72040
rect 523830 71984 523835 72040
rect 521916 71982 523835 71984
rect 523769 71979 523835 71982
rect -960 64562 480 64652
rect 3509 64562 3575 64565
rect -960 64560 3575 64562
rect -960 64504 3514 64560
rect 3570 64504 3575 64560
rect -960 64502 3575 64504
rect -960 64412 480 64502
rect 3509 64499 3575 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 59353 59122 59419 59125
rect 59353 59120 62100 59122
rect 59353 59064 59358 59120
rect 59414 59064 62100 59120
rect 59353 59062 62100 59064
rect 59353 59059 59419 59062
rect 523861 58714 523927 58717
rect 521916 58712 523927 58714
rect 521916 58656 523866 58712
rect 523922 58656 523927 58712
rect 521916 58654 523927 58656
rect 523861 58651 523927 58654
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3601 50146 3667 50149
rect -960 50144 3667 50146
rect -960 50088 3606 50144
rect 3662 50088 3667 50144
rect -960 50086 3667 50088
rect -960 49996 480 50086
rect 3601 50083 3667 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3325 35866 3391 35869
rect -960 35864 3391 35866
rect -960 35808 3330 35864
rect 3386 35808 3391 35864
rect -960 35806 3391 35808
rect -960 35716 480 35806
rect 3325 35803 3391 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3417 21450 3483 21453
rect -960 21448 3483 21450
rect -960 21392 3422 21448
rect 3478 21392 3483 21448
rect -960 21390 3483 21392
rect -960 21300 480 21390
rect 3417 21387 3483 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3509 7170 3575 7173
rect -960 7168 3575 7170
rect -960 7112 3514 7168
rect 3570 7112 3575 7168
rect -960 7110 3575 7112
rect -960 7020 480 7110
rect 3509 7107 3575 7110
rect 583520 5796 584960 6036
rect 485681 3634 485747 3637
rect 546493 3634 546559 3637
rect 485681 3632 546559 3634
rect 485681 3576 485686 3632
rect 485742 3576 546498 3632
rect 546554 3576 546559 3632
rect 485681 3574 546559 3576
rect 485681 3571 485747 3574
rect 546493 3571 546559 3574
rect 85481 3498 85547 3501
rect 146845 3498 146911 3501
rect 85481 3496 146911 3498
rect 85481 3440 85486 3496
rect 85542 3440 146850 3496
rect 146906 3440 146911 3496
rect 85481 3438 146911 3440
rect 85481 3435 85547 3438
rect 146845 3435 146911 3438
rect 364241 3498 364307 3501
rect 425145 3498 425211 3501
rect 364241 3496 425211 3498
rect 364241 3440 364246 3496
rect 364302 3440 425150 3496
rect 425206 3440 425211 3496
rect 364241 3438 425211 3440
rect 364241 3435 364307 3438
rect 425145 3435 425211 3438
rect 449801 3498 449867 3501
rect 510797 3498 510863 3501
rect 449801 3496 510863 3498
rect 449801 3440 449806 3496
rect 449862 3440 510802 3496
rect 510858 3440 510863 3496
rect 449801 3438 510863 3440
rect 449801 3435 449867 3438
rect 510797 3435 510863 3438
rect 92381 3362 92447 3365
rect 153929 3362 153995 3365
rect 92381 3360 153995 3362
rect 92381 3304 92386 3360
rect 92442 3304 153934 3360
rect 153990 3304 153995 3360
rect 92381 3302 153995 3304
rect 92381 3299 92447 3302
rect 153929 3299 153995 3302
rect 339401 3362 339467 3365
rect 400213 3362 400279 3365
rect 339401 3360 400279 3362
rect 339401 3304 339406 3360
rect 339462 3304 400218 3360
rect 400274 3304 400279 3360
rect 339401 3302 400279 3304
rect 339401 3299 339467 3302
rect 400213 3299 400279 3302
rect 407021 3362 407087 3365
rect 467925 3362 467991 3365
rect 407021 3360 467991 3362
rect 407021 3304 407026 3360
rect 407082 3304 467930 3360
rect 467986 3304 467991 3360
rect 407021 3302 467991 3304
rect 407021 3299 407087 3302
rect 467925 3299 467991 3302
rect 520181 3362 520247 3365
rect 580993 3362 581059 3365
rect 520181 3360 581059 3362
rect 520181 3304 520186 3360
rect 520242 3304 580998 3360
rect 581054 3304 581059 3360
rect 520181 3302 581059 3304
rect 520181 3299 520247 3302
rect 580993 3299 581059 3302
<< metal4 >>
rect -4876 707718 -4276 707740
rect -4876 707482 -4694 707718
rect -4458 707482 -4276 707718
rect -4876 707398 -4276 707482
rect -4876 707162 -4694 707398
rect -4458 707162 -4276 707398
rect -4876 672054 -4276 707162
rect -4876 671818 -4694 672054
rect -4458 671818 -4276 672054
rect -4876 671734 -4276 671818
rect -4876 671498 -4694 671734
rect -4458 671498 -4276 671734
rect -4876 636054 -4276 671498
rect -4876 635818 -4694 636054
rect -4458 635818 -4276 636054
rect -4876 635734 -4276 635818
rect -4876 635498 -4694 635734
rect -4458 635498 -4276 635734
rect -4876 600054 -4276 635498
rect -4876 599818 -4694 600054
rect -4458 599818 -4276 600054
rect -4876 599734 -4276 599818
rect -4876 599498 -4694 599734
rect -4458 599498 -4276 599734
rect -4876 564054 -4276 599498
rect -4876 563818 -4694 564054
rect -4458 563818 -4276 564054
rect -4876 563734 -4276 563818
rect -4876 563498 -4694 563734
rect -4458 563498 -4276 563734
rect -4876 528054 -4276 563498
rect -4876 527818 -4694 528054
rect -4458 527818 -4276 528054
rect -4876 527734 -4276 527818
rect -4876 527498 -4694 527734
rect -4458 527498 -4276 527734
rect -4876 492054 -4276 527498
rect -4876 491818 -4694 492054
rect -4458 491818 -4276 492054
rect -4876 491734 -4276 491818
rect -4876 491498 -4694 491734
rect -4458 491498 -4276 491734
rect -4876 456054 -4276 491498
rect -4876 455818 -4694 456054
rect -4458 455818 -4276 456054
rect -4876 455734 -4276 455818
rect -4876 455498 -4694 455734
rect -4458 455498 -4276 455734
rect -4876 420054 -4276 455498
rect -4876 419818 -4694 420054
rect -4458 419818 -4276 420054
rect -4876 419734 -4276 419818
rect -4876 419498 -4694 419734
rect -4458 419498 -4276 419734
rect -4876 384054 -4276 419498
rect -4876 383818 -4694 384054
rect -4458 383818 -4276 384054
rect -4876 383734 -4276 383818
rect -4876 383498 -4694 383734
rect -4458 383498 -4276 383734
rect -4876 348054 -4276 383498
rect -4876 347818 -4694 348054
rect -4458 347818 -4276 348054
rect -4876 347734 -4276 347818
rect -4876 347498 -4694 347734
rect -4458 347498 -4276 347734
rect -4876 312054 -4276 347498
rect -4876 311818 -4694 312054
rect -4458 311818 -4276 312054
rect -4876 311734 -4276 311818
rect -4876 311498 -4694 311734
rect -4458 311498 -4276 311734
rect -4876 276054 -4276 311498
rect -4876 275818 -4694 276054
rect -4458 275818 -4276 276054
rect -4876 275734 -4276 275818
rect -4876 275498 -4694 275734
rect -4458 275498 -4276 275734
rect -4876 240054 -4276 275498
rect -4876 239818 -4694 240054
rect -4458 239818 -4276 240054
rect -4876 239734 -4276 239818
rect -4876 239498 -4694 239734
rect -4458 239498 -4276 239734
rect -4876 204054 -4276 239498
rect -4876 203818 -4694 204054
rect -4458 203818 -4276 204054
rect -4876 203734 -4276 203818
rect -4876 203498 -4694 203734
rect -4458 203498 -4276 203734
rect -4876 168054 -4276 203498
rect -4876 167818 -4694 168054
rect -4458 167818 -4276 168054
rect -4876 167734 -4276 167818
rect -4876 167498 -4694 167734
rect -4458 167498 -4276 167734
rect -4876 132054 -4276 167498
rect -4876 131818 -4694 132054
rect -4458 131818 -4276 132054
rect -4876 131734 -4276 131818
rect -4876 131498 -4694 131734
rect -4458 131498 -4276 131734
rect -4876 96054 -4276 131498
rect -4876 95818 -4694 96054
rect -4458 95818 -4276 96054
rect -4876 95734 -4276 95818
rect -4876 95498 -4694 95734
rect -4458 95498 -4276 95734
rect -4876 60054 -4276 95498
rect -4876 59818 -4694 60054
rect -4458 59818 -4276 60054
rect -4876 59734 -4276 59818
rect -4876 59498 -4694 59734
rect -4458 59498 -4276 59734
rect -4876 24054 -4276 59498
rect -4876 23818 -4694 24054
rect -4458 23818 -4276 24054
rect -4876 23734 -4276 23818
rect -4876 23498 -4694 23734
rect -4458 23498 -4276 23734
rect -4876 -3226 -4276 23498
rect -3916 706758 -3316 706780
rect -3916 706522 -3734 706758
rect -3498 706522 -3316 706758
rect -3916 706438 -3316 706522
rect -3916 706202 -3734 706438
rect -3498 706202 -3316 706438
rect -3916 690054 -3316 706202
rect 4404 706758 5004 707740
rect 4404 706522 4586 706758
rect 4822 706522 5004 706758
rect 4404 706438 5004 706522
rect 4404 706202 4586 706438
rect 4822 706202 5004 706438
rect -3916 689818 -3734 690054
rect -3498 689818 -3316 690054
rect -3916 689734 -3316 689818
rect -3916 689498 -3734 689734
rect -3498 689498 -3316 689734
rect -3916 654054 -3316 689498
rect -3916 653818 -3734 654054
rect -3498 653818 -3316 654054
rect -3916 653734 -3316 653818
rect -3916 653498 -3734 653734
rect -3498 653498 -3316 653734
rect -3916 618054 -3316 653498
rect -3916 617818 -3734 618054
rect -3498 617818 -3316 618054
rect -3916 617734 -3316 617818
rect -3916 617498 -3734 617734
rect -3498 617498 -3316 617734
rect -3916 582054 -3316 617498
rect -3916 581818 -3734 582054
rect -3498 581818 -3316 582054
rect -3916 581734 -3316 581818
rect -3916 581498 -3734 581734
rect -3498 581498 -3316 581734
rect -3916 546054 -3316 581498
rect -3916 545818 -3734 546054
rect -3498 545818 -3316 546054
rect -3916 545734 -3316 545818
rect -3916 545498 -3734 545734
rect -3498 545498 -3316 545734
rect -3916 510054 -3316 545498
rect -3916 509818 -3734 510054
rect -3498 509818 -3316 510054
rect -3916 509734 -3316 509818
rect -3916 509498 -3734 509734
rect -3498 509498 -3316 509734
rect -3916 474054 -3316 509498
rect -3916 473818 -3734 474054
rect -3498 473818 -3316 474054
rect -3916 473734 -3316 473818
rect -3916 473498 -3734 473734
rect -3498 473498 -3316 473734
rect -3916 438054 -3316 473498
rect -3916 437818 -3734 438054
rect -3498 437818 -3316 438054
rect -3916 437734 -3316 437818
rect -3916 437498 -3734 437734
rect -3498 437498 -3316 437734
rect -3916 402054 -3316 437498
rect -3916 401818 -3734 402054
rect -3498 401818 -3316 402054
rect -3916 401734 -3316 401818
rect -3916 401498 -3734 401734
rect -3498 401498 -3316 401734
rect -3916 366054 -3316 401498
rect -3916 365818 -3734 366054
rect -3498 365818 -3316 366054
rect -3916 365734 -3316 365818
rect -3916 365498 -3734 365734
rect -3498 365498 -3316 365734
rect -3916 330054 -3316 365498
rect -3916 329818 -3734 330054
rect -3498 329818 -3316 330054
rect -3916 329734 -3316 329818
rect -3916 329498 -3734 329734
rect -3498 329498 -3316 329734
rect -3916 294054 -3316 329498
rect -3916 293818 -3734 294054
rect -3498 293818 -3316 294054
rect -3916 293734 -3316 293818
rect -3916 293498 -3734 293734
rect -3498 293498 -3316 293734
rect -3916 258054 -3316 293498
rect -3916 257818 -3734 258054
rect -3498 257818 -3316 258054
rect -3916 257734 -3316 257818
rect -3916 257498 -3734 257734
rect -3498 257498 -3316 257734
rect -3916 222054 -3316 257498
rect -3916 221818 -3734 222054
rect -3498 221818 -3316 222054
rect -3916 221734 -3316 221818
rect -3916 221498 -3734 221734
rect -3498 221498 -3316 221734
rect -3916 186054 -3316 221498
rect -3916 185818 -3734 186054
rect -3498 185818 -3316 186054
rect -3916 185734 -3316 185818
rect -3916 185498 -3734 185734
rect -3498 185498 -3316 185734
rect -3916 150054 -3316 185498
rect -3916 149818 -3734 150054
rect -3498 149818 -3316 150054
rect -3916 149734 -3316 149818
rect -3916 149498 -3734 149734
rect -3498 149498 -3316 149734
rect -3916 114054 -3316 149498
rect -3916 113818 -3734 114054
rect -3498 113818 -3316 114054
rect -3916 113734 -3316 113818
rect -3916 113498 -3734 113734
rect -3498 113498 -3316 113734
rect -3916 78054 -3316 113498
rect -3916 77818 -3734 78054
rect -3498 77818 -3316 78054
rect -3916 77734 -3316 77818
rect -3916 77498 -3734 77734
rect -3498 77498 -3316 77734
rect -3916 42054 -3316 77498
rect -3916 41818 -3734 42054
rect -3498 41818 -3316 42054
rect -3916 41734 -3316 41818
rect -3916 41498 -3734 41734
rect -3498 41498 -3316 41734
rect -3916 6054 -3316 41498
rect -3916 5818 -3734 6054
rect -3498 5818 -3316 6054
rect -3916 5734 -3316 5818
rect -3916 5498 -3734 5734
rect -3498 5498 -3316 5734
rect -3916 -2266 -3316 5498
rect -2956 705798 -2356 705820
rect -2956 705562 -2774 705798
rect -2538 705562 -2356 705798
rect -2956 705478 -2356 705562
rect -2956 705242 -2774 705478
rect -2538 705242 -2356 705478
rect -2956 668454 -2356 705242
rect -2956 668218 -2774 668454
rect -2538 668218 -2356 668454
rect -2956 668134 -2356 668218
rect -2956 667898 -2774 668134
rect -2538 667898 -2356 668134
rect -2956 632454 -2356 667898
rect -2956 632218 -2774 632454
rect -2538 632218 -2356 632454
rect -2956 632134 -2356 632218
rect -2956 631898 -2774 632134
rect -2538 631898 -2356 632134
rect -2956 596454 -2356 631898
rect -2956 596218 -2774 596454
rect -2538 596218 -2356 596454
rect -2956 596134 -2356 596218
rect -2956 595898 -2774 596134
rect -2538 595898 -2356 596134
rect -2956 560454 -2356 595898
rect -2956 560218 -2774 560454
rect -2538 560218 -2356 560454
rect -2956 560134 -2356 560218
rect -2956 559898 -2774 560134
rect -2538 559898 -2356 560134
rect -2956 524454 -2356 559898
rect -2956 524218 -2774 524454
rect -2538 524218 -2356 524454
rect -2956 524134 -2356 524218
rect -2956 523898 -2774 524134
rect -2538 523898 -2356 524134
rect -2956 488454 -2356 523898
rect -2956 488218 -2774 488454
rect -2538 488218 -2356 488454
rect -2956 488134 -2356 488218
rect -2956 487898 -2774 488134
rect -2538 487898 -2356 488134
rect -2956 452454 -2356 487898
rect -2956 452218 -2774 452454
rect -2538 452218 -2356 452454
rect -2956 452134 -2356 452218
rect -2956 451898 -2774 452134
rect -2538 451898 -2356 452134
rect -2956 416454 -2356 451898
rect -2956 416218 -2774 416454
rect -2538 416218 -2356 416454
rect -2956 416134 -2356 416218
rect -2956 415898 -2774 416134
rect -2538 415898 -2356 416134
rect -2956 380454 -2356 415898
rect -2956 380218 -2774 380454
rect -2538 380218 -2356 380454
rect -2956 380134 -2356 380218
rect -2956 379898 -2774 380134
rect -2538 379898 -2356 380134
rect -2956 344454 -2356 379898
rect -2956 344218 -2774 344454
rect -2538 344218 -2356 344454
rect -2956 344134 -2356 344218
rect -2956 343898 -2774 344134
rect -2538 343898 -2356 344134
rect -2956 308454 -2356 343898
rect -2956 308218 -2774 308454
rect -2538 308218 -2356 308454
rect -2956 308134 -2356 308218
rect -2956 307898 -2774 308134
rect -2538 307898 -2356 308134
rect -2956 272454 -2356 307898
rect -2956 272218 -2774 272454
rect -2538 272218 -2356 272454
rect -2956 272134 -2356 272218
rect -2956 271898 -2774 272134
rect -2538 271898 -2356 272134
rect -2956 236454 -2356 271898
rect -2956 236218 -2774 236454
rect -2538 236218 -2356 236454
rect -2956 236134 -2356 236218
rect -2956 235898 -2774 236134
rect -2538 235898 -2356 236134
rect -2956 200454 -2356 235898
rect -2956 200218 -2774 200454
rect -2538 200218 -2356 200454
rect -2956 200134 -2356 200218
rect -2956 199898 -2774 200134
rect -2538 199898 -2356 200134
rect -2956 164454 -2356 199898
rect -2956 164218 -2774 164454
rect -2538 164218 -2356 164454
rect -2956 164134 -2356 164218
rect -2956 163898 -2774 164134
rect -2538 163898 -2356 164134
rect -2956 128454 -2356 163898
rect -2956 128218 -2774 128454
rect -2538 128218 -2356 128454
rect -2956 128134 -2356 128218
rect -2956 127898 -2774 128134
rect -2538 127898 -2356 128134
rect -2956 92454 -2356 127898
rect -2956 92218 -2774 92454
rect -2538 92218 -2356 92454
rect -2956 92134 -2356 92218
rect -2956 91898 -2774 92134
rect -2538 91898 -2356 92134
rect -2956 56454 -2356 91898
rect -2956 56218 -2774 56454
rect -2538 56218 -2356 56454
rect -2956 56134 -2356 56218
rect -2956 55898 -2774 56134
rect -2538 55898 -2356 56134
rect -2956 20454 -2356 55898
rect -2956 20218 -2774 20454
rect -2538 20218 -2356 20454
rect -2956 20134 -2356 20218
rect -2956 19898 -2774 20134
rect -2538 19898 -2356 20134
rect -2956 -1306 -2356 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705820
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2956 -1542 -2774 -1306
rect -2538 -1542 -2356 -1306
rect -2956 -1626 -2356 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 -2356 -1626
rect -2956 -1884 -2356 -1862
rect 804 -1884 1404 -902
rect 4404 690054 5004 706202
rect 22404 707718 23004 707740
rect 22404 707482 22586 707718
rect 22822 707482 23004 707718
rect 22404 707398 23004 707482
rect 22404 707162 22586 707398
rect 22822 707162 23004 707398
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3916 -2502 -3734 -2266
rect -3498 -2502 -3316 -2266
rect -3916 -2586 -3316 -2502
rect -3916 -2822 -3734 -2586
rect -3498 -2822 -3316 -2586
rect -3916 -2844 -3316 -2822
rect 4404 -2266 5004 5498
rect 18804 705798 19404 705820
rect 18804 705562 18986 705798
rect 19222 705562 19404 705798
rect 18804 705478 19404 705562
rect 18804 705242 18986 705478
rect 19222 705242 19404 705478
rect 18804 668454 19404 705242
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1306 19404 19898
rect 18804 -1542 18986 -1306
rect 19222 -1542 19404 -1306
rect 18804 -1626 19404 -1542
rect 18804 -1862 18986 -1626
rect 19222 -1862 19404 -1626
rect 18804 -1884 19404 -1862
rect 22404 672054 23004 707162
rect 40404 706758 41004 707740
rect 40404 706522 40586 706758
rect 40822 706522 41004 706758
rect 40404 706438 41004 706522
rect 40404 706202 40586 706438
rect 40822 706202 41004 706438
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 4404 -2502 4586 -2266
rect 4822 -2502 5004 -2266
rect 4404 -2586 5004 -2502
rect 4404 -2822 4586 -2586
rect 4822 -2822 5004 -2586
rect -4876 -3462 -4694 -3226
rect -4458 -3462 -4276 -3226
rect -4876 -3546 -4276 -3462
rect -4876 -3782 -4694 -3546
rect -4458 -3782 -4276 -3546
rect -4876 -3804 -4276 -3782
rect 4404 -3804 5004 -2822
rect 22404 -3226 23004 23498
rect 36804 704838 37404 705820
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1884 37404 -902
rect 40404 690054 41004 706202
rect 58404 707718 59004 707740
rect 58404 707482 58586 707718
rect 58822 707482 59004 707718
rect 58404 707398 59004 707482
rect 58404 707162 58586 707398
rect 58822 707162 59004 707398
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 22404 -3462 22586 -3226
rect 22822 -3462 23004 -3226
rect 22404 -3546 23004 -3462
rect 22404 -3782 22586 -3546
rect 22822 -3782 23004 -3546
rect 22404 -3804 23004 -3782
rect 40404 -2266 41004 5498
rect 54804 705798 55404 705820
rect 54804 705562 54986 705798
rect 55222 705562 55404 705798
rect 54804 705478 55404 705562
rect 54804 705242 54986 705478
rect 55222 705242 55404 705478
rect 54804 668454 55404 705242
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1306 55404 19898
rect 54804 -1542 54986 -1306
rect 55222 -1542 55404 -1306
rect 54804 -1626 55404 -1542
rect 54804 -1862 54986 -1626
rect 55222 -1862 55404 -1626
rect 54804 -1884 55404 -1862
rect 58404 672054 59004 707162
rect 76404 706758 77004 707740
rect 76404 706522 76586 706758
rect 76822 706522 77004 706758
rect 76404 706438 77004 706522
rect 76404 706202 76586 706438
rect 76822 706202 77004 706438
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 72804 704838 73404 705820
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 652000 73404 685898
rect 76404 690054 77004 706202
rect 94404 707718 95004 707740
rect 94404 707482 94586 707718
rect 94822 707482 95004 707718
rect 94404 707398 95004 707482
rect 94404 707162 94586 707398
rect 94822 707162 95004 707398
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 652000 77004 653498
rect 90804 705798 91404 705820
rect 90804 705562 90986 705798
rect 91222 705562 91404 705798
rect 90804 705478 91404 705562
rect 90804 705242 90986 705478
rect 91222 705242 91404 705478
rect 90804 668454 91404 705242
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 652000 91404 667898
rect 94404 672054 95004 707162
rect 112404 706758 113004 707740
rect 112404 706522 112586 706758
rect 112822 706522 113004 706758
rect 112404 706438 113004 706522
rect 112404 706202 112586 706438
rect 112822 706202 113004 706438
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 652000 95004 671498
rect 108804 704838 109404 705820
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 652000 109404 685898
rect 112404 690054 113004 706202
rect 130404 707718 131004 707740
rect 130404 707482 130586 707718
rect 130822 707482 131004 707718
rect 130404 707398 131004 707482
rect 130404 707162 130586 707398
rect 130822 707162 131004 707398
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 652000 113004 653498
rect 126804 705798 127404 705820
rect 126804 705562 126986 705798
rect 127222 705562 127404 705798
rect 126804 705478 127404 705562
rect 126804 705242 126986 705478
rect 127222 705242 127404 705478
rect 126804 668454 127404 705242
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 652000 127404 667898
rect 130404 672054 131004 707162
rect 148404 706758 149004 707740
rect 148404 706522 148586 706758
rect 148822 706522 149004 706758
rect 148404 706438 149004 706522
rect 148404 706202 148586 706438
rect 148822 706202 149004 706438
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 652000 131004 671498
rect 144804 704838 145404 705820
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 652000 145404 685898
rect 148404 690054 149004 706202
rect 166404 707718 167004 707740
rect 166404 707482 166586 707718
rect 166822 707482 167004 707718
rect 166404 707398 167004 707482
rect 166404 707162 166586 707398
rect 166822 707162 167004 707398
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 652000 149004 653498
rect 162804 705798 163404 705820
rect 162804 705562 162986 705798
rect 163222 705562 163404 705798
rect 162804 705478 163404 705562
rect 162804 705242 162986 705478
rect 163222 705242 163404 705478
rect 162804 668454 163404 705242
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 652000 163404 667898
rect 166404 672054 167004 707162
rect 184404 706758 185004 707740
rect 184404 706522 184586 706758
rect 184822 706522 185004 706758
rect 184404 706438 185004 706522
rect 184404 706202 184586 706438
rect 184822 706202 185004 706438
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 652000 167004 671498
rect 180804 704838 181404 705820
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 652000 181404 685898
rect 184404 690054 185004 706202
rect 202404 707718 203004 707740
rect 202404 707482 202586 707718
rect 202822 707482 203004 707718
rect 202404 707398 203004 707482
rect 202404 707162 202586 707398
rect 202822 707162 203004 707398
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 652000 185004 653498
rect 198804 705798 199404 705820
rect 198804 705562 198986 705798
rect 199222 705562 199404 705798
rect 198804 705478 199404 705562
rect 198804 705242 198986 705478
rect 199222 705242 199404 705478
rect 198804 668454 199404 705242
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 652000 199404 667898
rect 202404 672054 203004 707162
rect 220404 706758 221004 707740
rect 220404 706522 220586 706758
rect 220822 706522 221004 706758
rect 220404 706438 221004 706522
rect 220404 706202 220586 706438
rect 220822 706202 221004 706438
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 652000 203004 671498
rect 216804 704838 217404 705820
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 652000 217404 685898
rect 220404 690054 221004 706202
rect 238404 707718 239004 707740
rect 238404 707482 238586 707718
rect 238822 707482 239004 707718
rect 238404 707398 239004 707482
rect 238404 707162 238586 707398
rect 238822 707162 239004 707398
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 652000 221004 653498
rect 234804 705798 235404 705820
rect 234804 705562 234986 705798
rect 235222 705562 235404 705798
rect 234804 705478 235404 705562
rect 234804 705242 234986 705478
rect 235222 705242 235404 705478
rect 234804 668454 235404 705242
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 652000 235404 667898
rect 238404 672054 239004 707162
rect 256404 706758 257004 707740
rect 256404 706522 256586 706758
rect 256822 706522 257004 706758
rect 256404 706438 257004 706522
rect 256404 706202 256586 706438
rect 256822 706202 257004 706438
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 652000 239004 671498
rect 252804 704838 253404 705820
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 652000 253404 685898
rect 256404 690054 257004 706202
rect 274404 707718 275004 707740
rect 274404 707482 274586 707718
rect 274822 707482 275004 707718
rect 274404 707398 275004 707482
rect 274404 707162 274586 707398
rect 274822 707162 275004 707398
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 652000 257004 653498
rect 270804 705798 271404 705820
rect 270804 705562 270986 705798
rect 271222 705562 271404 705798
rect 270804 705478 271404 705562
rect 270804 705242 270986 705478
rect 271222 705242 271404 705478
rect 270804 668454 271404 705242
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 652000 271404 667898
rect 274404 672054 275004 707162
rect 292404 706758 293004 707740
rect 292404 706522 292586 706758
rect 292822 706522 293004 706758
rect 292404 706438 293004 706522
rect 292404 706202 292586 706438
rect 292822 706202 293004 706438
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 652000 275004 671498
rect 288804 704838 289404 705820
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 652000 289404 685898
rect 292404 690054 293004 706202
rect 310404 707718 311004 707740
rect 310404 707482 310586 707718
rect 310822 707482 311004 707718
rect 310404 707398 311004 707482
rect 310404 707162 310586 707398
rect 310822 707162 311004 707398
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 652000 293004 653498
rect 306804 705798 307404 705820
rect 306804 705562 306986 705798
rect 307222 705562 307404 705798
rect 306804 705478 307404 705562
rect 306804 705242 306986 705478
rect 307222 705242 307404 705478
rect 306804 668454 307404 705242
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 652000 307404 667898
rect 310404 672054 311004 707162
rect 328404 706758 329004 707740
rect 328404 706522 328586 706758
rect 328822 706522 329004 706758
rect 328404 706438 329004 706522
rect 328404 706202 328586 706438
rect 328822 706202 329004 706438
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 652000 311004 671498
rect 324804 704838 325404 705820
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 652000 325404 685898
rect 328404 690054 329004 706202
rect 346404 707718 347004 707740
rect 346404 707482 346586 707718
rect 346822 707482 347004 707718
rect 346404 707398 347004 707482
rect 346404 707162 346586 707398
rect 346822 707162 347004 707398
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 652000 329004 653498
rect 342804 705798 343404 705820
rect 342804 705562 342986 705798
rect 343222 705562 343404 705798
rect 342804 705478 343404 705562
rect 342804 705242 342986 705478
rect 343222 705242 343404 705478
rect 342804 668454 343404 705242
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 652000 343404 667898
rect 346404 672054 347004 707162
rect 364404 706758 365004 707740
rect 364404 706522 364586 706758
rect 364822 706522 365004 706758
rect 364404 706438 365004 706522
rect 364404 706202 364586 706438
rect 364822 706202 365004 706438
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 652000 347004 671498
rect 360804 704838 361404 705820
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 652000 361404 685898
rect 364404 690054 365004 706202
rect 382404 707718 383004 707740
rect 382404 707482 382586 707718
rect 382822 707482 383004 707718
rect 382404 707398 383004 707482
rect 382404 707162 382586 707398
rect 382822 707162 383004 707398
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 652000 365004 653498
rect 378804 705798 379404 705820
rect 378804 705562 378986 705798
rect 379222 705562 379404 705798
rect 378804 705478 379404 705562
rect 378804 705242 378986 705478
rect 379222 705242 379404 705478
rect 378804 668454 379404 705242
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 652000 379404 667898
rect 382404 672054 383004 707162
rect 400404 706758 401004 707740
rect 400404 706522 400586 706758
rect 400822 706522 401004 706758
rect 400404 706438 401004 706522
rect 400404 706202 400586 706438
rect 400822 706202 401004 706438
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 652000 383004 671498
rect 396804 704838 397404 705820
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 652000 397404 685898
rect 400404 690054 401004 706202
rect 418404 707718 419004 707740
rect 418404 707482 418586 707718
rect 418822 707482 419004 707718
rect 418404 707398 419004 707482
rect 418404 707162 418586 707398
rect 418822 707162 419004 707398
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 652000 401004 653498
rect 414804 705798 415404 705820
rect 414804 705562 414986 705798
rect 415222 705562 415404 705798
rect 414804 705478 415404 705562
rect 414804 705242 414986 705478
rect 415222 705242 415404 705478
rect 414804 668454 415404 705242
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 652000 415404 667898
rect 418404 672054 419004 707162
rect 436404 706758 437004 707740
rect 436404 706522 436586 706758
rect 436822 706522 437004 706758
rect 436404 706438 437004 706522
rect 436404 706202 436586 706438
rect 436822 706202 437004 706438
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 652000 419004 671498
rect 432804 704838 433404 705820
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 652000 433404 685898
rect 436404 690054 437004 706202
rect 454404 707718 455004 707740
rect 454404 707482 454586 707718
rect 454822 707482 455004 707718
rect 454404 707398 455004 707482
rect 454404 707162 454586 707398
rect 454822 707162 455004 707398
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 652000 437004 653498
rect 450804 705798 451404 705820
rect 450804 705562 450986 705798
rect 451222 705562 451404 705798
rect 450804 705478 451404 705562
rect 450804 705242 450986 705478
rect 451222 705242 451404 705478
rect 450804 668454 451404 705242
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 652000 451404 667898
rect 454404 672054 455004 707162
rect 472404 706758 473004 707740
rect 472404 706522 472586 706758
rect 472822 706522 473004 706758
rect 472404 706438 473004 706522
rect 472404 706202 472586 706438
rect 472822 706202 473004 706438
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 652000 455004 671498
rect 468804 704838 469404 705820
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 652000 469404 685898
rect 472404 690054 473004 706202
rect 490404 707718 491004 707740
rect 490404 707482 490586 707718
rect 490822 707482 491004 707718
rect 490404 707398 491004 707482
rect 490404 707162 490586 707398
rect 490822 707162 491004 707398
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 652000 473004 653498
rect 486804 705798 487404 705820
rect 486804 705562 486986 705798
rect 487222 705562 487404 705798
rect 486804 705478 487404 705562
rect 486804 705242 486986 705478
rect 487222 705242 487404 705478
rect 486804 668454 487404 705242
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 652000 487404 667898
rect 490404 672054 491004 707162
rect 508404 706758 509004 707740
rect 508404 706522 508586 706758
rect 508822 706522 509004 706758
rect 508404 706438 509004 706522
rect 508404 706202 508586 706438
rect 508822 706202 509004 706438
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 652000 491004 671498
rect 504804 704838 505404 705820
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 652000 505404 685898
rect 508404 690054 509004 706202
rect 526404 707718 527004 707740
rect 526404 707482 526586 707718
rect 526822 707482 527004 707718
rect 526404 707398 527004 707482
rect 526404 707162 526586 707398
rect 526822 707162 527004 707398
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 652000 509004 653498
rect 522804 705798 523404 705820
rect 522804 705562 522986 705798
rect 523222 705562 523404 705798
rect 522804 705478 523404 705562
rect 522804 705242 522986 705478
rect 523222 705242 523404 705478
rect 522804 668454 523404 705242
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 81568 636054 81888 636076
rect 81568 635818 81610 636054
rect 81846 635818 81888 636054
rect 81568 635734 81888 635818
rect 81568 635498 81610 635734
rect 81846 635498 81888 635734
rect 81568 635476 81888 635498
rect 81568 632454 81888 632476
rect 81568 632218 81610 632454
rect 81846 632218 81888 632454
rect 81568 632134 81888 632218
rect 81568 631898 81610 632134
rect 81846 631898 81888 632134
rect 81568 631876 81888 631898
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 66208 618054 66528 618076
rect 66208 617818 66250 618054
rect 66486 617818 66528 618054
rect 66208 617734 66528 617818
rect 66208 617498 66250 617734
rect 66486 617498 66528 617734
rect 66208 617476 66528 617498
rect 66208 614454 66528 614476
rect 66208 614218 66250 614454
rect 66486 614218 66528 614454
rect 66208 614134 66528 614218
rect 66208 613898 66250 614134
rect 66486 613898 66528 614134
rect 66208 613876 66528 613898
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 81568 600054 81888 600076
rect 81568 599818 81610 600054
rect 81846 599818 81888 600054
rect 81568 599734 81888 599818
rect 81568 599498 81610 599734
rect 81846 599498 81888 599734
rect 81568 599476 81888 599498
rect 81568 596454 81888 596476
rect 81568 596218 81610 596454
rect 81846 596218 81888 596454
rect 81568 596134 81888 596218
rect 81568 595898 81610 596134
rect 81846 595898 81888 596134
rect 81568 595876 81888 595898
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 66208 582054 66528 582076
rect 66208 581818 66250 582054
rect 66486 581818 66528 582054
rect 66208 581734 66528 581818
rect 66208 581498 66250 581734
rect 66486 581498 66528 581734
rect 66208 581476 66528 581498
rect 66208 578454 66528 578476
rect 66208 578218 66250 578454
rect 66486 578218 66528 578454
rect 66208 578134 66528 578218
rect 66208 577898 66250 578134
rect 66486 577898 66528 578134
rect 66208 577876 66528 577898
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 81568 564054 81888 564076
rect 81568 563818 81610 564054
rect 81846 563818 81888 564054
rect 81568 563734 81888 563818
rect 81568 563498 81610 563734
rect 81846 563498 81888 563734
rect 81568 563476 81888 563498
rect 81568 560454 81888 560476
rect 81568 560218 81610 560454
rect 81846 560218 81888 560454
rect 81568 560134 81888 560218
rect 81568 559898 81610 560134
rect 81846 559898 81888 560134
rect 81568 559876 81888 559898
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 66208 546054 66528 546076
rect 66208 545818 66250 546054
rect 66486 545818 66528 546054
rect 66208 545734 66528 545818
rect 66208 545498 66250 545734
rect 66486 545498 66528 545734
rect 66208 545476 66528 545498
rect 66208 542454 66528 542476
rect 66208 542218 66250 542454
rect 66486 542218 66528 542454
rect 66208 542134 66528 542218
rect 66208 541898 66250 542134
rect 66486 541898 66528 542134
rect 66208 541876 66528 541898
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 81568 528054 81888 528076
rect 81568 527818 81610 528054
rect 81846 527818 81888 528054
rect 81568 527734 81888 527818
rect 81568 527498 81610 527734
rect 81846 527498 81888 527734
rect 81568 527476 81888 527498
rect 81568 524454 81888 524476
rect 81568 524218 81610 524454
rect 81846 524218 81888 524454
rect 81568 524134 81888 524218
rect 81568 523898 81610 524134
rect 81846 523898 81888 524134
rect 81568 523876 81888 523898
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 66208 510054 66528 510076
rect 66208 509818 66250 510054
rect 66486 509818 66528 510054
rect 66208 509734 66528 509818
rect 66208 509498 66250 509734
rect 66486 509498 66528 509734
rect 66208 509476 66528 509498
rect 66208 506454 66528 506476
rect 66208 506218 66250 506454
rect 66486 506218 66528 506454
rect 66208 506134 66528 506218
rect 66208 505898 66250 506134
rect 66486 505898 66528 506134
rect 66208 505876 66528 505898
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 81568 492054 81888 492076
rect 81568 491818 81610 492054
rect 81846 491818 81888 492054
rect 81568 491734 81888 491818
rect 81568 491498 81610 491734
rect 81846 491498 81888 491734
rect 81568 491476 81888 491498
rect 81568 488454 81888 488476
rect 81568 488218 81610 488454
rect 81846 488218 81888 488454
rect 81568 488134 81888 488218
rect 81568 487898 81610 488134
rect 81846 487898 81888 488134
rect 81568 487876 81888 487898
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 66208 474054 66528 474076
rect 66208 473818 66250 474054
rect 66486 473818 66528 474054
rect 66208 473734 66528 473818
rect 66208 473498 66250 473734
rect 66486 473498 66528 473734
rect 66208 473476 66528 473498
rect 66208 470454 66528 470476
rect 66208 470218 66250 470454
rect 66486 470218 66528 470454
rect 66208 470134 66528 470218
rect 66208 469898 66250 470134
rect 66486 469898 66528 470134
rect 66208 469876 66528 469898
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 81568 456054 81888 456076
rect 81568 455818 81610 456054
rect 81846 455818 81888 456054
rect 81568 455734 81888 455818
rect 81568 455498 81610 455734
rect 81846 455498 81888 455734
rect 81568 455476 81888 455498
rect 81568 452454 81888 452476
rect 81568 452218 81610 452454
rect 81846 452218 81888 452454
rect 81568 452134 81888 452218
rect 81568 451898 81610 452134
rect 81846 451898 81888 452134
rect 81568 451876 81888 451898
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 66208 438054 66528 438076
rect 66208 437818 66250 438054
rect 66486 437818 66528 438054
rect 66208 437734 66528 437818
rect 66208 437498 66250 437734
rect 66486 437498 66528 437734
rect 66208 437476 66528 437498
rect 66208 434454 66528 434476
rect 66208 434218 66250 434454
rect 66486 434218 66528 434454
rect 66208 434134 66528 434218
rect 66208 433898 66250 434134
rect 66486 433898 66528 434134
rect 66208 433876 66528 433898
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 81568 420054 81888 420076
rect 81568 419818 81610 420054
rect 81846 419818 81888 420054
rect 81568 419734 81888 419818
rect 81568 419498 81610 419734
rect 81846 419498 81888 419734
rect 81568 419476 81888 419498
rect 81568 416454 81888 416476
rect 81568 416218 81610 416454
rect 81846 416218 81888 416454
rect 81568 416134 81888 416218
rect 81568 415898 81610 416134
rect 81846 415898 81888 416134
rect 81568 415876 81888 415898
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 66208 402054 66528 402076
rect 66208 401818 66250 402054
rect 66486 401818 66528 402054
rect 66208 401734 66528 401818
rect 66208 401498 66250 401734
rect 66486 401498 66528 401734
rect 66208 401476 66528 401498
rect 66208 398454 66528 398476
rect 66208 398218 66250 398454
rect 66486 398218 66528 398454
rect 66208 398134 66528 398218
rect 66208 397898 66250 398134
rect 66486 397898 66528 398134
rect 66208 397876 66528 397898
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 81568 384054 81888 384076
rect 81568 383818 81610 384054
rect 81846 383818 81888 384054
rect 81568 383734 81888 383818
rect 81568 383498 81610 383734
rect 81846 383498 81888 383734
rect 81568 383476 81888 383498
rect 81568 380454 81888 380476
rect 81568 380218 81610 380454
rect 81846 380218 81888 380454
rect 81568 380134 81888 380218
rect 81568 379898 81610 380134
rect 81846 379898 81888 380134
rect 81568 379876 81888 379898
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 66208 366054 66528 366076
rect 66208 365818 66250 366054
rect 66486 365818 66528 366054
rect 66208 365734 66528 365818
rect 66208 365498 66250 365734
rect 66486 365498 66528 365734
rect 66208 365476 66528 365498
rect 66208 362454 66528 362476
rect 66208 362218 66250 362454
rect 66486 362218 66528 362454
rect 66208 362134 66528 362218
rect 66208 361898 66250 362134
rect 66486 361898 66528 362134
rect 66208 361876 66528 361898
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 81568 348054 81888 348076
rect 81568 347818 81610 348054
rect 81846 347818 81888 348054
rect 81568 347734 81888 347818
rect 81568 347498 81610 347734
rect 81846 347498 81888 347734
rect 81568 347476 81888 347498
rect 81568 344454 81888 344476
rect 81568 344218 81610 344454
rect 81846 344218 81888 344454
rect 81568 344134 81888 344218
rect 81568 343898 81610 344134
rect 81846 343898 81888 344134
rect 81568 343876 81888 343898
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 66208 330054 66528 330076
rect 66208 329818 66250 330054
rect 66486 329818 66528 330054
rect 66208 329734 66528 329818
rect 66208 329498 66250 329734
rect 66486 329498 66528 329734
rect 66208 329476 66528 329498
rect 66208 326454 66528 326476
rect 66208 326218 66250 326454
rect 66486 326218 66528 326454
rect 66208 326134 66528 326218
rect 66208 325898 66250 326134
rect 66486 325898 66528 326134
rect 66208 325876 66528 325898
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 81568 312054 81888 312076
rect 81568 311818 81610 312054
rect 81846 311818 81888 312054
rect 81568 311734 81888 311818
rect 81568 311498 81610 311734
rect 81846 311498 81888 311734
rect 81568 311476 81888 311498
rect 81568 308454 81888 308476
rect 81568 308218 81610 308454
rect 81846 308218 81888 308454
rect 81568 308134 81888 308218
rect 81568 307898 81610 308134
rect 81846 307898 81888 308134
rect 81568 307876 81888 307898
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 66208 294054 66528 294076
rect 66208 293818 66250 294054
rect 66486 293818 66528 294054
rect 66208 293734 66528 293818
rect 66208 293498 66250 293734
rect 66486 293498 66528 293734
rect 66208 293476 66528 293498
rect 66208 290454 66528 290476
rect 66208 290218 66250 290454
rect 66486 290218 66528 290454
rect 66208 290134 66528 290218
rect 66208 289898 66250 290134
rect 66486 289898 66528 290134
rect 66208 289876 66528 289898
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 81568 276054 81888 276076
rect 81568 275818 81610 276054
rect 81846 275818 81888 276054
rect 81568 275734 81888 275818
rect 81568 275498 81610 275734
rect 81846 275498 81888 275734
rect 81568 275476 81888 275498
rect 81568 272454 81888 272476
rect 81568 272218 81610 272454
rect 81846 272218 81888 272454
rect 81568 272134 81888 272218
rect 81568 271898 81610 272134
rect 81846 271898 81888 272134
rect 81568 271876 81888 271898
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 66208 258054 66528 258076
rect 66208 257818 66250 258054
rect 66486 257818 66528 258054
rect 66208 257734 66528 257818
rect 66208 257498 66250 257734
rect 66486 257498 66528 257734
rect 66208 257476 66528 257498
rect 66208 254454 66528 254476
rect 66208 254218 66250 254454
rect 66486 254218 66528 254454
rect 66208 254134 66528 254218
rect 66208 253898 66250 254134
rect 66486 253898 66528 254134
rect 66208 253876 66528 253898
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 81568 240054 81888 240076
rect 81568 239818 81610 240054
rect 81846 239818 81888 240054
rect 81568 239734 81888 239818
rect 81568 239498 81610 239734
rect 81846 239498 81888 239734
rect 81568 239476 81888 239498
rect 81568 236454 81888 236476
rect 81568 236218 81610 236454
rect 81846 236218 81888 236454
rect 81568 236134 81888 236218
rect 81568 235898 81610 236134
rect 81846 235898 81888 236134
rect 81568 235876 81888 235898
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 66208 222054 66528 222076
rect 66208 221818 66250 222054
rect 66486 221818 66528 222054
rect 66208 221734 66528 221818
rect 66208 221498 66250 221734
rect 66486 221498 66528 221734
rect 66208 221476 66528 221498
rect 66208 218454 66528 218476
rect 66208 218218 66250 218454
rect 66486 218218 66528 218454
rect 66208 218134 66528 218218
rect 66208 217898 66250 218134
rect 66486 217898 66528 218134
rect 66208 217876 66528 217898
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 81568 204054 81888 204076
rect 81568 203818 81610 204054
rect 81846 203818 81888 204054
rect 81568 203734 81888 203818
rect 81568 203498 81610 203734
rect 81846 203498 81888 203734
rect 81568 203476 81888 203498
rect 81568 200454 81888 200476
rect 81568 200218 81610 200454
rect 81846 200218 81888 200454
rect 81568 200134 81888 200218
rect 81568 199898 81610 200134
rect 81846 199898 81888 200134
rect 81568 199876 81888 199898
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 66208 186054 66528 186076
rect 66208 185818 66250 186054
rect 66486 185818 66528 186054
rect 66208 185734 66528 185818
rect 66208 185498 66250 185734
rect 66486 185498 66528 185734
rect 66208 185476 66528 185498
rect 66208 182454 66528 182476
rect 66208 182218 66250 182454
rect 66486 182218 66528 182454
rect 66208 182134 66528 182218
rect 66208 181898 66250 182134
rect 66486 181898 66528 182134
rect 66208 181876 66528 181898
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 81568 168054 81888 168076
rect 81568 167818 81610 168054
rect 81846 167818 81888 168054
rect 81568 167734 81888 167818
rect 81568 167498 81610 167734
rect 81846 167498 81888 167734
rect 81568 167476 81888 167498
rect 81568 164454 81888 164476
rect 81568 164218 81610 164454
rect 81846 164218 81888 164454
rect 81568 164134 81888 164218
rect 81568 163898 81610 164134
rect 81846 163898 81888 164134
rect 81568 163876 81888 163898
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 66208 150054 66528 150076
rect 66208 149818 66250 150054
rect 66486 149818 66528 150054
rect 66208 149734 66528 149818
rect 66208 149498 66250 149734
rect 66486 149498 66528 149734
rect 66208 149476 66528 149498
rect 66208 146454 66528 146476
rect 66208 146218 66250 146454
rect 66486 146218 66528 146454
rect 66208 146134 66528 146218
rect 66208 145898 66250 146134
rect 66486 145898 66528 146134
rect 66208 145876 66528 145898
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 81568 132054 81888 132076
rect 81568 131818 81610 132054
rect 81846 131818 81888 132054
rect 81568 131734 81888 131818
rect 81568 131498 81610 131734
rect 81846 131498 81888 131734
rect 81568 131476 81888 131498
rect 81568 128454 81888 128476
rect 81568 128218 81610 128454
rect 81846 128218 81888 128454
rect 81568 128134 81888 128218
rect 81568 127898 81610 128134
rect 81846 127898 81888 128134
rect 81568 127876 81888 127898
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 66208 114054 66528 114076
rect 66208 113818 66250 114054
rect 66486 113818 66528 114054
rect 66208 113734 66528 113818
rect 66208 113498 66250 113734
rect 66486 113498 66528 113734
rect 66208 113476 66528 113498
rect 66208 110454 66528 110476
rect 66208 110218 66250 110454
rect 66486 110218 66528 110454
rect 66208 110134 66528 110218
rect 66208 109898 66250 110134
rect 66486 109898 66528 110134
rect 66208 109876 66528 109898
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 81568 96054 81888 96076
rect 81568 95818 81610 96054
rect 81846 95818 81888 96054
rect 81568 95734 81888 95818
rect 81568 95498 81610 95734
rect 81846 95498 81888 95734
rect 81568 95476 81888 95498
rect 81568 92454 81888 92476
rect 81568 92218 81610 92454
rect 81846 92218 81888 92454
rect 81568 92134 81888 92218
rect 81568 91898 81610 92134
rect 81846 91898 81888 92134
rect 81568 91876 81888 91898
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 66208 78054 66528 78076
rect 66208 77818 66250 78054
rect 66486 77818 66528 78054
rect 66208 77734 66528 77818
rect 66208 77498 66250 77734
rect 66486 77498 66528 77734
rect 66208 77476 66528 77498
rect 66208 74454 66528 74476
rect 66208 74218 66250 74454
rect 66486 74218 66528 74454
rect 66208 74134 66528 74218
rect 66208 73898 66250 74134
rect 66486 73898 66528 74134
rect 66208 73876 66528 73898
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 81568 60054 81888 60076
rect 81568 59818 81610 60054
rect 81846 59818 81888 60054
rect 81568 59734 81888 59818
rect 81568 59498 81610 59734
rect 81846 59498 81888 59734
rect 81568 59476 81888 59498
rect 81568 56454 81888 56476
rect 81568 56218 81610 56454
rect 81846 56218 81888 56454
rect 81568 56134 81888 56218
rect 81568 55898 81610 56134
rect 81846 55898 81888 56134
rect 81568 55876 81888 55898
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 40404 -2502 40586 -2266
rect 40822 -2502 41004 -2266
rect 40404 -2586 41004 -2502
rect 40404 -2822 40586 -2586
rect 40822 -2822 41004 -2586
rect 40404 -3804 41004 -2822
rect 58404 -3226 59004 23498
rect 72804 38454 73404 52000
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1884 73404 -902
rect 76404 42054 77004 52000
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 58404 -3462 58586 -3226
rect 58822 -3462 59004 -3226
rect 58404 -3546 59004 -3462
rect 58404 -3782 58586 -3546
rect 58822 -3782 59004 -3546
rect 58404 -3804 59004 -3782
rect 76404 -2266 77004 5498
rect 90804 20454 91404 52000
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1306 91404 19898
rect 90804 -1542 90986 -1306
rect 91222 -1542 91404 -1306
rect 90804 -1626 91404 -1542
rect 90804 -1862 90986 -1626
rect 91222 -1862 91404 -1626
rect 90804 -1884 91404 -1862
rect 94404 24054 95004 52000
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 76404 -2502 76586 -2266
rect 76822 -2502 77004 -2266
rect 76404 -2586 77004 -2502
rect 76404 -2822 76586 -2586
rect 76822 -2822 77004 -2586
rect 76404 -3804 77004 -2822
rect 94404 -3226 95004 23498
rect 108804 38454 109404 52000
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1884 109404 -902
rect 112404 42054 113004 52000
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 94404 -3462 94586 -3226
rect 94822 -3462 95004 -3226
rect 94404 -3546 95004 -3462
rect 94404 -3782 94586 -3546
rect 94822 -3782 95004 -3546
rect 94404 -3804 95004 -3782
rect 112404 -2266 113004 5498
rect 126804 20454 127404 52000
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1306 127404 19898
rect 126804 -1542 126986 -1306
rect 127222 -1542 127404 -1306
rect 126804 -1626 127404 -1542
rect 126804 -1862 126986 -1626
rect 127222 -1862 127404 -1626
rect 126804 -1884 127404 -1862
rect 130404 24054 131004 52000
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 112404 -2502 112586 -2266
rect 112822 -2502 113004 -2266
rect 112404 -2586 113004 -2502
rect 112404 -2822 112586 -2586
rect 112822 -2822 113004 -2586
rect 112404 -3804 113004 -2822
rect 130404 -3226 131004 23498
rect 144804 38454 145404 52000
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1884 145404 -902
rect 148404 42054 149004 52000
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 130404 -3462 130586 -3226
rect 130822 -3462 131004 -3226
rect 130404 -3546 131004 -3462
rect 130404 -3782 130586 -3546
rect 130822 -3782 131004 -3546
rect 130404 -3804 131004 -3782
rect 148404 -2266 149004 5498
rect 162804 20454 163404 52000
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1306 163404 19898
rect 162804 -1542 162986 -1306
rect 163222 -1542 163404 -1306
rect 162804 -1626 163404 -1542
rect 162804 -1862 162986 -1626
rect 163222 -1862 163404 -1626
rect 162804 -1884 163404 -1862
rect 166404 24054 167004 52000
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 148404 -2502 148586 -2266
rect 148822 -2502 149004 -2266
rect 148404 -2586 149004 -2502
rect 148404 -2822 148586 -2586
rect 148822 -2822 149004 -2586
rect 148404 -3804 149004 -2822
rect 166404 -3226 167004 23498
rect 180804 38454 181404 52000
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1884 181404 -902
rect 184404 42054 185004 52000
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 166404 -3462 166586 -3226
rect 166822 -3462 167004 -3226
rect 166404 -3546 167004 -3462
rect 166404 -3782 166586 -3546
rect 166822 -3782 167004 -3546
rect 166404 -3804 167004 -3782
rect 184404 -2266 185004 5498
rect 198804 20454 199404 52000
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1306 199404 19898
rect 198804 -1542 198986 -1306
rect 199222 -1542 199404 -1306
rect 198804 -1626 199404 -1542
rect 198804 -1862 198986 -1626
rect 199222 -1862 199404 -1626
rect 198804 -1884 199404 -1862
rect 202404 24054 203004 52000
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 184404 -2502 184586 -2266
rect 184822 -2502 185004 -2266
rect 184404 -2586 185004 -2502
rect 184404 -2822 184586 -2586
rect 184822 -2822 185004 -2586
rect 184404 -3804 185004 -2822
rect 202404 -3226 203004 23498
rect 216804 38454 217404 52000
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1884 217404 -902
rect 220404 42054 221004 52000
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 202404 -3462 202586 -3226
rect 202822 -3462 203004 -3226
rect 202404 -3546 203004 -3462
rect 202404 -3782 202586 -3546
rect 202822 -3782 203004 -3546
rect 202404 -3804 203004 -3782
rect 220404 -2266 221004 5498
rect 234804 20454 235404 52000
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1306 235404 19898
rect 234804 -1542 234986 -1306
rect 235222 -1542 235404 -1306
rect 234804 -1626 235404 -1542
rect 234804 -1862 234986 -1626
rect 235222 -1862 235404 -1626
rect 234804 -1884 235404 -1862
rect 238404 24054 239004 52000
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 220404 -2502 220586 -2266
rect 220822 -2502 221004 -2266
rect 220404 -2586 221004 -2502
rect 220404 -2822 220586 -2586
rect 220822 -2822 221004 -2586
rect 220404 -3804 221004 -2822
rect 238404 -3226 239004 23498
rect 252804 38454 253404 52000
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1884 253404 -902
rect 256404 42054 257004 52000
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 238404 -3462 238586 -3226
rect 238822 -3462 239004 -3226
rect 238404 -3546 239004 -3462
rect 238404 -3782 238586 -3546
rect 238822 -3782 239004 -3546
rect 238404 -3804 239004 -3782
rect 256404 -2266 257004 5498
rect 270804 20454 271404 52000
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1306 271404 19898
rect 270804 -1542 270986 -1306
rect 271222 -1542 271404 -1306
rect 270804 -1626 271404 -1542
rect 270804 -1862 270986 -1626
rect 271222 -1862 271404 -1626
rect 270804 -1884 271404 -1862
rect 274404 24054 275004 52000
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 256404 -2502 256586 -2266
rect 256822 -2502 257004 -2266
rect 256404 -2586 257004 -2502
rect 256404 -2822 256586 -2586
rect 256822 -2822 257004 -2586
rect 256404 -3804 257004 -2822
rect 274404 -3226 275004 23498
rect 288804 38454 289404 52000
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1884 289404 -902
rect 292404 42054 293004 52000
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 274404 -3462 274586 -3226
rect 274822 -3462 275004 -3226
rect 274404 -3546 275004 -3462
rect 274404 -3782 274586 -3546
rect 274822 -3782 275004 -3546
rect 274404 -3804 275004 -3782
rect 292404 -2266 293004 5498
rect 306804 20454 307404 52000
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1306 307404 19898
rect 306804 -1542 306986 -1306
rect 307222 -1542 307404 -1306
rect 306804 -1626 307404 -1542
rect 306804 -1862 306986 -1626
rect 307222 -1862 307404 -1626
rect 306804 -1884 307404 -1862
rect 310404 24054 311004 52000
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 292404 -2502 292586 -2266
rect 292822 -2502 293004 -2266
rect 292404 -2586 293004 -2502
rect 292404 -2822 292586 -2586
rect 292822 -2822 293004 -2586
rect 292404 -3804 293004 -2822
rect 310404 -3226 311004 23498
rect 324804 38454 325404 52000
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1884 325404 -902
rect 328404 42054 329004 52000
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 310404 -3462 310586 -3226
rect 310822 -3462 311004 -3226
rect 310404 -3546 311004 -3462
rect 310404 -3782 310586 -3546
rect 310822 -3782 311004 -3546
rect 310404 -3804 311004 -3782
rect 328404 -2266 329004 5498
rect 342804 20454 343404 52000
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1306 343404 19898
rect 342804 -1542 342986 -1306
rect 343222 -1542 343404 -1306
rect 342804 -1626 343404 -1542
rect 342804 -1862 342986 -1626
rect 343222 -1862 343404 -1626
rect 342804 -1884 343404 -1862
rect 346404 24054 347004 52000
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 328404 -2502 328586 -2266
rect 328822 -2502 329004 -2266
rect 328404 -2586 329004 -2502
rect 328404 -2822 328586 -2586
rect 328822 -2822 329004 -2586
rect 328404 -3804 329004 -2822
rect 346404 -3226 347004 23498
rect 360804 38454 361404 52000
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1884 361404 -902
rect 364404 42054 365004 52000
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 346404 -3462 346586 -3226
rect 346822 -3462 347004 -3226
rect 346404 -3546 347004 -3462
rect 346404 -3782 346586 -3546
rect 346822 -3782 347004 -3546
rect 346404 -3804 347004 -3782
rect 364404 -2266 365004 5498
rect 378804 20454 379404 52000
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1306 379404 19898
rect 378804 -1542 378986 -1306
rect 379222 -1542 379404 -1306
rect 378804 -1626 379404 -1542
rect 378804 -1862 378986 -1626
rect 379222 -1862 379404 -1626
rect 378804 -1884 379404 -1862
rect 382404 24054 383004 52000
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 364404 -2502 364586 -2266
rect 364822 -2502 365004 -2266
rect 364404 -2586 365004 -2502
rect 364404 -2822 364586 -2586
rect 364822 -2822 365004 -2586
rect 364404 -3804 365004 -2822
rect 382404 -3226 383004 23498
rect 396804 38454 397404 52000
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1884 397404 -902
rect 400404 42054 401004 52000
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 382404 -3462 382586 -3226
rect 382822 -3462 383004 -3226
rect 382404 -3546 383004 -3462
rect 382404 -3782 382586 -3546
rect 382822 -3782 383004 -3546
rect 382404 -3804 383004 -3782
rect 400404 -2266 401004 5498
rect 414804 20454 415404 52000
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1306 415404 19898
rect 414804 -1542 414986 -1306
rect 415222 -1542 415404 -1306
rect 414804 -1626 415404 -1542
rect 414804 -1862 414986 -1626
rect 415222 -1862 415404 -1626
rect 414804 -1884 415404 -1862
rect 418404 24054 419004 52000
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 400404 -2502 400586 -2266
rect 400822 -2502 401004 -2266
rect 400404 -2586 401004 -2502
rect 400404 -2822 400586 -2586
rect 400822 -2822 401004 -2586
rect 400404 -3804 401004 -2822
rect 418404 -3226 419004 23498
rect 432804 38454 433404 52000
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1884 433404 -902
rect 436404 42054 437004 52000
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 418404 -3462 418586 -3226
rect 418822 -3462 419004 -3226
rect 418404 -3546 419004 -3462
rect 418404 -3782 418586 -3546
rect 418822 -3782 419004 -3546
rect 418404 -3804 419004 -3782
rect 436404 -2266 437004 5498
rect 450804 20454 451404 52000
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1306 451404 19898
rect 450804 -1542 450986 -1306
rect 451222 -1542 451404 -1306
rect 450804 -1626 451404 -1542
rect 450804 -1862 450986 -1626
rect 451222 -1862 451404 -1626
rect 450804 -1884 451404 -1862
rect 454404 24054 455004 52000
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 436404 -2502 436586 -2266
rect 436822 -2502 437004 -2266
rect 436404 -2586 437004 -2502
rect 436404 -2822 436586 -2586
rect 436822 -2822 437004 -2586
rect 436404 -3804 437004 -2822
rect 454404 -3226 455004 23498
rect 468804 38454 469404 52000
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1884 469404 -902
rect 472404 42054 473004 52000
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 454404 -3462 454586 -3226
rect 454822 -3462 455004 -3226
rect 454404 -3546 455004 -3462
rect 454404 -3782 454586 -3546
rect 454822 -3782 455004 -3546
rect 454404 -3804 455004 -3782
rect 472404 -2266 473004 5498
rect 486804 20454 487404 52000
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1306 487404 19898
rect 486804 -1542 486986 -1306
rect 487222 -1542 487404 -1306
rect 486804 -1626 487404 -1542
rect 486804 -1862 486986 -1626
rect 487222 -1862 487404 -1626
rect 486804 -1884 487404 -1862
rect 490404 24054 491004 52000
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 472404 -2502 472586 -2266
rect 472822 -2502 473004 -2266
rect 472404 -2586 473004 -2502
rect 472404 -2822 472586 -2586
rect 472822 -2822 473004 -2586
rect 472404 -3804 473004 -2822
rect 490404 -3226 491004 23498
rect 504804 38454 505404 52000
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1884 505404 -902
rect 508404 42054 509004 52000
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 490404 -3462 490586 -3226
rect 490822 -3462 491004 -3226
rect 490404 -3546 491004 -3462
rect 490404 -3782 490586 -3546
rect 490822 -3782 491004 -3546
rect 490404 -3804 491004 -3782
rect 508404 -2266 509004 5498
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1306 523404 19898
rect 522804 -1542 522986 -1306
rect 523222 -1542 523404 -1306
rect 522804 -1626 523404 -1542
rect 522804 -1862 522986 -1626
rect 523222 -1862 523404 -1626
rect 522804 -1884 523404 -1862
rect 526404 672054 527004 707162
rect 544404 706758 545004 707740
rect 544404 706522 544586 706758
rect 544822 706522 545004 706758
rect 544404 706438 545004 706522
rect 544404 706202 544586 706438
rect 544822 706202 545004 706438
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 508404 -2502 508586 -2266
rect 508822 -2502 509004 -2266
rect 508404 -2586 509004 -2502
rect 508404 -2822 508586 -2586
rect 508822 -2822 509004 -2586
rect 508404 -3804 509004 -2822
rect 526404 -3226 527004 23498
rect 540804 704838 541404 705820
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1884 541404 -902
rect 544404 690054 545004 706202
rect 562404 707718 563004 707740
rect 562404 707482 562586 707718
rect 562822 707482 563004 707718
rect 562404 707398 563004 707482
rect 562404 707162 562586 707398
rect 562822 707162 563004 707398
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 526404 -3462 526586 -3226
rect 526822 -3462 527004 -3226
rect 526404 -3546 527004 -3462
rect 526404 -3782 526586 -3546
rect 526822 -3782 527004 -3546
rect 526404 -3804 527004 -3782
rect 544404 -2266 545004 5498
rect 558804 705798 559404 705820
rect 558804 705562 558986 705798
rect 559222 705562 559404 705798
rect 558804 705478 559404 705562
rect 558804 705242 558986 705478
rect 559222 705242 559404 705478
rect 558804 668454 559404 705242
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1306 559404 19898
rect 558804 -1542 558986 -1306
rect 559222 -1542 559404 -1306
rect 558804 -1626 559404 -1542
rect 558804 -1862 558986 -1626
rect 559222 -1862 559404 -1626
rect 558804 -1884 559404 -1862
rect 562404 672054 563004 707162
rect 580404 706758 581004 707740
rect 588200 707718 588800 707740
rect 588200 707482 588382 707718
rect 588618 707482 588800 707718
rect 588200 707398 588800 707482
rect 588200 707162 588382 707398
rect 588618 707162 588800 707398
rect 580404 706522 580586 706758
rect 580822 706522 581004 706758
rect 580404 706438 581004 706522
rect 580404 706202 580586 706438
rect 580822 706202 581004 706438
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 544404 -2502 544586 -2266
rect 544822 -2502 545004 -2266
rect 544404 -2586 545004 -2502
rect 544404 -2822 544586 -2586
rect 544822 -2822 545004 -2586
rect 544404 -3804 545004 -2822
rect 562404 -3226 563004 23498
rect 576804 704838 577404 705820
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1884 577404 -902
rect 580404 690054 581004 706202
rect 587240 706758 587840 706780
rect 587240 706522 587422 706758
rect 587658 706522 587840 706758
rect 587240 706438 587840 706522
rect 587240 706202 587422 706438
rect 587658 706202 587840 706438
rect 586280 705798 586880 705820
rect 586280 705562 586462 705798
rect 586698 705562 586880 705798
rect 586280 705478 586880 705562
rect 586280 705242 586462 705478
rect 586698 705242 586880 705478
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 562404 -3462 562586 -3226
rect 562822 -3462 563004 -3226
rect 562404 -3546 563004 -3462
rect 562404 -3782 562586 -3546
rect 562822 -3782 563004 -3546
rect 562404 -3804 563004 -3782
rect 580404 -2266 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586280 668454 586880 705242
rect 586280 668218 586462 668454
rect 586698 668218 586880 668454
rect 586280 668134 586880 668218
rect 586280 667898 586462 668134
rect 586698 667898 586880 668134
rect 586280 632454 586880 667898
rect 586280 632218 586462 632454
rect 586698 632218 586880 632454
rect 586280 632134 586880 632218
rect 586280 631898 586462 632134
rect 586698 631898 586880 632134
rect 586280 596454 586880 631898
rect 586280 596218 586462 596454
rect 586698 596218 586880 596454
rect 586280 596134 586880 596218
rect 586280 595898 586462 596134
rect 586698 595898 586880 596134
rect 586280 560454 586880 595898
rect 586280 560218 586462 560454
rect 586698 560218 586880 560454
rect 586280 560134 586880 560218
rect 586280 559898 586462 560134
rect 586698 559898 586880 560134
rect 586280 524454 586880 559898
rect 586280 524218 586462 524454
rect 586698 524218 586880 524454
rect 586280 524134 586880 524218
rect 586280 523898 586462 524134
rect 586698 523898 586880 524134
rect 586280 488454 586880 523898
rect 586280 488218 586462 488454
rect 586698 488218 586880 488454
rect 586280 488134 586880 488218
rect 586280 487898 586462 488134
rect 586698 487898 586880 488134
rect 586280 452454 586880 487898
rect 586280 452218 586462 452454
rect 586698 452218 586880 452454
rect 586280 452134 586880 452218
rect 586280 451898 586462 452134
rect 586698 451898 586880 452134
rect 586280 416454 586880 451898
rect 586280 416218 586462 416454
rect 586698 416218 586880 416454
rect 586280 416134 586880 416218
rect 586280 415898 586462 416134
rect 586698 415898 586880 416134
rect 586280 380454 586880 415898
rect 586280 380218 586462 380454
rect 586698 380218 586880 380454
rect 586280 380134 586880 380218
rect 586280 379898 586462 380134
rect 586698 379898 586880 380134
rect 586280 344454 586880 379898
rect 586280 344218 586462 344454
rect 586698 344218 586880 344454
rect 586280 344134 586880 344218
rect 586280 343898 586462 344134
rect 586698 343898 586880 344134
rect 586280 308454 586880 343898
rect 586280 308218 586462 308454
rect 586698 308218 586880 308454
rect 586280 308134 586880 308218
rect 586280 307898 586462 308134
rect 586698 307898 586880 308134
rect 586280 272454 586880 307898
rect 586280 272218 586462 272454
rect 586698 272218 586880 272454
rect 586280 272134 586880 272218
rect 586280 271898 586462 272134
rect 586698 271898 586880 272134
rect 586280 236454 586880 271898
rect 586280 236218 586462 236454
rect 586698 236218 586880 236454
rect 586280 236134 586880 236218
rect 586280 235898 586462 236134
rect 586698 235898 586880 236134
rect 586280 200454 586880 235898
rect 586280 200218 586462 200454
rect 586698 200218 586880 200454
rect 586280 200134 586880 200218
rect 586280 199898 586462 200134
rect 586698 199898 586880 200134
rect 586280 164454 586880 199898
rect 586280 164218 586462 164454
rect 586698 164218 586880 164454
rect 586280 164134 586880 164218
rect 586280 163898 586462 164134
rect 586698 163898 586880 164134
rect 586280 128454 586880 163898
rect 586280 128218 586462 128454
rect 586698 128218 586880 128454
rect 586280 128134 586880 128218
rect 586280 127898 586462 128134
rect 586698 127898 586880 128134
rect 586280 92454 586880 127898
rect 586280 92218 586462 92454
rect 586698 92218 586880 92454
rect 586280 92134 586880 92218
rect 586280 91898 586462 92134
rect 586698 91898 586880 92134
rect 586280 56454 586880 91898
rect 586280 56218 586462 56454
rect 586698 56218 586880 56454
rect 586280 56134 586880 56218
rect 586280 55898 586462 56134
rect 586698 55898 586880 56134
rect 586280 20454 586880 55898
rect 586280 20218 586462 20454
rect 586698 20218 586880 20454
rect 586280 20134 586880 20218
rect 586280 19898 586462 20134
rect 586698 19898 586880 20134
rect 586280 -1306 586880 19898
rect 586280 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect 586280 -1626 586880 -1542
rect 586280 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect 586280 -1884 586880 -1862
rect 587240 690054 587840 706202
rect 587240 689818 587422 690054
rect 587658 689818 587840 690054
rect 587240 689734 587840 689818
rect 587240 689498 587422 689734
rect 587658 689498 587840 689734
rect 587240 654054 587840 689498
rect 587240 653818 587422 654054
rect 587658 653818 587840 654054
rect 587240 653734 587840 653818
rect 587240 653498 587422 653734
rect 587658 653498 587840 653734
rect 587240 618054 587840 653498
rect 587240 617818 587422 618054
rect 587658 617818 587840 618054
rect 587240 617734 587840 617818
rect 587240 617498 587422 617734
rect 587658 617498 587840 617734
rect 587240 582054 587840 617498
rect 587240 581818 587422 582054
rect 587658 581818 587840 582054
rect 587240 581734 587840 581818
rect 587240 581498 587422 581734
rect 587658 581498 587840 581734
rect 587240 546054 587840 581498
rect 587240 545818 587422 546054
rect 587658 545818 587840 546054
rect 587240 545734 587840 545818
rect 587240 545498 587422 545734
rect 587658 545498 587840 545734
rect 587240 510054 587840 545498
rect 587240 509818 587422 510054
rect 587658 509818 587840 510054
rect 587240 509734 587840 509818
rect 587240 509498 587422 509734
rect 587658 509498 587840 509734
rect 587240 474054 587840 509498
rect 587240 473818 587422 474054
rect 587658 473818 587840 474054
rect 587240 473734 587840 473818
rect 587240 473498 587422 473734
rect 587658 473498 587840 473734
rect 587240 438054 587840 473498
rect 587240 437818 587422 438054
rect 587658 437818 587840 438054
rect 587240 437734 587840 437818
rect 587240 437498 587422 437734
rect 587658 437498 587840 437734
rect 587240 402054 587840 437498
rect 587240 401818 587422 402054
rect 587658 401818 587840 402054
rect 587240 401734 587840 401818
rect 587240 401498 587422 401734
rect 587658 401498 587840 401734
rect 587240 366054 587840 401498
rect 587240 365818 587422 366054
rect 587658 365818 587840 366054
rect 587240 365734 587840 365818
rect 587240 365498 587422 365734
rect 587658 365498 587840 365734
rect 587240 330054 587840 365498
rect 587240 329818 587422 330054
rect 587658 329818 587840 330054
rect 587240 329734 587840 329818
rect 587240 329498 587422 329734
rect 587658 329498 587840 329734
rect 587240 294054 587840 329498
rect 587240 293818 587422 294054
rect 587658 293818 587840 294054
rect 587240 293734 587840 293818
rect 587240 293498 587422 293734
rect 587658 293498 587840 293734
rect 587240 258054 587840 293498
rect 587240 257818 587422 258054
rect 587658 257818 587840 258054
rect 587240 257734 587840 257818
rect 587240 257498 587422 257734
rect 587658 257498 587840 257734
rect 587240 222054 587840 257498
rect 587240 221818 587422 222054
rect 587658 221818 587840 222054
rect 587240 221734 587840 221818
rect 587240 221498 587422 221734
rect 587658 221498 587840 221734
rect 587240 186054 587840 221498
rect 587240 185818 587422 186054
rect 587658 185818 587840 186054
rect 587240 185734 587840 185818
rect 587240 185498 587422 185734
rect 587658 185498 587840 185734
rect 587240 150054 587840 185498
rect 587240 149818 587422 150054
rect 587658 149818 587840 150054
rect 587240 149734 587840 149818
rect 587240 149498 587422 149734
rect 587658 149498 587840 149734
rect 587240 114054 587840 149498
rect 587240 113818 587422 114054
rect 587658 113818 587840 114054
rect 587240 113734 587840 113818
rect 587240 113498 587422 113734
rect 587658 113498 587840 113734
rect 587240 78054 587840 113498
rect 587240 77818 587422 78054
rect 587658 77818 587840 78054
rect 587240 77734 587840 77818
rect 587240 77498 587422 77734
rect 587658 77498 587840 77734
rect 587240 42054 587840 77498
rect 587240 41818 587422 42054
rect 587658 41818 587840 42054
rect 587240 41734 587840 41818
rect 587240 41498 587422 41734
rect 587658 41498 587840 41734
rect 587240 6054 587840 41498
rect 587240 5818 587422 6054
rect 587658 5818 587840 6054
rect 587240 5734 587840 5818
rect 587240 5498 587422 5734
rect 587658 5498 587840 5734
rect 580404 -2502 580586 -2266
rect 580822 -2502 581004 -2266
rect 580404 -2586 581004 -2502
rect 580404 -2822 580586 -2586
rect 580822 -2822 581004 -2586
rect 580404 -3804 581004 -2822
rect 587240 -2266 587840 5498
rect 587240 -2502 587422 -2266
rect 587658 -2502 587840 -2266
rect 587240 -2586 587840 -2502
rect 587240 -2822 587422 -2586
rect 587658 -2822 587840 -2586
rect 587240 -2844 587840 -2822
rect 588200 672054 588800 707162
rect 588200 671818 588382 672054
rect 588618 671818 588800 672054
rect 588200 671734 588800 671818
rect 588200 671498 588382 671734
rect 588618 671498 588800 671734
rect 588200 636054 588800 671498
rect 588200 635818 588382 636054
rect 588618 635818 588800 636054
rect 588200 635734 588800 635818
rect 588200 635498 588382 635734
rect 588618 635498 588800 635734
rect 588200 600054 588800 635498
rect 588200 599818 588382 600054
rect 588618 599818 588800 600054
rect 588200 599734 588800 599818
rect 588200 599498 588382 599734
rect 588618 599498 588800 599734
rect 588200 564054 588800 599498
rect 588200 563818 588382 564054
rect 588618 563818 588800 564054
rect 588200 563734 588800 563818
rect 588200 563498 588382 563734
rect 588618 563498 588800 563734
rect 588200 528054 588800 563498
rect 588200 527818 588382 528054
rect 588618 527818 588800 528054
rect 588200 527734 588800 527818
rect 588200 527498 588382 527734
rect 588618 527498 588800 527734
rect 588200 492054 588800 527498
rect 588200 491818 588382 492054
rect 588618 491818 588800 492054
rect 588200 491734 588800 491818
rect 588200 491498 588382 491734
rect 588618 491498 588800 491734
rect 588200 456054 588800 491498
rect 588200 455818 588382 456054
rect 588618 455818 588800 456054
rect 588200 455734 588800 455818
rect 588200 455498 588382 455734
rect 588618 455498 588800 455734
rect 588200 420054 588800 455498
rect 588200 419818 588382 420054
rect 588618 419818 588800 420054
rect 588200 419734 588800 419818
rect 588200 419498 588382 419734
rect 588618 419498 588800 419734
rect 588200 384054 588800 419498
rect 588200 383818 588382 384054
rect 588618 383818 588800 384054
rect 588200 383734 588800 383818
rect 588200 383498 588382 383734
rect 588618 383498 588800 383734
rect 588200 348054 588800 383498
rect 588200 347818 588382 348054
rect 588618 347818 588800 348054
rect 588200 347734 588800 347818
rect 588200 347498 588382 347734
rect 588618 347498 588800 347734
rect 588200 312054 588800 347498
rect 588200 311818 588382 312054
rect 588618 311818 588800 312054
rect 588200 311734 588800 311818
rect 588200 311498 588382 311734
rect 588618 311498 588800 311734
rect 588200 276054 588800 311498
rect 588200 275818 588382 276054
rect 588618 275818 588800 276054
rect 588200 275734 588800 275818
rect 588200 275498 588382 275734
rect 588618 275498 588800 275734
rect 588200 240054 588800 275498
rect 588200 239818 588382 240054
rect 588618 239818 588800 240054
rect 588200 239734 588800 239818
rect 588200 239498 588382 239734
rect 588618 239498 588800 239734
rect 588200 204054 588800 239498
rect 588200 203818 588382 204054
rect 588618 203818 588800 204054
rect 588200 203734 588800 203818
rect 588200 203498 588382 203734
rect 588618 203498 588800 203734
rect 588200 168054 588800 203498
rect 588200 167818 588382 168054
rect 588618 167818 588800 168054
rect 588200 167734 588800 167818
rect 588200 167498 588382 167734
rect 588618 167498 588800 167734
rect 588200 132054 588800 167498
rect 588200 131818 588382 132054
rect 588618 131818 588800 132054
rect 588200 131734 588800 131818
rect 588200 131498 588382 131734
rect 588618 131498 588800 131734
rect 588200 96054 588800 131498
rect 588200 95818 588382 96054
rect 588618 95818 588800 96054
rect 588200 95734 588800 95818
rect 588200 95498 588382 95734
rect 588618 95498 588800 95734
rect 588200 60054 588800 95498
rect 588200 59818 588382 60054
rect 588618 59818 588800 60054
rect 588200 59734 588800 59818
rect 588200 59498 588382 59734
rect 588618 59498 588800 59734
rect 588200 24054 588800 59498
rect 588200 23818 588382 24054
rect 588618 23818 588800 24054
rect 588200 23734 588800 23818
rect 588200 23498 588382 23734
rect 588618 23498 588800 23734
rect 588200 -3226 588800 23498
rect 588200 -3462 588382 -3226
rect 588618 -3462 588800 -3226
rect 588200 -3546 588800 -3462
rect 588200 -3782 588382 -3546
rect 588618 -3782 588800 -3546
rect 588200 -3804 588800 -3782
<< via4 >>
rect -4694 707482 -4458 707718
rect -4694 707162 -4458 707398
rect -4694 671818 -4458 672054
rect -4694 671498 -4458 671734
rect -4694 635818 -4458 636054
rect -4694 635498 -4458 635734
rect -4694 599818 -4458 600054
rect -4694 599498 -4458 599734
rect -4694 563818 -4458 564054
rect -4694 563498 -4458 563734
rect -4694 527818 -4458 528054
rect -4694 527498 -4458 527734
rect -4694 491818 -4458 492054
rect -4694 491498 -4458 491734
rect -4694 455818 -4458 456054
rect -4694 455498 -4458 455734
rect -4694 419818 -4458 420054
rect -4694 419498 -4458 419734
rect -4694 383818 -4458 384054
rect -4694 383498 -4458 383734
rect -4694 347818 -4458 348054
rect -4694 347498 -4458 347734
rect -4694 311818 -4458 312054
rect -4694 311498 -4458 311734
rect -4694 275818 -4458 276054
rect -4694 275498 -4458 275734
rect -4694 239818 -4458 240054
rect -4694 239498 -4458 239734
rect -4694 203818 -4458 204054
rect -4694 203498 -4458 203734
rect -4694 167818 -4458 168054
rect -4694 167498 -4458 167734
rect -4694 131818 -4458 132054
rect -4694 131498 -4458 131734
rect -4694 95818 -4458 96054
rect -4694 95498 -4458 95734
rect -4694 59818 -4458 60054
rect -4694 59498 -4458 59734
rect -4694 23818 -4458 24054
rect -4694 23498 -4458 23734
rect -3734 706522 -3498 706758
rect -3734 706202 -3498 706438
rect 4586 706522 4822 706758
rect 4586 706202 4822 706438
rect -3734 689818 -3498 690054
rect -3734 689498 -3498 689734
rect -3734 653818 -3498 654054
rect -3734 653498 -3498 653734
rect -3734 617818 -3498 618054
rect -3734 617498 -3498 617734
rect -3734 581818 -3498 582054
rect -3734 581498 -3498 581734
rect -3734 545818 -3498 546054
rect -3734 545498 -3498 545734
rect -3734 509818 -3498 510054
rect -3734 509498 -3498 509734
rect -3734 473818 -3498 474054
rect -3734 473498 -3498 473734
rect -3734 437818 -3498 438054
rect -3734 437498 -3498 437734
rect -3734 401818 -3498 402054
rect -3734 401498 -3498 401734
rect -3734 365818 -3498 366054
rect -3734 365498 -3498 365734
rect -3734 329818 -3498 330054
rect -3734 329498 -3498 329734
rect -3734 293818 -3498 294054
rect -3734 293498 -3498 293734
rect -3734 257818 -3498 258054
rect -3734 257498 -3498 257734
rect -3734 221818 -3498 222054
rect -3734 221498 -3498 221734
rect -3734 185818 -3498 186054
rect -3734 185498 -3498 185734
rect -3734 149818 -3498 150054
rect -3734 149498 -3498 149734
rect -3734 113818 -3498 114054
rect -3734 113498 -3498 113734
rect -3734 77818 -3498 78054
rect -3734 77498 -3498 77734
rect -3734 41818 -3498 42054
rect -3734 41498 -3498 41734
rect -3734 5818 -3498 6054
rect -3734 5498 -3498 5734
rect -2774 705562 -2538 705798
rect -2774 705242 -2538 705478
rect -2774 668218 -2538 668454
rect -2774 667898 -2538 668134
rect -2774 632218 -2538 632454
rect -2774 631898 -2538 632134
rect -2774 596218 -2538 596454
rect -2774 595898 -2538 596134
rect -2774 560218 -2538 560454
rect -2774 559898 -2538 560134
rect -2774 524218 -2538 524454
rect -2774 523898 -2538 524134
rect -2774 488218 -2538 488454
rect -2774 487898 -2538 488134
rect -2774 452218 -2538 452454
rect -2774 451898 -2538 452134
rect -2774 416218 -2538 416454
rect -2774 415898 -2538 416134
rect -2774 380218 -2538 380454
rect -2774 379898 -2538 380134
rect -2774 344218 -2538 344454
rect -2774 343898 -2538 344134
rect -2774 308218 -2538 308454
rect -2774 307898 -2538 308134
rect -2774 272218 -2538 272454
rect -2774 271898 -2538 272134
rect -2774 236218 -2538 236454
rect -2774 235898 -2538 236134
rect -2774 200218 -2538 200454
rect -2774 199898 -2538 200134
rect -2774 164218 -2538 164454
rect -2774 163898 -2538 164134
rect -2774 128218 -2538 128454
rect -2774 127898 -2538 128134
rect -2774 92218 -2538 92454
rect -2774 91898 -2538 92134
rect -2774 56218 -2538 56454
rect -2774 55898 -2538 56134
rect -2774 20218 -2538 20454
rect -2774 19898 -2538 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2774 -1542 -2538 -1306
rect -2774 -1862 -2538 -1626
rect 22586 707482 22822 707718
rect 22586 707162 22822 707398
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3734 -2502 -3498 -2266
rect -3734 -2822 -3498 -2586
rect 18986 705562 19222 705798
rect 18986 705242 19222 705478
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1542 19222 -1306
rect 18986 -1862 19222 -1626
rect 40586 706522 40822 706758
rect 40586 706202 40822 706438
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 4586 -2502 4822 -2266
rect 4586 -2822 4822 -2586
rect -4694 -3462 -4458 -3226
rect -4694 -3782 -4458 -3546
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 58586 707482 58822 707718
rect 58586 707162 58822 707398
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 22586 -3462 22822 -3226
rect 22586 -3782 22822 -3546
rect 54986 705562 55222 705798
rect 54986 705242 55222 705478
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1542 55222 -1306
rect 54986 -1862 55222 -1626
rect 76586 706522 76822 706758
rect 76586 706202 76822 706438
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 94586 707482 94822 707718
rect 94586 707162 94822 707398
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 90986 705562 91222 705798
rect 90986 705242 91222 705478
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 112586 706522 112822 706758
rect 112586 706202 112822 706438
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 130586 707482 130822 707718
rect 130586 707162 130822 707398
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 126986 705562 127222 705798
rect 126986 705242 127222 705478
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 148586 706522 148822 706758
rect 148586 706202 148822 706438
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 166586 707482 166822 707718
rect 166586 707162 166822 707398
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 162986 705562 163222 705798
rect 162986 705242 163222 705478
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 184586 706522 184822 706758
rect 184586 706202 184822 706438
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 202586 707482 202822 707718
rect 202586 707162 202822 707398
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 198986 705562 199222 705798
rect 198986 705242 199222 705478
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 220586 706522 220822 706758
rect 220586 706202 220822 706438
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 238586 707482 238822 707718
rect 238586 707162 238822 707398
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 234986 705562 235222 705798
rect 234986 705242 235222 705478
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 256586 706522 256822 706758
rect 256586 706202 256822 706438
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 274586 707482 274822 707718
rect 274586 707162 274822 707398
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 270986 705562 271222 705798
rect 270986 705242 271222 705478
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 292586 706522 292822 706758
rect 292586 706202 292822 706438
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 310586 707482 310822 707718
rect 310586 707162 310822 707398
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 306986 705562 307222 705798
rect 306986 705242 307222 705478
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 328586 706522 328822 706758
rect 328586 706202 328822 706438
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 346586 707482 346822 707718
rect 346586 707162 346822 707398
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 342986 705562 343222 705798
rect 342986 705242 343222 705478
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 364586 706522 364822 706758
rect 364586 706202 364822 706438
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 382586 707482 382822 707718
rect 382586 707162 382822 707398
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 378986 705562 379222 705798
rect 378986 705242 379222 705478
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 400586 706522 400822 706758
rect 400586 706202 400822 706438
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 418586 707482 418822 707718
rect 418586 707162 418822 707398
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 414986 705562 415222 705798
rect 414986 705242 415222 705478
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 436586 706522 436822 706758
rect 436586 706202 436822 706438
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 454586 707482 454822 707718
rect 454586 707162 454822 707398
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 450986 705562 451222 705798
rect 450986 705242 451222 705478
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 472586 706522 472822 706758
rect 472586 706202 472822 706438
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 490586 707482 490822 707718
rect 490586 707162 490822 707398
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 486986 705562 487222 705798
rect 486986 705242 487222 705478
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 508586 706522 508822 706758
rect 508586 706202 508822 706438
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 526586 707482 526822 707718
rect 526586 707162 526822 707398
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 522986 705562 523222 705798
rect 522986 705242 523222 705478
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 81610 635818 81846 636054
rect 81610 635498 81846 635734
rect 81610 632218 81846 632454
rect 81610 631898 81846 632134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 66250 617818 66486 618054
rect 66250 617498 66486 617734
rect 66250 614218 66486 614454
rect 66250 613898 66486 614134
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 81610 599818 81846 600054
rect 81610 599498 81846 599734
rect 81610 596218 81846 596454
rect 81610 595898 81846 596134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 66250 581818 66486 582054
rect 66250 581498 66486 581734
rect 66250 578218 66486 578454
rect 66250 577898 66486 578134
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 81610 563818 81846 564054
rect 81610 563498 81846 563734
rect 81610 560218 81846 560454
rect 81610 559898 81846 560134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 66250 545818 66486 546054
rect 66250 545498 66486 545734
rect 66250 542218 66486 542454
rect 66250 541898 66486 542134
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 81610 527818 81846 528054
rect 81610 527498 81846 527734
rect 81610 524218 81846 524454
rect 81610 523898 81846 524134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 66250 509818 66486 510054
rect 66250 509498 66486 509734
rect 66250 506218 66486 506454
rect 66250 505898 66486 506134
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 81610 491818 81846 492054
rect 81610 491498 81846 491734
rect 81610 488218 81846 488454
rect 81610 487898 81846 488134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 66250 473818 66486 474054
rect 66250 473498 66486 473734
rect 66250 470218 66486 470454
rect 66250 469898 66486 470134
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 81610 455818 81846 456054
rect 81610 455498 81846 455734
rect 81610 452218 81846 452454
rect 81610 451898 81846 452134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 66250 437818 66486 438054
rect 66250 437498 66486 437734
rect 66250 434218 66486 434454
rect 66250 433898 66486 434134
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 81610 419818 81846 420054
rect 81610 419498 81846 419734
rect 81610 416218 81846 416454
rect 81610 415898 81846 416134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 66250 401818 66486 402054
rect 66250 401498 66486 401734
rect 66250 398218 66486 398454
rect 66250 397898 66486 398134
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 81610 383818 81846 384054
rect 81610 383498 81846 383734
rect 81610 380218 81846 380454
rect 81610 379898 81846 380134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 66250 365818 66486 366054
rect 66250 365498 66486 365734
rect 66250 362218 66486 362454
rect 66250 361898 66486 362134
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 81610 347818 81846 348054
rect 81610 347498 81846 347734
rect 81610 344218 81846 344454
rect 81610 343898 81846 344134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 66250 329818 66486 330054
rect 66250 329498 66486 329734
rect 66250 326218 66486 326454
rect 66250 325898 66486 326134
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 81610 311818 81846 312054
rect 81610 311498 81846 311734
rect 81610 308218 81846 308454
rect 81610 307898 81846 308134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 66250 293818 66486 294054
rect 66250 293498 66486 293734
rect 66250 290218 66486 290454
rect 66250 289898 66486 290134
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 81610 275818 81846 276054
rect 81610 275498 81846 275734
rect 81610 272218 81846 272454
rect 81610 271898 81846 272134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 66250 257818 66486 258054
rect 66250 257498 66486 257734
rect 66250 254218 66486 254454
rect 66250 253898 66486 254134
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 81610 239818 81846 240054
rect 81610 239498 81846 239734
rect 81610 236218 81846 236454
rect 81610 235898 81846 236134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 66250 221818 66486 222054
rect 66250 221498 66486 221734
rect 66250 218218 66486 218454
rect 66250 217898 66486 218134
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 81610 203818 81846 204054
rect 81610 203498 81846 203734
rect 81610 200218 81846 200454
rect 81610 199898 81846 200134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 66250 185818 66486 186054
rect 66250 185498 66486 185734
rect 66250 182218 66486 182454
rect 66250 181898 66486 182134
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 81610 167818 81846 168054
rect 81610 167498 81846 167734
rect 81610 164218 81846 164454
rect 81610 163898 81846 164134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 66250 149818 66486 150054
rect 66250 149498 66486 149734
rect 66250 146218 66486 146454
rect 66250 145898 66486 146134
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 81610 131818 81846 132054
rect 81610 131498 81846 131734
rect 81610 128218 81846 128454
rect 81610 127898 81846 128134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 66250 113818 66486 114054
rect 66250 113498 66486 113734
rect 66250 110218 66486 110454
rect 66250 109898 66486 110134
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 81610 95818 81846 96054
rect 81610 95498 81846 95734
rect 81610 92218 81846 92454
rect 81610 91898 81846 92134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 66250 77818 66486 78054
rect 66250 77498 66486 77734
rect 66250 74218 66486 74454
rect 66250 73898 66486 74134
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 81610 59818 81846 60054
rect 81610 59498 81846 59734
rect 81610 56218 81846 56454
rect 81610 55898 81846 56134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 40586 -2502 40822 -2266
rect 40586 -2822 40822 -2586
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 58586 -3462 58822 -3226
rect 58586 -3782 58822 -3546
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1542 91222 -1306
rect 90986 -1862 91222 -1626
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 76586 -2502 76822 -2266
rect 76586 -2822 76822 -2586
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 94586 -3462 94822 -3226
rect 94586 -3782 94822 -3546
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1542 127222 -1306
rect 126986 -1862 127222 -1626
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 112586 -2502 112822 -2266
rect 112586 -2822 112822 -2586
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 130586 -3462 130822 -3226
rect 130586 -3782 130822 -3546
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1542 163222 -1306
rect 162986 -1862 163222 -1626
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 148586 -2502 148822 -2266
rect 148586 -2822 148822 -2586
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 166586 -3462 166822 -3226
rect 166586 -3782 166822 -3546
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1542 199222 -1306
rect 198986 -1862 199222 -1626
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 184586 -2502 184822 -2266
rect 184586 -2822 184822 -2586
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 202586 -3462 202822 -3226
rect 202586 -3782 202822 -3546
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1542 235222 -1306
rect 234986 -1862 235222 -1626
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 220586 -2502 220822 -2266
rect 220586 -2822 220822 -2586
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 238586 -3462 238822 -3226
rect 238586 -3782 238822 -3546
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1542 271222 -1306
rect 270986 -1862 271222 -1626
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 256586 -2502 256822 -2266
rect 256586 -2822 256822 -2586
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 274586 -3462 274822 -3226
rect 274586 -3782 274822 -3546
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1542 307222 -1306
rect 306986 -1862 307222 -1626
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 292586 -2502 292822 -2266
rect 292586 -2822 292822 -2586
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 310586 -3462 310822 -3226
rect 310586 -3782 310822 -3546
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1542 343222 -1306
rect 342986 -1862 343222 -1626
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 328586 -2502 328822 -2266
rect 328586 -2822 328822 -2586
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 346586 -3462 346822 -3226
rect 346586 -3782 346822 -3546
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1542 379222 -1306
rect 378986 -1862 379222 -1626
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 364586 -2502 364822 -2266
rect 364586 -2822 364822 -2586
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 382586 -3462 382822 -3226
rect 382586 -3782 382822 -3546
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1542 415222 -1306
rect 414986 -1862 415222 -1626
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 400586 -2502 400822 -2266
rect 400586 -2822 400822 -2586
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 418586 -3462 418822 -3226
rect 418586 -3782 418822 -3546
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1542 451222 -1306
rect 450986 -1862 451222 -1626
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 436586 -2502 436822 -2266
rect 436586 -2822 436822 -2586
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 454586 -3462 454822 -3226
rect 454586 -3782 454822 -3546
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1542 487222 -1306
rect 486986 -1862 487222 -1626
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 472586 -2502 472822 -2266
rect 472586 -2822 472822 -2586
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 490586 -3462 490822 -3226
rect 490586 -3782 490822 -3546
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1542 523222 -1306
rect 522986 -1862 523222 -1626
rect 544586 706522 544822 706758
rect 544586 706202 544822 706438
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 508586 -2502 508822 -2266
rect 508586 -2822 508822 -2586
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 562586 707482 562822 707718
rect 562586 707162 562822 707398
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 526586 -3462 526822 -3226
rect 526586 -3782 526822 -3546
rect 558986 705562 559222 705798
rect 558986 705242 559222 705478
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1542 559222 -1306
rect 558986 -1862 559222 -1626
rect 588382 707482 588618 707718
rect 588382 707162 588618 707398
rect 580586 706522 580822 706758
rect 580586 706202 580822 706438
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 544586 -2502 544822 -2266
rect 544586 -2822 544822 -2586
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587422 706522 587658 706758
rect 587422 706202 587658 706438
rect 586462 705562 586698 705798
rect 586462 705242 586698 705478
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 562586 -3462 562822 -3226
rect 562586 -3782 562822 -3546
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586462 668218 586698 668454
rect 586462 667898 586698 668134
rect 586462 632218 586698 632454
rect 586462 631898 586698 632134
rect 586462 596218 586698 596454
rect 586462 595898 586698 596134
rect 586462 560218 586698 560454
rect 586462 559898 586698 560134
rect 586462 524218 586698 524454
rect 586462 523898 586698 524134
rect 586462 488218 586698 488454
rect 586462 487898 586698 488134
rect 586462 452218 586698 452454
rect 586462 451898 586698 452134
rect 586462 416218 586698 416454
rect 586462 415898 586698 416134
rect 586462 380218 586698 380454
rect 586462 379898 586698 380134
rect 586462 344218 586698 344454
rect 586462 343898 586698 344134
rect 586462 308218 586698 308454
rect 586462 307898 586698 308134
rect 586462 272218 586698 272454
rect 586462 271898 586698 272134
rect 586462 236218 586698 236454
rect 586462 235898 586698 236134
rect 586462 200218 586698 200454
rect 586462 199898 586698 200134
rect 586462 164218 586698 164454
rect 586462 163898 586698 164134
rect 586462 128218 586698 128454
rect 586462 127898 586698 128134
rect 586462 92218 586698 92454
rect 586462 91898 586698 92134
rect 586462 56218 586698 56454
rect 586462 55898 586698 56134
rect 586462 20218 586698 20454
rect 586462 19898 586698 20134
rect 586462 -1542 586698 -1306
rect 586462 -1862 586698 -1626
rect 587422 689818 587658 690054
rect 587422 689498 587658 689734
rect 587422 653818 587658 654054
rect 587422 653498 587658 653734
rect 587422 617818 587658 618054
rect 587422 617498 587658 617734
rect 587422 581818 587658 582054
rect 587422 581498 587658 581734
rect 587422 545818 587658 546054
rect 587422 545498 587658 545734
rect 587422 509818 587658 510054
rect 587422 509498 587658 509734
rect 587422 473818 587658 474054
rect 587422 473498 587658 473734
rect 587422 437818 587658 438054
rect 587422 437498 587658 437734
rect 587422 401818 587658 402054
rect 587422 401498 587658 401734
rect 587422 365818 587658 366054
rect 587422 365498 587658 365734
rect 587422 329818 587658 330054
rect 587422 329498 587658 329734
rect 587422 293818 587658 294054
rect 587422 293498 587658 293734
rect 587422 257818 587658 258054
rect 587422 257498 587658 257734
rect 587422 221818 587658 222054
rect 587422 221498 587658 221734
rect 587422 185818 587658 186054
rect 587422 185498 587658 185734
rect 587422 149818 587658 150054
rect 587422 149498 587658 149734
rect 587422 113818 587658 114054
rect 587422 113498 587658 113734
rect 587422 77818 587658 78054
rect 587422 77498 587658 77734
rect 587422 41818 587658 42054
rect 587422 41498 587658 41734
rect 587422 5818 587658 6054
rect 587422 5498 587658 5734
rect 580586 -2502 580822 -2266
rect 580586 -2822 580822 -2586
rect 587422 -2502 587658 -2266
rect 587422 -2822 587658 -2586
rect 588382 671818 588618 672054
rect 588382 671498 588618 671734
rect 588382 635818 588618 636054
rect 588382 635498 588618 635734
rect 588382 599818 588618 600054
rect 588382 599498 588618 599734
rect 588382 563818 588618 564054
rect 588382 563498 588618 563734
rect 588382 527818 588618 528054
rect 588382 527498 588618 527734
rect 588382 491818 588618 492054
rect 588382 491498 588618 491734
rect 588382 455818 588618 456054
rect 588382 455498 588618 455734
rect 588382 419818 588618 420054
rect 588382 419498 588618 419734
rect 588382 383818 588618 384054
rect 588382 383498 588618 383734
rect 588382 347818 588618 348054
rect 588382 347498 588618 347734
rect 588382 311818 588618 312054
rect 588382 311498 588618 311734
rect 588382 275818 588618 276054
rect 588382 275498 588618 275734
rect 588382 239818 588618 240054
rect 588382 239498 588618 239734
rect 588382 203818 588618 204054
rect 588382 203498 588618 203734
rect 588382 167818 588618 168054
rect 588382 167498 588618 167734
rect 588382 131818 588618 132054
rect 588382 131498 588618 131734
rect 588382 95818 588618 96054
rect 588382 95498 588618 95734
rect 588382 59818 588618 60054
rect 588382 59498 588618 59734
rect 588382 23818 588618 24054
rect 588382 23498 588618 23734
rect 588382 -3462 588618 -3226
rect 588382 -3782 588618 -3546
<< metal5 >>
rect -4876 707740 -4276 707742
rect 22404 707740 23004 707742
rect 58404 707740 59004 707742
rect 94404 707740 95004 707742
rect 130404 707740 131004 707742
rect 166404 707740 167004 707742
rect 202404 707740 203004 707742
rect 238404 707740 239004 707742
rect 274404 707740 275004 707742
rect 310404 707740 311004 707742
rect 346404 707740 347004 707742
rect 382404 707740 383004 707742
rect 418404 707740 419004 707742
rect 454404 707740 455004 707742
rect 490404 707740 491004 707742
rect 526404 707740 527004 707742
rect 562404 707740 563004 707742
rect 588200 707740 588800 707742
rect -4876 707718 588800 707740
rect -4876 707482 -4694 707718
rect -4458 707482 22586 707718
rect 22822 707482 58586 707718
rect 58822 707482 94586 707718
rect 94822 707482 130586 707718
rect 130822 707482 166586 707718
rect 166822 707482 202586 707718
rect 202822 707482 238586 707718
rect 238822 707482 274586 707718
rect 274822 707482 310586 707718
rect 310822 707482 346586 707718
rect 346822 707482 382586 707718
rect 382822 707482 418586 707718
rect 418822 707482 454586 707718
rect 454822 707482 490586 707718
rect 490822 707482 526586 707718
rect 526822 707482 562586 707718
rect 562822 707482 588382 707718
rect 588618 707482 588800 707718
rect -4876 707398 588800 707482
rect -4876 707162 -4694 707398
rect -4458 707162 22586 707398
rect 22822 707162 58586 707398
rect 58822 707162 94586 707398
rect 94822 707162 130586 707398
rect 130822 707162 166586 707398
rect 166822 707162 202586 707398
rect 202822 707162 238586 707398
rect 238822 707162 274586 707398
rect 274822 707162 310586 707398
rect 310822 707162 346586 707398
rect 346822 707162 382586 707398
rect 382822 707162 418586 707398
rect 418822 707162 454586 707398
rect 454822 707162 490586 707398
rect 490822 707162 526586 707398
rect 526822 707162 562586 707398
rect 562822 707162 588382 707398
rect 588618 707162 588800 707398
rect -4876 707140 588800 707162
rect -4876 707138 -4276 707140
rect 22404 707138 23004 707140
rect 58404 707138 59004 707140
rect 94404 707138 95004 707140
rect 130404 707138 131004 707140
rect 166404 707138 167004 707140
rect 202404 707138 203004 707140
rect 238404 707138 239004 707140
rect 274404 707138 275004 707140
rect 310404 707138 311004 707140
rect 346404 707138 347004 707140
rect 382404 707138 383004 707140
rect 418404 707138 419004 707140
rect 454404 707138 455004 707140
rect 490404 707138 491004 707140
rect 526404 707138 527004 707140
rect 562404 707138 563004 707140
rect 588200 707138 588800 707140
rect -3916 706780 -3316 706782
rect 4404 706780 5004 706782
rect 40404 706780 41004 706782
rect 76404 706780 77004 706782
rect 112404 706780 113004 706782
rect 148404 706780 149004 706782
rect 184404 706780 185004 706782
rect 220404 706780 221004 706782
rect 256404 706780 257004 706782
rect 292404 706780 293004 706782
rect 328404 706780 329004 706782
rect 364404 706780 365004 706782
rect 400404 706780 401004 706782
rect 436404 706780 437004 706782
rect 472404 706780 473004 706782
rect 508404 706780 509004 706782
rect 544404 706780 545004 706782
rect 580404 706780 581004 706782
rect 587240 706780 587840 706782
rect -3916 706758 587840 706780
rect -3916 706522 -3734 706758
rect -3498 706522 4586 706758
rect 4822 706522 40586 706758
rect 40822 706522 76586 706758
rect 76822 706522 112586 706758
rect 112822 706522 148586 706758
rect 148822 706522 184586 706758
rect 184822 706522 220586 706758
rect 220822 706522 256586 706758
rect 256822 706522 292586 706758
rect 292822 706522 328586 706758
rect 328822 706522 364586 706758
rect 364822 706522 400586 706758
rect 400822 706522 436586 706758
rect 436822 706522 472586 706758
rect 472822 706522 508586 706758
rect 508822 706522 544586 706758
rect 544822 706522 580586 706758
rect 580822 706522 587422 706758
rect 587658 706522 587840 706758
rect -3916 706438 587840 706522
rect -3916 706202 -3734 706438
rect -3498 706202 4586 706438
rect 4822 706202 40586 706438
rect 40822 706202 76586 706438
rect 76822 706202 112586 706438
rect 112822 706202 148586 706438
rect 148822 706202 184586 706438
rect 184822 706202 220586 706438
rect 220822 706202 256586 706438
rect 256822 706202 292586 706438
rect 292822 706202 328586 706438
rect 328822 706202 364586 706438
rect 364822 706202 400586 706438
rect 400822 706202 436586 706438
rect 436822 706202 472586 706438
rect 472822 706202 508586 706438
rect 508822 706202 544586 706438
rect 544822 706202 580586 706438
rect 580822 706202 587422 706438
rect 587658 706202 587840 706438
rect -3916 706180 587840 706202
rect -3916 706178 -3316 706180
rect 4404 706178 5004 706180
rect 40404 706178 41004 706180
rect 76404 706178 77004 706180
rect 112404 706178 113004 706180
rect 148404 706178 149004 706180
rect 184404 706178 185004 706180
rect 220404 706178 221004 706180
rect 256404 706178 257004 706180
rect 292404 706178 293004 706180
rect 328404 706178 329004 706180
rect 364404 706178 365004 706180
rect 400404 706178 401004 706180
rect 436404 706178 437004 706180
rect 472404 706178 473004 706180
rect 508404 706178 509004 706180
rect 544404 706178 545004 706180
rect 580404 706178 581004 706180
rect 587240 706178 587840 706180
rect -2956 705820 -2356 705822
rect 18804 705820 19404 705822
rect 54804 705820 55404 705822
rect 90804 705820 91404 705822
rect 126804 705820 127404 705822
rect 162804 705820 163404 705822
rect 198804 705820 199404 705822
rect 234804 705820 235404 705822
rect 270804 705820 271404 705822
rect 306804 705820 307404 705822
rect 342804 705820 343404 705822
rect 378804 705820 379404 705822
rect 414804 705820 415404 705822
rect 450804 705820 451404 705822
rect 486804 705820 487404 705822
rect 522804 705820 523404 705822
rect 558804 705820 559404 705822
rect 586280 705820 586880 705822
rect -2956 705798 586880 705820
rect -2956 705562 -2774 705798
rect -2538 705562 18986 705798
rect 19222 705562 54986 705798
rect 55222 705562 90986 705798
rect 91222 705562 126986 705798
rect 127222 705562 162986 705798
rect 163222 705562 198986 705798
rect 199222 705562 234986 705798
rect 235222 705562 270986 705798
rect 271222 705562 306986 705798
rect 307222 705562 342986 705798
rect 343222 705562 378986 705798
rect 379222 705562 414986 705798
rect 415222 705562 450986 705798
rect 451222 705562 486986 705798
rect 487222 705562 522986 705798
rect 523222 705562 558986 705798
rect 559222 705562 586462 705798
rect 586698 705562 586880 705798
rect -2956 705478 586880 705562
rect -2956 705242 -2774 705478
rect -2538 705242 18986 705478
rect 19222 705242 54986 705478
rect 55222 705242 90986 705478
rect 91222 705242 126986 705478
rect 127222 705242 162986 705478
rect 163222 705242 198986 705478
rect 199222 705242 234986 705478
rect 235222 705242 270986 705478
rect 271222 705242 306986 705478
rect 307222 705242 342986 705478
rect 343222 705242 378986 705478
rect 379222 705242 414986 705478
rect 415222 705242 450986 705478
rect 451222 705242 486986 705478
rect 487222 705242 522986 705478
rect 523222 705242 558986 705478
rect 559222 705242 586462 705478
rect 586698 705242 586880 705478
rect -2956 705220 586880 705242
rect -2956 705218 -2356 705220
rect 18804 705218 19404 705220
rect 54804 705218 55404 705220
rect 90804 705218 91404 705220
rect 126804 705218 127404 705220
rect 162804 705218 163404 705220
rect 198804 705218 199404 705220
rect 234804 705218 235404 705220
rect 270804 705218 271404 705220
rect 306804 705218 307404 705220
rect 342804 705218 343404 705220
rect 378804 705218 379404 705220
rect 414804 705218 415404 705220
rect 450804 705218 451404 705220
rect 486804 705218 487404 705220
rect 522804 705218 523404 705220
rect 558804 705218 559404 705220
rect 586280 705218 586880 705220
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -3916 690076 -3316 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587240 690076 587840 690078
rect -4876 690054 588800 690076
rect -4876 689818 -3734 690054
rect -3498 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587422 690054
rect 587658 689818 588800 690054
rect -4876 689734 588800 689818
rect -4876 689498 -3734 689734
rect -3498 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587422 689734
rect 587658 689498 588800 689734
rect -4876 689476 588800 689498
rect -3916 689474 -3316 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587240 689474 587840 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2956 686454 586880 686476
rect -2956 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586880 686454
rect -2956 686134 586880 686218
rect -2956 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586880 686134
rect -2956 685876 586880 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -4876 672076 -4276 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588200 672076 588800 672078
rect -4876 672054 588800 672076
rect -4876 671818 -4694 672054
rect -4458 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588382 672054
rect 588618 671818 588800 672054
rect -4876 671734 588800 671818
rect -4876 671498 -4694 671734
rect -4458 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588382 671734
rect 588618 671498 588800 671734
rect -4876 671476 588800 671498
rect -4876 671474 -4276 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588200 671474 588800 671476
rect -2956 668476 -2356 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586280 668476 586880 668478
rect -2956 668454 586880 668476
rect -2956 668218 -2774 668454
rect -2538 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586462 668454
rect 586698 668218 586880 668454
rect -2956 668134 586880 668218
rect -2956 667898 -2774 668134
rect -2538 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586462 668134
rect 586698 667898 586880 668134
rect -2956 667876 586880 667898
rect -2956 667874 -2356 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586280 667874 586880 667876
rect -3916 654076 -3316 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587240 654076 587840 654078
rect -4876 654054 588800 654076
rect -4876 653818 -3734 654054
rect -3498 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587422 654054
rect 587658 653818 588800 654054
rect -4876 653734 588800 653818
rect -4876 653498 -3734 653734
rect -3498 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587422 653734
rect 587658 653498 588800 653734
rect -4876 653476 588800 653498
rect -3916 653474 -3316 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587240 653474 587840 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2956 650454 586880 650476
rect -2956 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586880 650454
rect -2956 650134 586880 650218
rect -2956 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586880 650134
rect -2956 649876 586880 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -4876 636076 -4276 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 81568 636076 81888 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588200 636076 588800 636078
rect -4876 636054 588800 636076
rect -4876 635818 -4694 636054
rect -4458 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 81610 636054
rect 81846 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588382 636054
rect 588618 635818 588800 636054
rect -4876 635734 588800 635818
rect -4876 635498 -4694 635734
rect -4458 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 81610 635734
rect 81846 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588382 635734
rect 588618 635498 588800 635734
rect -4876 635476 588800 635498
rect -4876 635474 -4276 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 81568 635474 81888 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588200 635474 588800 635476
rect -2956 632476 -2356 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 81568 632476 81888 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586280 632476 586880 632478
rect -2956 632454 586880 632476
rect -2956 632218 -2774 632454
rect -2538 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 81610 632454
rect 81846 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586462 632454
rect 586698 632218 586880 632454
rect -2956 632134 586880 632218
rect -2956 631898 -2774 632134
rect -2538 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 81610 632134
rect 81846 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586462 632134
rect 586698 631898 586880 632134
rect -2956 631876 586880 631898
rect -2956 631874 -2356 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 81568 631874 81888 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586280 631874 586880 631876
rect -3916 618076 -3316 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 66208 618076 66528 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587240 618076 587840 618078
rect -4876 618054 588800 618076
rect -4876 617818 -3734 618054
rect -3498 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 66250 618054
rect 66486 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587422 618054
rect 587658 617818 588800 618054
rect -4876 617734 588800 617818
rect -4876 617498 -3734 617734
rect -3498 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 66250 617734
rect 66486 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587422 617734
rect 587658 617498 588800 617734
rect -4876 617476 588800 617498
rect -3916 617474 -3316 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 66208 617474 66528 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587240 617474 587840 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 66208 614476 66528 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2956 614454 586880 614476
rect -2956 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 66250 614454
rect 66486 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586880 614454
rect -2956 614134 586880 614218
rect -2956 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 66250 614134
rect 66486 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586880 614134
rect -2956 613876 586880 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 66208 613874 66528 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -4876 600076 -4276 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 81568 600076 81888 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588200 600076 588800 600078
rect -4876 600054 588800 600076
rect -4876 599818 -4694 600054
rect -4458 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 81610 600054
rect 81846 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588382 600054
rect 588618 599818 588800 600054
rect -4876 599734 588800 599818
rect -4876 599498 -4694 599734
rect -4458 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 81610 599734
rect 81846 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588382 599734
rect 588618 599498 588800 599734
rect -4876 599476 588800 599498
rect -4876 599474 -4276 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 81568 599474 81888 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588200 599474 588800 599476
rect -2956 596476 -2356 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 81568 596476 81888 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586280 596476 586880 596478
rect -2956 596454 586880 596476
rect -2956 596218 -2774 596454
rect -2538 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 81610 596454
rect 81846 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586462 596454
rect 586698 596218 586880 596454
rect -2956 596134 586880 596218
rect -2956 595898 -2774 596134
rect -2538 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 81610 596134
rect 81846 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586462 596134
rect 586698 595898 586880 596134
rect -2956 595876 586880 595898
rect -2956 595874 -2356 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 81568 595874 81888 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586280 595874 586880 595876
rect -3916 582076 -3316 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 66208 582076 66528 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587240 582076 587840 582078
rect -4876 582054 588800 582076
rect -4876 581818 -3734 582054
rect -3498 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 66250 582054
rect 66486 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587422 582054
rect 587658 581818 588800 582054
rect -4876 581734 588800 581818
rect -4876 581498 -3734 581734
rect -3498 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 66250 581734
rect 66486 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587422 581734
rect 587658 581498 588800 581734
rect -4876 581476 588800 581498
rect -3916 581474 -3316 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 66208 581474 66528 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587240 581474 587840 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 66208 578476 66528 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2956 578454 586880 578476
rect -2956 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 66250 578454
rect 66486 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586880 578454
rect -2956 578134 586880 578218
rect -2956 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 66250 578134
rect 66486 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586880 578134
rect -2956 577876 586880 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 66208 577874 66528 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -4876 564076 -4276 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 81568 564076 81888 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588200 564076 588800 564078
rect -4876 564054 588800 564076
rect -4876 563818 -4694 564054
rect -4458 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 81610 564054
rect 81846 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588382 564054
rect 588618 563818 588800 564054
rect -4876 563734 588800 563818
rect -4876 563498 -4694 563734
rect -4458 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 81610 563734
rect 81846 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588382 563734
rect 588618 563498 588800 563734
rect -4876 563476 588800 563498
rect -4876 563474 -4276 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 81568 563474 81888 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588200 563474 588800 563476
rect -2956 560476 -2356 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 81568 560476 81888 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586280 560476 586880 560478
rect -2956 560454 586880 560476
rect -2956 560218 -2774 560454
rect -2538 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 81610 560454
rect 81846 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586462 560454
rect 586698 560218 586880 560454
rect -2956 560134 586880 560218
rect -2956 559898 -2774 560134
rect -2538 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 81610 560134
rect 81846 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586462 560134
rect 586698 559898 586880 560134
rect -2956 559876 586880 559898
rect -2956 559874 -2356 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 81568 559874 81888 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586280 559874 586880 559876
rect -3916 546076 -3316 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 66208 546076 66528 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587240 546076 587840 546078
rect -4876 546054 588800 546076
rect -4876 545818 -3734 546054
rect -3498 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 66250 546054
rect 66486 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587422 546054
rect 587658 545818 588800 546054
rect -4876 545734 588800 545818
rect -4876 545498 -3734 545734
rect -3498 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 66250 545734
rect 66486 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587422 545734
rect 587658 545498 588800 545734
rect -4876 545476 588800 545498
rect -3916 545474 -3316 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 66208 545474 66528 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587240 545474 587840 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 66208 542476 66528 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2956 542454 586880 542476
rect -2956 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 66250 542454
rect 66486 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586880 542454
rect -2956 542134 586880 542218
rect -2956 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 66250 542134
rect 66486 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586880 542134
rect -2956 541876 586880 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 66208 541874 66528 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -4876 528076 -4276 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 81568 528076 81888 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588200 528076 588800 528078
rect -4876 528054 588800 528076
rect -4876 527818 -4694 528054
rect -4458 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 81610 528054
rect 81846 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588382 528054
rect 588618 527818 588800 528054
rect -4876 527734 588800 527818
rect -4876 527498 -4694 527734
rect -4458 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 81610 527734
rect 81846 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588382 527734
rect 588618 527498 588800 527734
rect -4876 527476 588800 527498
rect -4876 527474 -4276 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 81568 527474 81888 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588200 527474 588800 527476
rect -2956 524476 -2356 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 81568 524476 81888 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586280 524476 586880 524478
rect -2956 524454 586880 524476
rect -2956 524218 -2774 524454
rect -2538 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 81610 524454
rect 81846 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586462 524454
rect 586698 524218 586880 524454
rect -2956 524134 586880 524218
rect -2956 523898 -2774 524134
rect -2538 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 81610 524134
rect 81846 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586462 524134
rect 586698 523898 586880 524134
rect -2956 523876 586880 523898
rect -2956 523874 -2356 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 81568 523874 81888 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586280 523874 586880 523876
rect -3916 510076 -3316 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 66208 510076 66528 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587240 510076 587840 510078
rect -4876 510054 588800 510076
rect -4876 509818 -3734 510054
rect -3498 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 66250 510054
rect 66486 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587422 510054
rect 587658 509818 588800 510054
rect -4876 509734 588800 509818
rect -4876 509498 -3734 509734
rect -3498 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 66250 509734
rect 66486 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587422 509734
rect 587658 509498 588800 509734
rect -4876 509476 588800 509498
rect -3916 509474 -3316 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 66208 509474 66528 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587240 509474 587840 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 66208 506476 66528 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2956 506454 586880 506476
rect -2956 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 66250 506454
rect 66486 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586880 506454
rect -2956 506134 586880 506218
rect -2956 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 66250 506134
rect 66486 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586880 506134
rect -2956 505876 586880 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 66208 505874 66528 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -4876 492076 -4276 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 81568 492076 81888 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588200 492076 588800 492078
rect -4876 492054 588800 492076
rect -4876 491818 -4694 492054
rect -4458 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 81610 492054
rect 81846 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588382 492054
rect 588618 491818 588800 492054
rect -4876 491734 588800 491818
rect -4876 491498 -4694 491734
rect -4458 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 81610 491734
rect 81846 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588382 491734
rect 588618 491498 588800 491734
rect -4876 491476 588800 491498
rect -4876 491474 -4276 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 81568 491474 81888 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588200 491474 588800 491476
rect -2956 488476 -2356 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 81568 488476 81888 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586280 488476 586880 488478
rect -2956 488454 586880 488476
rect -2956 488218 -2774 488454
rect -2538 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 81610 488454
rect 81846 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586462 488454
rect 586698 488218 586880 488454
rect -2956 488134 586880 488218
rect -2956 487898 -2774 488134
rect -2538 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 81610 488134
rect 81846 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586462 488134
rect 586698 487898 586880 488134
rect -2956 487876 586880 487898
rect -2956 487874 -2356 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 81568 487874 81888 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586280 487874 586880 487876
rect -3916 474076 -3316 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 66208 474076 66528 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587240 474076 587840 474078
rect -4876 474054 588800 474076
rect -4876 473818 -3734 474054
rect -3498 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 66250 474054
rect 66486 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587422 474054
rect 587658 473818 588800 474054
rect -4876 473734 588800 473818
rect -4876 473498 -3734 473734
rect -3498 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 66250 473734
rect 66486 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587422 473734
rect 587658 473498 588800 473734
rect -4876 473476 588800 473498
rect -3916 473474 -3316 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 66208 473474 66528 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587240 473474 587840 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 66208 470476 66528 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2956 470454 586880 470476
rect -2956 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 66250 470454
rect 66486 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586880 470454
rect -2956 470134 586880 470218
rect -2956 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 66250 470134
rect 66486 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586880 470134
rect -2956 469876 586880 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 66208 469874 66528 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -4876 456076 -4276 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 81568 456076 81888 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588200 456076 588800 456078
rect -4876 456054 588800 456076
rect -4876 455818 -4694 456054
rect -4458 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 81610 456054
rect 81846 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588382 456054
rect 588618 455818 588800 456054
rect -4876 455734 588800 455818
rect -4876 455498 -4694 455734
rect -4458 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 81610 455734
rect 81846 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588382 455734
rect 588618 455498 588800 455734
rect -4876 455476 588800 455498
rect -4876 455474 -4276 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 81568 455474 81888 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588200 455474 588800 455476
rect -2956 452476 -2356 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 81568 452476 81888 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586280 452476 586880 452478
rect -2956 452454 586880 452476
rect -2956 452218 -2774 452454
rect -2538 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 81610 452454
rect 81846 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586462 452454
rect 586698 452218 586880 452454
rect -2956 452134 586880 452218
rect -2956 451898 -2774 452134
rect -2538 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 81610 452134
rect 81846 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586462 452134
rect 586698 451898 586880 452134
rect -2956 451876 586880 451898
rect -2956 451874 -2356 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 81568 451874 81888 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586280 451874 586880 451876
rect -3916 438076 -3316 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 66208 438076 66528 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587240 438076 587840 438078
rect -4876 438054 588800 438076
rect -4876 437818 -3734 438054
rect -3498 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 66250 438054
rect 66486 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587422 438054
rect 587658 437818 588800 438054
rect -4876 437734 588800 437818
rect -4876 437498 -3734 437734
rect -3498 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 66250 437734
rect 66486 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587422 437734
rect 587658 437498 588800 437734
rect -4876 437476 588800 437498
rect -3916 437474 -3316 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 66208 437474 66528 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587240 437474 587840 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 66208 434476 66528 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2956 434454 586880 434476
rect -2956 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 66250 434454
rect 66486 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586880 434454
rect -2956 434134 586880 434218
rect -2956 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 66250 434134
rect 66486 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586880 434134
rect -2956 433876 586880 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 66208 433874 66528 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -4876 420076 -4276 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 81568 420076 81888 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588200 420076 588800 420078
rect -4876 420054 588800 420076
rect -4876 419818 -4694 420054
rect -4458 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 81610 420054
rect 81846 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588382 420054
rect 588618 419818 588800 420054
rect -4876 419734 588800 419818
rect -4876 419498 -4694 419734
rect -4458 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 81610 419734
rect 81846 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588382 419734
rect 588618 419498 588800 419734
rect -4876 419476 588800 419498
rect -4876 419474 -4276 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 81568 419474 81888 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588200 419474 588800 419476
rect -2956 416476 -2356 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 81568 416476 81888 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586280 416476 586880 416478
rect -2956 416454 586880 416476
rect -2956 416218 -2774 416454
rect -2538 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 81610 416454
rect 81846 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586462 416454
rect 586698 416218 586880 416454
rect -2956 416134 586880 416218
rect -2956 415898 -2774 416134
rect -2538 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 81610 416134
rect 81846 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586462 416134
rect 586698 415898 586880 416134
rect -2956 415876 586880 415898
rect -2956 415874 -2356 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 81568 415874 81888 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586280 415874 586880 415876
rect -3916 402076 -3316 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 66208 402076 66528 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587240 402076 587840 402078
rect -4876 402054 588800 402076
rect -4876 401818 -3734 402054
rect -3498 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 66250 402054
rect 66486 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587422 402054
rect 587658 401818 588800 402054
rect -4876 401734 588800 401818
rect -4876 401498 -3734 401734
rect -3498 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 66250 401734
rect 66486 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587422 401734
rect 587658 401498 588800 401734
rect -4876 401476 588800 401498
rect -3916 401474 -3316 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 66208 401474 66528 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587240 401474 587840 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 66208 398476 66528 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2956 398454 586880 398476
rect -2956 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 66250 398454
rect 66486 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586880 398454
rect -2956 398134 586880 398218
rect -2956 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 66250 398134
rect 66486 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586880 398134
rect -2956 397876 586880 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 66208 397874 66528 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -4876 384076 -4276 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 81568 384076 81888 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588200 384076 588800 384078
rect -4876 384054 588800 384076
rect -4876 383818 -4694 384054
rect -4458 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 81610 384054
rect 81846 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588382 384054
rect 588618 383818 588800 384054
rect -4876 383734 588800 383818
rect -4876 383498 -4694 383734
rect -4458 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 81610 383734
rect 81846 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588382 383734
rect 588618 383498 588800 383734
rect -4876 383476 588800 383498
rect -4876 383474 -4276 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 81568 383474 81888 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588200 383474 588800 383476
rect -2956 380476 -2356 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 81568 380476 81888 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586280 380476 586880 380478
rect -2956 380454 586880 380476
rect -2956 380218 -2774 380454
rect -2538 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 81610 380454
rect 81846 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586462 380454
rect 586698 380218 586880 380454
rect -2956 380134 586880 380218
rect -2956 379898 -2774 380134
rect -2538 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 81610 380134
rect 81846 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586462 380134
rect 586698 379898 586880 380134
rect -2956 379876 586880 379898
rect -2956 379874 -2356 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 81568 379874 81888 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586280 379874 586880 379876
rect -3916 366076 -3316 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 66208 366076 66528 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587240 366076 587840 366078
rect -4876 366054 588800 366076
rect -4876 365818 -3734 366054
rect -3498 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 66250 366054
rect 66486 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587422 366054
rect 587658 365818 588800 366054
rect -4876 365734 588800 365818
rect -4876 365498 -3734 365734
rect -3498 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 66250 365734
rect 66486 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587422 365734
rect 587658 365498 588800 365734
rect -4876 365476 588800 365498
rect -3916 365474 -3316 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 66208 365474 66528 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587240 365474 587840 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 66208 362476 66528 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2956 362454 586880 362476
rect -2956 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 66250 362454
rect 66486 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586880 362454
rect -2956 362134 586880 362218
rect -2956 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 66250 362134
rect 66486 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586880 362134
rect -2956 361876 586880 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 66208 361874 66528 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -4876 348076 -4276 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 81568 348076 81888 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588200 348076 588800 348078
rect -4876 348054 588800 348076
rect -4876 347818 -4694 348054
rect -4458 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 81610 348054
rect 81846 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588382 348054
rect 588618 347818 588800 348054
rect -4876 347734 588800 347818
rect -4876 347498 -4694 347734
rect -4458 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 81610 347734
rect 81846 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588382 347734
rect 588618 347498 588800 347734
rect -4876 347476 588800 347498
rect -4876 347474 -4276 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 81568 347474 81888 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588200 347474 588800 347476
rect -2956 344476 -2356 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 81568 344476 81888 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586280 344476 586880 344478
rect -2956 344454 586880 344476
rect -2956 344218 -2774 344454
rect -2538 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 81610 344454
rect 81846 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586462 344454
rect 586698 344218 586880 344454
rect -2956 344134 586880 344218
rect -2956 343898 -2774 344134
rect -2538 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 81610 344134
rect 81846 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586462 344134
rect 586698 343898 586880 344134
rect -2956 343876 586880 343898
rect -2956 343874 -2356 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 81568 343874 81888 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586280 343874 586880 343876
rect -3916 330076 -3316 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 66208 330076 66528 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587240 330076 587840 330078
rect -4876 330054 588800 330076
rect -4876 329818 -3734 330054
rect -3498 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 66250 330054
rect 66486 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587422 330054
rect 587658 329818 588800 330054
rect -4876 329734 588800 329818
rect -4876 329498 -3734 329734
rect -3498 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 66250 329734
rect 66486 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587422 329734
rect 587658 329498 588800 329734
rect -4876 329476 588800 329498
rect -3916 329474 -3316 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 66208 329474 66528 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587240 329474 587840 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 66208 326476 66528 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2956 326454 586880 326476
rect -2956 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 66250 326454
rect 66486 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586880 326454
rect -2956 326134 586880 326218
rect -2956 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 66250 326134
rect 66486 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586880 326134
rect -2956 325876 586880 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 66208 325874 66528 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -4876 312076 -4276 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 81568 312076 81888 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588200 312076 588800 312078
rect -4876 312054 588800 312076
rect -4876 311818 -4694 312054
rect -4458 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 81610 312054
rect 81846 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588382 312054
rect 588618 311818 588800 312054
rect -4876 311734 588800 311818
rect -4876 311498 -4694 311734
rect -4458 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 81610 311734
rect 81846 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588382 311734
rect 588618 311498 588800 311734
rect -4876 311476 588800 311498
rect -4876 311474 -4276 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 81568 311474 81888 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588200 311474 588800 311476
rect -2956 308476 -2356 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 81568 308476 81888 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586280 308476 586880 308478
rect -2956 308454 586880 308476
rect -2956 308218 -2774 308454
rect -2538 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 81610 308454
rect 81846 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586462 308454
rect 586698 308218 586880 308454
rect -2956 308134 586880 308218
rect -2956 307898 -2774 308134
rect -2538 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 81610 308134
rect 81846 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586462 308134
rect 586698 307898 586880 308134
rect -2956 307876 586880 307898
rect -2956 307874 -2356 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 81568 307874 81888 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586280 307874 586880 307876
rect -3916 294076 -3316 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 66208 294076 66528 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587240 294076 587840 294078
rect -4876 294054 588800 294076
rect -4876 293818 -3734 294054
rect -3498 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 66250 294054
rect 66486 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587422 294054
rect 587658 293818 588800 294054
rect -4876 293734 588800 293818
rect -4876 293498 -3734 293734
rect -3498 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 66250 293734
rect 66486 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587422 293734
rect 587658 293498 588800 293734
rect -4876 293476 588800 293498
rect -3916 293474 -3316 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 66208 293474 66528 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587240 293474 587840 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 66208 290476 66528 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2956 290454 586880 290476
rect -2956 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 66250 290454
rect 66486 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586880 290454
rect -2956 290134 586880 290218
rect -2956 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 66250 290134
rect 66486 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586880 290134
rect -2956 289876 586880 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 66208 289874 66528 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -4876 276076 -4276 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 81568 276076 81888 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588200 276076 588800 276078
rect -4876 276054 588800 276076
rect -4876 275818 -4694 276054
rect -4458 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 81610 276054
rect 81846 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588382 276054
rect 588618 275818 588800 276054
rect -4876 275734 588800 275818
rect -4876 275498 -4694 275734
rect -4458 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 81610 275734
rect 81846 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588382 275734
rect 588618 275498 588800 275734
rect -4876 275476 588800 275498
rect -4876 275474 -4276 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 81568 275474 81888 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588200 275474 588800 275476
rect -2956 272476 -2356 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 81568 272476 81888 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586280 272476 586880 272478
rect -2956 272454 586880 272476
rect -2956 272218 -2774 272454
rect -2538 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 81610 272454
rect 81846 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586462 272454
rect 586698 272218 586880 272454
rect -2956 272134 586880 272218
rect -2956 271898 -2774 272134
rect -2538 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 81610 272134
rect 81846 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586462 272134
rect 586698 271898 586880 272134
rect -2956 271876 586880 271898
rect -2956 271874 -2356 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 81568 271874 81888 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586280 271874 586880 271876
rect -3916 258076 -3316 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 66208 258076 66528 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587240 258076 587840 258078
rect -4876 258054 588800 258076
rect -4876 257818 -3734 258054
rect -3498 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 66250 258054
rect 66486 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587422 258054
rect 587658 257818 588800 258054
rect -4876 257734 588800 257818
rect -4876 257498 -3734 257734
rect -3498 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 66250 257734
rect 66486 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587422 257734
rect 587658 257498 588800 257734
rect -4876 257476 588800 257498
rect -3916 257474 -3316 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 66208 257474 66528 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587240 257474 587840 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 66208 254476 66528 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2956 254454 586880 254476
rect -2956 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 66250 254454
rect 66486 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586880 254454
rect -2956 254134 586880 254218
rect -2956 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 66250 254134
rect 66486 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586880 254134
rect -2956 253876 586880 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 66208 253874 66528 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -4876 240076 -4276 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 81568 240076 81888 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588200 240076 588800 240078
rect -4876 240054 588800 240076
rect -4876 239818 -4694 240054
rect -4458 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 81610 240054
rect 81846 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588382 240054
rect 588618 239818 588800 240054
rect -4876 239734 588800 239818
rect -4876 239498 -4694 239734
rect -4458 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 81610 239734
rect 81846 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588382 239734
rect 588618 239498 588800 239734
rect -4876 239476 588800 239498
rect -4876 239474 -4276 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 81568 239474 81888 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588200 239474 588800 239476
rect -2956 236476 -2356 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 81568 236476 81888 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586280 236476 586880 236478
rect -2956 236454 586880 236476
rect -2956 236218 -2774 236454
rect -2538 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 81610 236454
rect 81846 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586462 236454
rect 586698 236218 586880 236454
rect -2956 236134 586880 236218
rect -2956 235898 -2774 236134
rect -2538 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 81610 236134
rect 81846 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586462 236134
rect 586698 235898 586880 236134
rect -2956 235876 586880 235898
rect -2956 235874 -2356 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 81568 235874 81888 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586280 235874 586880 235876
rect -3916 222076 -3316 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 66208 222076 66528 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587240 222076 587840 222078
rect -4876 222054 588800 222076
rect -4876 221818 -3734 222054
rect -3498 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 66250 222054
rect 66486 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587422 222054
rect 587658 221818 588800 222054
rect -4876 221734 588800 221818
rect -4876 221498 -3734 221734
rect -3498 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 66250 221734
rect 66486 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587422 221734
rect 587658 221498 588800 221734
rect -4876 221476 588800 221498
rect -3916 221474 -3316 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 66208 221474 66528 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587240 221474 587840 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 66208 218476 66528 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2956 218454 586880 218476
rect -2956 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 66250 218454
rect 66486 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586880 218454
rect -2956 218134 586880 218218
rect -2956 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 66250 218134
rect 66486 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586880 218134
rect -2956 217876 586880 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 66208 217874 66528 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -4876 204076 -4276 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 81568 204076 81888 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588200 204076 588800 204078
rect -4876 204054 588800 204076
rect -4876 203818 -4694 204054
rect -4458 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 81610 204054
rect 81846 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588382 204054
rect 588618 203818 588800 204054
rect -4876 203734 588800 203818
rect -4876 203498 -4694 203734
rect -4458 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 81610 203734
rect 81846 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588382 203734
rect 588618 203498 588800 203734
rect -4876 203476 588800 203498
rect -4876 203474 -4276 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 81568 203474 81888 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588200 203474 588800 203476
rect -2956 200476 -2356 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 81568 200476 81888 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586280 200476 586880 200478
rect -2956 200454 586880 200476
rect -2956 200218 -2774 200454
rect -2538 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 81610 200454
rect 81846 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586462 200454
rect 586698 200218 586880 200454
rect -2956 200134 586880 200218
rect -2956 199898 -2774 200134
rect -2538 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 81610 200134
rect 81846 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586462 200134
rect 586698 199898 586880 200134
rect -2956 199876 586880 199898
rect -2956 199874 -2356 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 81568 199874 81888 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586280 199874 586880 199876
rect -3916 186076 -3316 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 66208 186076 66528 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587240 186076 587840 186078
rect -4876 186054 588800 186076
rect -4876 185818 -3734 186054
rect -3498 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 66250 186054
rect 66486 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587422 186054
rect 587658 185818 588800 186054
rect -4876 185734 588800 185818
rect -4876 185498 -3734 185734
rect -3498 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 66250 185734
rect 66486 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587422 185734
rect 587658 185498 588800 185734
rect -4876 185476 588800 185498
rect -3916 185474 -3316 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 66208 185474 66528 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587240 185474 587840 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 66208 182476 66528 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2956 182454 586880 182476
rect -2956 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 66250 182454
rect 66486 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586880 182454
rect -2956 182134 586880 182218
rect -2956 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 66250 182134
rect 66486 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586880 182134
rect -2956 181876 586880 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 66208 181874 66528 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -4876 168076 -4276 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 81568 168076 81888 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588200 168076 588800 168078
rect -4876 168054 588800 168076
rect -4876 167818 -4694 168054
rect -4458 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 81610 168054
rect 81846 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588382 168054
rect 588618 167818 588800 168054
rect -4876 167734 588800 167818
rect -4876 167498 -4694 167734
rect -4458 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 81610 167734
rect 81846 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588382 167734
rect 588618 167498 588800 167734
rect -4876 167476 588800 167498
rect -4876 167474 -4276 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 81568 167474 81888 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588200 167474 588800 167476
rect -2956 164476 -2356 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 81568 164476 81888 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586280 164476 586880 164478
rect -2956 164454 586880 164476
rect -2956 164218 -2774 164454
rect -2538 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 81610 164454
rect 81846 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586462 164454
rect 586698 164218 586880 164454
rect -2956 164134 586880 164218
rect -2956 163898 -2774 164134
rect -2538 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 81610 164134
rect 81846 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586462 164134
rect 586698 163898 586880 164134
rect -2956 163876 586880 163898
rect -2956 163874 -2356 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 81568 163874 81888 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586280 163874 586880 163876
rect -3916 150076 -3316 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 66208 150076 66528 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587240 150076 587840 150078
rect -4876 150054 588800 150076
rect -4876 149818 -3734 150054
rect -3498 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 66250 150054
rect 66486 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587422 150054
rect 587658 149818 588800 150054
rect -4876 149734 588800 149818
rect -4876 149498 -3734 149734
rect -3498 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 66250 149734
rect 66486 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587422 149734
rect 587658 149498 588800 149734
rect -4876 149476 588800 149498
rect -3916 149474 -3316 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 66208 149474 66528 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587240 149474 587840 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 66208 146476 66528 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2956 146454 586880 146476
rect -2956 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 66250 146454
rect 66486 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586880 146454
rect -2956 146134 586880 146218
rect -2956 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 66250 146134
rect 66486 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586880 146134
rect -2956 145876 586880 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 66208 145874 66528 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -4876 132076 -4276 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 81568 132076 81888 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588200 132076 588800 132078
rect -4876 132054 588800 132076
rect -4876 131818 -4694 132054
rect -4458 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 81610 132054
rect 81846 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588382 132054
rect 588618 131818 588800 132054
rect -4876 131734 588800 131818
rect -4876 131498 -4694 131734
rect -4458 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 81610 131734
rect 81846 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588382 131734
rect 588618 131498 588800 131734
rect -4876 131476 588800 131498
rect -4876 131474 -4276 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 81568 131474 81888 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588200 131474 588800 131476
rect -2956 128476 -2356 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 81568 128476 81888 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586280 128476 586880 128478
rect -2956 128454 586880 128476
rect -2956 128218 -2774 128454
rect -2538 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 81610 128454
rect 81846 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586462 128454
rect 586698 128218 586880 128454
rect -2956 128134 586880 128218
rect -2956 127898 -2774 128134
rect -2538 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 81610 128134
rect 81846 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586462 128134
rect 586698 127898 586880 128134
rect -2956 127876 586880 127898
rect -2956 127874 -2356 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 81568 127874 81888 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586280 127874 586880 127876
rect -3916 114076 -3316 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 66208 114076 66528 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587240 114076 587840 114078
rect -4876 114054 588800 114076
rect -4876 113818 -3734 114054
rect -3498 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 66250 114054
rect 66486 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587422 114054
rect 587658 113818 588800 114054
rect -4876 113734 588800 113818
rect -4876 113498 -3734 113734
rect -3498 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 66250 113734
rect 66486 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587422 113734
rect 587658 113498 588800 113734
rect -4876 113476 588800 113498
rect -3916 113474 -3316 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 66208 113474 66528 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587240 113474 587840 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 66208 110476 66528 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2956 110454 586880 110476
rect -2956 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 66250 110454
rect 66486 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586880 110454
rect -2956 110134 586880 110218
rect -2956 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 66250 110134
rect 66486 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586880 110134
rect -2956 109876 586880 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 66208 109874 66528 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -4876 96076 -4276 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 81568 96076 81888 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588200 96076 588800 96078
rect -4876 96054 588800 96076
rect -4876 95818 -4694 96054
rect -4458 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 81610 96054
rect 81846 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588382 96054
rect 588618 95818 588800 96054
rect -4876 95734 588800 95818
rect -4876 95498 -4694 95734
rect -4458 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 81610 95734
rect 81846 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588382 95734
rect 588618 95498 588800 95734
rect -4876 95476 588800 95498
rect -4876 95474 -4276 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 81568 95474 81888 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588200 95474 588800 95476
rect -2956 92476 -2356 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 81568 92476 81888 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586280 92476 586880 92478
rect -2956 92454 586880 92476
rect -2956 92218 -2774 92454
rect -2538 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 81610 92454
rect 81846 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586462 92454
rect 586698 92218 586880 92454
rect -2956 92134 586880 92218
rect -2956 91898 -2774 92134
rect -2538 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 81610 92134
rect 81846 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586462 92134
rect 586698 91898 586880 92134
rect -2956 91876 586880 91898
rect -2956 91874 -2356 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 81568 91874 81888 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586280 91874 586880 91876
rect -3916 78076 -3316 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 66208 78076 66528 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587240 78076 587840 78078
rect -4876 78054 588800 78076
rect -4876 77818 -3734 78054
rect -3498 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 66250 78054
rect 66486 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587422 78054
rect 587658 77818 588800 78054
rect -4876 77734 588800 77818
rect -4876 77498 -3734 77734
rect -3498 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 66250 77734
rect 66486 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587422 77734
rect 587658 77498 588800 77734
rect -4876 77476 588800 77498
rect -3916 77474 -3316 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 66208 77474 66528 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587240 77474 587840 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 66208 74476 66528 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2956 74454 586880 74476
rect -2956 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 66250 74454
rect 66486 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586880 74454
rect -2956 74134 586880 74218
rect -2956 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 66250 74134
rect 66486 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586880 74134
rect -2956 73876 586880 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 66208 73874 66528 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -4876 60076 -4276 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 81568 60076 81888 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588200 60076 588800 60078
rect -4876 60054 588800 60076
rect -4876 59818 -4694 60054
rect -4458 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 81610 60054
rect 81846 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588382 60054
rect 588618 59818 588800 60054
rect -4876 59734 588800 59818
rect -4876 59498 -4694 59734
rect -4458 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 81610 59734
rect 81846 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588382 59734
rect 588618 59498 588800 59734
rect -4876 59476 588800 59498
rect -4876 59474 -4276 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 81568 59474 81888 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588200 59474 588800 59476
rect -2956 56476 -2356 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 81568 56476 81888 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586280 56476 586880 56478
rect -2956 56454 586880 56476
rect -2956 56218 -2774 56454
rect -2538 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 81610 56454
rect 81846 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586462 56454
rect 586698 56218 586880 56454
rect -2956 56134 586880 56218
rect -2956 55898 -2774 56134
rect -2538 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 81610 56134
rect 81846 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586462 56134
rect 586698 55898 586880 56134
rect -2956 55876 586880 55898
rect -2956 55874 -2356 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 81568 55874 81888 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586280 55874 586880 55876
rect -3916 42076 -3316 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587240 42076 587840 42078
rect -4876 42054 588800 42076
rect -4876 41818 -3734 42054
rect -3498 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587422 42054
rect 587658 41818 588800 42054
rect -4876 41734 588800 41818
rect -4876 41498 -3734 41734
rect -3498 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587422 41734
rect 587658 41498 588800 41734
rect -4876 41476 588800 41498
rect -3916 41474 -3316 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587240 41474 587840 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2956 38454 586880 38476
rect -2956 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586880 38454
rect -2956 38134 586880 38218
rect -2956 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586880 38134
rect -2956 37876 586880 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -4876 24076 -4276 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588200 24076 588800 24078
rect -4876 24054 588800 24076
rect -4876 23818 -4694 24054
rect -4458 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588382 24054
rect 588618 23818 588800 24054
rect -4876 23734 588800 23818
rect -4876 23498 -4694 23734
rect -4458 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588382 23734
rect 588618 23498 588800 23734
rect -4876 23476 588800 23498
rect -4876 23474 -4276 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588200 23474 588800 23476
rect -2956 20476 -2356 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586280 20476 586880 20478
rect -2956 20454 586880 20476
rect -2956 20218 -2774 20454
rect -2538 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586462 20454
rect 586698 20218 586880 20454
rect -2956 20134 586880 20218
rect -2956 19898 -2774 20134
rect -2538 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586462 20134
rect 586698 19898 586880 20134
rect -2956 19876 586880 19898
rect -2956 19874 -2356 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586280 19874 586880 19876
rect -3916 6076 -3316 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587240 6076 587840 6078
rect -4876 6054 588800 6076
rect -4876 5818 -3734 6054
rect -3498 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587422 6054
rect 587658 5818 588800 6054
rect -4876 5734 588800 5818
rect -4876 5498 -3734 5734
rect -3498 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587422 5734
rect 587658 5498 588800 5734
rect -4876 5476 588800 5498
rect -3916 5474 -3316 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587240 5474 587840 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2956 2454 586880 2476
rect -2956 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586880 2454
rect -2956 2134 586880 2218
rect -2956 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586880 2134
rect -2956 1876 586880 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2956 -1284 -2356 -1282
rect 18804 -1284 19404 -1282
rect 54804 -1284 55404 -1282
rect 90804 -1284 91404 -1282
rect 126804 -1284 127404 -1282
rect 162804 -1284 163404 -1282
rect 198804 -1284 199404 -1282
rect 234804 -1284 235404 -1282
rect 270804 -1284 271404 -1282
rect 306804 -1284 307404 -1282
rect 342804 -1284 343404 -1282
rect 378804 -1284 379404 -1282
rect 414804 -1284 415404 -1282
rect 450804 -1284 451404 -1282
rect 486804 -1284 487404 -1282
rect 522804 -1284 523404 -1282
rect 558804 -1284 559404 -1282
rect 586280 -1284 586880 -1282
rect -2956 -1306 586880 -1284
rect -2956 -1542 -2774 -1306
rect -2538 -1542 18986 -1306
rect 19222 -1542 54986 -1306
rect 55222 -1542 90986 -1306
rect 91222 -1542 126986 -1306
rect 127222 -1542 162986 -1306
rect 163222 -1542 198986 -1306
rect 199222 -1542 234986 -1306
rect 235222 -1542 270986 -1306
rect 271222 -1542 306986 -1306
rect 307222 -1542 342986 -1306
rect 343222 -1542 378986 -1306
rect 379222 -1542 414986 -1306
rect 415222 -1542 450986 -1306
rect 451222 -1542 486986 -1306
rect 487222 -1542 522986 -1306
rect 523222 -1542 558986 -1306
rect 559222 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect -2956 -1626 586880 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 18986 -1626
rect 19222 -1862 54986 -1626
rect 55222 -1862 90986 -1626
rect 91222 -1862 126986 -1626
rect 127222 -1862 162986 -1626
rect 163222 -1862 198986 -1626
rect 199222 -1862 234986 -1626
rect 235222 -1862 270986 -1626
rect 271222 -1862 306986 -1626
rect 307222 -1862 342986 -1626
rect 343222 -1862 378986 -1626
rect 379222 -1862 414986 -1626
rect 415222 -1862 450986 -1626
rect 451222 -1862 486986 -1626
rect 487222 -1862 522986 -1626
rect 523222 -1862 558986 -1626
rect 559222 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect -2956 -1884 586880 -1862
rect -2956 -1886 -2356 -1884
rect 18804 -1886 19404 -1884
rect 54804 -1886 55404 -1884
rect 90804 -1886 91404 -1884
rect 126804 -1886 127404 -1884
rect 162804 -1886 163404 -1884
rect 198804 -1886 199404 -1884
rect 234804 -1886 235404 -1884
rect 270804 -1886 271404 -1884
rect 306804 -1886 307404 -1884
rect 342804 -1886 343404 -1884
rect 378804 -1886 379404 -1884
rect 414804 -1886 415404 -1884
rect 450804 -1886 451404 -1884
rect 486804 -1886 487404 -1884
rect 522804 -1886 523404 -1884
rect 558804 -1886 559404 -1884
rect 586280 -1886 586880 -1884
rect -3916 -2244 -3316 -2242
rect 4404 -2244 5004 -2242
rect 40404 -2244 41004 -2242
rect 76404 -2244 77004 -2242
rect 112404 -2244 113004 -2242
rect 148404 -2244 149004 -2242
rect 184404 -2244 185004 -2242
rect 220404 -2244 221004 -2242
rect 256404 -2244 257004 -2242
rect 292404 -2244 293004 -2242
rect 328404 -2244 329004 -2242
rect 364404 -2244 365004 -2242
rect 400404 -2244 401004 -2242
rect 436404 -2244 437004 -2242
rect 472404 -2244 473004 -2242
rect 508404 -2244 509004 -2242
rect 544404 -2244 545004 -2242
rect 580404 -2244 581004 -2242
rect 587240 -2244 587840 -2242
rect -3916 -2266 587840 -2244
rect -3916 -2502 -3734 -2266
rect -3498 -2502 4586 -2266
rect 4822 -2502 40586 -2266
rect 40822 -2502 76586 -2266
rect 76822 -2502 112586 -2266
rect 112822 -2502 148586 -2266
rect 148822 -2502 184586 -2266
rect 184822 -2502 220586 -2266
rect 220822 -2502 256586 -2266
rect 256822 -2502 292586 -2266
rect 292822 -2502 328586 -2266
rect 328822 -2502 364586 -2266
rect 364822 -2502 400586 -2266
rect 400822 -2502 436586 -2266
rect 436822 -2502 472586 -2266
rect 472822 -2502 508586 -2266
rect 508822 -2502 544586 -2266
rect 544822 -2502 580586 -2266
rect 580822 -2502 587422 -2266
rect 587658 -2502 587840 -2266
rect -3916 -2586 587840 -2502
rect -3916 -2822 -3734 -2586
rect -3498 -2822 4586 -2586
rect 4822 -2822 40586 -2586
rect 40822 -2822 76586 -2586
rect 76822 -2822 112586 -2586
rect 112822 -2822 148586 -2586
rect 148822 -2822 184586 -2586
rect 184822 -2822 220586 -2586
rect 220822 -2822 256586 -2586
rect 256822 -2822 292586 -2586
rect 292822 -2822 328586 -2586
rect 328822 -2822 364586 -2586
rect 364822 -2822 400586 -2586
rect 400822 -2822 436586 -2586
rect 436822 -2822 472586 -2586
rect 472822 -2822 508586 -2586
rect 508822 -2822 544586 -2586
rect 544822 -2822 580586 -2586
rect 580822 -2822 587422 -2586
rect 587658 -2822 587840 -2586
rect -3916 -2844 587840 -2822
rect -3916 -2846 -3316 -2844
rect 4404 -2846 5004 -2844
rect 40404 -2846 41004 -2844
rect 76404 -2846 77004 -2844
rect 112404 -2846 113004 -2844
rect 148404 -2846 149004 -2844
rect 184404 -2846 185004 -2844
rect 220404 -2846 221004 -2844
rect 256404 -2846 257004 -2844
rect 292404 -2846 293004 -2844
rect 328404 -2846 329004 -2844
rect 364404 -2846 365004 -2844
rect 400404 -2846 401004 -2844
rect 436404 -2846 437004 -2844
rect 472404 -2846 473004 -2844
rect 508404 -2846 509004 -2844
rect 544404 -2846 545004 -2844
rect 580404 -2846 581004 -2844
rect 587240 -2846 587840 -2844
rect -4876 -3204 -4276 -3202
rect 22404 -3204 23004 -3202
rect 58404 -3204 59004 -3202
rect 94404 -3204 95004 -3202
rect 130404 -3204 131004 -3202
rect 166404 -3204 167004 -3202
rect 202404 -3204 203004 -3202
rect 238404 -3204 239004 -3202
rect 274404 -3204 275004 -3202
rect 310404 -3204 311004 -3202
rect 346404 -3204 347004 -3202
rect 382404 -3204 383004 -3202
rect 418404 -3204 419004 -3202
rect 454404 -3204 455004 -3202
rect 490404 -3204 491004 -3202
rect 526404 -3204 527004 -3202
rect 562404 -3204 563004 -3202
rect 588200 -3204 588800 -3202
rect -4876 -3226 588800 -3204
rect -4876 -3462 -4694 -3226
rect -4458 -3462 22586 -3226
rect 22822 -3462 58586 -3226
rect 58822 -3462 94586 -3226
rect 94822 -3462 130586 -3226
rect 130822 -3462 166586 -3226
rect 166822 -3462 202586 -3226
rect 202822 -3462 238586 -3226
rect 238822 -3462 274586 -3226
rect 274822 -3462 310586 -3226
rect 310822 -3462 346586 -3226
rect 346822 -3462 382586 -3226
rect 382822 -3462 418586 -3226
rect 418822 -3462 454586 -3226
rect 454822 -3462 490586 -3226
rect 490822 -3462 526586 -3226
rect 526822 -3462 562586 -3226
rect 562822 -3462 588382 -3226
rect 588618 -3462 588800 -3226
rect -4876 -3546 588800 -3462
rect -4876 -3782 -4694 -3546
rect -4458 -3782 22586 -3546
rect 22822 -3782 58586 -3546
rect 58822 -3782 94586 -3546
rect 94822 -3782 130586 -3546
rect 130822 -3782 166586 -3546
rect 166822 -3782 202586 -3546
rect 202822 -3782 238586 -3546
rect 238822 -3782 274586 -3546
rect 274822 -3782 310586 -3546
rect 310822 -3782 346586 -3546
rect 346822 -3782 382586 -3546
rect 382822 -3782 418586 -3546
rect 418822 -3782 454586 -3546
rect 454822 -3782 490586 -3546
rect 490822 -3782 526586 -3546
rect 526822 -3782 562586 -3546
rect 562822 -3782 588382 -3546
rect 588618 -3782 588800 -3546
rect -4876 -3804 588800 -3782
rect -4876 -3806 -4276 -3804
rect 22404 -3806 23004 -3804
rect 58404 -3806 59004 -3804
rect 94404 -3806 95004 -3804
rect 130404 -3806 131004 -3804
rect 166404 -3806 167004 -3804
rect 202404 -3806 203004 -3804
rect 238404 -3806 239004 -3804
rect 274404 -3806 275004 -3804
rect 310404 -3806 311004 -3804
rect 346404 -3806 347004 -3804
rect 382404 -3806 383004 -3804
rect 418404 -3806 419004 -3804
rect 454404 -3806 455004 -3804
rect 490404 -3806 491004 -3804
rect 526404 -3806 527004 -3804
rect 562404 -3806 563004 -3804
rect 588200 -3806 588800 -3804
use ghazi_top_dffram_csv  mprj
timestamp 1608008999
transform 1 0 62000 0 1 52000
box 0 0 460000 600000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2956 -1884 586880 -1284 8 vssd1
port 637 nsew default input
rlabel metal5 s -3916 -2844 587840 -2244 8 vccd2
port 638 nsew default input
rlabel metal5 s -4876 -3804 588800 -3204 8 vssd2
port 639 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
