magic
tech sky130A
magscale 1 2
timestamp 1608285900
<< locali >>
rect 8125 685899 8159 695453
rect 72525 683247 72559 692733
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72709 678895 72743 683077
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 72801 656931 72835 666485
rect 219081 656931 219115 666485
rect 398849 37315 398883 37961
rect 407221 37315 407255 46869
rect 443193 37315 443227 46869
rect 450001 37315 450035 46869
rect 535469 37315 535503 46869
rect 516149 29019 516183 35173
rect 333989 9707 334023 19261
rect 345029 9707 345063 19261
rect 372629 9707 372663 19261
rect 394709 9707 394743 19261
rect 397469 9707 397503 19261
rect 398849 9707 398883 27557
rect 407221 12291 407255 27557
rect 443009 9707 443043 27557
rect 535469 9707 535503 27557
rect 336657 3655 336691 7021
rect 388395 5321 388579 5355
rect 388545 5219 388579 5321
rect 388453 4947 388487 5185
rect 405749 4539 405783 4709
rect 345029 3655 345063 4165
rect 340831 3621 340889 3655
rect 354597 3655 354631 4165
rect 357449 3655 357483 3825
rect 336841 3587 336875 3621
rect 336783 3553 336875 3587
rect 361221 3519 361255 3689
rect 367017 3587 367051 3825
rect 386279 3621 386337 3655
rect 369961 3519 369995 3553
rect 369961 3485 370053 3519
rect 183477 3247 183511 3417
rect 376769 3315 376803 3553
rect 412097 595 412131 9605
rect 413293 4811 413327 5253
rect 415317 4539 415351 4641
rect 420377 595 420411 9605
rect 422953 4811 422987 5253
rect 433625 4539 433659 4845
rect 480269 4743 480303 4913
rect 489837 4743 489871 4913
rect 499589 4743 499623 4913
rect 509157 4743 509191 4913
rect 514769 4743 514803 4913
rect 515689 4743 515723 4981
rect 428749 595 428783 2805
rect 435833 595 435867 2805
rect 516793 595 516827 9605
rect 520289 595 520323 9605
rect 524371 4981 524429 5015
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 692733 72559 692767
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 72525 683213 72559 683247
rect 154313 685797 154347 685831
rect 72709 683077 72743 683111
rect 72709 678861 72743 678895
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 284033 676209 284067 676243
rect 72801 666485 72835 666519
rect 72801 656897 72835 656931
rect 219081 666485 219115 666519
rect 219081 656897 219115 656931
rect 407221 46869 407255 46903
rect 398849 37961 398883 37995
rect 398849 37281 398883 37315
rect 407221 37281 407255 37315
rect 443193 46869 443227 46903
rect 443193 37281 443227 37315
rect 450001 46869 450035 46903
rect 450001 37281 450035 37315
rect 535469 46869 535503 46903
rect 535469 37281 535503 37315
rect 516149 35173 516183 35207
rect 516149 28985 516183 29019
rect 398849 27557 398883 27591
rect 333989 19261 334023 19295
rect 333989 9673 334023 9707
rect 345029 19261 345063 19295
rect 345029 9673 345063 9707
rect 372629 19261 372663 19295
rect 372629 9673 372663 9707
rect 394709 19261 394743 19295
rect 394709 9673 394743 9707
rect 397469 19261 397503 19295
rect 397469 9673 397503 9707
rect 407221 27557 407255 27591
rect 407221 12257 407255 12291
rect 443009 27557 443043 27591
rect 398849 9673 398883 9707
rect 443009 9673 443043 9707
rect 535469 27557 535503 27591
rect 535469 9673 535503 9707
rect 412097 9605 412131 9639
rect 336657 7021 336691 7055
rect 388361 5321 388395 5355
rect 388453 5185 388487 5219
rect 388545 5185 388579 5219
rect 388453 4913 388487 4947
rect 405749 4709 405783 4743
rect 405749 4505 405783 4539
rect 345029 4165 345063 4199
rect 336657 3621 336691 3655
rect 336841 3621 336875 3655
rect 340797 3621 340831 3655
rect 340889 3621 340923 3655
rect 345029 3621 345063 3655
rect 354597 4165 354631 4199
rect 354597 3621 354631 3655
rect 357449 3825 357483 3859
rect 367017 3825 367051 3859
rect 357449 3621 357483 3655
rect 361221 3689 361255 3723
rect 336749 3553 336783 3587
rect 386245 3621 386279 3655
rect 386337 3621 386371 3655
rect 367017 3553 367051 3587
rect 369961 3553 369995 3587
rect 361221 3485 361255 3519
rect 376769 3553 376803 3587
rect 370053 3485 370087 3519
rect 183477 3417 183511 3451
rect 376769 3281 376803 3315
rect 183477 3213 183511 3247
rect 420377 9605 420411 9639
rect 413293 5253 413327 5287
rect 413293 4777 413327 4811
rect 415317 4641 415351 4675
rect 415317 4505 415351 4539
rect 412097 561 412131 595
rect 516793 9605 516827 9639
rect 422953 5253 422987 5287
rect 515689 4981 515723 5015
rect 480269 4913 480303 4947
rect 422953 4777 422987 4811
rect 433625 4845 433659 4879
rect 480269 4709 480303 4743
rect 489837 4913 489871 4947
rect 489837 4709 489871 4743
rect 499589 4913 499623 4947
rect 499589 4709 499623 4743
rect 509157 4913 509191 4947
rect 509157 4709 509191 4743
rect 514769 4913 514803 4947
rect 514769 4709 514803 4743
rect 515689 4709 515723 4743
rect 433625 4505 433659 4539
rect 420377 561 420411 595
rect 428749 2805 428783 2839
rect 428749 561 428783 595
rect 435833 2805 435867 2839
rect 435833 561 435867 595
rect 516793 561 516827 595
rect 520289 9605 520323 9639
rect 524337 4981 524371 5015
rect 524429 4981 524463 5015
rect 520289 561 520323 595
<< metal1 >>
rect 411162 700408 411168 700460
rect 411220 700448 411226 700460
rect 429838 700448 429844 700460
rect 411220 700420 429844 700448
rect 411220 700408 411226 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 463602 700408 463608 700460
rect 463660 700448 463666 700460
rect 494790 700448 494796 700460
rect 463660 700420 494796 700448
rect 463660 700408 463666 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 514662 700408 514668 700460
rect 514720 700448 514726 700460
rect 559650 700448 559656 700460
rect 514720 700420 559656 700448
rect 514720 700408 514726 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 394602 700340 394608 700392
rect 394660 700380 394666 700392
rect 413646 700380 413652 700392
rect 394660 700352 413652 700380
rect 394660 700340 394666 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 445662 700340 445668 700392
rect 445720 700380 445726 700392
rect 478506 700380 478512 700392
rect 445720 700352 478512 700380
rect 445720 700340 445726 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 496722 700340 496728 700392
rect 496780 700380 496786 700392
rect 543458 700380 543464 700392
rect 496780 700352 543464 700380
rect 496780 700340 496786 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 343542 700272 343548 700324
rect 343600 700312 343606 700324
rect 348786 700312 348792 700324
rect 343600 700284 348792 700312
rect 343600 700272 343606 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 378042 700272 378048 700324
rect 378100 700312 378106 700324
rect 397454 700312 397460 700324
rect 378100 700284 397460 700312
rect 378100 700272 378106 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 429102 700272 429108 700324
rect 429160 700312 429166 700324
rect 462314 700312 462320 700324
rect 429160 700284 462320 700312
rect 429160 700272 429166 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 480162 700272 480168 700324
rect 480220 700312 480226 700324
rect 527174 700312 527180 700324
rect 480220 700284 527180 700312
rect 480220 700272 480226 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 326982 699660 326988 699712
rect 327040 699700 327046 699712
rect 332502 699700 332508 699712
rect 327040 699672 332508 699700
rect 327040 699660 327046 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 360102 699660 360108 699712
rect 360160 699700 360166 699712
rect 364978 699700 364984 699712
rect 360160 699672 364984 699700
rect 360160 699660 360166 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 523770 696940 523776 696992
rect 523828 696980 523834 696992
rect 580166 696980 580172 696992
rect 523828 696952 580172 696980
rect 523828 696940 523834 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 692767 72571 692773
rect 72513 692733 72525 692767
rect 72559 692764 72571 692767
rect 72694 692764 72700 692776
rect 72559 692736 72700 692764
rect 72559 692733 72571 692736
rect 72513 692727 72571 692733
rect 72694 692724 72700 692736
rect 72752 692724 72758 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 523678 685856 523684 685908
rect 523736 685896 523742 685908
rect 580166 685896 580172 685908
rect 523736 685868 580172 685896
rect 523736 685856 523742 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 683244 72516 683256
rect 72471 683216 72516 683244
rect 72510 683204 72516 683216
rect 72568 683204 72574 683256
rect 72510 683068 72516 683120
rect 72568 683108 72574 683120
rect 72697 683111 72755 683117
rect 72697 683108 72709 683111
rect 72568 683080 72709 683108
rect 72568 683068 72574 683080
rect 72697 683077 72709 683080
rect 72743 683077 72755 683111
rect 72697 683071 72755 683077
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 219066 679028 219072 679040
rect 218992 679000 219072 679028
rect 218992 678972 219020 679000
rect 219066 678988 219072 679000
rect 219124 678988 219130 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 218974 678920 218980 678972
rect 219032 678920 219038 678972
rect 72694 678892 72700 678904
rect 72655 678864 72700 678892
rect 72694 678852 72700 678864
rect 72752 678852 72758 678904
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 72694 669264 72700 669316
rect 72752 669304 72758 669316
rect 72878 669304 72884 669316
rect 72752 669276 72884 669304
rect 72752 669264 72758 669276
rect 72878 669264 72884 669276
rect 72936 669264 72942 669316
rect 218974 669264 218980 669316
rect 219032 669304 219038 669316
rect 219158 669304 219164 669316
rect 219032 669276 219164 669304
rect 219032 669264 219038 669276
rect 219158 669264 219164 669276
rect 219216 669264 219222 669316
rect 72789 666519 72847 666525
rect 72789 666485 72801 666519
rect 72835 666516 72847 666519
rect 72878 666516 72884 666528
rect 72835 666488 72884 666516
rect 72835 666485 72847 666488
rect 72789 666479 72847 666485
rect 72878 666476 72884 666488
rect 72936 666476 72942 666528
rect 219069 666519 219127 666525
rect 219069 666485 219081 666519
rect 219115 666516 219127 666519
rect 219158 666516 219164 666528
rect 219115 666488 219164 666516
rect 219115 666485 219127 666488
rect 219069 666479 219127 666485
rect 219158 666476 219164 666488
rect 219216 666476 219222 666528
rect 72786 656928 72792 656940
rect 72747 656900 72792 656928
rect 72786 656888 72792 656900
rect 72844 656888 72850 656940
rect 219066 656928 219072 656940
rect 219027 656900 219072 656928
rect 219066 656888 219072 656900
rect 219124 656888 219130 656940
rect 377122 655460 377128 655512
rect 377180 655500 377186 655512
rect 378042 655500 378048 655512
rect 377180 655472 378048 655500
rect 377180 655460 377186 655472
rect 378042 655460 378048 655472
rect 378100 655460 378106 655512
rect 428182 655460 428188 655512
rect 428240 655500 428246 655512
rect 429102 655500 429108 655512
rect 428240 655472 429108 655500
rect 428240 655460 428246 655472
rect 429102 655460 429108 655472
rect 429160 655460 429166 655512
rect 462314 655460 462320 655512
rect 462372 655500 462378 655512
rect 463602 655500 463608 655512
rect 462372 655472 463608 655500
rect 462372 655460 462378 655472
rect 463602 655460 463608 655472
rect 463660 655460 463666 655512
rect 479334 655460 479340 655512
rect 479392 655500 479398 655512
rect 480162 655500 480168 655512
rect 479392 655472 480168 655500
rect 479392 655460 479398 655472
rect 480162 655460 480168 655472
rect 480220 655460 480226 655512
rect 513374 655256 513380 655308
rect 513432 655296 513438 655308
rect 514662 655296 514668 655308
rect 513432 655268 514668 655296
rect 513432 655256 513438 655268
rect 514662 655256 514668 655268
rect 514720 655256 514726 655308
rect 325970 655120 325976 655172
rect 326028 655160 326034 655172
rect 326982 655160 326988 655172
rect 326028 655132 326988 655160
rect 326028 655120 326034 655132
rect 326982 655120 326988 655132
rect 327040 655120 327046 655172
rect 72786 654984 72792 655036
rect 72844 655024 72850 655036
rect 121546 655024 121552 655036
rect 72844 654996 121552 655024
rect 72844 654984 72850 654996
rect 121546 654984 121552 654996
rect 121604 654984 121610 655036
rect 137738 654984 137744 655036
rect 137796 655024 137802 655036
rect 172698 655024 172704 655036
rect 137796 654996 172704 655024
rect 137796 654984 137802 654996
rect 172698 654984 172704 654996
rect 172756 654984 172762 655036
rect 41322 654916 41328 654968
rect 41380 654956 41386 654968
rect 104526 654956 104532 654968
rect 41380 654928 104532 654956
rect 41380 654916 41386 654928
rect 104526 654916 104532 654928
rect 104584 654916 104590 654968
rect 154298 654916 154304 654968
rect 154356 654956 154362 654968
rect 189718 654956 189724 654968
rect 154356 654928 189724 654956
rect 154356 654916 154362 654928
rect 189718 654916 189724 654928
rect 189776 654916 189782 654968
rect 219066 654916 219072 654968
rect 219124 654956 219130 654968
rect 240778 654956 240784 654968
rect 219124 654928 240784 654956
rect 219124 654916 219130 654928
rect 240778 654916 240784 654928
rect 240836 654916 240842 654968
rect 24762 654848 24768 654900
rect 24820 654888 24826 654900
rect 87506 654888 87512 654900
rect 24820 654860 87512 654888
rect 24820 654848 24826 654860
rect 87506 654848 87512 654860
rect 87564 654848 87570 654900
rect 106182 654848 106188 654900
rect 106240 654888 106246 654900
rect 155586 654888 155592 654900
rect 106240 654860 155592 654888
rect 106240 654848 106246 654860
rect 155586 654848 155592 654860
rect 155644 654848 155650 654900
rect 202782 654848 202788 654900
rect 202840 654888 202846 654900
rect 223758 654888 223764 654900
rect 202840 654860 223764 654888
rect 202840 654848 202846 654860
rect 223758 654848 223764 654860
rect 223816 654848 223822 654900
rect 8018 654780 8024 654832
rect 8076 654820 8082 654832
rect 70486 654820 70492 654832
rect 8076 654792 70492 654820
rect 8076 654780 8082 654792
rect 70486 654780 70492 654792
rect 70544 654780 70550 654832
rect 89622 654780 89628 654832
rect 89680 654820 89686 654832
rect 138566 654820 138572 654832
rect 89680 654792 138572 654820
rect 89680 654780 89686 654792
rect 138566 654780 138572 654792
rect 138624 654780 138630 654832
rect 171042 654780 171048 654832
rect 171100 654820 171106 654832
rect 206738 654820 206744 654832
rect 171100 654792 206744 654820
rect 171100 654780 171106 654792
rect 206738 654780 206744 654792
rect 206796 654780 206802 654832
rect 235902 654780 235908 654832
rect 235960 654820 235966 654832
rect 257890 654820 257896 654832
rect 235960 654792 257896 654820
rect 235960 654780 235966 654792
rect 257890 654780 257896 654792
rect 257948 654780 257954 654832
rect 267642 654780 267648 654832
rect 267700 654820 267706 654832
rect 274910 654820 274916 654832
rect 267700 654792 274916 654820
rect 267700 654780 267706 654792
rect 274910 654780 274916 654792
rect 274968 654780 274974 654832
rect 284018 654780 284024 654832
rect 284076 654820 284082 654832
rect 291930 654820 291936 654832
rect 284076 654792 291936 654820
rect 284076 654780 284082 654792
rect 291930 654780 291936 654792
rect 291988 654780 291994 654832
rect 300762 654100 300768 654152
rect 300820 654140 300826 654152
rect 308950 654140 308956 654152
rect 300820 654112 308956 654140
rect 300820 654100 300826 654112
rect 308950 654100 308956 654112
rect 309008 654100 309014 654152
rect 3510 645804 3516 645856
rect 3568 645844 3574 645856
rect 59354 645844 59360 645856
rect 3568 645816 59360 645844
rect 3568 645804 3574 645816
rect 59354 645804 59360 645816
rect 59412 645804 59418 645856
rect 523770 638936 523776 638988
rect 523828 638976 523834 638988
rect 580166 638976 580172 638988
rect 523828 638948 580172 638976
rect 523828 638936 523834 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 3418 630572 3424 630624
rect 3476 630612 3482 630624
rect 59354 630612 59360 630624
rect 3476 630584 59360 630612
rect 3476 630572 3482 630584
rect 59354 630572 59360 630584
rect 59412 630572 59418 630624
rect 524322 619556 524328 619608
rect 524380 619596 524386 619608
rect 580258 619596 580264 619608
rect 524380 619568 580264 619596
rect 524380 619556 524386 619568
rect 580258 619556 580264 619568
rect 580316 619556 580322 619608
rect 3602 616768 3608 616820
rect 3660 616808 3666 616820
rect 59354 616808 59360 616820
rect 3660 616780 59360 616808
rect 3660 616768 3666 616780
rect 59354 616768 59360 616780
rect 59412 616768 59418 616820
rect 523126 605752 523132 605804
rect 523184 605792 523190 605804
rect 580442 605792 580448 605804
rect 523184 605764 580448 605792
rect 523184 605752 523190 605764
rect 580442 605752 580448 605764
rect 580500 605752 580506 605804
rect 3510 603032 3516 603084
rect 3568 603072 3574 603084
rect 59354 603072 59360 603084
rect 3568 603044 59360 603072
rect 3568 603032 3574 603044
rect 59354 603032 59360 603044
rect 59412 603032 59418 603084
rect 523678 592016 523684 592068
rect 523736 592056 523742 592068
rect 579798 592056 579804 592068
rect 523736 592028 579804 592056
rect 523736 592016 523742 592028
rect 579798 592016 579804 592028
rect 579856 592016 579862 592068
rect 3418 587800 3424 587852
rect 3476 587840 3482 587852
rect 59354 587840 59360 587852
rect 3476 587812 59360 587840
rect 3476 587800 3482 587812
rect 59354 587800 59360 587812
rect 59412 587800 59418 587852
rect 524322 579572 524328 579624
rect 524380 579612 524386 579624
rect 580350 579612 580356 579624
rect 524380 579584 580356 579612
rect 524380 579572 524386 579584
rect 580350 579572 580356 579584
rect 580408 579572 580414 579624
rect 3510 573996 3516 574048
rect 3568 574036 3574 574048
rect 59354 574036 59360 574048
rect 3568 574008 59360 574036
rect 3568 573996 3574 574008
rect 59354 573996 59360 574008
rect 59412 573996 59418 574048
rect 523126 565768 523132 565820
rect 523184 565808 523190 565820
rect 580442 565808 580448 565820
rect 523184 565780 580448 565808
rect 523184 565768 523190 565780
rect 580442 565768 580448 565780
rect 580500 565768 580506 565820
rect 3418 560192 3424 560244
rect 3476 560232 3482 560244
rect 59354 560232 59360 560244
rect 3476 560204 59360 560232
rect 3476 560192 3482 560204
rect 59354 560192 59360 560204
rect 59412 560192 59418 560244
rect 523770 556180 523776 556232
rect 523828 556220 523834 556232
rect 580166 556220 580172 556232
rect 523828 556192 580172 556220
rect 523828 556180 523834 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 523494 545096 523500 545148
rect 523552 545136 523558 545148
rect 580166 545136 580172 545148
rect 523552 545108 580172 545136
rect 523552 545096 523558 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 3418 545028 3424 545080
rect 3476 545068 3482 545080
rect 59354 545068 59360 545080
rect 3476 545040 59360 545068
rect 3476 545028 3482 545040
rect 59354 545028 59360 545040
rect 59412 545028 59418 545080
rect 523678 539520 523684 539572
rect 523736 539560 523742 539572
rect 580258 539560 580264 539572
rect 523736 539532 580264 539560
rect 523736 539520 523742 539532
rect 580258 539520 580264 539532
rect 580316 539520 580322 539572
rect 3418 531224 3424 531276
rect 3476 531264 3482 531276
rect 59354 531264 59360 531276
rect 3476 531236 59360 531264
rect 3476 531224 3482 531236
rect 59354 531224 59360 531236
rect 59412 531224 59418 531276
rect 3418 516128 3424 516180
rect 3476 516168 3482 516180
rect 59354 516168 59360 516180
rect 3476 516140 59360 516168
rect 3476 516128 3482 516140
rect 59354 516128 59360 516140
rect 59412 516128 59418 516180
rect 523770 509260 523776 509312
rect 523828 509300 523834 509312
rect 580166 509300 580172 509312
rect 523828 509272 580172 509300
rect 523828 509260 523834 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 59354 501004 59360 501016
rect 3384 500976 59360 501004
rect 3384 500964 3390 500976
rect 59354 500964 59360 500976
rect 59412 500964 59418 501016
rect 523678 499468 523684 499520
rect 523736 499508 523742 499520
rect 580258 499508 580264 499520
rect 523736 499480 580264 499508
rect 523736 499468 523742 499480
rect 580258 499468 580264 499480
rect 580316 499468 580322 499520
rect 523678 498176 523684 498228
rect 523736 498216 523742 498228
rect 580166 498216 580172 498228
rect 523736 498188 580172 498216
rect 523736 498176 523742 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3418 487160 3424 487212
rect 3476 487200 3482 487212
rect 59354 487200 59360 487212
rect 3476 487172 59360 487200
rect 3476 487160 3482 487172
rect 59354 487160 59360 487172
rect 59412 487160 59418 487212
rect 3418 473356 3424 473408
rect 3476 473396 3482 473408
rect 59354 473396 59360 473408
rect 3476 473368 59360 473396
rect 3476 473356 3482 473368
rect 59354 473356 59360 473368
rect 59412 473356 59418 473408
rect 523678 462340 523684 462392
rect 523736 462380 523742 462392
rect 580166 462380 580172 462392
rect 523736 462352 580172 462380
rect 523736 462340 523742 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 524322 459484 524328 459536
rect 524380 459524 524386 459536
rect 580258 459524 580264 459536
rect 524380 459496 580264 459524
rect 524380 459484 524386 459496
rect 580258 459484 580264 459496
rect 580316 459484 580322 459536
rect 3510 458192 3516 458244
rect 3568 458232 3574 458244
rect 59354 458232 59360 458244
rect 3568 458204 59360 458232
rect 3568 458192 3574 458204
rect 59354 458192 59360 458204
rect 59412 458192 59418 458244
rect 523770 451256 523776 451308
rect 523828 451296 523834 451308
rect 580166 451296 580172 451308
rect 523828 451268 580172 451296
rect 523828 451256 523834 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 3418 444388 3424 444440
rect 3476 444428 3482 444440
rect 59354 444428 59360 444440
rect 3476 444400 59360 444428
rect 3476 444388 3482 444400
rect 59354 444388 59360 444400
rect 59412 444388 59418 444440
rect 523678 438880 523684 438932
rect 523736 438920 523742 438932
rect 580166 438920 580172 438932
rect 523736 438892 580172 438920
rect 523736 438880 523742 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3602 429156 3608 429208
rect 3660 429196 3666 429208
rect 59354 429196 59360 429208
rect 3660 429168 59360 429196
rect 3660 429156 3666 429168
rect 59354 429156 59360 429168
rect 59412 429156 59418 429208
rect 3418 415420 3424 415472
rect 3476 415460 3482 415472
rect 59354 415460 59360 415472
rect 3476 415432 59360 415460
rect 3476 415420 3482 415432
rect 59354 415420 59360 415432
rect 59412 415420 59418 415472
rect 523678 415420 523684 415472
rect 523736 415460 523742 415472
rect 580166 415460 580172 415472
rect 523736 415432 580172 415460
rect 523736 415420 523742 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 523770 404336 523776 404388
rect 523828 404376 523834 404388
rect 580166 404376 580172 404388
rect 523828 404348 580172 404376
rect 523828 404336 523834 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 401616 3516 401668
rect 3568 401656 3574 401668
rect 59354 401656 59360 401668
rect 3568 401628 59360 401656
rect 3568 401616 3574 401628
rect 59354 401616 59360 401628
rect 59412 401616 59418 401668
rect 523678 391960 523684 392012
rect 523736 392000 523742 392012
rect 580166 392000 580172 392012
rect 523736 391972 580172 392000
rect 523736 391960 523742 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 3602 372580 3608 372632
rect 3660 372620 3666 372632
rect 59354 372620 59360 372632
rect 3660 372592 59360 372620
rect 3660 372580 3666 372592
rect 59354 372580 59360 372592
rect 59412 372580 59418 372632
rect 524230 368500 524236 368552
rect 524288 368540 524294 368552
rect 580166 368540 580172 368552
rect 524288 368512 580172 368540
rect 524288 368500 524294 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 3510 358776 3516 358828
rect 3568 358816 3574 358828
rect 59354 358816 59360 358828
rect 3568 358788 59360 358816
rect 3568 358776 3574 358788
rect 59354 358776 59360 358788
rect 59412 358776 59418 358828
rect 523678 357416 523684 357468
rect 523736 357456 523742 357468
rect 580166 357456 580172 357468
rect 523736 357428 580172 357456
rect 523736 357416 523742 357428
rect 580166 357416 580172 357428
rect 580224 357416 580230 357468
rect 523770 345040 523776 345092
rect 523828 345080 523834 345092
rect 580166 345080 580172 345092
rect 523828 345052 580172 345080
rect 523828 345040 523834 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 3326 338036 3332 338088
rect 3384 338076 3390 338088
rect 60090 338076 60096 338088
rect 3384 338048 60096 338076
rect 3384 338036 3390 338048
rect 60090 338036 60096 338048
rect 60148 338036 60154 338088
rect 3418 329808 3424 329860
rect 3476 329848 3482 329860
rect 59354 329848 59360 329860
rect 3476 329820 59360 329848
rect 3476 329808 3482 329820
rect 59354 329808 59360 329820
rect 59412 329808 59418 329860
rect 524322 322872 524328 322924
rect 524380 322912 524386 322924
rect 580166 322912 580172 322924
rect 524380 322884 580172 322912
rect 524380 322872 524386 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 3602 316004 3608 316056
rect 3660 316044 3666 316056
rect 59354 316044 59360 316056
rect 3660 316016 59360 316044
rect 3660 316004 3666 316016
rect 59354 316004 59360 316016
rect 59412 316004 59418 316056
rect 524322 311788 524328 311840
rect 524380 311828 524386 311840
rect 580166 311828 580172 311840
rect 524380 311800 580172 311828
rect 524380 311788 524386 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 524322 298732 524328 298784
rect 524380 298772 524386 298784
rect 580166 298772 580172 298784
rect 524380 298744 580172 298772
rect 524380 298732 524386 298744
rect 580166 298732 580172 298744
rect 580224 298732 580230 298784
rect 3050 295264 3056 295316
rect 3108 295304 3114 295316
rect 59998 295304 60004 295316
rect 3108 295276 60004 295304
rect 3108 295264 3114 295276
rect 59998 295264 60004 295276
rect 60056 295264 60062 295316
rect 3510 287036 3516 287088
rect 3568 287076 3574 287088
rect 59354 287076 59360 287088
rect 3568 287048 59360 287076
rect 3568 287036 3574 287048
rect 59354 287036 59360 287048
rect 59412 287036 59418 287088
rect 523678 275952 523684 276004
rect 523736 275992 523742 276004
rect 580166 275992 580172 276004
rect 523736 275964 580172 275992
rect 523736 275952 523742 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 3418 273232 3424 273284
rect 3476 273272 3482 273284
rect 59354 273272 59360 273284
rect 3476 273244 59360 273272
rect 3476 273232 3482 273244
rect 59354 273232 59360 273244
rect 59412 273232 59418 273284
rect 523678 264868 523684 264920
rect 523736 264908 523742 264920
rect 580166 264908 580172 264920
rect 523736 264880 580172 264908
rect 523736 264868 523742 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 3142 252492 3148 252544
rect 3200 252532 3206 252544
rect 60090 252532 60096 252544
rect 3200 252504 60096 252532
rect 3200 252492 3206 252504
rect 60090 252492 60096 252504
rect 60148 252492 60154 252544
rect 523678 252492 523684 252544
rect 523736 252532 523742 252544
rect 579798 252532 579804 252544
rect 523736 252504 579804 252532
rect 523736 252492 523742 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 3602 244264 3608 244316
rect 3660 244304 3666 244316
rect 59354 244304 59360 244316
rect 3660 244276 59360 244304
rect 3660 244264 3666 244276
rect 59354 244264 59360 244276
rect 59412 244264 59418 244316
rect 3694 229100 3700 229152
rect 3752 229140 3758 229152
rect 59354 229140 59360 229152
rect 3752 229112 59360 229140
rect 3752 229100 3758 229112
rect 59354 229100 59360 229112
rect 59412 229100 59418 229152
rect 523678 229032 523684 229084
rect 523736 229072 523742 229084
rect 580166 229072 580172 229084
rect 523736 229044 580172 229072
rect 523736 229032 523742 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 523770 217948 523776 218000
rect 523828 217988 523834 218000
rect 580166 217988 580172 218000
rect 523828 217960 580172 217988
rect 523828 217948 523834 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 3142 208292 3148 208344
rect 3200 208332 3206 208344
rect 59998 208332 60004 208344
rect 3200 208304 60004 208332
rect 3200 208292 3206 208304
rect 59998 208292 60004 208304
rect 60056 208292 60062 208344
rect 523862 205572 523868 205624
rect 523920 205612 523926 205624
rect 579798 205612 579804 205624
rect 523920 205584 579804 205612
rect 523920 205572 523926 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 3510 201492 3516 201544
rect 3568 201532 3574 201544
rect 59354 201532 59360 201544
rect 3568 201504 59360 201532
rect 3568 201492 3574 201504
rect 59354 201492 59360 201504
rect 59412 201492 59418 201544
rect 3602 186328 3608 186380
rect 3660 186368 3666 186380
rect 59354 186368 59360 186380
rect 3660 186340 59360 186368
rect 3660 186328 3666 186340
rect 59354 186328 59360 186340
rect 59412 186328 59418 186380
rect 523678 182112 523684 182164
rect 523736 182152 523742 182164
rect 580166 182152 580172 182164
rect 523736 182124 580172 182152
rect 523736 182112 523742 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 523770 171028 523776 171080
rect 523828 171068 523834 171080
rect 580166 171068 580172 171080
rect 523828 171040 580172 171068
rect 523828 171028 523834 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 3418 165520 3424 165572
rect 3476 165560 3482 165572
rect 60090 165560 60096 165572
rect 3476 165532 60096 165560
rect 3476 165520 3482 165532
rect 60090 165520 60096 165532
rect 60148 165520 60154 165572
rect 3418 158720 3424 158772
rect 3476 158760 3482 158772
rect 59354 158760 59360 158772
rect 3476 158732 59360 158760
rect 3476 158720 3482 158732
rect 59354 158720 59360 158732
rect 59412 158720 59418 158772
rect 523862 158652 523868 158704
rect 523920 158692 523926 158704
rect 579798 158692 579804 158704
rect 523920 158664 579804 158692
rect 523920 158652 523926 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 3694 143556 3700 143608
rect 3752 143596 3758 143608
rect 59354 143596 59360 143608
rect 3752 143568 59360 143596
rect 3752 143556 3758 143568
rect 59354 143556 59360 143568
rect 59412 143556 59418 143608
rect 523678 135192 523684 135244
rect 523736 135232 523742 135244
rect 580166 135232 580172 135244
rect 523736 135204 580172 135232
rect 523736 135192 523742 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 523770 124108 523776 124160
rect 523828 124148 523834 124160
rect 580166 124148 580172 124160
rect 523828 124120 580172 124148
rect 523828 124108 523834 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 2958 122748 2964 122800
rect 3016 122788 3022 122800
rect 59998 122788 60004 122800
rect 3016 122760 60004 122788
rect 3016 122748 3022 122760
rect 59998 122748 60004 122760
rect 60056 122748 60062 122800
rect 3510 115948 3516 116000
rect 3568 115988 3574 116000
rect 59354 115988 59360 116000
rect 3568 115960 59360 115988
rect 3568 115948 3574 115960
rect 59354 115948 59360 115960
rect 59412 115948 59418 116000
rect 523862 111732 523868 111784
rect 523920 111772 523926 111784
rect 579798 111772 579804 111784
rect 523920 111744 579804 111772
rect 523920 111732 523926 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3602 100716 3608 100768
rect 3660 100756 3666 100768
rect 59354 100756 59360 100768
rect 3660 100728 59360 100756
rect 3660 100716 3666 100728
rect 59354 100716 59360 100728
rect 59412 100716 59418 100768
rect 523678 88272 523684 88324
rect 523736 88312 523742 88324
rect 580166 88312 580172 88324
rect 523736 88284 580172 88312
rect 523736 88272 523742 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 3050 79976 3056 80028
rect 3108 80016 3114 80028
rect 60090 80016 60096 80028
rect 3108 79988 60096 80016
rect 3108 79976 3114 79988
rect 60090 79976 60096 79988
rect 60148 79976 60154 80028
rect 523770 77188 523776 77240
rect 523828 77228 523834 77240
rect 580166 77228 580172 77240
rect 523828 77200 580172 77228
rect 523828 77188 523834 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 3418 73176 3424 73228
rect 3476 73216 3482 73228
rect 59354 73216 59360 73228
rect 3476 73188 59360 73216
rect 3476 73176 3482 73188
rect 59354 73176 59360 73188
rect 59412 73176 59418 73228
rect 523862 64812 523868 64864
rect 523920 64852 523926 64864
rect 579798 64852 579804 64864
rect 523920 64824 579804 64852
rect 523920 64812 523926 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 3510 57944 3516 57996
rect 3568 57984 3574 57996
rect 59354 57984 59360 57996
rect 3568 57956 59360 57984
rect 3568 57944 3574 57956
rect 59354 57944 59360 57956
rect 59412 57944 59418 57996
rect 81618 49444 81624 49496
rect 81676 49484 81682 49496
rect 142246 49484 142252 49496
rect 81676 49456 142252 49484
rect 81676 49444 81682 49456
rect 142246 49444 142252 49456
rect 142304 49444 142310 49496
rect 167362 49444 167368 49496
rect 167420 49484 167426 49496
rect 227898 49484 227904 49496
rect 167420 49456 227904 49484
rect 167420 49444 167426 49456
rect 227898 49444 227904 49456
rect 227956 49444 227962 49496
rect 110230 49376 110236 49428
rect 110288 49416 110294 49428
rect 171226 49416 171232 49428
rect 110288 49388 171232 49416
rect 110288 49376 110294 49388
rect 171226 49376 171232 49388
rect 171284 49376 171290 49428
rect 403342 49376 403348 49428
rect 403400 49416 403406 49428
rect 463786 49416 463792 49428
rect 403400 49388 463792 49416
rect 403400 49376 403406 49388
rect 463786 49376 463792 49388
rect 463844 49376 463850 49428
rect 138842 49308 138848 49360
rect 138900 49348 138906 49360
rect 200206 49348 200212 49360
rect 138900 49320 200212 49348
rect 138900 49308 138906 49320
rect 200206 49308 200212 49320
rect 200264 49308 200270 49360
rect 210326 49308 210332 49360
rect 210384 49348 210390 49360
rect 270494 49348 270500 49360
rect 210384 49320 270500 49348
rect 210384 49308 210390 49320
rect 270494 49308 270500 49320
rect 270552 49308 270558 49360
rect 396166 49308 396172 49360
rect 396224 49348 396230 49360
rect 456886 49348 456892 49360
rect 396224 49320 456892 49348
rect 396224 49308 396230 49320
rect 456886 49308 456892 49320
rect 456944 49308 456950 49360
rect 95878 49240 95884 49292
rect 95936 49280 95942 49292
rect 157426 49280 157432 49292
rect 95936 49252 157432 49280
rect 95936 49240 95942 49252
rect 157426 49240 157432 49252
rect 157484 49240 157490 49292
rect 174538 49240 174544 49292
rect 174596 49280 174602 49292
rect 236178 49280 236184 49292
rect 174596 49252 236184 49280
rect 174596 49240 174602 49252
rect 236178 49240 236184 49252
rect 236236 49240 236242 49292
rect 253198 49240 253204 49292
rect 253256 49280 253262 49292
rect 313458 49280 313464 49292
rect 253256 49252 313464 49280
rect 253256 49240 253262 49252
rect 313458 49240 313464 49252
rect 313516 49240 313522 49292
rect 367646 49240 367652 49292
rect 367704 49280 367710 49292
rect 427906 49280 427912 49292
rect 367704 49252 427912 49280
rect 367704 49240 367710 49252
rect 427906 49240 427912 49252
rect 427964 49240 427970 49292
rect 131666 49172 131672 49224
rect 131724 49212 131730 49224
rect 193398 49212 193404 49224
rect 131724 49184 193404 49212
rect 131724 49172 131730 49184
rect 193398 49172 193404 49184
rect 193456 49172 193462 49224
rect 217410 49172 217416 49224
rect 217468 49212 217474 49224
rect 278958 49212 278964 49224
rect 217468 49184 278964 49212
rect 217468 49172 217474 49184
rect 278958 49172 278964 49184
rect 279016 49172 279022 49224
rect 374730 49172 374736 49224
rect 374788 49212 374794 49224
rect 434806 49212 434812 49224
rect 374788 49184 434812 49212
rect 374788 49172 374794 49184
rect 434806 49172 434812 49184
rect 434864 49172 434870 49224
rect 482002 49172 482008 49224
rect 482060 49212 482066 49224
rect 542354 49212 542360 49224
rect 482060 49184 542360 49212
rect 482060 49172 482066 49184
rect 542354 49172 542360 49184
rect 542412 49172 542418 49224
rect 103054 49104 103060 49156
rect 103112 49144 103118 49156
rect 164326 49144 164332 49156
rect 103112 49116 164332 49144
rect 103112 49104 103118 49116
rect 164326 49104 164332 49116
rect 164384 49104 164390 49156
rect 181714 49104 181720 49156
rect 181772 49144 181778 49156
rect 242986 49144 242992 49156
rect 181772 49116 242992 49144
rect 181772 49104 181778 49116
rect 242986 49104 242992 49116
rect 243044 49104 243050 49156
rect 260374 49104 260380 49156
rect 260432 49144 260438 49156
rect 321738 49144 321744 49156
rect 260432 49116 321744 49144
rect 260432 49104 260438 49116
rect 321738 49104 321744 49116
rect 321796 49104 321802 49156
rect 346118 49104 346124 49156
rect 346176 49144 346182 49156
rect 407206 49144 407212 49156
rect 346176 49116 407212 49144
rect 346176 49104 346182 49116
rect 407206 49104 407212 49116
rect 407264 49104 407270 49156
rect 474826 49104 474832 49156
rect 474884 49144 474890 49156
rect 535454 49144 535460 49156
rect 474884 49116 535460 49144
rect 474884 49104 474890 49116
rect 535454 49104 535460 49116
rect 535512 49104 535518 49156
rect 88702 49036 88708 49088
rect 88760 49076 88766 49088
rect 150618 49076 150624 49088
rect 88760 49048 150624 49076
rect 88760 49036 88766 49048
rect 150618 49036 150624 49048
rect 150676 49036 150682 49088
rect 188890 49036 188896 49088
rect 188948 49076 188954 49088
rect 249886 49076 249892 49088
rect 188948 49048 249892 49076
rect 188948 49036 188954 49048
rect 249886 49036 249892 49048
rect 249944 49036 249950 49088
rect 267458 49036 267464 49088
rect 267516 49076 267522 49088
rect 328546 49076 328552 49088
rect 267516 49048 328552 49076
rect 267516 49036 267522 49048
rect 328546 49036 328552 49048
rect 328604 49036 328610 49088
rect 344922 49036 344928 49088
rect 344980 49076 344986 49088
rect 351178 49076 351184 49088
rect 344980 49048 351184 49076
rect 344980 49036 344986 49048
rect 351178 49036 351184 49048
rect 351236 49036 351242 49088
rect 389082 49036 389088 49088
rect 389140 49076 389146 49088
rect 449986 49076 449992 49088
rect 389140 49048 449992 49076
rect 389140 49036 389146 49048
rect 449986 49036 449992 49048
rect 450044 49036 450050 49088
rect 489178 49036 489184 49088
rect 489236 49076 489242 49088
rect 549254 49076 549260 49088
rect 489236 49048 549260 49076
rect 489236 49036 489242 49048
rect 549254 49036 549260 49048
rect 549312 49036 549318 49088
rect 67266 48968 67272 49020
rect 67324 49008 67330 49020
rect 128446 49008 128452 49020
rect 67324 48980 128452 49008
rect 67324 48968 67330 48980
rect 128446 48968 128452 48980
rect 128504 48968 128510 49020
rect 145926 48968 145932 49020
rect 145984 49008 145990 49020
rect 207106 49008 207112 49020
rect 145984 48980 207112 49008
rect 145984 48968 145990 48980
rect 207106 48968 207112 48980
rect 207164 48968 207170 49020
rect 224586 48968 224592 49020
rect 224644 49008 224650 49020
rect 285766 49008 285772 49020
rect 224644 48980 285772 49008
rect 224644 48968 224650 48980
rect 285766 48968 285772 48980
rect 285824 48968 285830 49020
rect 318702 48968 318708 49020
rect 318760 49008 318766 49020
rect 345658 49008 345664 49020
rect 318760 48980 345664 49008
rect 318760 48968 318766 48980
rect 345658 48968 345664 48980
rect 345716 48968 345722 49020
rect 354490 48968 354496 49020
rect 354548 49008 354554 49020
rect 367738 49008 367744 49020
rect 354548 48980 367744 49008
rect 354548 48968 354554 48980
rect 367738 48968 367744 48980
rect 367796 48968 367802 49020
rect 381906 48968 381912 49020
rect 381964 49008 381970 49020
rect 443178 49008 443184 49020
rect 381964 48980 443184 49008
rect 381964 48968 381970 48980
rect 443178 48968 443184 48980
rect 443236 48968 443242 49020
rect 467742 48968 467748 49020
rect 467800 49008 467806 49020
rect 528554 49008 528560 49020
rect 467800 48980 528560 49008
rect 467800 48968 467806 48980
rect 528554 48968 528560 48980
rect 528612 48968 528618 49020
rect 379514 48832 379520 48884
rect 379572 48872 379578 48884
rect 380802 48872 380808 48884
rect 379572 48844 380808 48872
rect 379572 48832 379578 48844
rect 380802 48832 380808 48844
rect 380860 48832 380866 48884
rect 66070 48764 66076 48816
rect 66128 48804 66134 48816
rect 66898 48804 66904 48816
rect 66128 48776 66904 48804
rect 66128 48764 66134 48776
rect 66898 48764 66904 48776
rect 66956 48764 66962 48816
rect 70854 48764 70860 48816
rect 70912 48804 70918 48816
rect 71682 48804 71688 48816
rect 70912 48776 71688 48804
rect 70912 48764 70918 48776
rect 71682 48764 71688 48776
rect 71740 48764 71746 48816
rect 72050 48764 72056 48816
rect 72108 48804 72114 48816
rect 73062 48804 73068 48816
rect 72108 48776 73068 48804
rect 72108 48764 72114 48776
rect 73062 48764 73068 48776
rect 73120 48764 73126 48816
rect 73246 48764 73252 48816
rect 73304 48804 73310 48816
rect 74350 48804 74356 48816
rect 73304 48776 74356 48804
rect 73304 48764 73310 48776
rect 74350 48764 74356 48776
rect 74408 48764 74414 48816
rect 89898 48764 89904 48816
rect 89956 48804 89962 48816
rect 91002 48804 91008 48816
rect 89956 48776 91008 48804
rect 89956 48764 89962 48776
rect 91002 48764 91008 48776
rect 91060 48764 91066 48816
rect 91094 48764 91100 48816
rect 91152 48804 91158 48816
rect 92290 48804 92296 48816
rect 91152 48776 92296 48804
rect 91152 48764 91158 48776
rect 92290 48764 92296 48776
rect 92348 48764 92354 48816
rect 97074 48764 97080 48816
rect 97132 48804 97138 48816
rect 97902 48804 97908 48816
rect 97132 48776 97908 48804
rect 97132 48764 97138 48776
rect 97902 48764 97908 48776
rect 97960 48764 97966 48816
rect 98270 48764 98276 48816
rect 98328 48804 98334 48816
rect 99282 48804 99288 48816
rect 98328 48776 99288 48804
rect 98328 48764 98334 48776
rect 99282 48764 99288 48776
rect 99340 48764 99346 48816
rect 99466 48764 99472 48816
rect 99524 48804 99530 48816
rect 100662 48804 100668 48816
rect 99524 48776 100668 48804
rect 99524 48764 99530 48776
rect 100662 48764 100668 48776
rect 100720 48764 100726 48816
rect 105446 48764 105452 48816
rect 105504 48804 105510 48816
rect 106182 48804 106188 48816
rect 105504 48776 106188 48804
rect 105504 48764 105510 48776
rect 106182 48764 106188 48776
rect 106240 48764 106246 48816
rect 106642 48764 106648 48816
rect 106700 48804 106706 48816
rect 107562 48804 107568 48816
rect 106700 48776 107568 48804
rect 106700 48764 106706 48776
rect 107562 48764 107568 48776
rect 107620 48764 107626 48816
rect 107838 48764 107844 48816
rect 107896 48804 107902 48816
rect 108942 48804 108948 48816
rect 107896 48776 108948 48804
rect 107896 48764 107902 48776
rect 108942 48764 108948 48776
rect 109000 48764 109006 48816
rect 109034 48764 109040 48816
rect 109092 48804 109098 48816
rect 110322 48804 110328 48816
rect 109092 48776 110328 48804
rect 109092 48764 109098 48776
rect 110322 48764 110328 48776
rect 110380 48764 110386 48816
rect 113726 48764 113732 48816
rect 113784 48804 113790 48816
rect 114462 48804 114468 48816
rect 113784 48776 114468 48804
rect 113784 48764 113790 48776
rect 114462 48764 114468 48776
rect 114520 48764 114526 48816
rect 114922 48764 114928 48816
rect 114980 48804 114986 48816
rect 115842 48804 115848 48816
rect 114980 48776 115848 48804
rect 114980 48764 114986 48776
rect 115842 48764 115848 48776
rect 115900 48764 115906 48816
rect 116118 48764 116124 48816
rect 116176 48804 116182 48816
rect 117222 48804 117228 48816
rect 116176 48776 117228 48804
rect 116176 48764 116182 48776
rect 117222 48764 117228 48776
rect 117280 48764 117286 48816
rect 117314 48764 117320 48816
rect 117372 48804 117378 48816
rect 118602 48804 118608 48816
rect 117372 48776 118608 48804
rect 117372 48764 117378 48776
rect 118602 48764 118608 48776
rect 118660 48764 118666 48816
rect 124490 48764 124496 48816
rect 124548 48804 124554 48816
rect 125502 48804 125508 48816
rect 124548 48776 125508 48804
rect 124548 48764 124554 48776
rect 125502 48764 125508 48776
rect 125560 48764 125566 48816
rect 132862 48764 132868 48816
rect 132920 48804 132926 48816
rect 133782 48804 133788 48816
rect 132920 48776 133788 48804
rect 132920 48764 132926 48776
rect 133782 48764 133788 48776
rect 133840 48764 133846 48816
rect 134058 48764 134064 48816
rect 134116 48804 134122 48816
rect 135162 48804 135168 48816
rect 134116 48776 135168 48804
rect 134116 48764 134122 48776
rect 135162 48764 135168 48776
rect 135220 48764 135226 48816
rect 135254 48764 135260 48816
rect 135312 48804 135318 48816
rect 136542 48804 136548 48816
rect 135312 48776 136548 48804
rect 135312 48764 135318 48776
rect 136542 48764 136548 48776
rect 136600 48764 136606 48816
rect 141142 48764 141148 48816
rect 141200 48804 141206 48816
rect 142062 48804 142068 48816
rect 141200 48776 142068 48804
rect 141200 48764 141206 48776
rect 142062 48764 142068 48776
rect 142120 48764 142126 48816
rect 142338 48764 142344 48816
rect 142396 48804 142402 48816
rect 143442 48804 143448 48816
rect 142396 48776 143448 48804
rect 142396 48764 142402 48776
rect 143442 48764 143448 48776
rect 143500 48764 143506 48816
rect 143534 48764 143540 48816
rect 143592 48804 143598 48816
rect 144822 48804 144828 48816
rect 143592 48776 144828 48804
rect 143592 48764 143598 48776
rect 144822 48764 144828 48776
rect 144880 48764 144886 48816
rect 149514 48764 149520 48816
rect 149572 48804 149578 48816
rect 150342 48804 150348 48816
rect 149572 48776 150348 48804
rect 149572 48764 149578 48776
rect 150342 48764 150348 48776
rect 150400 48764 150406 48816
rect 150710 48764 150716 48816
rect 150768 48804 150774 48816
rect 151722 48804 151728 48816
rect 150768 48776 151728 48804
rect 150768 48764 150774 48776
rect 151722 48764 151728 48776
rect 151780 48764 151786 48816
rect 159082 48764 159088 48816
rect 159140 48804 159146 48816
rect 160002 48804 160008 48816
rect 159140 48776 160008 48804
rect 159140 48764 159146 48776
rect 160002 48764 160008 48776
rect 160060 48764 160066 48816
rect 160278 48764 160284 48816
rect 160336 48804 160342 48816
rect 161382 48804 161388 48816
rect 160336 48776 161388 48804
rect 160336 48764 160342 48776
rect 161382 48764 161388 48776
rect 161440 48764 161446 48816
rect 161474 48764 161480 48816
rect 161532 48804 161538 48816
rect 162762 48804 162768 48816
rect 161532 48776 162768 48804
rect 161532 48764 161538 48776
rect 162762 48764 162768 48776
rect 162820 48764 162826 48816
rect 166166 48764 166172 48816
rect 166224 48804 166230 48816
rect 166902 48804 166908 48816
rect 166224 48776 166908 48804
rect 166224 48764 166230 48776
rect 166902 48764 166908 48776
rect 166960 48764 166966 48816
rect 168558 48764 168564 48816
rect 168616 48804 168622 48816
rect 169662 48804 169668 48816
rect 168616 48776 169668 48804
rect 168616 48764 168622 48776
rect 169662 48764 169668 48776
rect 169720 48764 169726 48816
rect 169754 48764 169760 48816
rect 169812 48804 169818 48816
rect 170950 48804 170956 48816
rect 169812 48776 170956 48804
rect 169812 48764 169818 48776
rect 170950 48764 170956 48776
rect 171008 48764 171014 48816
rect 175734 48764 175740 48816
rect 175792 48804 175798 48816
rect 176562 48804 176568 48816
rect 175792 48776 176568 48804
rect 175792 48764 175798 48776
rect 176562 48764 176568 48776
rect 176620 48764 176626 48816
rect 178126 48764 178132 48816
rect 178184 48804 178190 48816
rect 179322 48804 179328 48816
rect 178184 48776 179328 48804
rect 178184 48764 178190 48776
rect 179322 48764 179328 48776
rect 179380 48764 179386 48816
rect 185302 48764 185308 48816
rect 185360 48804 185366 48816
rect 186222 48804 186228 48816
rect 185360 48776 186228 48804
rect 185360 48764 185366 48776
rect 186222 48764 186228 48776
rect 186280 48764 186286 48816
rect 187694 48764 187700 48816
rect 187752 48804 187758 48816
rect 188982 48804 188988 48816
rect 187752 48776 188988 48804
rect 187752 48764 187758 48776
rect 188982 48764 188988 48776
rect 189040 48764 189046 48816
rect 193582 48764 193588 48816
rect 193640 48804 193646 48816
rect 194502 48804 194508 48816
rect 193640 48776 194508 48804
rect 193640 48764 193646 48776
rect 194502 48764 194508 48776
rect 194560 48764 194566 48816
rect 194778 48764 194784 48816
rect 194836 48804 194842 48816
rect 195882 48804 195888 48816
rect 194836 48776 195888 48804
rect 194836 48764 194842 48776
rect 195882 48764 195888 48776
rect 195940 48764 195946 48816
rect 203150 48764 203156 48816
rect 203208 48804 203214 48816
rect 204162 48804 204168 48816
rect 203208 48776 204168 48804
rect 203208 48764 203214 48776
rect 204162 48764 204168 48776
rect 204220 48764 204226 48816
rect 204346 48764 204352 48816
rect 204404 48804 204410 48816
rect 205450 48804 205456 48816
rect 204404 48776 205456 48804
rect 204404 48764 204410 48776
rect 205450 48764 205456 48776
rect 205508 48764 205514 48816
rect 211522 48764 211528 48816
rect 211580 48804 211586 48816
rect 212442 48804 212448 48816
rect 211580 48776 212448 48804
rect 211580 48764 211586 48776
rect 212442 48764 212448 48776
rect 212500 48764 212506 48816
rect 212718 48764 212724 48816
rect 212776 48804 212782 48816
rect 213822 48804 213828 48816
rect 212776 48776 213828 48804
rect 212776 48764 212782 48776
rect 213822 48764 213828 48776
rect 213880 48764 213886 48816
rect 213914 48764 213920 48816
rect 213972 48804 213978 48816
rect 215202 48804 215208 48816
rect 213972 48776 215208 48804
rect 213972 48764 213978 48776
rect 215202 48764 215208 48776
rect 215260 48764 215266 48816
rect 218606 48764 218612 48816
rect 218664 48804 218670 48816
rect 219342 48804 219348 48816
rect 218664 48776 219348 48804
rect 218664 48764 218670 48776
rect 219342 48764 219348 48776
rect 219400 48764 219406 48816
rect 219802 48764 219808 48816
rect 219860 48804 219866 48816
rect 220722 48804 220728 48816
rect 219860 48776 220728 48804
rect 219860 48764 219866 48776
rect 220722 48764 220728 48776
rect 220780 48764 220786 48816
rect 220998 48764 221004 48816
rect 221056 48804 221062 48816
rect 222102 48804 222108 48816
rect 221056 48776 222108 48804
rect 221056 48764 221062 48776
rect 222102 48764 222108 48776
rect 222160 48764 222166 48816
rect 222194 48764 222200 48816
rect 222252 48804 222258 48816
rect 223482 48804 223488 48816
rect 222252 48776 223488 48804
rect 222252 48764 222258 48776
rect 223482 48764 223488 48776
rect 223540 48764 223546 48816
rect 228174 48764 228180 48816
rect 228232 48804 228238 48816
rect 229002 48804 229008 48816
rect 228232 48776 229008 48804
rect 228232 48764 228238 48776
rect 229002 48764 229008 48776
rect 229060 48764 229066 48816
rect 229370 48764 229376 48816
rect 229428 48804 229434 48816
rect 230382 48804 230388 48816
rect 229428 48776 230388 48804
rect 229428 48764 229434 48776
rect 230382 48764 230388 48776
rect 230440 48764 230446 48816
rect 237742 48764 237748 48816
rect 237800 48804 237806 48816
rect 238662 48804 238668 48816
rect 237800 48776 238668 48804
rect 237800 48764 237806 48776
rect 238662 48764 238668 48776
rect 238720 48764 238726 48816
rect 238938 48764 238944 48816
rect 238996 48804 239002 48816
rect 240042 48804 240048 48816
rect 238996 48776 240048 48804
rect 238996 48764 239002 48776
rect 240042 48764 240048 48776
rect 240100 48764 240106 48816
rect 240134 48764 240140 48816
rect 240192 48804 240198 48816
rect 241422 48804 241428 48816
rect 240192 48776 241428 48804
rect 240192 48764 240198 48776
rect 241422 48764 241428 48776
rect 241480 48764 241486 48816
rect 246022 48764 246028 48816
rect 246080 48804 246086 48816
rect 246942 48804 246948 48816
rect 246080 48776 246948 48804
rect 246080 48764 246086 48776
rect 246942 48764 246948 48776
rect 247000 48764 247006 48816
rect 247218 48764 247224 48816
rect 247276 48804 247282 48816
rect 248322 48804 248328 48816
rect 247276 48776 248328 48804
rect 247276 48764 247282 48776
rect 248322 48764 248328 48776
rect 248380 48764 248386 48816
rect 248414 48764 248420 48816
rect 248472 48804 248478 48816
rect 249610 48804 249616 48816
rect 248472 48776 249616 48804
rect 248472 48764 248478 48776
rect 249610 48764 249616 48776
rect 249668 48764 249674 48816
rect 254394 48764 254400 48816
rect 254452 48804 254458 48816
rect 255222 48804 255228 48816
rect 254452 48776 255228 48804
rect 254452 48764 254458 48776
rect 255222 48764 255228 48776
rect 255280 48764 255286 48816
rect 255590 48764 255596 48816
rect 255648 48804 255654 48816
rect 256602 48804 256608 48816
rect 255648 48776 256608 48804
rect 255648 48764 255654 48776
rect 256602 48764 256608 48776
rect 256660 48764 256666 48816
rect 256786 48764 256792 48816
rect 256844 48804 256850 48816
rect 257982 48804 257988 48816
rect 256844 48776 257988 48804
rect 256844 48764 256850 48776
rect 257982 48764 257988 48776
rect 258040 48764 258046 48816
rect 263962 48764 263968 48816
rect 264020 48804 264026 48816
rect 264882 48804 264888 48816
rect 264020 48776 264888 48804
rect 264020 48764 264026 48776
rect 264882 48764 264888 48776
rect 264940 48764 264946 48816
rect 265158 48764 265164 48816
rect 265216 48804 265222 48816
rect 266262 48804 266268 48816
rect 265216 48776 266268 48804
rect 265216 48764 265222 48776
rect 266262 48764 266268 48776
rect 266320 48764 266326 48816
rect 266354 48764 266360 48816
rect 266412 48804 266418 48816
rect 267642 48804 267648 48816
rect 266412 48776 267648 48804
rect 266412 48764 266418 48776
rect 267642 48764 267648 48776
rect 267700 48764 267706 48816
rect 272242 48764 272248 48816
rect 272300 48804 272306 48816
rect 273162 48804 273168 48816
rect 272300 48776 273168 48804
rect 272300 48764 272306 48776
rect 273162 48764 273168 48776
rect 273220 48764 273226 48816
rect 273438 48764 273444 48816
rect 273496 48804 273502 48816
rect 274542 48804 274548 48816
rect 273496 48776 274548 48804
rect 273496 48764 273502 48776
rect 274542 48764 274548 48776
rect 274600 48764 274606 48816
rect 274634 48764 274640 48816
rect 274692 48804 274698 48816
rect 275830 48804 275836 48816
rect 274692 48776 275836 48804
rect 274692 48764 274698 48776
rect 275830 48764 275836 48776
rect 275888 48764 275894 48816
rect 280614 48764 280620 48816
rect 280672 48804 280678 48816
rect 281442 48804 281448 48816
rect 280672 48776 281448 48804
rect 280672 48764 280678 48776
rect 281442 48764 281448 48776
rect 281500 48764 281506 48816
rect 281810 48764 281816 48816
rect 281868 48804 281874 48816
rect 282822 48804 282828 48816
rect 281868 48776 282828 48804
rect 281868 48764 281874 48776
rect 282822 48764 282828 48776
rect 282880 48764 282886 48816
rect 283006 48764 283012 48816
rect 283064 48804 283070 48816
rect 284202 48804 284208 48816
rect 283064 48776 284208 48804
rect 283064 48764 283070 48776
rect 284202 48764 284208 48776
rect 284260 48764 284266 48816
rect 291378 48764 291384 48816
rect 291436 48804 291442 48816
rect 292482 48804 292488 48816
rect 291436 48776 292488 48804
rect 291436 48764 291442 48776
rect 292482 48764 292488 48776
rect 292540 48764 292546 48816
rect 292574 48764 292580 48816
rect 292632 48804 292638 48816
rect 293862 48804 293868 48816
rect 292632 48776 293868 48804
rect 292632 48764 292638 48776
rect 293862 48764 293868 48776
rect 293920 48764 293926 48816
rect 299658 48764 299664 48816
rect 299716 48804 299722 48816
rect 300762 48804 300768 48816
rect 299716 48776 300768 48804
rect 299716 48764 299722 48776
rect 300762 48764 300768 48776
rect 300820 48764 300826 48816
rect 300854 48764 300860 48816
rect 300912 48804 300918 48816
rect 302142 48804 302148 48816
rect 300912 48776 302148 48804
rect 300912 48764 300918 48776
rect 302142 48764 302148 48776
rect 302200 48764 302206 48816
rect 306834 48764 306840 48816
rect 306892 48804 306898 48816
rect 307662 48804 307668 48816
rect 306892 48776 307668 48804
rect 306892 48764 306898 48776
rect 307662 48764 307668 48776
rect 307720 48764 307726 48816
rect 309226 48764 309232 48816
rect 309284 48804 309290 48816
rect 310330 48804 310336 48816
rect 309284 48776 310336 48804
rect 309284 48764 309290 48776
rect 310330 48764 310336 48776
rect 310388 48764 310394 48816
rect 323486 48764 323492 48816
rect 323544 48804 323550 48816
rect 324222 48804 324228 48816
rect 323544 48776 324228 48804
rect 323544 48764 323550 48776
rect 324222 48764 324228 48776
rect 324280 48764 324286 48816
rect 324682 48764 324688 48816
rect 324740 48804 324746 48816
rect 325602 48804 325608 48816
rect 324740 48776 325608 48804
rect 324740 48764 324746 48776
rect 325602 48764 325608 48776
rect 325660 48764 325666 48816
rect 325878 48764 325884 48816
rect 325936 48804 325942 48816
rect 326982 48804 326988 48816
rect 325936 48776 326988 48804
rect 325936 48764 325942 48776
rect 326982 48764 326988 48776
rect 327040 48764 327046 48816
rect 327074 48764 327080 48816
rect 327132 48804 327138 48816
rect 328270 48804 328276 48816
rect 327132 48776 328276 48804
rect 327132 48764 327138 48776
rect 328270 48764 328276 48776
rect 328328 48764 328334 48816
rect 333054 48764 333060 48816
rect 333112 48804 333118 48816
rect 333882 48804 333888 48816
rect 333112 48776 333888 48804
rect 333112 48764 333118 48776
rect 333882 48764 333888 48776
rect 333940 48764 333946 48816
rect 334250 48764 334256 48816
rect 334308 48804 334314 48816
rect 335262 48804 335268 48816
rect 334308 48776 335268 48804
rect 334308 48764 334314 48776
rect 335262 48764 335268 48776
rect 335320 48764 335326 48816
rect 335446 48764 335452 48816
rect 335504 48804 335510 48816
rect 336642 48804 336648 48816
rect 335504 48776 336648 48804
rect 335504 48764 335510 48776
rect 336642 48764 336648 48776
rect 336700 48764 336706 48816
rect 342622 48764 342628 48816
rect 342680 48804 342686 48816
rect 343542 48804 343548 48816
rect 342680 48776 343548 48804
rect 342680 48764 342686 48776
rect 343542 48764 343548 48776
rect 343600 48764 343606 48816
rect 343726 48764 343732 48816
rect 343784 48804 343790 48816
rect 344922 48804 344928 48816
rect 343784 48776 344928 48804
rect 343784 48764 343790 48776
rect 344922 48764 344928 48776
rect 344980 48764 344986 48816
rect 350902 48764 350908 48816
rect 350960 48804 350966 48816
rect 351822 48804 351828 48816
rect 350960 48776 351828 48804
rect 350960 48764 350966 48776
rect 351822 48764 351828 48776
rect 351880 48764 351886 48816
rect 352098 48764 352104 48816
rect 352156 48804 352162 48816
rect 353202 48804 353208 48816
rect 352156 48776 353208 48804
rect 352156 48764 352162 48776
rect 353202 48764 353208 48776
rect 353260 48764 353266 48816
rect 353294 48764 353300 48816
rect 353352 48804 353358 48816
rect 354582 48804 354588 48816
rect 353352 48776 354588 48804
rect 353352 48764 353358 48776
rect 354582 48764 354588 48776
rect 354640 48764 354646 48816
rect 359274 48764 359280 48816
rect 359332 48804 359338 48816
rect 360102 48804 360108 48816
rect 359332 48776 360108 48804
rect 359332 48764 359338 48776
rect 360102 48764 360108 48776
rect 360160 48764 360166 48816
rect 360470 48764 360476 48816
rect 360528 48804 360534 48816
rect 361482 48804 361488 48816
rect 360528 48776 361488 48804
rect 360528 48764 360534 48776
rect 361482 48764 361488 48776
rect 361540 48764 361546 48816
rect 361666 48764 361672 48816
rect 361724 48804 361730 48816
rect 362862 48804 362868 48816
rect 361724 48776 362868 48804
rect 361724 48764 361730 48776
rect 362862 48764 362868 48776
rect 362920 48764 362926 48816
rect 377122 48764 377128 48816
rect 377180 48804 377186 48816
rect 378042 48804 378048 48816
rect 377180 48776 378048 48804
rect 377180 48764 377186 48776
rect 378042 48764 378048 48776
rect 378100 48764 378106 48816
rect 378318 48764 378324 48816
rect 378376 48804 378382 48816
rect 379422 48804 379428 48816
rect 378376 48776 379428 48804
rect 378376 48764 378382 48776
rect 379422 48764 379428 48776
rect 379480 48764 379486 48816
rect 380710 48764 380716 48816
rect 380768 48804 380774 48816
rect 381538 48804 381544 48816
rect 380768 48776 381544 48804
rect 380768 48764 380774 48776
rect 381538 48764 381544 48776
rect 381596 48764 381602 48816
rect 386690 48764 386696 48816
rect 386748 48804 386754 48816
rect 387702 48804 387708 48816
rect 386748 48776 387708 48804
rect 386748 48764 386754 48776
rect 387702 48764 387708 48776
rect 387760 48764 387766 48816
rect 387886 48764 387892 48816
rect 387944 48804 387950 48816
rect 389082 48804 389088 48816
rect 387944 48776 389088 48804
rect 387944 48764 387950 48776
rect 389082 48764 389088 48776
rect 389140 48764 389146 48816
rect 394970 48764 394976 48816
rect 395028 48804 395034 48816
rect 395982 48804 395988 48816
rect 395028 48776 395988 48804
rect 395028 48764 395034 48776
rect 395982 48764 395988 48776
rect 396040 48764 396046 48816
rect 404538 48764 404544 48816
rect 404596 48804 404602 48816
rect 405642 48804 405648 48816
rect 404596 48776 405648 48804
rect 404596 48764 404602 48776
rect 405642 48764 405648 48776
rect 405700 48764 405706 48816
rect 411714 48764 411720 48816
rect 411772 48804 411778 48816
rect 412542 48804 412548 48816
rect 411772 48776 412548 48804
rect 411772 48764 411778 48776
rect 412542 48764 412548 48776
rect 412600 48764 412606 48816
rect 412910 48764 412916 48816
rect 412968 48804 412974 48816
rect 413922 48804 413928 48816
rect 412968 48776 413928 48804
rect 412968 48764 412974 48776
rect 413922 48764 413928 48776
rect 413980 48764 413986 48816
rect 414106 48764 414112 48816
rect 414164 48804 414170 48816
rect 415302 48804 415308 48816
rect 414164 48776 415308 48804
rect 414164 48764 414170 48776
rect 415302 48764 415308 48776
rect 415360 48764 415366 48816
rect 420086 48764 420092 48816
rect 420144 48804 420150 48816
rect 420822 48804 420828 48816
rect 420144 48776 420828 48804
rect 420144 48764 420150 48776
rect 420822 48764 420828 48776
rect 420880 48764 420886 48816
rect 421190 48764 421196 48816
rect 421248 48804 421254 48816
rect 422202 48804 422208 48816
rect 421248 48776 422208 48804
rect 421248 48764 421254 48776
rect 422202 48764 422208 48776
rect 422260 48764 422266 48816
rect 428366 48764 428372 48816
rect 428424 48804 428430 48816
rect 429102 48804 429108 48816
rect 428424 48776 429108 48804
rect 428424 48764 428430 48776
rect 429102 48764 429108 48776
rect 429160 48764 429166 48816
rect 429562 48764 429568 48816
rect 429620 48804 429626 48816
rect 430482 48804 430488 48816
rect 429620 48776 430488 48804
rect 429620 48764 429626 48776
rect 430482 48764 430488 48776
rect 430540 48764 430546 48816
rect 430758 48764 430764 48816
rect 430816 48804 430822 48816
rect 431862 48804 431868 48816
rect 430816 48776 431868 48804
rect 430816 48764 430822 48776
rect 431862 48764 431868 48776
rect 431920 48764 431926 48816
rect 431954 48764 431960 48816
rect 432012 48804 432018 48816
rect 433150 48804 433156 48816
rect 432012 48776 433156 48804
rect 432012 48764 432018 48776
rect 433150 48764 433156 48776
rect 433208 48764 433214 48816
rect 437934 48764 437940 48816
rect 437992 48804 437998 48816
rect 438762 48804 438768 48816
rect 437992 48776 438768 48804
rect 437992 48764 437998 48776
rect 438762 48764 438768 48776
rect 438820 48764 438826 48816
rect 439130 48764 439136 48816
rect 439188 48804 439194 48816
rect 440142 48804 440148 48816
rect 439188 48776 440148 48804
rect 439188 48764 439194 48776
rect 440142 48764 440148 48776
rect 440200 48764 440206 48816
rect 440326 48764 440332 48816
rect 440384 48804 440390 48816
rect 441522 48804 441528 48816
rect 440384 48776 441528 48804
rect 440384 48764 440390 48776
rect 441522 48764 441528 48776
rect 441580 48764 441586 48816
rect 446214 48764 446220 48816
rect 446272 48804 446278 48816
rect 447042 48804 447048 48816
rect 446272 48776 447048 48804
rect 446272 48764 446278 48776
rect 447042 48764 447048 48776
rect 447100 48764 447106 48816
rect 447410 48764 447416 48816
rect 447468 48804 447474 48816
rect 448422 48804 448428 48816
rect 447468 48776 448428 48804
rect 447468 48764 447474 48776
rect 448422 48764 448428 48776
rect 448480 48764 448486 48816
rect 448606 48764 448612 48816
rect 448664 48804 448670 48816
rect 449710 48804 449716 48816
rect 448664 48776 449716 48804
rect 448664 48764 448670 48776
rect 449710 48764 449716 48776
rect 449768 48764 449774 48816
rect 455782 48764 455788 48816
rect 455840 48804 455846 48816
rect 456702 48804 456708 48816
rect 455840 48776 456708 48804
rect 455840 48764 455846 48776
rect 456702 48764 456708 48776
rect 456760 48764 456766 48816
rect 456978 48764 456984 48816
rect 457036 48804 457042 48816
rect 458082 48804 458088 48816
rect 457036 48776 458088 48804
rect 457036 48764 457042 48776
rect 458082 48764 458088 48776
rect 458140 48764 458146 48816
rect 458174 48764 458180 48816
rect 458232 48804 458238 48816
rect 459462 48804 459468 48816
rect 458232 48776 459468 48804
rect 458232 48764 458238 48776
rect 459462 48764 459468 48776
rect 459520 48764 459526 48816
rect 464154 48764 464160 48816
rect 464212 48804 464218 48816
rect 464982 48804 464988 48816
rect 464212 48776 464988 48804
rect 464212 48764 464218 48776
rect 464982 48764 464988 48776
rect 465040 48764 465046 48816
rect 465350 48764 465356 48816
rect 465408 48804 465414 48816
rect 466362 48804 466368 48816
rect 465408 48776 466368 48804
rect 465408 48764 465414 48776
rect 466362 48764 466368 48776
rect 466420 48764 466426 48816
rect 466546 48764 466552 48816
rect 466604 48804 466610 48816
rect 467742 48804 467748 48816
rect 466604 48776 467748 48804
rect 466604 48764 466610 48776
rect 467742 48764 467748 48776
rect 467800 48764 467806 48816
rect 472434 48764 472440 48816
rect 472492 48804 472498 48816
rect 473262 48804 473268 48816
rect 472492 48776 473268 48804
rect 472492 48764 472498 48776
rect 473262 48764 473268 48776
rect 473320 48764 473326 48816
rect 473630 48764 473636 48816
rect 473688 48804 473694 48816
rect 474642 48804 474648 48816
rect 473688 48776 474648 48804
rect 473688 48764 473694 48776
rect 474642 48764 474648 48776
rect 474700 48764 474706 48816
rect 480806 48764 480812 48816
rect 480864 48804 480870 48816
rect 481542 48804 481548 48816
rect 480864 48776 481548 48804
rect 480864 48764 480870 48776
rect 481542 48764 481548 48776
rect 481600 48764 481606 48816
rect 483198 48764 483204 48816
rect 483256 48804 483262 48816
rect 484302 48804 484308 48816
rect 483256 48776 484308 48804
rect 483256 48764 483262 48776
rect 484302 48764 484308 48776
rect 484360 48764 484366 48816
rect 484394 48764 484400 48816
rect 484452 48804 484458 48816
rect 485590 48804 485596 48816
rect 484452 48776 485596 48804
rect 484452 48764 484458 48776
rect 485590 48764 485596 48776
rect 485648 48764 485654 48816
rect 490374 48764 490380 48816
rect 490432 48804 490438 48816
rect 491202 48804 491208 48816
rect 490432 48776 491208 48804
rect 490432 48764 490438 48776
rect 491202 48764 491208 48776
rect 491260 48764 491266 48816
rect 491570 48764 491576 48816
rect 491628 48804 491634 48816
rect 492582 48804 492588 48816
rect 491628 48776 492588 48804
rect 491628 48764 491634 48776
rect 492582 48764 492588 48776
rect 492640 48764 492646 48816
rect 492766 48764 492772 48816
rect 492824 48804 492830 48816
rect 493962 48804 493968 48816
rect 492824 48776 493968 48804
rect 492824 48764 492830 48776
rect 493962 48764 493968 48776
rect 494020 48764 494026 48816
rect 498654 48764 498660 48816
rect 498712 48804 498718 48816
rect 499482 48804 499488 48816
rect 498712 48776 499488 48804
rect 498712 48764 498718 48776
rect 499482 48764 499488 48776
rect 499540 48764 499546 48816
rect 499850 48764 499856 48816
rect 499908 48804 499914 48816
rect 500862 48804 500868 48816
rect 499908 48776 500868 48804
rect 499908 48764 499914 48776
rect 500862 48764 500868 48776
rect 500920 48764 500926 48816
rect 508222 48764 508228 48816
rect 508280 48804 508286 48816
rect 509142 48804 509148 48816
rect 508280 48776 509148 48804
rect 508280 48764 508286 48776
rect 509142 48764 509148 48776
rect 509200 48764 509206 48816
rect 509418 48764 509424 48816
rect 509476 48804 509482 48816
rect 510522 48804 510528 48816
rect 509476 48776 510528 48804
rect 509476 48764 509482 48776
rect 510522 48764 510528 48776
rect 510580 48764 510586 48816
rect 516594 48764 516600 48816
rect 516652 48804 516658 48816
rect 517422 48804 517428 48816
rect 516652 48776 517428 48804
rect 516652 48764 516658 48776
rect 517422 48764 517428 48776
rect 517480 48764 517486 48816
rect 517790 48764 517796 48816
rect 517848 48804 517854 48816
rect 518802 48804 518808 48816
rect 517848 48776 518808 48804
rect 517848 48764 517854 48776
rect 518802 48764 518808 48776
rect 518860 48764 518866 48816
rect 518986 48764 518992 48816
rect 519044 48804 519050 48816
rect 520090 48804 520096 48816
rect 519044 48776 520096 48804
rect 519044 48764 519050 48776
rect 520090 48764 520096 48776
rect 520148 48764 520154 48816
rect 64874 48696 64880 48748
rect 64932 48736 64938 48748
rect 66162 48736 66168 48748
rect 64932 48708 66168 48736
rect 64932 48696 64938 48708
rect 66162 48696 66168 48708
rect 66220 48696 66226 48748
rect 123294 48696 123300 48748
rect 123352 48736 123358 48748
rect 124122 48736 124128 48748
rect 123352 48708 124128 48736
rect 123352 48696 123358 48708
rect 124122 48696 124128 48708
rect 124180 48696 124186 48748
rect 157886 48696 157892 48748
rect 157944 48736 157950 48748
rect 158622 48736 158628 48748
rect 157944 48708 158628 48736
rect 157944 48696 157950 48708
rect 158622 48696 158628 48708
rect 158680 48696 158686 48748
rect 271046 48696 271052 48748
rect 271104 48736 271110 48748
rect 272518 48736 272524 48748
rect 271104 48708 272524 48736
rect 271104 48696 271110 48708
rect 272518 48696 272524 48708
rect 272576 48696 272582 48748
rect 315206 48696 315212 48748
rect 315264 48736 315270 48748
rect 315942 48736 315948 48748
rect 315264 48708 315948 48736
rect 315264 48696 315270 48708
rect 315942 48696 315948 48708
rect 316000 48696 316006 48748
rect 385494 48696 385500 48748
rect 385552 48736 385558 48748
rect 386322 48736 386328 48748
rect 385552 48708 386328 48736
rect 385552 48696 385558 48708
rect 386322 48696 386328 48708
rect 386380 48696 386386 48748
rect 125686 48628 125692 48680
rect 125744 48668 125750 48680
rect 126882 48668 126888 48680
rect 125744 48640 126888 48668
rect 125744 48628 125750 48640
rect 126882 48628 126888 48640
rect 126940 48628 126946 48680
rect 186498 48628 186504 48680
rect 186556 48668 186562 48680
rect 187602 48668 187608 48680
rect 186556 48640 187608 48668
rect 186556 48628 186562 48640
rect 187602 48628 187608 48640
rect 187660 48628 187666 48680
rect 230566 48628 230572 48680
rect 230624 48668 230630 48680
rect 231670 48668 231676 48680
rect 230624 48640 231676 48668
rect 230624 48628 230630 48640
rect 231670 48628 231676 48640
rect 231728 48628 231734 48680
rect 308030 48560 308036 48612
rect 308088 48600 308094 48612
rect 309042 48600 309048 48612
rect 308088 48572 309048 48600
rect 308088 48560 308094 48572
rect 309042 48560 309048 48572
rect 309100 48560 309106 48612
rect 368842 48560 368848 48612
rect 368900 48600 368906 48612
rect 369762 48600 369768 48612
rect 368900 48572 369768 48600
rect 368900 48560 368906 48572
rect 369762 48560 369768 48572
rect 369820 48560 369826 48612
rect 375926 48560 375932 48612
rect 375984 48600 375990 48612
rect 376662 48600 376668 48612
rect 375984 48572 376668 48600
rect 375984 48560 375990 48572
rect 376662 48560 376668 48572
rect 376720 48560 376726 48612
rect 195974 48492 195980 48544
rect 196032 48532 196038 48544
rect 197262 48532 197268 48544
rect 196032 48504 197268 48532
rect 196032 48492 196038 48504
rect 197262 48492 197268 48504
rect 197320 48492 197326 48544
rect 405734 48492 405740 48544
rect 405792 48532 405798 48544
rect 406930 48532 406936 48544
rect 405792 48504 406936 48532
rect 405792 48492 405798 48504
rect 406930 48492 406936 48504
rect 406988 48492 406994 48544
rect 510614 48492 510620 48544
rect 510672 48532 510678 48544
rect 511902 48532 511908 48544
rect 510672 48504 511908 48532
rect 510672 48492 510678 48504
rect 511902 48492 511908 48504
rect 511960 48492 511966 48544
rect 82814 48424 82820 48476
rect 82872 48464 82878 48476
rect 84010 48464 84016 48476
rect 82872 48436 84016 48464
rect 82872 48424 82878 48436
rect 84010 48424 84016 48436
rect 84068 48424 84074 48476
rect 176930 48424 176936 48476
rect 176988 48464 176994 48476
rect 177942 48464 177948 48476
rect 176988 48436 177948 48464
rect 176988 48424 176994 48436
rect 177942 48424 177948 48436
rect 178000 48424 178006 48476
rect 290182 48424 290188 48476
rect 290240 48464 290246 48476
rect 291102 48464 291108 48476
rect 290240 48436 291108 48464
rect 290240 48424 290246 48436
rect 291102 48424 291108 48436
rect 291160 48424 291166 48476
rect 298462 48424 298468 48476
rect 298520 48464 298526 48476
rect 299382 48464 299388 48476
rect 298520 48436 299388 48464
rect 298520 48424 298526 48436
rect 299382 48424 299388 48436
rect 299440 48424 299446 48476
rect 317598 48288 317604 48340
rect 317656 48328 317662 48340
rect 318702 48328 318708 48340
rect 317656 48300 318708 48328
rect 317656 48288 317662 48300
rect 318702 48288 318708 48300
rect 318760 48288 318766 48340
rect 422386 48288 422392 48340
rect 422444 48328 422450 48340
rect 423582 48328 423588 48340
rect 422444 48300 423588 48328
rect 422444 48288 422450 48300
rect 423582 48288 423588 48300
rect 423640 48288 423646 48340
rect 151906 47608 151912 47660
rect 151964 47648 151970 47660
rect 212534 47648 212540 47660
rect 151964 47620 212540 47648
rect 151964 47608 151970 47620
rect 212534 47608 212540 47620
rect 212592 47608 212598 47660
rect 262766 47608 262772 47660
rect 262824 47648 262830 47660
rect 322934 47648 322940 47660
rect 262824 47620 322940 47648
rect 262824 47608 262830 47620
rect 322934 47608 322940 47620
rect 322992 47608 322998 47660
rect 84102 47540 84108 47592
rect 84160 47580 84166 47592
rect 144914 47580 144920 47592
rect 84160 47552 144920 47580
rect 84160 47540 84166 47552
rect 144914 47540 144920 47552
rect 144972 47540 144978 47592
rect 205542 47540 205548 47592
rect 205600 47580 205606 47592
rect 266354 47580 266360 47592
rect 205600 47552 266360 47580
rect 205600 47540 205606 47552
rect 266354 47540 266360 47552
rect 266412 47540 266418 47592
rect 316402 47540 316408 47592
rect 316460 47580 316466 47592
rect 376754 47580 376760 47592
rect 316460 47552 376760 47580
rect 316460 47540 316466 47552
rect 376754 47540 376760 47552
rect 376812 47540 376818 47592
rect 433242 47540 433248 47592
rect 433300 47580 433306 47592
rect 494054 47580 494060 47592
rect 433300 47552 494060 47580
rect 433300 47540 433306 47552
rect 494054 47540 494060 47552
rect 494112 47540 494118 47592
rect 501046 47540 501052 47592
rect 501104 47580 501110 47592
rect 561674 47580 561680 47592
rect 501104 47552 561680 47580
rect 501104 47540 501110 47552
rect 561674 47540 561680 47552
rect 561732 47540 561738 47592
rect 407206 46900 407212 46912
rect 407167 46872 407212 46900
rect 407206 46860 407212 46872
rect 407264 46860 407270 46912
rect 443178 46900 443184 46912
rect 443139 46872 443184 46900
rect 443178 46860 443184 46872
rect 443236 46860 443242 46912
rect 449986 46900 449992 46912
rect 449947 46872 449992 46900
rect 449986 46860 449992 46872
rect 450044 46860 450050 46912
rect 535454 46900 535460 46912
rect 535415 46872 535460 46900
rect 535454 46860 535460 46872
rect 535512 46860 535518 46912
rect 201954 46248 201960 46300
rect 202012 46288 202018 46300
rect 262214 46288 262220 46300
rect 202012 46260 262220 46288
rect 202012 46248 202018 46260
rect 262214 46248 262220 46260
rect 262272 46248 262278 46300
rect 312814 46248 312820 46300
rect 312872 46288 312878 46300
rect 374086 46288 374092 46300
rect 312872 46260 374092 46288
rect 312872 46248 312878 46260
rect 374086 46248 374092 46260
rect 374144 46248 374150 46300
rect 80422 46180 80428 46232
rect 80480 46220 80486 46232
rect 140774 46220 140780 46232
rect 80480 46192 140780 46220
rect 80480 46180 80486 46192
rect 140774 46180 140780 46192
rect 140832 46180 140838 46232
rect 148318 46180 148324 46232
rect 148376 46220 148382 46232
rect 209866 46220 209872 46232
rect 148376 46192 209872 46220
rect 148376 46180 148382 46192
rect 209866 46180 209872 46192
rect 209924 46180 209930 46232
rect 259178 46180 259184 46232
rect 259236 46220 259242 46232
rect 320174 46220 320180 46232
rect 259236 46192 320180 46220
rect 259236 46180 259242 46192
rect 320174 46180 320180 46192
rect 320232 46180 320238 46232
rect 369946 46180 369952 46232
rect 370004 46220 370010 46232
rect 430574 46220 430580 46232
rect 370004 46192 430580 46220
rect 370004 46180 370010 46192
rect 430574 46180 430580 46192
rect 430632 46180 430638 46232
rect 450998 46180 451004 46232
rect 451056 46220 451062 46232
rect 511994 46220 512000 46232
rect 451056 46192 512000 46220
rect 451056 46180 451062 46192
rect 511994 46180 512000 46192
rect 512052 46180 512058 46232
rect 515398 46180 515404 46232
rect 515456 46220 515462 46232
rect 575474 46220 575480 46232
rect 515456 46192 575480 46220
rect 515456 46180 515462 46192
rect 575474 46180 575480 46192
rect 575532 46180 575538 46232
rect 256602 44956 256608 45008
rect 256660 44996 256666 45008
rect 316034 44996 316040 45008
rect 256660 44968 316040 44996
rect 256660 44956 256666 44968
rect 316034 44956 316040 44968
rect 316092 44956 316098 45008
rect 198642 44888 198648 44940
rect 198700 44928 198706 44940
rect 259454 44928 259460 44940
rect 198700 44900 259460 44928
rect 198700 44888 198706 44900
rect 259454 44888 259460 44900
rect 259512 44888 259518 44940
rect 77202 44820 77208 44872
rect 77260 44860 77266 44872
rect 138014 44860 138020 44872
rect 77260 44832 138020 44860
rect 77260 44820 77266 44832
rect 138014 44820 138020 44832
rect 138072 44820 138078 44872
rect 144730 44820 144736 44872
rect 144788 44860 144794 44872
rect 205634 44860 205640 44872
rect 144788 44832 205640 44860
rect 144788 44820 144794 44832
rect 205634 44820 205640 44832
rect 205692 44820 205698 44872
rect 310330 44820 310336 44872
rect 310388 44860 310394 44872
rect 369854 44860 369860 44872
rect 310388 44832 369860 44860
rect 310388 44820 310394 44832
rect 369854 44820 369860 44832
rect 369912 44820 369918 44872
rect 415210 44820 415216 44872
rect 415268 44860 415274 44872
rect 476114 44860 476120 44872
rect 415268 44832 476120 44860
rect 415268 44820 415274 44832
rect 476114 44820 476120 44832
rect 476172 44820 476178 44872
rect 493870 44820 493876 44872
rect 493928 44860 493934 44872
rect 554774 44860 554780 44872
rect 493928 44832 554780 44860
rect 493928 44820 493934 44832
rect 554774 44820 554780 44832
rect 554832 44820 554838 44872
rect 195882 43460 195888 43512
rect 195940 43500 195946 43512
rect 255314 43500 255320 43512
rect 195940 43472 255320 43500
rect 195940 43460 195946 43472
rect 255314 43460 255320 43472
rect 255372 43460 255378 43512
rect 302050 43460 302056 43512
rect 302108 43500 302114 43512
rect 362954 43500 362960 43512
rect 302108 43472 362960 43500
rect 302108 43460 302114 43472
rect 362954 43460 362960 43472
rect 363012 43460 363018 43512
rect 409782 43460 409788 43512
rect 409840 43500 409846 43512
rect 469214 43500 469220 43512
rect 409840 43472 469220 43500
rect 409840 43460 409846 43472
rect 469214 43460 469220 43472
rect 469272 43460 469278 43512
rect 74350 43392 74356 43444
rect 74408 43432 74414 43444
rect 133874 43432 133880 43444
rect 74408 43404 133880 43432
rect 74408 43392 74414 43404
rect 133874 43392 133880 43404
rect 133932 43392 133938 43444
rect 142062 43392 142068 43444
rect 142120 43432 142126 43444
rect 201494 43432 201500 43444
rect 142120 43404 201500 43432
rect 142120 43392 142126 43404
rect 201494 43392 201500 43404
rect 201552 43392 201558 43444
rect 249610 43392 249616 43444
rect 249668 43432 249674 43444
rect 309134 43432 309140 43444
rect 249668 43404 309140 43432
rect 249668 43392 249674 43404
rect 309134 43392 309140 43404
rect 309192 43392 309198 43444
rect 362770 43392 362776 43444
rect 362828 43432 362834 43444
rect 423674 43432 423680 43444
rect 362828 43404 423680 43432
rect 362828 43392 362834 43404
rect 423674 43392 423680 43404
rect 423732 43392 423738 43444
rect 511810 43392 511816 43444
rect 511868 43432 511874 43444
rect 571426 43432 571432 43444
rect 511868 43404 571432 43432
rect 511868 43392 511874 43404
rect 571426 43392 571432 43404
rect 571484 43392 571490 43444
rect 135162 42100 135168 42152
rect 135220 42140 135226 42152
rect 194594 42140 194600 42152
rect 135220 42112 194600 42140
rect 135220 42100 135226 42112
rect 194594 42100 194600 42112
rect 194652 42100 194658 42152
rect 245562 42100 245568 42152
rect 245620 42140 245626 42152
rect 304994 42140 305000 42152
rect 245620 42112 305000 42140
rect 245620 42100 245626 42112
rect 304994 42100 305000 42112
rect 305052 42100 305058 42152
rect 360102 42100 360108 42152
rect 360160 42140 360166 42152
rect 419534 42140 419540 42152
rect 360160 42112 419540 42140
rect 360160 42100 360166 42112
rect 419534 42100 419540 42112
rect 419592 42100 419598 42152
rect 70302 42032 70308 42084
rect 70360 42072 70366 42084
rect 131114 42072 131120 42084
rect 70360 42044 131120 42072
rect 70360 42032 70366 42044
rect 131114 42032 131120 42044
rect 131172 42032 131178 42084
rect 191742 42032 191748 42084
rect 191800 42072 191806 42084
rect 252646 42072 252652 42084
rect 191800 42044 252652 42072
rect 191800 42032 191806 42044
rect 252646 42032 252652 42044
rect 252704 42032 252710 42084
rect 299382 42032 299388 42084
rect 299440 42072 299446 42084
rect 358814 42072 358820 42084
rect 299440 42044 358820 42072
rect 299440 42032 299446 42044
rect 358814 42032 358820 42044
rect 358872 42032 358878 42084
rect 406930 42032 406936 42084
rect 406988 42072 406994 42084
rect 466454 42072 466460 42084
rect 406988 42044 466460 42072
rect 406988 42032 406994 42044
rect 466454 42032 466460 42044
rect 466512 42032 466518 42084
rect 520090 42032 520096 42084
rect 520148 42072 520154 42084
rect 579614 42072 579620 42084
rect 520148 42044 579620 42072
rect 520148 42032 520154 42044
rect 579614 42032 579620 42044
rect 579672 42032 579678 42084
rect 523678 41352 523684 41404
rect 523736 41392 523742 41404
rect 580166 41392 580172 41404
rect 523736 41364 580172 41392
rect 523736 41352 523742 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 188982 40740 188988 40792
rect 189040 40780 189046 40792
rect 248414 40780 248420 40792
rect 189040 40752 248420 40780
rect 189040 40740 189046 40752
rect 248414 40740 248420 40752
rect 248472 40740 248478 40792
rect 292482 40740 292488 40792
rect 292540 40780 292546 40792
rect 351914 40780 351920 40792
rect 292540 40752 351920 40780
rect 292540 40740 292546 40752
rect 351914 40740 351920 40752
rect 351972 40740 351978 40792
rect 402882 40740 402888 40792
rect 402940 40780 402946 40792
rect 462314 40780 462320 40792
rect 402940 40752 462320 40780
rect 402940 40740 402946 40752
rect 462314 40740 462320 40752
rect 462372 40740 462378 40792
rect 131022 40672 131028 40724
rect 131080 40712 131086 40724
rect 191834 40712 191840 40724
rect 131080 40684 191840 40712
rect 131080 40672 131086 40684
rect 191834 40672 191840 40684
rect 191892 40672 191898 40724
rect 241330 40672 241336 40724
rect 241388 40712 241394 40724
rect 302234 40712 302240 40724
rect 241388 40684 302240 40712
rect 241388 40672 241394 40684
rect 302234 40672 302240 40684
rect 302292 40672 302298 40724
rect 349062 40672 349068 40724
rect 349120 40712 349126 40724
rect 408494 40712 408500 40724
rect 349120 40684 408500 40712
rect 349120 40672 349126 40684
rect 408494 40672 408500 40684
rect 408552 40672 408558 40724
rect 424962 40672 424968 40724
rect 425020 40712 425026 40724
rect 485774 40712 485780 40724
rect 425020 40684 485780 40712
rect 425020 40672 425026 40684
rect 485774 40672 485780 40684
rect 485832 40672 485838 40724
rect 288342 39448 288348 39500
rect 288400 39488 288406 39500
rect 347774 39488 347780 39500
rect 288400 39460 347780 39488
rect 288400 39448 288406 39460
rect 347774 39448 347780 39460
rect 347832 39448 347838 39500
rect 184842 39380 184848 39432
rect 184900 39420 184906 39432
rect 244274 39420 244280 39432
rect 184900 39392 244280 39420
rect 184900 39380 184906 39392
rect 244274 39380 244280 39392
rect 244332 39380 244338 39432
rect 342162 39380 342168 39432
rect 342220 39420 342226 39432
rect 401594 39420 401600 39432
rect 342220 39392 401600 39420
rect 342220 39380 342226 39392
rect 401594 39380 401600 39392
rect 401652 39380 401658 39432
rect 126790 39312 126796 39364
rect 126848 39352 126854 39364
rect 187694 39352 187700 39364
rect 126848 39324 187700 39352
rect 126848 39312 126854 39324
rect 187694 39312 187700 39324
rect 187752 39312 187758 39364
rect 238662 39312 238668 39364
rect 238720 39352 238726 39364
rect 298094 39352 298100 39364
rect 238720 39324 298100 39352
rect 238720 39312 238726 39324
rect 298094 39312 298100 39324
rect 298152 39312 298158 39364
rect 398742 39312 398748 39364
rect 398800 39352 398806 39364
rect 459646 39352 459652 39364
rect 398800 39324 459652 39352
rect 398800 39312 398806 39324
rect 459646 39312 459652 39324
rect 459704 39312 459710 39364
rect 477402 39312 477408 39364
rect 477460 39352 477466 39364
rect 536834 39352 536840 39364
rect 477460 39324 536840 39352
rect 477460 39312 477466 39324
rect 536834 39312 536840 39324
rect 536892 39312 536898 39364
rect 369854 38564 369860 38616
rect 369912 38604 369918 38616
rect 369946 38604 369952 38616
rect 369912 38576 369952 38604
rect 369912 38564 369918 38576
rect 369946 38564 369952 38576
rect 370004 38564 370010 38616
rect 124122 37952 124128 38004
rect 124180 37992 124186 38004
rect 183554 37992 183560 38004
rect 124180 37964 183560 37992
rect 124180 37952 124186 37964
rect 183554 37952 183560 37964
rect 183612 37952 183618 38004
rect 234522 37952 234528 38004
rect 234580 37992 234586 38004
rect 295334 37992 295340 38004
rect 234580 37964 295340 37992
rect 234580 37952 234586 37964
rect 295334 37952 295340 37964
rect 295392 37952 295398 38004
rect 338022 37952 338028 38004
rect 338080 37992 338086 38004
rect 398837 37995 398895 38001
rect 398837 37992 398849 37995
rect 338080 37964 398849 37992
rect 338080 37952 338086 37964
rect 398837 37961 398849 37964
rect 398883 37961 398895 37995
rect 398837 37955 398895 37961
rect 420822 37952 420828 38004
rect 420880 37992 420886 38004
rect 480254 37992 480260 38004
rect 420880 37964 480260 37992
rect 420880 37952 420886 37964
rect 480254 37952 480260 37964
rect 480312 37952 480318 38004
rect 180702 37884 180708 37936
rect 180760 37924 180766 37936
rect 241514 37924 241520 37936
rect 180760 37896 241520 37924
rect 180760 37884 180766 37896
rect 241514 37884 241520 37896
rect 241572 37884 241578 37936
rect 284110 37884 284116 37936
rect 284168 37924 284174 37936
rect 345014 37924 345020 37936
rect 284168 37896 345020 37924
rect 284168 37884 284174 37896
rect 345014 37884 345020 37896
rect 345072 37884 345078 37936
rect 395982 37884 395988 37936
rect 396040 37924 396046 37936
rect 455414 37924 455420 37936
rect 396040 37896 455420 37924
rect 396040 37884 396046 37896
rect 455414 37884 455420 37896
rect 455472 37884 455478 37936
rect 485590 37884 485596 37936
rect 485648 37924 485654 37936
rect 545114 37924 545120 37936
rect 485648 37896 545120 37924
rect 485648 37884 485654 37896
rect 545114 37884 545120 37896
rect 545172 37884 545178 37936
rect 398834 37312 398840 37324
rect 398795 37284 398840 37312
rect 398834 37272 398840 37284
rect 398892 37272 398898 37324
rect 407206 37312 407212 37324
rect 407167 37284 407212 37312
rect 407206 37272 407212 37284
rect 407264 37272 407270 37324
rect 443178 37312 443184 37324
rect 443139 37284 443184 37312
rect 443178 37272 443184 37284
rect 443236 37272 443242 37324
rect 449986 37312 449992 37324
rect 449947 37284 449992 37312
rect 449986 37272 449992 37284
rect 450044 37272 450050 37324
rect 535454 37312 535460 37324
rect 535415 37284 535460 37312
rect 535454 37272 535460 37284
rect 535512 37272 535518 37324
rect 177942 36592 177948 36644
rect 178000 36632 178006 36644
rect 237374 36632 237380 36644
rect 178000 36604 237380 36632
rect 178000 36592 178006 36604
rect 237374 36592 237380 36604
rect 237432 36592 237438 36644
rect 281442 36592 281448 36644
rect 281500 36632 281506 36644
rect 340874 36632 340880 36644
rect 281500 36604 340880 36632
rect 281500 36592 281506 36604
rect 340874 36592 340880 36604
rect 340932 36592 340938 36644
rect 391842 36592 391848 36644
rect 391900 36632 391906 36644
rect 451274 36632 451280 36644
rect 391900 36604 451280 36632
rect 391900 36592 391906 36604
rect 451274 36592 451280 36604
rect 451332 36592 451338 36644
rect 119982 36524 119988 36576
rect 120040 36564 120046 36576
rect 180794 36564 180800 36576
rect 120040 36536 180800 36564
rect 120040 36524 120046 36536
rect 180794 36524 180800 36536
rect 180852 36524 180858 36576
rect 231670 36524 231676 36576
rect 231728 36564 231734 36576
rect 291194 36564 291200 36576
rect 231728 36536 291200 36564
rect 231728 36524 231734 36536
rect 291194 36524 291200 36536
rect 291252 36524 291258 36576
rect 335262 36524 335268 36576
rect 335320 36564 335326 36576
rect 394694 36564 394700 36576
rect 335320 36536 394700 36564
rect 335320 36524 335326 36536
rect 394694 36524 394700 36536
rect 394752 36524 394758 36576
rect 459370 36524 459376 36576
rect 459428 36564 459434 36576
rect 520366 36564 520372 36576
rect 459428 36536 520372 36564
rect 459428 36524 459434 36536
rect 520366 36524 520372 36536
rect 520424 36524 520430 36576
rect 3326 35844 3332 35896
rect 3384 35884 3390 35896
rect 59998 35884 60004 35896
rect 3384 35856 60004 35884
rect 3384 35844 3390 35856
rect 59998 35844 60004 35856
rect 60056 35844 60062 35896
rect 117222 35232 117228 35284
rect 117280 35272 117286 35284
rect 176654 35272 176660 35284
rect 117280 35244 176660 35272
rect 117280 35232 117286 35244
rect 176654 35232 176660 35244
rect 176712 35232 176718 35284
rect 227622 35232 227628 35284
rect 227680 35272 227686 35284
rect 287054 35272 287060 35284
rect 227680 35244 287060 35272
rect 227680 35232 227686 35244
rect 287054 35232 287060 35244
rect 287112 35232 287118 35284
rect 331122 35232 331128 35284
rect 331180 35272 331186 35284
rect 390554 35272 390560 35284
rect 331180 35244 390560 35272
rect 331180 35232 331186 35244
rect 390554 35232 390560 35244
rect 390612 35232 390618 35284
rect 170950 35164 170956 35216
rect 171008 35204 171014 35216
rect 230474 35204 230480 35216
rect 171008 35176 230480 35204
rect 171008 35164 171014 35176
rect 230474 35164 230480 35176
rect 230532 35164 230538 35216
rect 277302 35164 277308 35216
rect 277360 35204 277366 35216
rect 338114 35204 338120 35216
rect 277360 35176 338120 35204
rect 277360 35164 277366 35176
rect 338114 35164 338120 35176
rect 338172 35164 338178 35216
rect 389082 35164 389088 35216
rect 389140 35204 389146 35216
rect 448514 35204 448520 35216
rect 389140 35176 448520 35204
rect 389140 35164 389146 35176
rect 448514 35164 448520 35176
rect 448572 35164 448578 35216
rect 456702 35164 456708 35216
rect 456760 35204 456766 35216
rect 516137 35207 516195 35213
rect 516137 35204 516149 35207
rect 456760 35176 516149 35204
rect 456760 35164 456766 35176
rect 516137 35173 516149 35176
rect 516183 35173 516195 35207
rect 516137 35167 516195 35173
rect 274542 33872 274548 33924
rect 274600 33912 274606 33924
rect 333974 33912 333980 33924
rect 274600 33884 333980 33912
rect 274600 33872 274606 33884
rect 333974 33872 333980 33884
rect 334032 33872 334038 33924
rect 113082 33804 113088 33856
rect 113140 33844 113146 33856
rect 173894 33844 173900 33856
rect 113140 33816 173900 33844
rect 113140 33804 113146 33816
rect 173894 33804 173900 33816
rect 173952 33804 173958 33856
rect 223390 33804 223396 33856
rect 223448 33844 223454 33856
rect 284294 33844 284300 33856
rect 223448 33816 284300 33844
rect 223448 33804 223454 33816
rect 284294 33804 284300 33816
rect 284352 33804 284358 33856
rect 166902 33736 166908 33788
rect 166960 33776 166966 33788
rect 227806 33776 227812 33788
rect 166960 33748 227812 33776
rect 166960 33736 166966 33748
rect 227806 33736 227812 33748
rect 227864 33736 227870 33788
rect 328270 33736 328276 33788
rect 328328 33776 328334 33788
rect 387794 33776 387800 33788
rect 328328 33748 387800 33776
rect 328328 33736 328334 33748
rect 387794 33736 387800 33748
rect 387852 33736 387858 33788
rect 441430 33736 441436 33788
rect 441488 33776 441494 33788
rect 502426 33776 502432 33788
rect 441488 33748 502432 33776
rect 441488 33736 441494 33748
rect 502426 33736 502432 33748
rect 502484 33736 502490 33788
rect 110322 32444 110328 32496
rect 110380 32484 110386 32496
rect 169754 32484 169760 32496
rect 110380 32456 169760 32484
rect 110380 32444 110386 32456
rect 169754 32444 169760 32456
rect 169812 32444 169818 32496
rect 220722 32444 220728 32496
rect 220780 32484 220786 32496
rect 280154 32484 280160 32496
rect 220780 32456 280160 32484
rect 220780 32444 220786 32456
rect 280154 32444 280160 32456
rect 280212 32444 280218 32496
rect 324222 32444 324228 32496
rect 324280 32484 324286 32496
rect 383654 32484 383660 32496
rect 324280 32456 383660 32484
rect 324280 32444 324286 32456
rect 383654 32444 383660 32456
rect 383712 32444 383718 32496
rect 162670 32376 162676 32428
rect 162728 32416 162734 32428
rect 223574 32416 223580 32428
rect 162728 32388 223580 32416
rect 162728 32376 162734 32388
rect 223574 32376 223580 32388
rect 223632 32376 223638 32428
rect 270402 32376 270408 32428
rect 270460 32416 270466 32428
rect 331214 32416 331220 32428
rect 270460 32388 331220 32416
rect 270460 32376 270466 32388
rect 331214 32376 331220 32388
rect 331272 32376 331278 32428
rect 384942 32376 384948 32428
rect 385000 32416 385006 32428
rect 444374 32416 444380 32428
rect 385000 32388 444380 32416
rect 385000 32376 385006 32388
rect 444374 32376 444380 32388
rect 444432 32376 444438 32428
rect 449710 32376 449716 32428
rect 449768 32416 449774 32428
rect 509234 32416 509240 32428
rect 449768 32388 509240 32416
rect 449768 32376 449774 32388
rect 509234 32376 509240 32388
rect 509292 32376 509298 32428
rect 510522 32376 510528 32428
rect 510580 32416 510586 32428
rect 569954 32416 569960 32428
rect 510580 32388 569960 32416
rect 510580 32376 510586 32388
rect 569954 32376 569960 32388
rect 570012 32376 570018 32428
rect 160002 31084 160008 31136
rect 160060 31124 160066 31136
rect 219434 31124 219440 31136
rect 160060 31096 219440 31124
rect 160060 31084 160066 31096
rect 219434 31084 219440 31096
rect 219492 31084 219498 31136
rect 267642 31084 267648 31136
rect 267700 31124 267706 31136
rect 327074 31124 327080 31136
rect 267700 31096 327080 31124
rect 267700 31084 267706 31096
rect 327074 31084 327080 31096
rect 327132 31084 327138 31136
rect 378042 31084 378048 31136
rect 378100 31124 378106 31136
rect 437474 31124 437480 31136
rect 378100 31096 437480 31124
rect 378100 31084 378106 31096
rect 437474 31084 437480 31096
rect 437532 31084 437538 31136
rect 106182 31016 106188 31068
rect 106240 31056 106246 31068
rect 167086 31056 167092 31068
rect 106240 31028 167092 31056
rect 106240 31016 106246 31028
rect 167086 31016 167092 31028
rect 167144 31016 167150 31068
rect 216582 31016 216588 31068
rect 216640 31056 216646 31068
rect 277394 31056 277400 31068
rect 216640 31028 277400 31056
rect 216640 31016 216646 31028
rect 277394 31016 277400 31028
rect 277452 31016 277458 31068
rect 320082 31016 320088 31068
rect 320140 31056 320146 31068
rect 380894 31056 380900 31068
rect 320140 31028 380900 31056
rect 320140 31016 320146 31028
rect 380894 31016 380900 31028
rect 380952 31016 380958 31068
rect 445662 31016 445668 31068
rect 445720 31056 445726 31068
rect 505094 31056 505100 31068
rect 445720 31028 505100 31056
rect 445720 31016 445726 31028
rect 505094 31016 505100 31028
rect 505152 31016 505158 31068
rect 506382 31016 506388 31068
rect 506440 31056 506446 31068
rect 565814 31056 565820 31068
rect 506440 31028 565820 31056
rect 506440 31016 506446 31028
rect 565814 31016 565820 31028
rect 565872 31016 565878 31068
rect 523770 30268 523776 30320
rect 523828 30308 523834 30320
rect 580166 30308 580172 30320
rect 523828 30280 580172 30308
rect 523828 30268 523834 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 213822 29724 213828 29776
rect 213880 29764 213886 29776
rect 273254 29764 273260 29776
rect 213880 29736 273260 29764
rect 213880 29724 213886 29736
rect 273254 29724 273260 29736
rect 273312 29724 273318 29776
rect 155862 29656 155868 29708
rect 155920 29696 155926 29708
rect 216674 29696 216680 29708
rect 155920 29668 216680 29696
rect 155920 29656 155926 29668
rect 216674 29656 216680 29668
rect 216732 29656 216738 29708
rect 306282 29656 306288 29708
rect 306340 29696 306346 29708
rect 365714 29696 365720 29708
rect 306340 29668 365720 29696
rect 306340 29656 306346 29668
rect 365714 29656 365720 29668
rect 365772 29656 365778 29708
rect 102042 29588 102048 29640
rect 102100 29628 102106 29640
rect 162854 29628 162860 29640
rect 102100 29600 162860 29628
rect 102100 29588 102106 29600
rect 162854 29588 162860 29600
rect 162912 29588 162918 29640
rect 252462 29588 252468 29640
rect 252520 29628 252526 29640
rect 313366 29628 313372 29640
rect 252520 29600 313372 29628
rect 252520 29588 252526 29600
rect 313366 29588 313372 29600
rect 313424 29588 313430 29640
rect 367002 29588 367008 29640
rect 367060 29628 367066 29640
rect 426434 29628 426440 29640
rect 367060 29600 426440 29628
rect 367060 29588 367066 29600
rect 426434 29588 426440 29600
rect 426492 29588 426498 29640
rect 438762 29588 438768 29640
rect 438820 29628 438826 29640
rect 498194 29628 498200 29640
rect 438820 29600 498200 29628
rect 438820 29588 438826 29600
rect 498194 29588 498200 29600
rect 498252 29588 498258 29640
rect 407206 29112 407212 29164
rect 407264 29112 407270 29164
rect 407224 29028 407252 29112
rect 407206 28976 407212 29028
rect 407264 28976 407270 29028
rect 516134 29016 516140 29028
rect 516095 28988 516140 29016
rect 516134 28976 516140 28988
rect 516192 28976 516198 29028
rect 272518 28296 272524 28348
rect 272576 28336 272582 28348
rect 331306 28336 331312 28348
rect 272576 28308 331312 28336
rect 272576 28296 272582 28308
rect 331306 28296 331312 28308
rect 331364 28296 331370 28348
rect 97902 28228 97908 28280
rect 97960 28268 97966 28280
rect 158806 28268 158812 28280
rect 97960 28240 158812 28268
rect 97960 28228 97966 28240
rect 158806 28228 158812 28240
rect 158864 28228 158870 28280
rect 165522 28228 165528 28280
rect 165580 28268 165586 28280
rect 226334 28268 226340 28280
rect 165580 28240 226340 28268
rect 165580 28228 165586 28240
rect 226334 28228 226340 28240
rect 226392 28228 226398 28280
rect 244182 28228 244188 28280
rect 244240 28268 244246 28280
rect 305086 28268 305092 28280
rect 244240 28240 305092 28268
rect 244240 28228 244246 28240
rect 305086 28228 305092 28240
rect 305144 28228 305150 28280
rect 322842 28228 322848 28280
rect 322900 28268 322906 28280
rect 382366 28268 382372 28280
rect 322900 28240 382372 28268
rect 322900 28228 322906 28240
rect 382366 28228 382372 28240
rect 382424 28228 382430 28280
rect 434622 28228 434628 28280
rect 434680 28268 434686 28280
rect 494146 28268 494152 28280
rect 434680 28240 494152 28268
rect 434680 28228 434686 28240
rect 494146 28228 494152 28240
rect 494204 28228 494210 28280
rect 495342 28228 495348 28280
rect 495400 28268 495406 28280
rect 554866 28268 554872 28280
rect 495400 28240 554872 28268
rect 495400 28228 495406 28240
rect 554866 28228 554872 28240
rect 554924 28228 554930 28280
rect 369854 27548 369860 27600
rect 369912 27588 369918 27600
rect 370498 27588 370504 27600
rect 369912 27560 370504 27588
rect 369912 27548 369918 27560
rect 370498 27548 370504 27560
rect 370556 27548 370562 27600
rect 398834 27588 398840 27600
rect 398795 27560 398840 27588
rect 398834 27548 398840 27560
rect 398892 27548 398898 27600
rect 407206 27588 407212 27600
rect 407167 27560 407212 27588
rect 407206 27548 407212 27560
rect 407264 27548 407270 27600
rect 442997 27591 443055 27597
rect 442997 27557 443009 27591
rect 443043 27588 443055 27591
rect 443178 27588 443184 27600
rect 443043 27560 443184 27588
rect 443043 27557 443055 27560
rect 442997 27551 443055 27557
rect 443178 27548 443184 27560
rect 443236 27548 443242 27600
rect 449986 27548 449992 27600
rect 450044 27588 450050 27600
rect 450354 27588 450360 27600
rect 450044 27560 450360 27588
rect 450044 27548 450050 27560
rect 450354 27548 450360 27560
rect 450412 27548 450418 27600
rect 535454 27588 535460 27600
rect 535415 27560 535460 27588
rect 535454 27548 535460 27560
rect 535512 27548 535518 27600
rect 275830 26936 275836 26988
rect 275888 26976 275894 26988
rect 335354 26976 335360 26988
rect 275888 26948 335360 26976
rect 275888 26936 275894 26948
rect 335354 26936 335360 26948
rect 335412 26936 335418 26988
rect 431862 26936 431868 26988
rect 431920 26976 431926 26988
rect 491294 26976 491300 26988
rect 431920 26948 491300 26976
rect 431920 26936 431926 26948
rect 491294 26936 491300 26948
rect 491352 26936 491358 26988
rect 93762 26868 93768 26920
rect 93820 26908 93826 26920
rect 154574 26908 154580 26920
rect 93820 26880 154580 26908
rect 93820 26868 93826 26880
rect 154574 26868 154580 26880
rect 154632 26868 154638 26920
rect 158622 26868 158628 26920
rect 158680 26908 158686 26920
rect 218146 26908 218152 26920
rect 158680 26880 218152 26908
rect 158680 26868 158686 26880
rect 218146 26868 218152 26880
rect 218204 26868 218210 26920
rect 237282 26868 237288 26920
rect 237340 26908 237346 26920
rect 296806 26908 296812 26920
rect 237340 26880 296812 26908
rect 237340 26868 237346 26880
rect 296806 26868 296812 26880
rect 296864 26868 296870 26920
rect 311802 26868 311808 26920
rect 311860 26908 311866 26920
rect 372614 26908 372620 26920
rect 311860 26880 372620 26908
rect 311860 26868 311866 26880
rect 372614 26868 372620 26880
rect 372672 26868 372678 26920
rect 373902 26868 373908 26920
rect 373960 26908 373966 26920
rect 433334 26908 433340 26920
rect 373960 26880 433340 26908
rect 373960 26868 373966 26880
rect 433334 26868 433340 26880
rect 433392 26868 433398 26920
rect 492582 26868 492588 26920
rect 492640 26908 492646 26920
rect 552014 26908 552020 26920
rect 492640 26880 552020 26908
rect 492640 26868 492646 26880
rect 552014 26868 552020 26880
rect 552072 26868 552078 26920
rect 353202 25576 353208 25628
rect 353260 25616 353266 25628
rect 412634 25616 412640 25628
rect 353260 25588 412640 25616
rect 353260 25576 353266 25588
rect 412634 25576 412640 25588
rect 412692 25576 412698 25628
rect 91002 25508 91008 25560
rect 91060 25548 91066 25560
rect 150526 25548 150532 25560
rect 91060 25520 150532 25548
rect 91060 25508 91066 25520
rect 150526 25508 150532 25520
rect 150584 25508 150590 25560
rect 154482 25508 154488 25560
rect 154540 25548 154546 25560
rect 215294 25548 215300 25560
rect 154540 25520 215300 25548
rect 154540 25508 154546 25520
rect 215294 25508 215300 25520
rect 215352 25508 215358 25560
rect 226242 25508 226248 25560
rect 226300 25548 226306 25560
rect 287146 25548 287152 25560
rect 226300 25520 287152 25548
rect 226300 25508 226306 25520
rect 287146 25508 287152 25520
rect 287204 25508 287210 25560
rect 293770 25508 293776 25560
rect 293828 25548 293834 25560
rect 354674 25548 354680 25560
rect 293828 25520 354680 25548
rect 293828 25508 293834 25520
rect 354674 25508 354680 25520
rect 354732 25508 354738 25560
rect 427722 25508 427728 25560
rect 427780 25548 427786 25560
rect 487154 25548 487160 25560
rect 427780 25520 487160 25548
rect 427780 25508 427786 25520
rect 487154 25508 487160 25520
rect 487212 25508 487218 25560
rect 488442 25508 488448 25560
rect 488500 25548 488506 25560
rect 547874 25548 547880 25560
rect 488500 25520 547880 25548
rect 488500 25508 488506 25520
rect 547874 25508 547880 25520
rect 547932 25508 547938 25560
rect 278682 24148 278688 24200
rect 278740 24188 278746 24200
rect 339494 24188 339500 24200
rect 278740 24160 339500 24188
rect 278740 24148 278746 24160
rect 339494 24148 339500 24160
rect 339552 24148 339558 24200
rect 86862 24080 86868 24132
rect 86920 24120 86926 24132
rect 147674 24120 147680 24132
rect 86920 24092 147680 24120
rect 86920 24080 86926 24092
rect 147674 24080 147680 24092
rect 147732 24080 147738 24132
rect 151722 24080 151728 24132
rect 151780 24120 151786 24132
rect 211154 24120 211160 24132
rect 151780 24092 211160 24120
rect 151780 24080 151786 24092
rect 211154 24080 211160 24092
rect 211212 24080 211218 24132
rect 215110 24080 215116 24132
rect 215168 24120 215174 24132
rect 276014 24120 276020 24132
rect 215168 24092 276020 24120
rect 215168 24080 215174 24092
rect 276014 24080 276020 24092
rect 276072 24080 276078 24132
rect 286962 24080 286968 24132
rect 287020 24120 287026 24132
rect 347866 24120 347872 24132
rect 287020 24092 347872 24120
rect 287020 24080 287026 24092
rect 347866 24080 347872 24092
rect 347924 24080 347930 24132
rect 351822 24080 351828 24132
rect 351880 24120 351886 24132
rect 411254 24120 411260 24132
rect 351880 24092 411260 24120
rect 351880 24080 351886 24092
rect 411254 24080 411260 24092
rect 411312 24080 411318 24132
rect 423490 24080 423496 24132
rect 423548 24120 423554 24132
rect 484394 24120 484400 24132
rect 423548 24092 484400 24120
rect 423548 24080 423554 24092
rect 484394 24080 484400 24092
rect 484452 24080 484458 24132
rect 499482 24080 499488 24132
rect 499540 24120 499546 24132
rect 558914 24120 558920 24132
rect 499540 24092 558920 24120
rect 499540 24080 499546 24092
rect 558914 24080 558920 24092
rect 558972 24080 558978 24132
rect 275922 22788 275928 22840
rect 275980 22828 275986 22840
rect 336734 22828 336740 22840
rect 275980 22800 336740 22828
rect 275980 22788 275986 22800
rect 336734 22788 336740 22800
rect 336792 22788 336798 22840
rect 344922 22788 344928 22840
rect 344980 22828 344986 22840
rect 404354 22828 404360 22840
rect 344980 22800 404360 22828
rect 344980 22788 344986 22800
rect 404354 22788 404360 22800
rect 404412 22788 404418 22840
rect 84010 22720 84016 22772
rect 84068 22760 84074 22772
rect 143534 22760 143540 22772
rect 84068 22732 143540 22760
rect 84068 22720 84074 22732
rect 143534 22720 143540 22732
rect 143592 22720 143598 22772
rect 147582 22720 147588 22772
rect 147640 22760 147646 22772
rect 208394 22760 208400 22772
rect 147640 22732 208400 22760
rect 147640 22720 147646 22732
rect 208394 22720 208400 22732
rect 208452 22720 208458 22772
rect 212442 22720 212448 22772
rect 212500 22760 212506 22772
rect 271874 22760 271880 22772
rect 212500 22732 271880 22760
rect 212500 22720 212506 22732
rect 271874 22720 271880 22732
rect 271932 22720 271938 22772
rect 285582 22720 285588 22772
rect 285640 22760 285646 22772
rect 346394 22760 346400 22772
rect 285640 22732 346400 22760
rect 285640 22720 285646 22732
rect 346394 22720 346400 22732
rect 346452 22720 346458 22772
rect 419442 22720 419448 22772
rect 419500 22760 419506 22772
rect 478874 22760 478880 22772
rect 419500 22732 478880 22760
rect 419500 22720 419506 22732
rect 478874 22720 478880 22732
rect 478932 22720 478938 22772
rect 79962 21360 79968 21412
rect 80020 21400 80026 21412
rect 140866 21400 140872 21412
rect 80020 21372 140872 21400
rect 80020 21360 80026 21372
rect 140866 21360 140872 21372
rect 140924 21360 140930 21412
rect 144822 21360 144828 21412
rect 144880 21400 144886 21412
rect 204254 21400 204260 21412
rect 144880 21372 204260 21400
rect 144880 21360 144886 21372
rect 204254 21360 204260 21372
rect 204312 21360 204318 21412
rect 205450 21360 205456 21412
rect 205508 21400 205514 21412
rect 264974 21400 264980 21412
rect 205508 21372 264980 21400
rect 205508 21360 205514 21372
rect 264974 21360 264980 21372
rect 265032 21360 265038 21412
rect 269022 21360 269028 21412
rect 269080 21400 269086 21412
rect 329834 21400 329840 21412
rect 269080 21372 329840 21400
rect 269080 21360 269086 21372
rect 329834 21360 329840 21372
rect 329892 21360 329898 21412
rect 336550 21360 336556 21412
rect 336608 21400 336614 21412
rect 397454 21400 397460 21412
rect 336608 21372 397460 21400
rect 336608 21360 336614 21372
rect 397454 21360 397460 21372
rect 397512 21360 397518 21412
rect 412542 21360 412548 21412
rect 412600 21400 412606 21412
rect 471974 21400 471980 21412
rect 412600 21372 471980 21400
rect 412600 21360 412606 21372
rect 471974 21360 471980 21372
rect 472032 21360 472038 21412
rect 474642 21360 474648 21412
rect 474700 21400 474706 21412
rect 534074 21400 534080 21412
rect 474700 21372 534080 21400
rect 474700 21360 474706 21372
rect 534074 21360 534080 21372
rect 534132 21360 534138 21412
rect 75822 19932 75828 19984
rect 75880 19972 75886 19984
rect 136634 19972 136640 19984
rect 75880 19944 136640 19972
rect 75880 19932 75886 19944
rect 136634 19932 136640 19944
rect 136692 19932 136698 19984
rect 140682 19932 140688 19984
rect 140740 19972 140746 19984
rect 201586 19972 201592 19984
rect 140740 19944 201592 19972
rect 140740 19932 140746 19944
rect 201586 19932 201592 19944
rect 201644 19932 201650 19984
rect 208302 19932 208308 19984
rect 208360 19972 208366 19984
rect 269114 19972 269120 19984
rect 208360 19944 269120 19972
rect 208360 19932 208366 19944
rect 269114 19932 269120 19944
rect 269172 19932 269178 19984
rect 273162 19932 273168 19984
rect 273220 19972 273226 19984
rect 332594 19972 332600 19984
rect 273220 19944 332600 19972
rect 273220 19932 273226 19944
rect 332594 19932 332600 19944
rect 332652 19932 332658 19984
rect 333882 19932 333888 19984
rect 333940 19972 333946 19984
rect 393314 19972 393320 19984
rect 333940 19944 393320 19972
rect 333940 19932 333946 19944
rect 393314 19932 393320 19944
rect 393372 19932 393378 19984
rect 408402 19932 408408 19984
rect 408460 19972 408466 19984
rect 467834 19972 467840 19984
rect 408460 19944 467840 19972
rect 408460 19932 408466 19944
rect 467834 19932 467840 19944
rect 467892 19932 467898 19984
rect 470502 19932 470508 19984
rect 470560 19972 470566 19984
rect 529934 19972 529940 19984
rect 470560 19944 529940 19972
rect 470560 19932 470566 19944
rect 529934 19932 529940 19944
rect 529992 19932 529998 19984
rect 333974 19292 333980 19304
rect 333935 19264 333980 19292
rect 333974 19252 333980 19264
rect 334032 19252 334038 19304
rect 345014 19292 345020 19304
rect 344975 19264 345020 19292
rect 345014 19252 345020 19264
rect 345072 19252 345078 19304
rect 372614 19292 372620 19304
rect 372575 19264 372620 19292
rect 372614 19252 372620 19264
rect 372672 19252 372678 19304
rect 394694 19292 394700 19304
rect 394655 19264 394700 19292
rect 394694 19252 394700 19264
rect 394752 19252 394758 19304
rect 397454 19292 397460 19304
rect 397415 19264 397460 19292
rect 397454 19252 397460 19264
rect 397512 19252 397518 19304
rect 515950 19252 515956 19304
rect 516008 19292 516014 19304
rect 516134 19292 516140 19304
rect 516008 19264 516140 19292
rect 516008 19252 516014 19264
rect 516134 19252 516140 19264
rect 516192 19252 516198 19304
rect 73062 18572 73068 18624
rect 73120 18612 73126 18624
rect 132586 18612 132592 18624
rect 73120 18584 132592 18612
rect 73120 18572 73126 18584
rect 132586 18572 132592 18584
rect 132644 18572 132650 18624
rect 136450 18572 136456 18624
rect 136508 18612 136514 18624
rect 197354 18612 197360 18624
rect 136508 18584 197360 18612
rect 136508 18572 136514 18584
rect 197354 18572 197360 18584
rect 197412 18572 197418 18624
rect 201402 18572 201408 18624
rect 201460 18612 201466 18624
rect 262306 18612 262312 18624
rect 201460 18584 262312 18612
rect 201460 18572 201466 18584
rect 262306 18572 262312 18584
rect 262364 18572 262370 18624
rect 266262 18572 266268 18624
rect 266320 18612 266326 18624
rect 325694 18612 325700 18624
rect 266320 18584 325700 18612
rect 266320 18572 266326 18584
rect 325694 18572 325700 18584
rect 325752 18572 325758 18624
rect 329742 18572 329748 18624
rect 329800 18612 329806 18624
rect 390646 18612 390652 18624
rect 329800 18584 390652 18612
rect 329800 18572 329806 18584
rect 390646 18572 390652 18584
rect 390704 18572 390710 18624
rect 405642 18572 405648 18624
rect 405700 18612 405706 18624
rect 465074 18612 465080 18624
rect 405700 18584 465080 18612
rect 405700 18572 405706 18584
rect 465074 18572 465080 18584
rect 465132 18572 465138 18624
rect 467742 18572 467748 18624
rect 467800 18612 467806 18624
rect 527266 18612 527272 18624
rect 467800 18584 527272 18612
rect 467800 18572 467806 18584
rect 527266 18572 527272 18584
rect 527324 18572 527330 18624
rect 523862 17892 523868 17944
rect 523920 17932 523926 17944
rect 580074 17932 580080 17944
rect 523920 17904 580080 17932
rect 523920 17892 523926 17904
rect 580074 17892 580080 17904
rect 580132 17892 580138 17944
rect 401502 17280 401508 17332
rect 401560 17320 401566 17332
rect 460934 17320 460940 17332
rect 401560 17292 460940 17320
rect 401560 17280 401566 17292
rect 460934 17280 460940 17292
rect 460992 17280 460998 17332
rect 129642 17212 129648 17264
rect 129700 17252 129706 17264
rect 190454 17252 190460 17264
rect 129700 17224 190460 17252
rect 129700 17212 129706 17224
rect 190454 17212 190460 17224
rect 190512 17212 190518 17264
rect 197170 17212 197176 17264
rect 197228 17252 197234 17264
rect 258074 17252 258080 17264
rect 197228 17224 258080 17252
rect 197228 17212 197234 17224
rect 258074 17212 258080 17224
rect 258132 17212 258138 17264
rect 262122 17212 262128 17264
rect 262180 17252 262186 17264
rect 321646 17252 321652 17264
rect 262180 17224 321652 17252
rect 262180 17212 262186 17224
rect 321646 17212 321652 17224
rect 321704 17212 321710 17264
rect 326982 17212 326988 17264
rect 327040 17252 327046 17264
rect 386414 17252 386420 17264
rect 327040 17224 386420 17252
rect 327040 17212 327046 17224
rect 386414 17212 386420 17224
rect 386472 17212 386478 17264
rect 452562 17212 452568 17264
rect 452620 17252 452626 17264
rect 512086 17252 512092 17264
rect 452620 17224 512092 17252
rect 452620 17212 452626 17224
rect 512086 17212 512092 17224
rect 512144 17212 512150 17264
rect 126882 15920 126888 15972
rect 126940 15960 126946 15972
rect 186314 15960 186320 15972
rect 126940 15932 186320 15960
rect 126940 15920 126946 15932
rect 186314 15920 186320 15932
rect 186372 15920 186378 15972
rect 315942 15920 315948 15972
rect 316000 15960 316006 15972
rect 375374 15960 375380 15972
rect 316000 15932 375380 15960
rect 316000 15920 316006 15932
rect 375374 15920 375380 15932
rect 375432 15920 375438 15972
rect 66898 15852 66904 15904
rect 66956 15892 66962 15904
rect 126974 15892 126980 15904
rect 66956 15864 126980 15892
rect 66956 15852 66962 15864
rect 126974 15852 126980 15864
rect 127032 15852 127038 15904
rect 194502 15852 194508 15904
rect 194560 15892 194566 15904
rect 253934 15892 253940 15904
rect 194560 15864 253940 15892
rect 194560 15852 194566 15864
rect 253934 15852 253940 15864
rect 253992 15852 253998 15904
rect 257890 15852 257896 15904
rect 257948 15892 257954 15904
rect 318794 15892 318800 15904
rect 257948 15864 318800 15892
rect 257948 15852 257954 15864
rect 318794 15852 318800 15864
rect 318852 15852 318858 15904
rect 397362 15852 397368 15904
rect 397420 15892 397426 15904
rect 458174 15892 458180 15904
rect 397420 15864 458180 15892
rect 397420 15852 397426 15864
rect 458174 15852 458180 15864
rect 458232 15852 458238 15904
rect 469122 15852 469128 15904
rect 469180 15892 469186 15904
rect 528646 15892 528652 15904
rect 469180 15864 528652 15892
rect 469180 15852 469186 15864
rect 528646 15852 528652 15864
rect 528704 15852 528710 15904
rect 248322 14492 248328 14544
rect 248380 14532 248386 14544
rect 307754 14532 307760 14544
rect 248380 14504 307760 14532
rect 248380 14492 248386 14504
rect 307754 14492 307760 14504
rect 307812 14492 307818 14544
rect 355962 14492 355968 14544
rect 356020 14532 356026 14544
rect 416866 14532 416872 14544
rect 356020 14504 416872 14532
rect 356020 14492 356026 14504
rect 416866 14492 416872 14504
rect 416924 14492 416930 14544
rect 448422 14492 448428 14544
rect 448480 14532 448486 14544
rect 507854 14532 507860 14544
rect 448480 14504 507860 14532
rect 448480 14492 448486 14504
rect 507854 14492 507860 14504
rect 507912 14492 507918 14544
rect 122742 14424 122748 14476
rect 122800 14464 122806 14476
rect 183646 14464 183652 14476
rect 122800 14436 183652 14464
rect 122800 14424 122806 14436
rect 183646 14424 183652 14436
rect 183704 14424 183710 14476
rect 187602 14424 187608 14476
rect 187660 14464 187666 14476
rect 247034 14464 247040 14476
rect 187660 14436 247040 14464
rect 187660 14424 187666 14436
rect 247034 14424 247040 14436
rect 247092 14424 247098 14476
rect 304902 14424 304908 14476
rect 304960 14464 304966 14476
rect 365806 14464 365812 14476
rect 304960 14436 365812 14464
rect 304960 14424 304966 14436
rect 365806 14424 365812 14436
rect 365864 14424 365870 14476
rect 413922 14424 413928 14476
rect 413980 14464 413986 14476
rect 473354 14464 473360 14476
rect 413980 14436 473360 14464
rect 413980 14424 413986 14436
rect 473354 14424 473360 14436
rect 473412 14424 473418 14476
rect 509142 14424 509148 14476
rect 509200 14464 509206 14476
rect 568574 14464 568580 14476
rect 509200 14436 568580 14464
rect 509200 14424 509206 14436
rect 568574 14424 568580 14436
rect 568632 14424 568638 14476
rect 309042 13132 309048 13184
rect 309100 13172 309106 13184
rect 368474 13172 368480 13184
rect 309100 13144 368480 13172
rect 309100 13132 309106 13144
rect 368474 13132 368480 13144
rect 368532 13132 368538 13184
rect 118510 13064 118516 13116
rect 118568 13104 118574 13116
rect 179414 13104 179420 13116
rect 118568 13076 179420 13104
rect 118568 13064 118574 13076
rect 179414 13064 179420 13076
rect 179472 13064 179478 13116
rect 183462 13064 183468 13116
rect 183520 13104 183526 13116
rect 244366 13104 244372 13116
rect 183520 13076 244372 13104
rect 183520 13064 183526 13076
rect 244366 13064 244372 13076
rect 244424 13064 244430 13116
rect 251082 13064 251088 13116
rect 251140 13104 251146 13116
rect 311894 13104 311900 13116
rect 251140 13076 311900 13104
rect 251140 13064 251146 13076
rect 311894 13064 311900 13076
rect 311952 13064 311958 13116
rect 381538 13064 381544 13116
rect 381596 13104 381602 13116
rect 441614 13104 441620 13116
rect 381596 13076 441620 13104
rect 381596 13064 381602 13076
rect 441614 13064 441620 13076
rect 441672 13064 441678 13116
rect 444282 13064 444288 13116
rect 444340 13104 444346 13116
rect 503714 13104 503720 13116
rect 444340 13076 503720 13104
rect 444340 13064 444346 13076
rect 503714 13064 503720 13076
rect 503772 13064 503778 13116
rect 505002 13064 505008 13116
rect 505060 13104 505066 13116
rect 564434 13104 564440 13116
rect 505060 13076 564440 13104
rect 505060 13064 505066 13076
rect 564434 13064 564440 13076
rect 564492 13064 564498 13116
rect 336734 12452 336740 12504
rect 336792 12452 336798 12504
rect 338114 12452 338120 12504
rect 338172 12452 338178 12504
rect 346394 12452 346400 12504
rect 346452 12452 346458 12504
rect 331306 12384 331312 12436
rect 331364 12424 331370 12436
rect 332410 12424 332416 12436
rect 331364 12396 332416 12424
rect 331364 12384 331370 12396
rect 332410 12384 332416 12396
rect 332468 12384 332474 12436
rect 332594 12384 332600 12436
rect 332652 12424 332658 12436
rect 333606 12424 333612 12436
rect 332652 12396 333612 12424
rect 332652 12384 332658 12396
rect 333606 12384 333612 12396
rect 333664 12384 333670 12436
rect 335354 12384 335360 12436
rect 335412 12424 335418 12436
rect 335906 12424 335912 12436
rect 335412 12396 335912 12424
rect 335412 12384 335418 12396
rect 335906 12384 335912 12396
rect 335964 12384 335970 12436
rect 336752 12356 336780 12452
rect 337102 12356 337108 12368
rect 336752 12328 337108 12356
rect 337102 12316 337108 12328
rect 337160 12316 337166 12368
rect 338132 12356 338160 12452
rect 340874 12384 340880 12436
rect 340932 12424 340938 12436
rect 341886 12424 341892 12436
rect 340932 12396 341892 12424
rect 340932 12384 340938 12396
rect 341886 12384 341892 12396
rect 341944 12384 341950 12436
rect 338298 12356 338304 12368
rect 338132 12328 338304 12356
rect 338298 12316 338304 12328
rect 338356 12316 338362 12368
rect 346412 12356 346440 12452
rect 351914 12384 351920 12436
rect 351972 12424 351978 12436
rect 352558 12424 352564 12436
rect 351972 12396 352564 12424
rect 351972 12384 351978 12396
rect 352558 12384 352564 12396
rect 352616 12384 352622 12436
rect 393314 12384 393320 12436
rect 393372 12424 393378 12436
rect 394234 12424 394240 12436
rect 393372 12396 394240 12424
rect 393372 12384 393378 12396
rect 394234 12384 394240 12396
rect 394292 12384 394298 12436
rect 401594 12384 401600 12436
rect 401652 12424 401658 12436
rect 402514 12424 402520 12436
rect 401652 12396 402520 12424
rect 401652 12384 401658 12396
rect 402514 12384 402520 12396
rect 402572 12384 402578 12436
rect 404354 12384 404360 12436
rect 404412 12424 404418 12436
rect 404906 12424 404912 12436
rect 404412 12396 404912 12424
rect 404412 12384 404418 12396
rect 404906 12384 404912 12396
rect 404964 12384 404970 12436
rect 448514 12384 448520 12436
rect 448572 12424 448578 12436
rect 448974 12424 448980 12436
rect 448572 12396 448980 12424
rect 448572 12384 448578 12396
rect 448974 12384 448980 12396
rect 449032 12384 449038 12436
rect 529934 12384 529940 12436
rect 529992 12424 529998 12436
rect 531038 12424 531044 12436
rect 529992 12396 531044 12424
rect 529992 12384 529998 12396
rect 531038 12384 531044 12396
rect 531096 12384 531102 12436
rect 534074 12384 534080 12436
rect 534132 12424 534138 12436
rect 534534 12424 534540 12436
rect 534132 12396 534540 12424
rect 534132 12384 534138 12396
rect 534534 12384 534540 12396
rect 534592 12384 534598 12436
rect 542354 12384 542360 12436
rect 542412 12424 542418 12436
rect 542906 12424 542912 12436
rect 542412 12396 542912 12424
rect 542412 12384 542418 12396
rect 542906 12384 542912 12396
rect 542964 12384 542970 12436
rect 346670 12356 346676 12368
rect 346412 12328 346676 12356
rect 346670 12316 346676 12328
rect 346728 12316 346734 12368
rect 407206 12288 407212 12300
rect 407167 12260 407212 12288
rect 407206 12248 407212 12260
rect 407264 12248 407270 12300
rect 351178 11772 351184 11824
rect 351236 11812 351242 11824
rect 406102 11812 406108 11824
rect 351236 11784 406108 11812
rect 351236 11772 351242 11784
rect 406102 11772 406108 11784
rect 406160 11772 406166 11824
rect 441522 11772 441528 11824
rect 441580 11812 441586 11824
rect 500954 11812 500960 11824
rect 441580 11784 500960 11812
rect 441580 11772 441586 11784
rect 500954 11772 500960 11784
rect 501012 11772 501018 11824
rect 115842 11704 115848 11756
rect 115900 11744 115906 11756
rect 175366 11744 175372 11756
rect 115900 11716 175372 11744
rect 115900 11704 115906 11716
rect 175366 11704 175372 11716
rect 175424 11704 175430 11756
rect 179230 11704 179236 11756
rect 179288 11744 179294 11756
rect 240134 11744 240140 11756
rect 179288 11716 240140 11744
rect 179288 11704 179294 11716
rect 240134 11704 240140 11716
rect 240192 11704 240198 11756
rect 241422 11704 241428 11756
rect 241480 11744 241486 11756
rect 300854 11744 300860 11756
rect 241480 11716 300860 11744
rect 241480 11704 241486 11716
rect 300854 11704 300860 11716
rect 300912 11704 300918 11756
rect 302142 11704 302148 11756
rect 302200 11744 302206 11756
rect 361574 11744 361580 11756
rect 302200 11716 361580 11744
rect 302200 11704 302206 11716
rect 361574 11704 361580 11716
rect 361632 11704 361638 11756
rect 416682 11704 416688 11756
rect 416740 11744 416746 11756
rect 477586 11744 477592 11756
rect 416740 11716 477592 11744
rect 416740 11704 416746 11716
rect 477586 11704 477592 11716
rect 477644 11704 477650 11756
rect 502150 11704 502156 11756
rect 502208 11744 502214 11756
rect 563146 11744 563152 11756
rect 502208 11716 563152 11744
rect 502208 11704 502214 11716
rect 563146 11704 563152 11716
rect 563204 11704 563210 11756
rect 176562 10344 176568 10396
rect 176620 10384 176626 10396
rect 236086 10384 236092 10396
rect 176620 10356 236092 10384
rect 176620 10344 176626 10356
rect 236086 10344 236092 10356
rect 236144 10344 236150 10396
rect 298002 10344 298008 10396
rect 298060 10384 298066 10396
rect 357434 10384 357440 10396
rect 298060 10356 357440 10384
rect 298060 10344 298066 10356
rect 357434 10344 357440 10356
rect 357492 10344 357498 10396
rect 111702 10276 111708 10328
rect 111760 10316 111766 10328
rect 172514 10316 172520 10328
rect 111760 10288 172520 10316
rect 111760 10276 111766 10288
rect 172514 10276 172520 10288
rect 172572 10276 172578 10328
rect 233142 10276 233148 10328
rect 233200 10316 233206 10328
rect 293954 10316 293960 10328
rect 233200 10288 293960 10316
rect 233200 10276 233206 10288
rect 293954 10276 293960 10288
rect 294012 10276 294018 10328
rect 303522 10276 303528 10328
rect 303580 10316 303586 10328
rect 364518 10316 364524 10328
rect 303580 10288 364524 10316
rect 303580 10276 303586 10288
rect 364518 10276 364524 10288
rect 364576 10276 364582 10328
rect 367738 10276 367744 10328
rect 367796 10316 367802 10328
rect 415394 10316 415400 10328
rect 367796 10288 415400 10316
rect 367796 10276 367802 10288
rect 415394 10276 415400 10288
rect 415452 10276 415458 10328
rect 437382 10276 437388 10328
rect 437440 10316 437446 10328
rect 496814 10316 496820 10328
rect 437440 10288 496820 10316
rect 437440 10276 437446 10288
rect 496814 10276 496820 10288
rect 496872 10276 496878 10328
rect 498102 10276 498108 10328
rect 498160 10316 498166 10328
rect 557534 10316 557540 10328
rect 498160 10288 557540 10316
rect 498160 10276 498166 10288
rect 557534 10276 557540 10288
rect 557592 10276 557598 10328
rect 333977 9707 334035 9713
rect 333977 9673 333989 9707
rect 334023 9704 334035 9707
rect 334710 9704 334716 9716
rect 334023 9676 334716 9704
rect 334023 9673 334035 9676
rect 333977 9667 334035 9673
rect 334710 9664 334716 9676
rect 334768 9664 334774 9716
rect 345017 9707 345075 9713
rect 345017 9673 345029 9707
rect 345063 9704 345075 9707
rect 345474 9704 345480 9716
rect 345063 9676 345480 9704
rect 345063 9673 345075 9676
rect 345017 9667 345075 9673
rect 345474 9664 345480 9676
rect 345532 9664 345538 9716
rect 372617 9707 372675 9713
rect 372617 9673 372629 9707
rect 372663 9704 372675 9707
rect 372890 9704 372896 9716
rect 372663 9676 372896 9704
rect 372663 9673 372675 9676
rect 372617 9667 372675 9673
rect 372890 9664 372896 9676
rect 372948 9664 372954 9716
rect 394697 9707 394755 9713
rect 394697 9673 394709 9707
rect 394743 9704 394755 9707
rect 395430 9704 395436 9716
rect 394743 9676 395436 9704
rect 394743 9673 394755 9676
rect 394697 9667 394755 9673
rect 395430 9664 395436 9676
rect 395488 9664 395494 9716
rect 397457 9707 397515 9713
rect 397457 9673 397469 9707
rect 397503 9704 397515 9707
rect 397822 9704 397828 9716
rect 397503 9676 397828 9704
rect 397503 9673 397515 9676
rect 397457 9667 397515 9673
rect 397822 9664 397828 9676
rect 397880 9664 397886 9716
rect 398837 9707 398895 9713
rect 398837 9673 398849 9707
rect 398883 9704 398895 9707
rect 399018 9704 399024 9716
rect 398883 9676 399024 9704
rect 398883 9673 398895 9676
rect 398837 9667 398895 9673
rect 399018 9664 399024 9676
rect 399076 9664 399082 9716
rect 442994 9704 443000 9716
rect 442955 9676 443000 9704
rect 442994 9664 443000 9676
rect 443052 9664 443058 9716
rect 535457 9707 535515 9713
rect 535457 9673 535469 9707
rect 535503 9704 535515 9707
rect 535730 9704 535736 9716
rect 535503 9676 535736 9704
rect 535503 9673 535515 9676
rect 535457 9667 535515 9673
rect 535730 9664 535736 9676
rect 535788 9664 535794 9716
rect 411254 9596 411260 9648
rect 411312 9636 411318 9648
rect 412085 9639 412143 9645
rect 412085 9636 412097 9639
rect 411312 9608 412097 9636
rect 411312 9596 411318 9608
rect 412085 9605 412097 9608
rect 412131 9605 412143 9639
rect 412085 9599 412143 9605
rect 419534 9596 419540 9648
rect 419592 9636 419598 9648
rect 420365 9639 420423 9645
rect 420365 9636 420377 9639
rect 419592 9608 420377 9636
rect 419592 9596 419598 9608
rect 420365 9605 420377 9608
rect 420411 9605 420423 9639
rect 420365 9599 420423 9605
rect 516134 9596 516140 9648
rect 516192 9636 516198 9648
rect 516781 9639 516839 9645
rect 516781 9636 516793 9639
rect 516192 9608 516793 9636
rect 516192 9596 516198 9608
rect 516781 9605 516793 9608
rect 516827 9605 516839 9639
rect 516781 9599 516839 9605
rect 520277 9639 520335 9645
rect 520277 9605 520289 9639
rect 520323 9636 520335 9639
rect 520366 9636 520372 9648
rect 520323 9608 520372 9636
rect 520323 9605 520335 9608
rect 520277 9599 520335 9605
rect 520366 9596 520372 9608
rect 520424 9596 520430 9648
rect 230382 8984 230388 9036
rect 230440 9024 230446 9036
rect 290734 9024 290740 9036
rect 230440 8996 290740 9024
rect 230440 8984 230446 8996
rect 290734 8984 290740 8996
rect 290792 8984 290798 9036
rect 291102 8984 291108 9036
rect 291160 9024 291166 9036
rect 351362 9024 351368 9036
rect 291160 8996 351368 9024
rect 291160 8984 291166 8996
rect 351362 8984 351368 8996
rect 351420 8984 351426 9036
rect 108942 8916 108948 8968
rect 109000 8956 109006 8968
rect 169386 8956 169392 8968
rect 109000 8928 169392 8956
rect 109000 8916 109006 8928
rect 169386 8916 169392 8928
rect 169444 8916 169450 8968
rect 172422 8916 172428 8968
rect 172480 8956 172486 8968
rect 233694 8956 233700 8968
rect 172480 8928 233700 8956
rect 172480 8916 172486 8928
rect 233694 8916 233700 8928
rect 233752 8916 233758 8968
rect 347682 8916 347688 8968
rect 347740 8956 347746 8968
rect 408678 8956 408684 8968
rect 347740 8928 408684 8956
rect 347740 8916 347746 8928
rect 408678 8916 408684 8928
rect 408736 8916 408742 8968
rect 430482 8916 430488 8968
rect 430540 8956 430546 8968
rect 490558 8956 490564 8968
rect 430540 8928 490564 8956
rect 430540 8916 430546 8928
rect 490558 8916 490564 8928
rect 490616 8916 490622 8968
rect 491202 8916 491208 8968
rect 491260 8956 491266 8968
rect 551186 8956 551192 8968
rect 491260 8928 551192 8956
rect 491260 8916 491266 8928
rect 551186 8916 551192 8928
rect 551244 8916 551250 8968
rect 104802 7624 104808 7676
rect 104860 7664 104866 7676
rect 165890 7664 165896 7676
rect 104860 7636 165896 7664
rect 104860 7624 104866 7636
rect 165890 7624 165896 7636
rect 165948 7624 165954 7676
rect 169662 7624 169668 7676
rect 169720 7664 169726 7676
rect 230106 7664 230112 7676
rect 169720 7636 230112 7664
rect 169720 7624 169726 7636
rect 230106 7624 230112 7636
rect 230164 7624 230170 7676
rect 340782 7624 340788 7676
rect 340840 7664 340846 7676
rect 401318 7664 401324 7676
rect 340840 7636 401324 7664
rect 340840 7624 340846 7636
rect 401318 7624 401324 7636
rect 401376 7624 401382 7676
rect 433334 7624 433340 7676
rect 433392 7664 433398 7676
rect 434622 7664 434628 7676
rect 433392 7636 434628 7664
rect 433392 7624 433398 7636
rect 434622 7624 434628 7636
rect 434680 7624 434686 7676
rect 451274 7624 451280 7676
rect 451332 7664 451338 7676
rect 452470 7664 452476 7676
rect 451332 7636 452476 7664
rect 451332 7624 451338 7636
rect 452470 7624 452476 7636
rect 452528 7624 452534 7676
rect 481542 7624 481548 7676
rect 481600 7664 481606 7676
rect 541710 7664 541716 7676
rect 481600 7636 541716 7664
rect 481600 7624 481606 7636
rect 541710 7624 541716 7636
rect 541768 7624 541774 7676
rect 137922 7556 137928 7608
rect 137980 7596 137986 7608
rect 199194 7596 199200 7608
rect 137980 7568 199200 7596
rect 137980 7556 137986 7568
rect 199194 7556 199200 7568
rect 199252 7556 199258 7608
rect 223482 7556 223488 7608
rect 223540 7596 223546 7608
rect 283650 7596 283656 7608
rect 223540 7568 283656 7596
rect 223540 7556 223546 7568
rect 283650 7556 283656 7568
rect 283708 7556 283714 7608
rect 284202 7556 284208 7608
rect 284260 7596 284266 7608
rect 344278 7596 344284 7608
rect 284260 7568 344284 7596
rect 284260 7556 284266 7568
rect 344278 7556 344284 7568
rect 344336 7556 344342 7608
rect 347774 7556 347780 7608
rect 347832 7596 347838 7608
rect 349062 7596 349068 7608
rect 347832 7568 349068 7596
rect 347832 7556 347838 7568
rect 349062 7556 349068 7568
rect 349120 7556 349126 7608
rect 365714 7556 365720 7608
rect 365772 7596 365778 7608
rect 366910 7596 366916 7608
rect 365772 7568 366916 7596
rect 365772 7556 365778 7568
rect 366910 7556 366916 7568
rect 366968 7556 366974 7608
rect 390554 7556 390560 7608
rect 390612 7596 390618 7608
rect 391842 7596 391848 7608
rect 390612 7568 391848 7596
rect 390612 7556 390618 7568
rect 391842 7556 391848 7568
rect 391900 7556 391906 7608
rect 408494 7556 408500 7608
rect 408552 7596 408558 7608
rect 409690 7596 409696 7608
rect 408552 7568 409696 7596
rect 408552 7556 408558 7568
rect 409690 7556 409696 7568
rect 409748 7556 409754 7608
rect 423582 7556 423588 7608
rect 423640 7596 423646 7608
rect 483474 7596 483480 7608
rect 423640 7568 483480 7596
rect 423640 7556 423646 7568
rect 483474 7556 483480 7568
rect 483532 7556 483538 7608
rect 528646 7556 528652 7608
rect 528704 7596 528710 7608
rect 529842 7596 529848 7608
rect 528704 7568 529848 7596
rect 528704 7556 528710 7568
rect 529842 7556 529848 7568
rect 529900 7556 529906 7608
rect 536834 7556 536840 7608
rect 536892 7596 536898 7608
rect 538122 7596 538128 7608
rect 536892 7568 538128 7596
rect 536892 7556 536898 7568
rect 538122 7556 538128 7568
rect 538180 7556 538186 7608
rect 328362 7012 328368 7064
rect 328420 7052 328426 7064
rect 336645 7055 336703 7061
rect 336645 7052 336657 7055
rect 328420 7024 336657 7052
rect 328420 7012 328426 7024
rect 336645 7021 336657 7024
rect 336691 7021 336703 7055
rect 336645 7015 336703 7021
rect 162762 6264 162768 6316
rect 162820 6304 162826 6316
rect 222930 6304 222936 6316
rect 162820 6276 222936 6304
rect 162820 6264 162826 6276
rect 222930 6264 222936 6276
rect 222988 6264 222994 6316
rect 219342 6196 219348 6248
rect 219400 6236 219406 6248
rect 279970 6236 279976 6248
rect 219400 6208 279976 6236
rect 219400 6196 219406 6208
rect 279970 6196 279976 6208
rect 280028 6196 280034 6248
rect 282822 6196 282828 6248
rect 282880 6236 282886 6248
rect 343082 6236 343088 6248
rect 282880 6208 343088 6236
rect 282880 6196 282886 6208
rect 343082 6196 343088 6208
rect 343140 6196 343146 6248
rect 100570 6128 100576 6180
rect 100628 6168 100634 6180
rect 162302 6168 162308 6180
rect 100628 6140 162308 6168
rect 100628 6128 100634 6140
rect 162302 6128 162308 6140
rect 162360 6128 162366 6180
rect 209682 6128 209688 6180
rect 209740 6168 209746 6180
rect 270586 6168 270592 6180
rect 209740 6140 270592 6168
rect 209740 6128 209746 6140
rect 270586 6128 270592 6140
rect 270644 6128 270650 6180
rect 280062 6128 280068 6180
rect 280120 6168 280126 6180
rect 340690 6168 340696 6180
rect 280120 6140 340696 6168
rect 280120 6128 280126 6140
rect 340690 6128 340696 6140
rect 340748 6128 340754 6180
rect 345658 6128 345664 6180
rect 345716 6168 345722 6180
rect 379974 6168 379980 6180
rect 345716 6140 379980 6168
rect 345716 6128 345722 6140
rect 379974 6128 379980 6140
rect 380032 6128 380038 6180
rect 426342 6128 426348 6180
rect 426400 6168 426406 6180
rect 486970 6168 486976 6180
rect 426400 6140 486976 6168
rect 426400 6128 426406 6140
rect 486970 6128 486976 6140
rect 487028 6128 487034 6180
rect 369762 5448 369768 5500
rect 369820 5488 369826 5500
rect 429930 5488 429936 5500
rect 369820 5460 429936 5488
rect 369820 5448 369826 5460
rect 429930 5448 429936 5460
rect 429988 5448 429994 5500
rect 358722 5380 358728 5432
rect 358780 5420 358786 5432
rect 419166 5420 419172 5432
rect 358780 5392 419172 5420
rect 358780 5380 358786 5392
rect 419166 5380 419172 5392
rect 419224 5380 419230 5432
rect 473262 5380 473268 5432
rect 473320 5420 473326 5432
rect 533430 5420 533436 5432
rect 473320 5392 533436 5420
rect 473320 5380 473326 5392
rect 533430 5380 533436 5392
rect 533488 5380 533494 5432
rect 387702 5312 387708 5364
rect 387760 5352 387766 5364
rect 388349 5355 388407 5361
rect 388349 5352 388361 5355
rect 387760 5324 388361 5352
rect 387760 5312 387766 5324
rect 388349 5321 388361 5324
rect 388395 5321 388407 5355
rect 388349 5315 388407 5321
rect 388456 5324 394004 5352
rect 380802 5244 380808 5296
rect 380860 5284 380866 5296
rect 388456 5284 388484 5324
rect 380860 5256 388484 5284
rect 393976 5284 394004 5324
rect 394602 5312 394608 5364
rect 394660 5352 394666 5364
rect 454862 5352 454868 5364
rect 394660 5324 454868 5352
rect 394660 5312 394666 5324
rect 454862 5312 454868 5324
rect 454920 5312 454926 5364
rect 463602 5312 463608 5364
rect 463660 5352 463666 5364
rect 523862 5352 523868 5364
rect 463660 5324 523868 5352
rect 463660 5312 463666 5324
rect 523862 5312 523868 5324
rect 523920 5312 523926 5364
rect 413281 5287 413339 5293
rect 413281 5284 413293 5287
rect 393976 5256 413293 5284
rect 380860 5244 380866 5256
rect 413281 5253 413293 5256
rect 413327 5253 413339 5287
rect 413281 5247 413339 5253
rect 422941 5287 422999 5293
rect 422941 5253 422953 5287
rect 422987 5284 422999 5287
rect 440602 5284 440608 5296
rect 422987 5256 440608 5284
rect 422987 5253 422999 5256
rect 422941 5247 422999 5253
rect 440602 5244 440608 5256
rect 440660 5244 440666 5296
rect 459462 5244 459468 5296
rect 459520 5284 459526 5296
rect 519078 5284 519084 5296
rect 459520 5256 519084 5284
rect 459520 5244 459526 5256
rect 519078 5244 519084 5256
rect 519136 5244 519142 5296
rect 383562 5176 383568 5228
rect 383620 5216 383626 5228
rect 388441 5219 388499 5225
rect 388441 5216 388453 5219
rect 383620 5188 388453 5216
rect 383620 5176 383626 5188
rect 388441 5185 388453 5188
rect 388487 5185 388499 5219
rect 388441 5179 388499 5185
rect 388533 5219 388591 5225
rect 388533 5185 388545 5219
rect 388579 5216 388591 5219
rect 447778 5216 447784 5228
rect 388579 5188 447784 5216
rect 388579 5185 388591 5188
rect 388533 5179 388591 5185
rect 447778 5176 447784 5188
rect 447836 5176 447842 5228
rect 462222 5176 462228 5228
rect 462280 5216 462286 5228
rect 522666 5216 522672 5228
rect 462280 5188 522672 5216
rect 462280 5176 462286 5188
rect 522666 5176 522672 5188
rect 522724 5176 522730 5228
rect 365622 5108 365628 5160
rect 365680 5148 365686 5160
rect 426342 5148 426348 5160
rect 365680 5120 426348 5148
rect 365680 5108 365686 5120
rect 426342 5108 426348 5120
rect 426400 5108 426406 5160
rect 484302 5108 484308 5160
rect 484360 5148 484366 5160
rect 544102 5148 544108 5160
rect 484360 5120 544108 5148
rect 484360 5108 484366 5120
rect 544102 5108 544108 5120
rect 544160 5108 544166 5160
rect 376662 5040 376668 5092
rect 376720 5080 376726 5092
rect 437014 5080 437020 5092
rect 376720 5052 437020 5080
rect 376720 5040 376726 5052
rect 437014 5040 437020 5052
rect 437072 5040 437078 5092
rect 466362 5040 466368 5092
rect 466420 5080 466426 5092
rect 526254 5080 526260 5092
rect 466420 5052 526260 5080
rect 466420 5040 466426 5052
rect 526254 5040 526260 5052
rect 526312 5040 526318 5092
rect 362862 4972 362868 5024
rect 362920 5012 362926 5024
rect 422754 5012 422760 5024
rect 362920 4984 422760 5012
rect 362920 4972 362926 4984
rect 422754 4972 422760 4984
rect 422812 4972 422818 5024
rect 455322 4972 455328 5024
rect 455380 5012 455386 5024
rect 515582 5012 515588 5024
rect 455380 4984 515588 5012
rect 455380 4972 455386 4984
rect 515582 4972 515588 4984
rect 515640 4972 515646 5024
rect 515677 5015 515735 5021
rect 515677 4981 515689 5015
rect 515723 5012 515735 5015
rect 524325 5015 524383 5021
rect 524325 5012 524337 5015
rect 515723 4984 524337 5012
rect 515723 4981 515735 4984
rect 515677 4975 515735 4981
rect 524325 4981 524337 4984
rect 524371 4981 524383 5015
rect 524325 4975 524383 4981
rect 524417 5015 524475 5021
rect 524417 4981 524429 5015
rect 524463 5012 524475 5015
rect 524463 4984 524644 5012
rect 524463 4981 524475 4984
rect 524417 4975 524475 4981
rect 133782 4904 133788 4956
rect 133840 4944 133846 4956
rect 194410 4944 194416 4956
rect 133840 4916 194416 4944
rect 133840 4904 133846 4916
rect 194410 4904 194416 4916
rect 194468 4904 194474 4956
rect 382366 4904 382372 4956
rect 382424 4944 382430 4956
rect 383562 4944 383568 4956
rect 382424 4916 383568 4944
rect 382424 4904 382430 4916
rect 383562 4904 383568 4916
rect 383620 4904 383626 4956
rect 388441 4947 388499 4953
rect 388441 4913 388453 4947
rect 388487 4944 388499 4947
rect 444190 4944 444196 4956
rect 388487 4916 444196 4944
rect 388487 4913 388499 4916
rect 388441 4907 388499 4913
rect 444190 4904 444196 4916
rect 444248 4904 444254 4956
rect 480162 4904 480168 4956
rect 480220 4944 480226 4956
rect 480257 4947 480315 4953
rect 480257 4944 480269 4947
rect 480220 4916 480269 4944
rect 480220 4904 480226 4916
rect 480257 4913 480269 4916
rect 480303 4913 480315 4947
rect 480257 4907 480315 4913
rect 489825 4947 489883 4953
rect 489825 4913 489837 4947
rect 489871 4944 489883 4947
rect 499577 4947 499635 4953
rect 499577 4944 499589 4947
rect 489871 4916 499589 4944
rect 489871 4913 489883 4916
rect 489825 4907 489883 4913
rect 499577 4913 499589 4916
rect 499623 4913 499635 4947
rect 499577 4907 499635 4913
rect 509145 4947 509203 4953
rect 509145 4913 509157 4947
rect 509191 4944 509203 4947
rect 514757 4947 514815 4953
rect 514757 4944 514769 4947
rect 509191 4916 514769 4944
rect 509191 4913 509203 4916
rect 509145 4907 509203 4913
rect 514757 4913 514769 4916
rect 514803 4913 514815 4947
rect 524616 4944 524644 4984
rect 540514 4944 540520 4956
rect 524616 4916 540520 4944
rect 514757 4907 514815 4913
rect 540514 4904 540520 4916
rect 540572 4904 540578 4956
rect 66162 4836 66168 4888
rect 66220 4876 66226 4888
rect 126606 4876 126612 4888
rect 66220 4848 126612 4876
rect 66220 4836 66226 4848
rect 126606 4836 126612 4848
rect 126664 4836 126670 4888
rect 190362 4836 190368 4888
rect 190420 4876 190426 4888
rect 251450 4876 251456 4888
rect 190420 4848 251456 4876
rect 190420 4836 190426 4848
rect 251450 4836 251456 4848
rect 251508 4836 251514 4888
rect 255222 4836 255228 4888
rect 255280 4876 255286 4888
rect 315758 4876 315764 4888
rect 255280 4848 315764 4876
rect 255280 4836 255286 4848
rect 315758 4836 315764 4848
rect 315816 4836 315822 4888
rect 372522 4836 372528 4888
rect 372580 4876 372586 4888
rect 433518 4876 433524 4888
rect 372580 4848 433524 4876
rect 372580 4836 372586 4848
rect 433518 4836 433524 4848
rect 433576 4836 433582 4888
rect 433613 4879 433671 4885
rect 433613 4845 433625 4879
rect 433659 4876 433671 4879
rect 433659 4848 439544 4876
rect 433659 4845 433671 4848
rect 433613 4839 433671 4845
rect 68922 4768 68928 4820
rect 68980 4808 68986 4820
rect 130194 4808 130200 4820
rect 68980 4780 130200 4808
rect 68980 4768 68986 4780
rect 130194 4768 130200 4780
rect 130252 4768 130258 4820
rect 173802 4768 173808 4820
rect 173860 4808 173866 4820
rect 234798 4808 234804 4820
rect 173860 4780 234804 4808
rect 173860 4768 173866 4780
rect 234798 4768 234804 4780
rect 234856 4768 234862 4820
rect 295242 4768 295248 4820
rect 295300 4808 295306 4820
rect 356146 4808 356152 4820
rect 295300 4780 356152 4808
rect 295300 4768 295306 4780
rect 356146 4768 356152 4780
rect 356204 4768 356210 4820
rect 413281 4811 413339 4817
rect 413281 4777 413293 4811
rect 413327 4808 413339 4811
rect 422941 4811 422999 4817
rect 422941 4808 422953 4811
rect 413327 4780 422953 4808
rect 413327 4777 413339 4780
rect 413281 4771 413339 4777
rect 422941 4777 422953 4780
rect 422987 4777 422999 4811
rect 422941 4771 422999 4777
rect 390462 4700 390468 4752
rect 390520 4740 390526 4752
rect 405737 4743 405795 4749
rect 405737 4740 405749 4743
rect 390520 4712 405749 4740
rect 390520 4700 390526 4712
rect 405737 4709 405749 4712
rect 405783 4709 405795 4743
rect 405737 4703 405795 4709
rect 415305 4675 415363 4681
rect 415305 4641 415317 4675
rect 415351 4672 415363 4675
rect 439516 4672 439544 4848
rect 487062 4836 487068 4888
rect 487120 4876 487126 4888
rect 547690 4876 547696 4888
rect 487120 4848 547696 4876
rect 487120 4836 487126 4848
rect 547690 4836 547696 4848
rect 547748 4836 547754 4888
rect 476022 4768 476028 4820
rect 476080 4808 476086 4820
rect 536926 4808 536932 4820
rect 476080 4780 536932 4808
rect 476080 4768 476086 4780
rect 536926 4768 536932 4780
rect 536984 4768 536990 4820
rect 480257 4743 480315 4749
rect 480257 4709 480269 4743
rect 480303 4740 480315 4743
rect 489825 4743 489883 4749
rect 489825 4740 489837 4743
rect 480303 4712 489837 4740
rect 480303 4709 480315 4712
rect 480257 4703 480315 4709
rect 489825 4709 489837 4712
rect 489871 4709 489883 4743
rect 489825 4703 489883 4709
rect 499577 4743 499635 4749
rect 499577 4709 499589 4743
rect 499623 4740 499635 4743
rect 509145 4743 509203 4749
rect 509145 4740 509157 4743
rect 499623 4712 509157 4740
rect 499623 4709 499635 4712
rect 499577 4703 499635 4709
rect 509145 4709 509157 4712
rect 509191 4709 509203 4743
rect 509145 4703 509203 4709
rect 514757 4743 514815 4749
rect 514757 4709 514769 4743
rect 514803 4740 514815 4743
rect 515677 4743 515735 4749
rect 515677 4740 515689 4743
rect 514803 4712 515689 4740
rect 514803 4709 514815 4712
rect 514757 4703 514815 4709
rect 515677 4709 515689 4712
rect 515723 4709 515735 4743
rect 515677 4703 515735 4709
rect 451274 4672 451280 4684
rect 415351 4644 416268 4672
rect 439516 4644 451280 4672
rect 415351 4641 415363 4644
rect 415305 4635 415363 4641
rect 405737 4539 405795 4545
rect 405737 4505 405749 4539
rect 405783 4536 405795 4539
rect 415305 4539 415363 4545
rect 415305 4536 415317 4539
rect 405783 4508 415317 4536
rect 405783 4505 405795 4508
rect 405737 4499 405795 4505
rect 415305 4505 415317 4508
rect 415351 4505 415363 4539
rect 416240 4536 416268 4644
rect 451274 4632 451280 4644
rect 451332 4632 451338 4684
rect 433613 4539 433671 4545
rect 433613 4536 433625 4539
rect 416240 4508 433625 4536
rect 415305 4499 415363 4505
rect 433613 4505 433625 4508
rect 433659 4505 433671 4539
rect 433613 4499 433671 4505
rect 345017 4199 345075 4205
rect 345017 4165 345029 4199
rect 345063 4196 345075 4199
rect 354585 4199 354643 4205
rect 354585 4196 354597 4199
rect 345063 4168 354597 4196
rect 345063 4165 345075 4168
rect 345017 4159 345075 4165
rect 354585 4165 354597 4168
rect 354631 4165 354643 4199
rect 354585 4159 354643 4165
rect 143442 4088 143448 4140
rect 143500 4128 143506 4140
rect 203886 4128 203892 4140
rect 143500 4100 203892 4128
rect 143500 4088 143506 4100
rect 203886 4088 203892 4100
rect 203944 4088 203950 4140
rect 246942 4088 246948 4140
rect 247000 4128 247006 4140
rect 307386 4128 307392 4140
rect 247000 4100 307392 4128
rect 247000 4088 247006 4100
rect 307386 4088 307392 4100
rect 307444 4088 307450 4140
rect 307662 4088 307668 4140
rect 307720 4128 307726 4140
rect 368014 4128 368020 4140
rect 307720 4100 368020 4128
rect 307720 4088 307726 4100
rect 368014 4088 368020 4100
rect 368072 4088 368078 4140
rect 379422 4088 379428 4140
rect 379480 4128 379486 4140
rect 439406 4128 439412 4140
rect 379480 4100 439412 4128
rect 379480 4088 379486 4100
rect 439406 4088 439412 4100
rect 439464 4088 439470 4140
rect 460842 4088 460848 4140
rect 460900 4128 460906 4140
rect 521470 4128 521476 4140
rect 460900 4100 521476 4128
rect 460900 4088 460906 4100
rect 521470 4088 521476 4100
rect 521528 4088 521534 4140
rect 521562 4088 521568 4140
rect 521620 4128 521626 4140
rect 582190 4128 582196 4140
rect 521620 4100 582196 4128
rect 521620 4088 521626 4100
rect 582190 4088 582196 4100
rect 582248 4088 582254 4140
rect 132586 4020 132592 4072
rect 132644 4060 132650 4072
rect 133782 4060 133788 4072
rect 132644 4032 133788 4060
rect 132644 4020 132650 4032
rect 133782 4020 133788 4032
rect 133840 4020 133846 4072
rect 150342 4020 150348 4072
rect 150400 4060 150406 4072
rect 211062 4060 211068 4072
rect 150400 4032 211068 4060
rect 150400 4020 150406 4032
rect 211062 4020 211068 4032
rect 211120 4020 211126 4072
rect 257982 4020 257988 4072
rect 258040 4060 258046 4072
rect 318058 4060 318064 4072
rect 258040 4032 318064 4060
rect 258040 4020 258046 4032
rect 318058 4020 318064 4032
rect 318116 4020 318122 4072
rect 336642 4020 336648 4072
rect 336700 4060 336706 4072
rect 396626 4060 396632 4072
rect 336700 4032 396632 4060
rect 336700 4020 336706 4032
rect 396626 4020 396632 4032
rect 396684 4020 396690 4072
rect 440142 4020 440148 4072
rect 440200 4060 440206 4072
rect 500126 4060 500132 4072
rect 440200 4032 500132 4060
rect 440200 4020 440206 4032
rect 500126 4020 500132 4032
rect 500184 4020 500190 4072
rect 518802 4020 518808 4072
rect 518860 4060 518866 4072
rect 578602 4060 578608 4072
rect 518860 4032 578608 4060
rect 518860 4020 518866 4032
rect 578602 4020 578608 4032
rect 578660 4020 578666 4072
rect 92290 3952 92296 4004
rect 92348 3992 92354 4004
rect 152734 3992 152740 4004
rect 92348 3964 152740 3992
rect 92348 3952 92354 3964
rect 152734 3952 152740 3964
rect 152792 3952 152798 4004
rect 161382 3952 161388 4004
rect 161440 3992 161446 4004
rect 221734 3992 221740 4004
rect 161440 3964 221740 3992
rect 161440 3952 161446 3964
rect 221734 3952 221740 3964
rect 221792 3952 221798 4004
rect 264882 3952 264888 4004
rect 264940 3992 264946 4004
rect 325234 3992 325240 4004
rect 264940 3964 325240 3992
rect 264940 3952 264946 3964
rect 325234 3952 325240 3964
rect 325292 3952 325298 4004
rect 343542 3952 343548 4004
rect 343600 3992 343606 4004
rect 403710 3992 403716 4004
rect 343600 3964 403716 3992
rect 343600 3952 343606 3964
rect 403710 3952 403716 3964
rect 403768 3952 403774 4004
rect 415302 3952 415308 4004
rect 415360 3992 415366 4004
rect 475102 3992 475108 4004
rect 415360 3964 475108 3992
rect 415360 3952 415366 3964
rect 475102 3952 475108 3964
rect 475160 3952 475166 4004
rect 496722 3952 496728 4004
rect 496780 3992 496786 4004
rect 557166 3992 557172 4004
rect 496780 3964 557172 3992
rect 496780 3952 496786 3964
rect 557166 3952 557172 3964
rect 557224 3952 557230 4004
rect 114462 3884 114468 3936
rect 114520 3924 114526 3936
rect 175274 3924 175280 3936
rect 114520 3896 175280 3924
rect 114520 3884 114526 3896
rect 175274 3884 175280 3896
rect 175332 3884 175338 3936
rect 215202 3884 215208 3936
rect 215260 3924 215266 3936
rect 275278 3924 275284 3936
rect 215260 3896 275284 3924
rect 215260 3884 215266 3896
rect 275278 3884 275284 3896
rect 275336 3884 275342 3936
rect 293862 3884 293868 3936
rect 293920 3924 293926 3936
rect 353754 3924 353760 3936
rect 293920 3896 353760 3924
rect 293920 3884 293926 3896
rect 353754 3884 353760 3896
rect 353812 3884 353818 3936
rect 393222 3884 393228 3936
rect 393280 3924 393286 3936
rect 453666 3924 453672 3936
rect 393280 3896 453672 3924
rect 393280 3884 393286 3896
rect 453666 3884 453672 3896
rect 453724 3884 453730 3936
rect 453942 3884 453948 3936
rect 454000 3924 454006 3936
rect 514386 3924 514392 3936
rect 454000 3896 514392 3924
rect 454000 3884 454006 3896
rect 514386 3884 514392 3896
rect 514444 3884 514450 3936
rect 514662 3884 514668 3936
rect 514720 3924 514726 3936
rect 575014 3924 575020 3936
rect 514720 3896 575020 3924
rect 514720 3884 514726 3896
rect 575014 3884 575020 3896
rect 575072 3884 575078 3936
rect 95142 3816 95148 3868
rect 95200 3856 95206 3868
rect 156322 3856 156328 3868
rect 95200 3828 156328 3856
rect 95200 3816 95206 3828
rect 156322 3816 156328 3828
rect 156380 3816 156386 3868
rect 201494 3816 201500 3868
rect 201552 3856 201558 3868
rect 202690 3856 202696 3868
rect 201552 3828 202696 3856
rect 201552 3816 201558 3828
rect 202690 3816 202696 3828
rect 202748 3816 202754 3868
rect 206922 3816 206928 3868
rect 206980 3856 206986 3868
rect 268102 3856 268108 3868
rect 206980 3828 268108 3856
rect 206980 3816 206986 3828
rect 268102 3816 268108 3828
rect 268160 3816 268166 3868
rect 289722 3816 289728 3868
rect 289780 3856 289786 3868
rect 350258 3856 350264 3868
rect 289780 3828 350264 3856
rect 289780 3816 289786 3828
rect 350258 3816 350264 3828
rect 350316 3816 350322 3868
rect 357437 3859 357495 3865
rect 357437 3825 357449 3859
rect 357483 3856 357495 3859
rect 367005 3859 367063 3865
rect 367005 3856 367017 3859
rect 357483 3828 367017 3856
rect 357483 3825 357495 3828
rect 357437 3819 357495 3825
rect 367005 3825 367017 3828
rect 367051 3825 367063 3859
rect 367005 3819 367063 3825
rect 386322 3816 386328 3868
rect 386380 3856 386386 3868
rect 446582 3856 446588 3868
rect 386380 3828 446588 3856
rect 386380 3816 386386 3828
rect 446582 3816 446588 3828
rect 446640 3816 446646 3868
rect 447042 3816 447048 3868
rect 447100 3856 447106 3868
rect 507210 3856 507216 3868
rect 447100 3828 507216 3856
rect 447100 3816 447106 3828
rect 507210 3816 507216 3828
rect 507268 3816 507274 3868
rect 511902 3816 511908 3868
rect 511960 3856 511966 3868
rect 571334 3856 571340 3868
rect 511960 3828 571340 3856
rect 511960 3816 511966 3828
rect 571334 3816 571340 3828
rect 571392 3816 571398 3868
rect 121362 3748 121368 3800
rect 121420 3788 121426 3800
rect 182542 3788 182548 3800
rect 121420 3760 182548 3788
rect 121420 3748 121426 3760
rect 182542 3748 182548 3760
rect 182600 3748 182606 3800
rect 200022 3748 200028 3800
rect 200080 3788 200086 3800
rect 261018 3788 261024 3800
rect 200080 3760 261024 3788
rect 200080 3748 200086 3760
rect 261018 3748 261024 3760
rect 261076 3748 261082 3800
rect 262214 3748 262220 3800
rect 262272 3788 262278 3800
rect 263410 3788 263416 3800
rect 262272 3760 263416 3788
rect 262272 3748 262278 3760
rect 263410 3748 263416 3760
rect 263468 3748 263474 3800
rect 296622 3748 296628 3800
rect 296680 3788 296686 3800
rect 357342 3788 357348 3800
rect 296680 3760 357348 3788
rect 296680 3748 296686 3760
rect 357342 3748 357348 3760
rect 357400 3748 357406 3800
rect 400122 3748 400128 3800
rect 400180 3788 400186 3800
rect 460842 3788 460848 3800
rect 400180 3760 460848 3788
rect 400180 3748 400186 3760
rect 460842 3748 460848 3760
rect 460900 3748 460906 3800
rect 507762 3748 507768 3800
rect 507820 3788 507826 3800
rect 567838 3788 567844 3800
rect 507820 3760 567844 3788
rect 507820 3748 507826 3760
rect 567838 3748 567844 3760
rect 567896 3748 567902 3800
rect 88242 3680 88248 3732
rect 88300 3720 88306 3732
rect 149238 3720 149244 3732
rect 88300 3692 149244 3720
rect 88300 3680 88306 3692
rect 149238 3680 149244 3692
rect 149296 3680 149302 3732
rect 153010 3680 153016 3732
rect 153068 3720 153074 3732
rect 214650 3720 214656 3732
rect 153068 3692 214656 3720
rect 153068 3680 153074 3692
rect 214650 3680 214656 3692
rect 214708 3680 214714 3732
rect 222102 3680 222108 3732
rect 222160 3720 222166 3732
rect 282454 3720 282460 3732
rect 222160 3692 282460 3720
rect 222160 3680 222166 3692
rect 282454 3680 282460 3692
rect 282512 3680 282518 3732
rect 300762 3680 300768 3732
rect 300820 3720 300826 3732
rect 360930 3720 360936 3732
rect 300820 3692 360936 3720
rect 300820 3680 300826 3692
rect 360930 3680 360936 3692
rect 360988 3680 360994 3732
rect 361209 3723 361267 3729
rect 361209 3689 361221 3723
rect 361255 3720 361267 3723
rect 371602 3720 371608 3732
rect 361255 3692 371608 3720
rect 361255 3689 361267 3692
rect 361209 3683 361267 3689
rect 371602 3680 371608 3692
rect 371660 3680 371666 3732
rect 411162 3680 411168 3732
rect 411220 3720 411226 3732
rect 471514 3720 471520 3732
rect 411220 3692 471520 3720
rect 411220 3680 411226 3692
rect 471514 3680 471520 3692
rect 471572 3680 471578 3732
rect 503622 3680 503628 3732
rect 503680 3720 503686 3732
rect 564342 3720 564348 3732
rect 503680 3692 564348 3720
rect 503680 3680 503686 3692
rect 564342 3680 564348 3692
rect 564400 3680 564406 3732
rect 78582 3612 78588 3664
rect 78640 3652 78646 3664
rect 139670 3652 139676 3664
rect 78640 3624 139676 3652
rect 78640 3612 78646 3624
rect 139670 3612 139676 3624
rect 139728 3612 139734 3664
rect 157242 3612 157248 3664
rect 157300 3652 157306 3664
rect 218054 3652 218060 3664
rect 157300 3624 218060 3652
rect 157300 3612 157306 3624
rect 218054 3612 218060 3624
rect 218112 3612 218118 3664
rect 242802 3612 242808 3664
rect 242860 3652 242866 3664
rect 242860 3624 245700 3652
rect 242860 3612 242866 3624
rect 71682 3544 71688 3596
rect 71740 3584 71746 3596
rect 132494 3584 132500 3596
rect 71740 3556 132500 3584
rect 71740 3544 71746 3556
rect 132494 3544 132500 3556
rect 132552 3544 132558 3596
rect 136082 3584 136088 3596
rect 132604 3556 136088 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 63494 3516 63500 3528
rect 1728 3488 63500 3516
rect 1728 3476 1734 3488
rect 63494 3476 63500 3488
rect 63552 3476 63558 3528
rect 74442 3476 74448 3528
rect 74500 3516 74506 3528
rect 132604 3516 132632 3556
rect 136082 3544 136088 3556
rect 136140 3544 136146 3596
rect 150526 3544 150532 3596
rect 150584 3584 150590 3596
rect 151538 3584 151544 3596
rect 150584 3556 151544 3584
rect 150584 3544 150590 3556
rect 151538 3544 151544 3556
rect 151596 3544 151602 3596
rect 164142 3544 164148 3596
rect 164200 3584 164206 3596
rect 225322 3584 225328 3596
rect 164200 3556 225328 3584
rect 164200 3544 164206 3556
rect 225322 3544 225328 3556
rect 225380 3544 225386 3596
rect 236086 3544 236092 3596
rect 236144 3584 236150 3596
rect 237190 3584 237196 3596
rect 236144 3556 237196 3584
rect 236144 3544 236150 3556
rect 237190 3544 237196 3556
rect 237248 3544 237254 3596
rect 244274 3544 244280 3596
rect 244332 3584 244338 3596
rect 245562 3584 245568 3596
rect 244332 3556 245568 3584
rect 244332 3544 244338 3556
rect 245562 3544 245568 3556
rect 245620 3544 245626 3596
rect 245672 3584 245700 3624
rect 249702 3612 249708 3664
rect 249760 3652 249766 3664
rect 310974 3652 310980 3664
rect 249760 3624 310980 3652
rect 249760 3612 249766 3624
rect 310974 3612 310980 3624
rect 311032 3612 311038 3664
rect 336645 3655 336703 3661
rect 311176 3624 314792 3652
rect 303798 3584 303804 3596
rect 245672 3556 303804 3584
rect 303798 3544 303804 3556
rect 303856 3544 303862 3596
rect 310422 3544 310428 3596
rect 310480 3584 310486 3596
rect 311176 3584 311204 3624
rect 310480 3556 311204 3584
rect 310480 3544 310486 3556
rect 314562 3544 314568 3596
rect 314620 3584 314626 3596
rect 314620 3556 314700 3584
rect 314620 3544 314626 3556
rect 74500 3488 132632 3516
rect 74500 3476 74506 3488
rect 140774 3476 140780 3528
rect 140832 3516 140838 3528
rect 142062 3516 142068 3528
rect 140832 3488 142068 3516
rect 140832 3476 140838 3488
rect 142062 3476 142068 3488
rect 142120 3476 142126 3528
rect 171042 3476 171048 3528
rect 171100 3516 171106 3528
rect 232498 3516 232504 3528
rect 171100 3488 232504 3516
rect 171100 3476 171106 3488
rect 232498 3476 232504 3488
rect 232556 3476 232562 3528
rect 235902 3476 235908 3528
rect 235960 3516 235966 3528
rect 296714 3516 296720 3528
rect 235960 3488 296720 3516
rect 235960 3476 235966 3488
rect 296714 3476 296720 3488
rect 296772 3476 296778 3528
rect 304994 3476 305000 3528
rect 305052 3516 305058 3528
rect 306190 3516 306196 3528
rect 305052 3488 306196 3516
rect 305052 3476 305058 3488
rect 306190 3476 306196 3488
rect 306248 3476 306254 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 62114 3448 62120 3460
rect 624 3420 62120 3448
rect 624 3408 630 3420
rect 62114 3408 62120 3420
rect 62172 3408 62178 3460
rect 128262 3408 128268 3460
rect 128320 3448 128326 3460
rect 183465 3451 183523 3457
rect 183465 3448 183477 3451
rect 128320 3420 183477 3448
rect 128320 3408 128326 3420
rect 183465 3417 183477 3420
rect 183511 3417 183523 3451
rect 183465 3411 183523 3417
rect 183554 3408 183560 3460
rect 183612 3448 183618 3460
rect 184842 3448 184848 3460
rect 183612 3420 184848 3448
rect 183612 3408 183618 3420
rect 184842 3408 184848 3420
rect 184900 3408 184906 3460
rect 218146 3408 218152 3460
rect 218204 3448 218210 3460
rect 219342 3448 219348 3460
rect 218204 3420 219348 3448
rect 218204 3408 218210 3420
rect 219342 3408 219348 3420
rect 219400 3408 219406 3460
rect 231762 3408 231768 3460
rect 231820 3448 231826 3460
rect 293126 3448 293132 3460
rect 231820 3420 293132 3448
rect 231820 3408 231826 3420
rect 293126 3408 293132 3420
rect 293184 3408 293190 3460
rect 136542 3340 136548 3392
rect 136600 3380 136606 3392
rect 196802 3380 196808 3392
rect 136600 3352 196808 3380
rect 136600 3340 136606 3352
rect 196802 3340 196808 3352
rect 196860 3340 196866 3392
rect 229002 3340 229008 3392
rect 229060 3380 229066 3392
rect 289538 3380 289544 3392
rect 229060 3352 289544 3380
rect 229060 3340 229066 3352
rect 289538 3340 289544 3352
rect 289596 3340 289602 3392
rect 125502 3272 125508 3324
rect 125560 3312 125566 3324
rect 186038 3312 186044 3324
rect 125560 3284 186044 3312
rect 125560 3272 125566 3284
rect 186038 3272 186044 3284
rect 186096 3272 186102 3324
rect 193122 3272 193128 3324
rect 193180 3312 193186 3324
rect 253842 3312 253848 3324
rect 193180 3284 253848 3312
rect 193180 3272 193186 3284
rect 253842 3272 253848 3284
rect 253900 3272 253906 3324
rect 270494 3272 270500 3324
rect 270552 3312 270558 3324
rect 271690 3312 271696 3324
rect 270552 3284 271696 3312
rect 270552 3272 270558 3284
rect 271690 3272 271696 3284
rect 271748 3272 271754 3324
rect 314672 3312 314700 3556
rect 314764 3516 314792 3624
rect 336645 3621 336657 3655
rect 336691 3652 336703 3655
rect 336829 3655 336887 3661
rect 336691 3624 336780 3652
rect 336691 3621 336703 3624
rect 336645 3615 336703 3621
rect 321646 3544 321652 3596
rect 321704 3584 321710 3596
rect 322842 3584 322848 3596
rect 321704 3556 322848 3584
rect 321704 3544 321710 3556
rect 322842 3544 322848 3556
rect 322900 3544 322906 3596
rect 336752 3593 336780 3624
rect 336829 3621 336841 3655
rect 336875 3652 336887 3655
rect 340785 3655 340843 3661
rect 340785 3652 340797 3655
rect 336875 3624 340797 3652
rect 336875 3621 336887 3624
rect 336829 3615 336887 3621
rect 340785 3621 340797 3624
rect 340831 3621 340843 3655
rect 340785 3615 340843 3621
rect 340877 3655 340935 3661
rect 340877 3621 340889 3655
rect 340923 3652 340935 3655
rect 345017 3655 345075 3661
rect 345017 3652 345029 3655
rect 340923 3624 345029 3652
rect 340923 3621 340935 3624
rect 340877 3615 340935 3621
rect 345017 3621 345029 3624
rect 345063 3621 345075 3655
rect 345017 3615 345075 3621
rect 354585 3655 354643 3661
rect 354585 3621 354597 3655
rect 354631 3652 354643 3655
rect 357437 3655 357495 3661
rect 357437 3652 357449 3655
rect 354631 3624 357449 3652
rect 354631 3621 354643 3624
rect 354585 3615 354643 3621
rect 357437 3621 357449 3624
rect 357483 3621 357495 3655
rect 357437 3615 357495 3621
rect 371142 3612 371148 3664
rect 371200 3652 371206 3664
rect 386233 3655 386291 3661
rect 386233 3652 386245 3655
rect 371200 3624 386245 3652
rect 371200 3612 371206 3624
rect 386233 3621 386245 3624
rect 386279 3621 386291 3655
rect 386233 3615 386291 3621
rect 386325 3655 386383 3661
rect 386325 3621 386337 3655
rect 386371 3652 386383 3655
rect 432322 3652 432328 3664
rect 386371 3624 432328 3652
rect 386371 3621 386383 3624
rect 386325 3615 386383 3621
rect 432322 3612 432328 3624
rect 432380 3612 432386 3664
rect 436002 3612 436008 3664
rect 436060 3652 436066 3664
rect 496538 3652 496544 3664
rect 436060 3624 496544 3652
rect 436060 3612 436066 3624
rect 496538 3612 496544 3624
rect 496596 3612 496602 3664
rect 500862 3612 500868 3664
rect 500920 3652 500926 3664
rect 560754 3652 560760 3664
rect 500920 3624 560760 3652
rect 500920 3612 500926 3624
rect 560754 3612 560760 3624
rect 560812 3612 560818 3664
rect 336737 3587 336795 3593
rect 336737 3553 336749 3587
rect 336783 3553 336795 3587
rect 336737 3547 336795 3553
rect 367005 3587 367063 3593
rect 367005 3553 367017 3587
rect 367051 3584 367063 3587
rect 369949 3587 370007 3593
rect 369949 3584 369961 3587
rect 367051 3556 369961 3584
rect 367051 3553 367063 3556
rect 367005 3547 367063 3553
rect 369949 3553 369961 3556
rect 369995 3553 370007 3587
rect 376757 3587 376815 3593
rect 376757 3584 376769 3587
rect 369949 3547 370007 3553
rect 376680 3556 376769 3584
rect 361209 3519 361267 3525
rect 361209 3516 361221 3519
rect 314764 3488 361221 3516
rect 361209 3485 361221 3488
rect 361255 3485 361267 3519
rect 361209 3479 361267 3485
rect 370041 3519 370099 3525
rect 370041 3485 370053 3519
rect 370087 3516 370099 3519
rect 376680 3516 376708 3556
rect 376757 3553 376769 3556
rect 376803 3553 376815 3587
rect 376757 3547 376815 3553
rect 422202 3544 422208 3596
rect 422260 3584 422266 3596
rect 482278 3584 482284 3596
rect 422260 3556 482284 3584
rect 422260 3544 422266 3556
rect 482278 3544 482284 3556
rect 482336 3544 482342 3596
rect 494146 3544 494152 3596
rect 494204 3584 494210 3596
rect 495342 3584 495348 3596
rect 494204 3556 495348 3584
rect 494204 3544 494210 3556
rect 495342 3544 495348 3556
rect 495400 3544 495406 3596
rect 517422 3544 517428 3596
rect 517480 3584 517486 3596
rect 577406 3584 577412 3596
rect 517480 3556 577412 3584
rect 517480 3544 517486 3556
rect 577406 3544 577412 3556
rect 577464 3544 577470 3596
rect 370087 3488 376708 3516
rect 370087 3485 370099 3488
rect 370041 3479 370099 3485
rect 418062 3476 418068 3528
rect 418120 3516 418126 3528
rect 478690 3516 478696 3528
rect 418120 3488 478696 3516
rect 418120 3476 418126 3488
rect 478690 3476 478696 3488
rect 478748 3476 478754 3528
rect 493962 3476 493968 3528
rect 494020 3516 494026 3528
rect 553578 3516 553584 3528
rect 494020 3488 553584 3516
rect 494020 3476 494026 3488
rect 553578 3476 553584 3488
rect 553636 3476 553642 3528
rect 571426 3476 571432 3528
rect 571484 3516 571490 3528
rect 572622 3516 572628 3528
rect 571484 3488 572628 3516
rect 571484 3476 571490 3488
rect 572622 3476 572628 3488
rect 572680 3476 572686 3528
rect 321462 3408 321468 3460
rect 321520 3448 321526 3460
rect 382274 3448 382280 3460
rect 321520 3420 382280 3448
rect 321520 3408 321526 3420
rect 382274 3408 382280 3420
rect 382332 3408 382338 3460
rect 429102 3408 429108 3460
rect 429160 3448 429166 3460
rect 489362 3448 489368 3460
rect 429160 3420 489368 3448
rect 429160 3408 429166 3420
rect 489362 3408 489368 3420
rect 489420 3408 489426 3460
rect 513282 3408 513288 3460
rect 513340 3448 513346 3460
rect 573818 3448 573824 3460
rect 513340 3420 573824 3448
rect 513340 3408 513346 3420
rect 573818 3408 573824 3420
rect 573876 3408 573882 3460
rect 332502 3340 332508 3392
rect 332560 3380 332566 3392
rect 393038 3380 393044 3392
rect 332560 3352 393044 3380
rect 332560 3340 332566 3352
rect 393038 3340 393044 3352
rect 393096 3340 393102 3392
rect 467834 3340 467840 3392
rect 467892 3380 467898 3392
rect 469122 3380 469128 3392
rect 467892 3352 469128 3380
rect 467892 3340 467898 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 478782 3340 478788 3392
rect 478840 3380 478846 3392
rect 539318 3380 539324 3392
rect 478840 3352 539324 3380
rect 478840 3340 478846 3352
rect 539318 3340 539324 3352
rect 539376 3340 539382 3392
rect 375190 3312 375196 3324
rect 314672 3284 375196 3312
rect 375190 3272 375196 3284
rect 375248 3272 375254 3324
rect 376757 3315 376815 3321
rect 376757 3281 376769 3315
rect 376803 3312 376815 3315
rect 389450 3312 389456 3324
rect 376803 3284 389456 3312
rect 376803 3281 376815 3284
rect 376757 3275 376815 3281
rect 389450 3272 389456 3284
rect 389508 3272 389514 3324
rect 464982 3272 464988 3324
rect 465040 3312 465046 3324
rect 525058 3312 525064 3324
rect 465040 3284 525064 3312
rect 465040 3272 465046 3284
rect 525058 3272 525064 3284
rect 525116 3272 525122 3324
rect 118602 3204 118608 3256
rect 118660 3244 118666 3256
rect 118660 3216 171824 3244
rect 118660 3204 118666 3216
rect 100662 3136 100668 3188
rect 100720 3176 100726 3188
rect 161106 3176 161112 3188
rect 100720 3148 161112 3176
rect 100720 3136 100726 3148
rect 161106 3136 161112 3148
rect 161164 3136 161170 3188
rect 171796 3176 171824 3216
rect 175366 3204 175372 3256
rect 175424 3244 175430 3256
rect 176562 3244 176568 3256
rect 175424 3216 176568 3244
rect 175424 3204 175430 3216
rect 176562 3204 176568 3216
rect 176620 3204 176626 3256
rect 183465 3247 183523 3253
rect 183465 3213 183477 3247
rect 183511 3244 183523 3247
rect 189626 3244 189632 3256
rect 183511 3216 189632 3244
rect 183511 3213 183523 3216
rect 183465 3207 183523 3213
rect 189626 3204 189632 3216
rect 189684 3204 189690 3256
rect 197262 3204 197268 3256
rect 197320 3244 197326 3256
rect 257430 3244 257436 3256
rect 197320 3216 257436 3244
rect 197320 3204 197326 3216
rect 257430 3204 257436 3216
rect 257488 3204 257494 3256
rect 318702 3204 318708 3256
rect 318760 3244 318766 3256
rect 378778 3244 378784 3256
rect 318760 3216 378784 3244
rect 318760 3204 318766 3216
rect 378778 3204 378784 3216
rect 378836 3204 378842 3256
rect 442902 3204 442908 3256
rect 442960 3244 442966 3256
rect 503622 3244 503628 3256
rect 442960 3216 503628 3244
rect 442960 3204 442966 3216
rect 503622 3204 503628 3216
rect 503680 3204 503686 3256
rect 178954 3176 178960 3188
rect 171796 3148 178960 3176
rect 178954 3136 178960 3148
rect 179012 3136 179018 3188
rect 179322 3136 179328 3188
rect 179380 3176 179386 3188
rect 239582 3176 239588 3188
rect 179380 3148 239588 3176
rect 179380 3136 179386 3148
rect 239582 3136 239588 3148
rect 239640 3136 239646 3188
rect 240042 3136 240048 3188
rect 240100 3176 240106 3188
rect 300302 3176 300308 3188
rect 240100 3148 300308 3176
rect 240100 3136 240106 3148
rect 300302 3136 300308 3148
rect 300360 3136 300366 3188
rect 350442 3136 350448 3188
rect 350500 3176 350506 3188
rect 410886 3176 410892 3188
rect 350500 3148 410892 3176
rect 350500 3136 350506 3148
rect 410886 3136 410892 3148
rect 410944 3136 410950 3188
rect 458082 3136 458088 3188
rect 458140 3176 458146 3188
rect 517882 3176 517888 3188
rect 458140 3148 517888 3176
rect 458140 3136 458146 3148
rect 517882 3136 517888 3148
rect 517940 3136 517946 3188
rect 99282 3068 99288 3120
rect 99340 3108 99346 3120
rect 159910 3108 159916 3120
rect 99340 3080 159916 3108
rect 99340 3068 99346 3080
rect 159910 3068 159916 3080
rect 159968 3068 159974 3120
rect 186222 3068 186228 3120
rect 186280 3108 186286 3120
rect 246758 3108 246764 3120
rect 186280 3080 246764 3108
rect 186280 3068 186286 3080
rect 246758 3068 246764 3080
rect 246816 3068 246822 3120
rect 354582 3068 354588 3120
rect 354640 3108 354646 3120
rect 414474 3108 414480 3120
rect 354640 3080 414480 3108
rect 354640 3068 354646 3080
rect 414474 3068 414480 3080
rect 414532 3068 414538 3120
rect 471882 3068 471888 3120
rect 471940 3108 471946 3120
rect 532234 3108 532240 3120
rect 471940 3080 532240 3108
rect 471940 3068 471946 3080
rect 532234 3068 532240 3080
rect 532292 3068 532298 3120
rect 107562 3000 107568 3052
rect 107620 3040 107626 3052
rect 168190 3040 168196 3052
rect 107620 3012 168196 3040
rect 107620 3000 107626 3012
rect 168190 3000 168196 3012
rect 168248 3000 168254 3052
rect 204162 3000 204168 3052
rect 204220 3040 204226 3052
rect 264606 3040 264612 3052
rect 204220 3012 264612 3040
rect 204220 3000 204226 3012
rect 264606 3000 264612 3012
rect 264664 3000 264670 3052
rect 361482 3000 361488 3052
rect 361540 3040 361546 3052
rect 421558 3040 421564 3052
rect 361540 3012 421564 3040
rect 361540 3000 361546 3012
rect 421558 3000 421564 3012
rect 421616 3000 421622 3052
rect 433150 3000 433156 3052
rect 433208 3040 433214 3052
rect 492950 3040 492956 3052
rect 433208 3012 492956 3040
rect 433208 3000 433214 3012
rect 492950 3000 492956 3012
rect 493008 3000 493014 3052
rect 357158 2932 357164 2984
rect 357216 2972 357222 2984
rect 417970 2972 417976 2984
rect 357216 2944 417976 2972
rect 357216 2932 357222 2944
rect 417970 2932 417976 2944
rect 418028 2932 418034 2984
rect 325602 2864 325608 2916
rect 325660 2904 325666 2916
rect 385862 2904 385868 2916
rect 325660 2876 385868 2904
rect 325660 2864 325666 2876
rect 385862 2864 385868 2876
rect 385920 2864 385926 2916
rect 368474 2796 368480 2848
rect 368532 2836 368538 2848
rect 368532 2808 369256 2836
rect 368532 2796 368538 2808
rect 369228 2780 369256 2808
rect 412634 2796 412640 2848
rect 412692 2836 412698 2848
rect 412692 2808 413324 2836
rect 412692 2796 412698 2808
rect 413296 2780 413324 2808
rect 423674 2796 423680 2848
rect 423732 2836 423738 2848
rect 423732 2808 423996 2836
rect 423732 2796 423738 2808
rect 423968 2780 423996 2808
rect 426434 2796 426440 2848
rect 426492 2836 426498 2848
rect 426492 2808 427584 2836
rect 426492 2796 426498 2808
rect 427556 2780 427584 2808
rect 427906 2796 427912 2848
rect 427964 2836 427970 2848
rect 428737 2839 428795 2845
rect 428737 2836 428749 2839
rect 427964 2808 428749 2836
rect 427964 2796 427970 2808
rect 428737 2805 428749 2808
rect 428783 2805 428795 2839
rect 428737 2799 428795 2805
rect 434806 2796 434812 2848
rect 434864 2836 434870 2848
rect 435821 2839 435879 2845
rect 435821 2836 435833 2839
rect 434864 2808 435833 2836
rect 434864 2796 434870 2808
rect 435821 2805 435833 2808
rect 435867 2805 435879 2839
rect 435821 2799 435879 2805
rect 437474 2796 437480 2848
rect 437532 2836 437538 2848
rect 437532 2808 438256 2836
rect 437532 2796 437538 2808
rect 438228 2780 438256 2808
rect 441614 2796 441620 2848
rect 441672 2836 441678 2848
rect 441672 2808 441844 2836
rect 441672 2796 441678 2808
rect 441816 2780 441844 2808
rect 444374 2796 444380 2848
rect 444432 2836 444438 2848
rect 444432 2808 445432 2836
rect 444432 2796 444438 2808
rect 445404 2780 445432 2808
rect 369210 2728 369216 2780
rect 369268 2728 369274 2780
rect 413278 2728 413284 2780
rect 413336 2728 413342 2780
rect 423950 2728 423956 2780
rect 424008 2728 424014 2780
rect 427538 2728 427544 2780
rect 427596 2728 427602 2780
rect 438210 2728 438216 2780
rect 438268 2728 438274 2780
rect 441798 2728 441804 2780
rect 441856 2728 441862 2780
rect 445386 2728 445392 2780
rect 445444 2728 445450 2780
rect 287054 2456 287060 2508
rect 287112 2496 287118 2508
rect 288342 2496 288348 2508
rect 287112 2468 288348 2496
rect 287112 2456 287118 2468
rect 288342 2456 288348 2468
rect 288400 2456 288406 2508
rect 354674 552 354680 604
rect 354732 592 354738 604
rect 354950 592 354956 604
rect 354732 564 354956 592
rect 354732 552 354738 564
rect 354950 552 354956 564
rect 355008 552 355014 604
rect 357434 552 357440 604
rect 357492 592 357498 604
rect 358538 592 358544 604
rect 357492 564 358544 592
rect 357492 552 357498 564
rect 358538 552 358544 564
rect 358596 552 358602 604
rect 358814 552 358820 604
rect 358872 592 358878 604
rect 359734 592 359740 604
rect 358872 564 359740 592
rect 358872 552 358878 564
rect 359734 552 359740 564
rect 359792 552 359798 604
rect 361574 552 361580 604
rect 361632 592 361638 604
rect 362126 592 362132 604
rect 361632 564 362132 592
rect 361632 552 361638 564
rect 362126 552 362132 564
rect 362184 552 362190 604
rect 370406 552 370412 604
rect 370464 592 370470 604
rect 370498 592 370504 604
rect 370464 564 370504 592
rect 370464 552 370470 564
rect 370498 552 370504 564
rect 370556 552 370562 604
rect 372798 552 372804 604
rect 372856 592 372862 604
rect 372890 592 372896 604
rect 372856 564 372896 592
rect 372856 552 372862 564
rect 372890 552 372896 564
rect 372948 552 372954 604
rect 375374 552 375380 604
rect 375432 592 375438 604
rect 376386 592 376392 604
rect 375432 564 376392 592
rect 375432 552 375438 564
rect 376386 552 376392 564
rect 376444 552 376450 604
rect 376754 552 376760 604
rect 376812 592 376818 604
rect 377582 592 377588 604
rect 376812 564 377588 592
rect 376812 552 376818 564
rect 377582 552 377588 564
rect 377640 552 377646 604
rect 383654 552 383660 604
rect 383712 592 383718 604
rect 384666 592 384672 604
rect 383712 564 384672 592
rect 383712 552 383718 564
rect 384666 552 384672 564
rect 384724 552 384730 604
rect 386414 552 386420 604
rect 386472 592 386478 604
rect 387058 592 387064 604
rect 386472 564 387064 592
rect 386472 552 386478 564
rect 387058 552 387064 564
rect 387116 552 387122 604
rect 387794 552 387800 604
rect 387852 592 387858 604
rect 388254 592 388260 604
rect 387852 564 388260 592
rect 387852 552 387858 564
rect 388254 552 388260 564
rect 388312 552 388318 604
rect 397822 552 397828 604
rect 397880 592 397886 604
rect 397914 592 397920 604
rect 397880 564 397920 592
rect 397880 552 397886 564
rect 397914 552 397920 564
rect 397972 552 397978 604
rect 412082 592 412088 604
rect 412043 564 412088 592
rect 412082 552 412088 564
rect 412140 552 412146 604
rect 420362 592 420368 604
rect 420323 564 420368 592
rect 420362 552 420368 564
rect 420420 552 420426 604
rect 428734 592 428740 604
rect 428695 564 428740 592
rect 428734 552 428740 564
rect 428792 552 428798 604
rect 430482 552 430488 604
rect 430540 592 430546 604
rect 431126 592 431132 604
rect 430540 564 431132 592
rect 430540 552 430546 564
rect 431126 552 431132 564
rect 431184 552 431190 604
rect 435818 592 435824 604
rect 435779 564 435824 592
rect 435818 552 435824 564
rect 435876 552 435882 604
rect 450170 552 450176 604
rect 450228 592 450234 604
rect 450354 592 450360 604
rect 450228 564 450360 592
rect 450228 552 450234 564
rect 450354 552 450360 564
rect 450412 552 450418 604
rect 455414 552 455420 604
rect 455472 592 455478 604
rect 456058 592 456064 604
rect 455472 564 456064 592
rect 455472 552 455478 564
rect 456058 552 456064 564
rect 456116 552 456122 604
rect 456886 552 456892 604
rect 456944 592 456950 604
rect 457254 592 457260 604
rect 456944 564 457260 592
rect 456944 552 456950 564
rect 457254 552 457260 564
rect 457312 552 457318 604
rect 471974 552 471980 604
rect 472032 592 472038 604
rect 472710 592 472716 604
rect 472032 564 472716 592
rect 472032 552 472038 564
rect 472710 552 472716 564
rect 472768 552 472774 604
rect 473354 552 473360 604
rect 473412 592 473418 604
rect 473906 592 473912 604
rect 473412 564 473912 592
rect 473412 552 473418 564
rect 473906 552 473912 564
rect 473964 552 473970 604
rect 478874 552 478880 604
rect 478932 592 478938 604
rect 479886 592 479892 604
rect 478932 564 479892 592
rect 478932 552 478938 564
rect 479886 552 479892 564
rect 479944 552 479950 604
rect 516778 592 516784 604
rect 516739 564 516784 592
rect 516778 552 516784 564
rect 516836 552 516842 604
rect 520274 592 520280 604
rect 520235 564 520280 592
rect 520274 552 520280 564
rect 520332 552 520338 604
rect 527266 552 527272 604
rect 527324 592 527330 604
rect 527450 592 527456 604
rect 527324 564 527456 592
rect 527324 552 527330 564
rect 527450 552 527456 564
rect 527508 552 527514 604
rect 579614 552 579620 604
rect 579672 592 579678 604
rect 579798 592 579804 604
rect 579672 564 579804 592
rect 579672 552 579678 564
rect 579798 552 579804 564
rect 579856 552 579862 604
<< via1 >>
rect 411168 700408 411220 700460
rect 429844 700408 429896 700460
rect 463608 700408 463660 700460
rect 494796 700408 494848 700460
rect 514668 700408 514720 700460
rect 559656 700408 559708 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 394608 700340 394660 700392
rect 413652 700340 413704 700392
rect 445668 700340 445720 700392
rect 478512 700340 478564 700392
rect 496728 700340 496780 700392
rect 543464 700340 543516 700392
rect 343548 700272 343600 700324
rect 348792 700272 348844 700324
rect 378048 700272 378100 700324
rect 397460 700272 397512 700324
rect 429108 700272 429160 700324
rect 462320 700272 462372 700324
rect 480168 700272 480220 700324
rect 527180 700272 527232 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 326988 699660 327040 699712
rect 332508 699660 332560 699712
rect 360108 699660 360160 699712
rect 364984 699660 365036 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 523776 696940 523828 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 692724 72752 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 523684 685856 523736 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 683247 72568 683256
rect 72516 683213 72525 683247
rect 72525 683213 72559 683247
rect 72559 683213 72568 683247
rect 72516 683204 72568 683213
rect 72516 683068 72568 683120
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 219072 678988 219124 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 218980 678920 219032 678972
rect 72700 678895 72752 678904
rect 72700 678861 72709 678895
rect 72709 678861 72743 678895
rect 72743 678861 72752 678895
rect 72700 678852 72752 678861
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 72700 669264 72752 669316
rect 72884 669264 72936 669316
rect 218980 669264 219032 669316
rect 219164 669264 219216 669316
rect 72884 666476 72936 666528
rect 219164 666476 219216 666528
rect 72792 656931 72844 656940
rect 72792 656897 72801 656931
rect 72801 656897 72835 656931
rect 72835 656897 72844 656931
rect 72792 656888 72844 656897
rect 219072 656931 219124 656940
rect 219072 656897 219081 656931
rect 219081 656897 219115 656931
rect 219115 656897 219124 656931
rect 219072 656888 219124 656897
rect 377128 655460 377180 655512
rect 378048 655460 378100 655512
rect 428188 655460 428240 655512
rect 429108 655460 429160 655512
rect 462320 655460 462372 655512
rect 463608 655460 463660 655512
rect 479340 655460 479392 655512
rect 480168 655460 480220 655512
rect 513380 655256 513432 655308
rect 514668 655256 514720 655308
rect 325976 655120 326028 655172
rect 326988 655120 327040 655172
rect 72792 654984 72844 655036
rect 121552 654984 121604 655036
rect 137744 654984 137796 655036
rect 172704 654984 172756 655036
rect 41328 654916 41380 654968
rect 104532 654916 104584 654968
rect 154304 654916 154356 654968
rect 189724 654916 189776 654968
rect 219072 654916 219124 654968
rect 240784 654916 240836 654968
rect 24768 654848 24820 654900
rect 87512 654848 87564 654900
rect 106188 654848 106240 654900
rect 155592 654848 155644 654900
rect 202788 654848 202840 654900
rect 223764 654848 223816 654900
rect 8024 654780 8076 654832
rect 70492 654780 70544 654832
rect 89628 654780 89680 654832
rect 138572 654780 138624 654832
rect 171048 654780 171100 654832
rect 206744 654780 206796 654832
rect 235908 654780 235960 654832
rect 257896 654780 257948 654832
rect 267648 654780 267700 654832
rect 274916 654780 274968 654832
rect 284024 654780 284076 654832
rect 291936 654780 291988 654832
rect 300768 654100 300820 654152
rect 308956 654100 309008 654152
rect 3516 645804 3568 645856
rect 59360 645804 59412 645856
rect 523776 638936 523828 638988
rect 580172 638936 580224 638988
rect 3424 630572 3476 630624
rect 59360 630572 59412 630624
rect 524328 619556 524380 619608
rect 580264 619556 580316 619608
rect 3608 616768 3660 616820
rect 59360 616768 59412 616820
rect 523132 605752 523184 605804
rect 580448 605752 580500 605804
rect 3516 603032 3568 603084
rect 59360 603032 59412 603084
rect 523684 592016 523736 592068
rect 579804 592016 579856 592068
rect 3424 587800 3476 587852
rect 59360 587800 59412 587852
rect 524328 579572 524380 579624
rect 580356 579572 580408 579624
rect 3516 573996 3568 574048
rect 59360 573996 59412 574048
rect 523132 565768 523184 565820
rect 580448 565768 580500 565820
rect 3424 560192 3476 560244
rect 59360 560192 59412 560244
rect 523776 556180 523828 556232
rect 580172 556180 580224 556232
rect 523500 545096 523552 545148
rect 580172 545096 580224 545148
rect 3424 545028 3476 545080
rect 59360 545028 59412 545080
rect 523684 539520 523736 539572
rect 580264 539520 580316 539572
rect 3424 531224 3476 531276
rect 59360 531224 59412 531276
rect 3424 516128 3476 516180
rect 59360 516128 59412 516180
rect 523776 509260 523828 509312
rect 580172 509260 580224 509312
rect 3332 500964 3384 501016
rect 59360 500964 59412 501016
rect 523684 499468 523736 499520
rect 580264 499468 580316 499520
rect 523684 498176 523736 498228
rect 580172 498176 580224 498228
rect 3424 487160 3476 487212
rect 59360 487160 59412 487212
rect 3424 473356 3476 473408
rect 59360 473356 59412 473408
rect 523684 462340 523736 462392
rect 580172 462340 580224 462392
rect 524328 459484 524380 459536
rect 580264 459484 580316 459536
rect 3516 458192 3568 458244
rect 59360 458192 59412 458244
rect 523776 451256 523828 451308
rect 580172 451256 580224 451308
rect 3424 444388 3476 444440
rect 59360 444388 59412 444440
rect 523684 438880 523736 438932
rect 580172 438880 580224 438932
rect 3608 429156 3660 429208
rect 59360 429156 59412 429208
rect 3424 415420 3476 415472
rect 59360 415420 59412 415472
rect 523684 415420 523736 415472
rect 580172 415420 580224 415472
rect 523776 404336 523828 404388
rect 580172 404336 580224 404388
rect 3516 401616 3568 401668
rect 59360 401616 59412 401668
rect 523684 391960 523736 392012
rect 580172 391960 580224 392012
rect 3608 372580 3660 372632
rect 59360 372580 59412 372632
rect 524236 368500 524288 368552
rect 580172 368500 580224 368552
rect 3516 358776 3568 358828
rect 59360 358776 59412 358828
rect 523684 357416 523736 357468
rect 580172 357416 580224 357468
rect 523776 345040 523828 345092
rect 580172 345040 580224 345092
rect 3332 338036 3384 338088
rect 60096 338036 60148 338088
rect 3424 329808 3476 329860
rect 59360 329808 59412 329860
rect 524328 322872 524380 322924
rect 580172 322872 580224 322924
rect 3608 316004 3660 316056
rect 59360 316004 59412 316056
rect 524328 311788 524380 311840
rect 580172 311788 580224 311840
rect 524328 298732 524380 298784
rect 580172 298732 580224 298784
rect 3056 295264 3108 295316
rect 60004 295264 60056 295316
rect 3516 287036 3568 287088
rect 59360 287036 59412 287088
rect 523684 275952 523736 276004
rect 580172 275952 580224 276004
rect 3424 273232 3476 273284
rect 59360 273232 59412 273284
rect 523684 264868 523736 264920
rect 580172 264868 580224 264920
rect 3148 252492 3200 252544
rect 60096 252492 60148 252544
rect 523684 252492 523736 252544
rect 579804 252492 579856 252544
rect 3608 244264 3660 244316
rect 59360 244264 59412 244316
rect 3700 229100 3752 229152
rect 59360 229100 59412 229152
rect 523684 229032 523736 229084
rect 580172 229032 580224 229084
rect 523776 217948 523828 218000
rect 580172 217948 580224 218000
rect 3148 208292 3200 208344
rect 60004 208292 60056 208344
rect 523868 205572 523920 205624
rect 579804 205572 579856 205624
rect 3516 201492 3568 201544
rect 59360 201492 59412 201544
rect 3608 186328 3660 186380
rect 59360 186328 59412 186380
rect 523684 182112 523736 182164
rect 580172 182112 580224 182164
rect 523776 171028 523828 171080
rect 580172 171028 580224 171080
rect 3424 165520 3476 165572
rect 60096 165520 60148 165572
rect 3424 158720 3476 158772
rect 59360 158720 59412 158772
rect 523868 158652 523920 158704
rect 579804 158652 579856 158704
rect 3700 143556 3752 143608
rect 59360 143556 59412 143608
rect 523684 135192 523736 135244
rect 580172 135192 580224 135244
rect 523776 124108 523828 124160
rect 580172 124108 580224 124160
rect 2964 122748 3016 122800
rect 60004 122748 60056 122800
rect 3516 115948 3568 116000
rect 59360 115948 59412 116000
rect 523868 111732 523920 111784
rect 579804 111732 579856 111784
rect 3608 100716 3660 100768
rect 59360 100716 59412 100768
rect 523684 88272 523736 88324
rect 580172 88272 580224 88324
rect 3056 79976 3108 80028
rect 60096 79976 60148 80028
rect 523776 77188 523828 77240
rect 580172 77188 580224 77240
rect 3424 73176 3476 73228
rect 59360 73176 59412 73228
rect 523868 64812 523920 64864
rect 579804 64812 579856 64864
rect 3516 57944 3568 57996
rect 59360 57944 59412 57996
rect 81624 49444 81676 49496
rect 142252 49444 142304 49496
rect 167368 49444 167420 49496
rect 227904 49444 227956 49496
rect 110236 49376 110288 49428
rect 171232 49376 171284 49428
rect 403348 49376 403400 49428
rect 463792 49376 463844 49428
rect 138848 49308 138900 49360
rect 200212 49308 200264 49360
rect 210332 49308 210384 49360
rect 270500 49308 270552 49360
rect 396172 49308 396224 49360
rect 456892 49308 456944 49360
rect 95884 49240 95936 49292
rect 157432 49240 157484 49292
rect 174544 49240 174596 49292
rect 236184 49240 236236 49292
rect 253204 49240 253256 49292
rect 313464 49240 313516 49292
rect 367652 49240 367704 49292
rect 427912 49240 427964 49292
rect 131672 49172 131724 49224
rect 193404 49172 193456 49224
rect 217416 49172 217468 49224
rect 278964 49172 279016 49224
rect 374736 49172 374788 49224
rect 434812 49172 434864 49224
rect 482008 49172 482060 49224
rect 542360 49172 542412 49224
rect 103060 49104 103112 49156
rect 164332 49104 164384 49156
rect 181720 49104 181772 49156
rect 242992 49104 243044 49156
rect 260380 49104 260432 49156
rect 321744 49104 321796 49156
rect 346124 49104 346176 49156
rect 407212 49104 407264 49156
rect 474832 49104 474884 49156
rect 535460 49104 535512 49156
rect 88708 49036 88760 49088
rect 150624 49036 150676 49088
rect 188896 49036 188948 49088
rect 249892 49036 249944 49088
rect 267464 49036 267516 49088
rect 328552 49036 328604 49088
rect 344928 49036 344980 49088
rect 351184 49036 351236 49088
rect 389088 49036 389140 49088
rect 449992 49036 450044 49088
rect 489184 49036 489236 49088
rect 549260 49036 549312 49088
rect 67272 48968 67324 49020
rect 128452 48968 128504 49020
rect 145932 48968 145984 49020
rect 207112 48968 207164 49020
rect 224592 48968 224644 49020
rect 285772 48968 285824 49020
rect 318708 48968 318760 49020
rect 345664 48968 345716 49020
rect 354496 48968 354548 49020
rect 367744 48968 367796 49020
rect 381912 48968 381964 49020
rect 443184 48968 443236 49020
rect 467748 48968 467800 49020
rect 528560 48968 528612 49020
rect 379520 48832 379572 48884
rect 380808 48832 380860 48884
rect 66076 48764 66128 48816
rect 66904 48764 66956 48816
rect 70860 48764 70912 48816
rect 71688 48764 71740 48816
rect 72056 48764 72108 48816
rect 73068 48764 73120 48816
rect 73252 48764 73304 48816
rect 74356 48764 74408 48816
rect 89904 48764 89956 48816
rect 91008 48764 91060 48816
rect 91100 48764 91152 48816
rect 92296 48764 92348 48816
rect 97080 48764 97132 48816
rect 97908 48764 97960 48816
rect 98276 48764 98328 48816
rect 99288 48764 99340 48816
rect 99472 48764 99524 48816
rect 100668 48764 100720 48816
rect 105452 48764 105504 48816
rect 106188 48764 106240 48816
rect 106648 48764 106700 48816
rect 107568 48764 107620 48816
rect 107844 48764 107896 48816
rect 108948 48764 109000 48816
rect 109040 48764 109092 48816
rect 110328 48764 110380 48816
rect 113732 48764 113784 48816
rect 114468 48764 114520 48816
rect 114928 48764 114980 48816
rect 115848 48764 115900 48816
rect 116124 48764 116176 48816
rect 117228 48764 117280 48816
rect 117320 48764 117372 48816
rect 118608 48764 118660 48816
rect 124496 48764 124548 48816
rect 125508 48764 125560 48816
rect 132868 48764 132920 48816
rect 133788 48764 133840 48816
rect 134064 48764 134116 48816
rect 135168 48764 135220 48816
rect 135260 48764 135312 48816
rect 136548 48764 136600 48816
rect 141148 48764 141200 48816
rect 142068 48764 142120 48816
rect 142344 48764 142396 48816
rect 143448 48764 143500 48816
rect 143540 48764 143592 48816
rect 144828 48764 144880 48816
rect 149520 48764 149572 48816
rect 150348 48764 150400 48816
rect 150716 48764 150768 48816
rect 151728 48764 151780 48816
rect 159088 48764 159140 48816
rect 160008 48764 160060 48816
rect 160284 48764 160336 48816
rect 161388 48764 161440 48816
rect 161480 48764 161532 48816
rect 162768 48764 162820 48816
rect 166172 48764 166224 48816
rect 166908 48764 166960 48816
rect 168564 48764 168616 48816
rect 169668 48764 169720 48816
rect 169760 48764 169812 48816
rect 170956 48764 171008 48816
rect 175740 48764 175792 48816
rect 176568 48764 176620 48816
rect 178132 48764 178184 48816
rect 179328 48764 179380 48816
rect 185308 48764 185360 48816
rect 186228 48764 186280 48816
rect 187700 48764 187752 48816
rect 188988 48764 189040 48816
rect 193588 48764 193640 48816
rect 194508 48764 194560 48816
rect 194784 48764 194836 48816
rect 195888 48764 195940 48816
rect 203156 48764 203208 48816
rect 204168 48764 204220 48816
rect 204352 48764 204404 48816
rect 205456 48764 205508 48816
rect 211528 48764 211580 48816
rect 212448 48764 212500 48816
rect 212724 48764 212776 48816
rect 213828 48764 213880 48816
rect 213920 48764 213972 48816
rect 215208 48764 215260 48816
rect 218612 48764 218664 48816
rect 219348 48764 219400 48816
rect 219808 48764 219860 48816
rect 220728 48764 220780 48816
rect 221004 48764 221056 48816
rect 222108 48764 222160 48816
rect 222200 48764 222252 48816
rect 223488 48764 223540 48816
rect 228180 48764 228232 48816
rect 229008 48764 229060 48816
rect 229376 48764 229428 48816
rect 230388 48764 230440 48816
rect 237748 48764 237800 48816
rect 238668 48764 238720 48816
rect 238944 48764 238996 48816
rect 240048 48764 240100 48816
rect 240140 48764 240192 48816
rect 241428 48764 241480 48816
rect 246028 48764 246080 48816
rect 246948 48764 247000 48816
rect 247224 48764 247276 48816
rect 248328 48764 248380 48816
rect 248420 48764 248472 48816
rect 249616 48764 249668 48816
rect 254400 48764 254452 48816
rect 255228 48764 255280 48816
rect 255596 48764 255648 48816
rect 256608 48764 256660 48816
rect 256792 48764 256844 48816
rect 257988 48764 258040 48816
rect 263968 48764 264020 48816
rect 264888 48764 264940 48816
rect 265164 48764 265216 48816
rect 266268 48764 266320 48816
rect 266360 48764 266412 48816
rect 267648 48764 267700 48816
rect 272248 48764 272300 48816
rect 273168 48764 273220 48816
rect 273444 48764 273496 48816
rect 274548 48764 274600 48816
rect 274640 48764 274692 48816
rect 275836 48764 275888 48816
rect 280620 48764 280672 48816
rect 281448 48764 281500 48816
rect 281816 48764 281868 48816
rect 282828 48764 282880 48816
rect 283012 48764 283064 48816
rect 284208 48764 284260 48816
rect 291384 48764 291436 48816
rect 292488 48764 292540 48816
rect 292580 48764 292632 48816
rect 293868 48764 293920 48816
rect 299664 48764 299716 48816
rect 300768 48764 300820 48816
rect 300860 48764 300912 48816
rect 302148 48764 302200 48816
rect 306840 48764 306892 48816
rect 307668 48764 307720 48816
rect 309232 48764 309284 48816
rect 310336 48764 310388 48816
rect 323492 48764 323544 48816
rect 324228 48764 324280 48816
rect 324688 48764 324740 48816
rect 325608 48764 325660 48816
rect 325884 48764 325936 48816
rect 326988 48764 327040 48816
rect 327080 48764 327132 48816
rect 328276 48764 328328 48816
rect 333060 48764 333112 48816
rect 333888 48764 333940 48816
rect 334256 48764 334308 48816
rect 335268 48764 335320 48816
rect 335452 48764 335504 48816
rect 336648 48764 336700 48816
rect 342628 48764 342680 48816
rect 343548 48764 343600 48816
rect 343732 48764 343784 48816
rect 344928 48764 344980 48816
rect 350908 48764 350960 48816
rect 351828 48764 351880 48816
rect 352104 48764 352156 48816
rect 353208 48764 353260 48816
rect 353300 48764 353352 48816
rect 354588 48764 354640 48816
rect 359280 48764 359332 48816
rect 360108 48764 360160 48816
rect 360476 48764 360528 48816
rect 361488 48764 361540 48816
rect 361672 48764 361724 48816
rect 362868 48764 362920 48816
rect 377128 48764 377180 48816
rect 378048 48764 378100 48816
rect 378324 48764 378376 48816
rect 379428 48764 379480 48816
rect 380716 48764 380768 48816
rect 381544 48764 381596 48816
rect 386696 48764 386748 48816
rect 387708 48764 387760 48816
rect 387892 48764 387944 48816
rect 389088 48764 389140 48816
rect 394976 48764 395028 48816
rect 395988 48764 396040 48816
rect 404544 48764 404596 48816
rect 405648 48764 405700 48816
rect 411720 48764 411772 48816
rect 412548 48764 412600 48816
rect 412916 48764 412968 48816
rect 413928 48764 413980 48816
rect 414112 48764 414164 48816
rect 415308 48764 415360 48816
rect 420092 48764 420144 48816
rect 420828 48764 420880 48816
rect 421196 48764 421248 48816
rect 422208 48764 422260 48816
rect 428372 48764 428424 48816
rect 429108 48764 429160 48816
rect 429568 48764 429620 48816
rect 430488 48764 430540 48816
rect 430764 48764 430816 48816
rect 431868 48764 431920 48816
rect 431960 48764 432012 48816
rect 433156 48764 433208 48816
rect 437940 48764 437992 48816
rect 438768 48764 438820 48816
rect 439136 48764 439188 48816
rect 440148 48764 440200 48816
rect 440332 48764 440384 48816
rect 441528 48764 441580 48816
rect 446220 48764 446272 48816
rect 447048 48764 447100 48816
rect 447416 48764 447468 48816
rect 448428 48764 448480 48816
rect 448612 48764 448664 48816
rect 449716 48764 449768 48816
rect 455788 48764 455840 48816
rect 456708 48764 456760 48816
rect 456984 48764 457036 48816
rect 458088 48764 458140 48816
rect 458180 48764 458232 48816
rect 459468 48764 459520 48816
rect 464160 48764 464212 48816
rect 464988 48764 465040 48816
rect 465356 48764 465408 48816
rect 466368 48764 466420 48816
rect 466552 48764 466604 48816
rect 467748 48764 467800 48816
rect 472440 48764 472492 48816
rect 473268 48764 473320 48816
rect 473636 48764 473688 48816
rect 474648 48764 474700 48816
rect 480812 48764 480864 48816
rect 481548 48764 481600 48816
rect 483204 48764 483256 48816
rect 484308 48764 484360 48816
rect 484400 48764 484452 48816
rect 485596 48764 485648 48816
rect 490380 48764 490432 48816
rect 491208 48764 491260 48816
rect 491576 48764 491628 48816
rect 492588 48764 492640 48816
rect 492772 48764 492824 48816
rect 493968 48764 494020 48816
rect 498660 48764 498712 48816
rect 499488 48764 499540 48816
rect 499856 48764 499908 48816
rect 500868 48764 500920 48816
rect 508228 48764 508280 48816
rect 509148 48764 509200 48816
rect 509424 48764 509476 48816
rect 510528 48764 510580 48816
rect 516600 48764 516652 48816
rect 517428 48764 517480 48816
rect 517796 48764 517848 48816
rect 518808 48764 518860 48816
rect 518992 48764 519044 48816
rect 520096 48764 520148 48816
rect 64880 48696 64932 48748
rect 66168 48696 66220 48748
rect 123300 48696 123352 48748
rect 124128 48696 124180 48748
rect 157892 48696 157944 48748
rect 158628 48696 158680 48748
rect 271052 48696 271104 48748
rect 272524 48696 272576 48748
rect 315212 48696 315264 48748
rect 315948 48696 316000 48748
rect 385500 48696 385552 48748
rect 386328 48696 386380 48748
rect 125692 48628 125744 48680
rect 126888 48628 126940 48680
rect 186504 48628 186556 48680
rect 187608 48628 187660 48680
rect 230572 48628 230624 48680
rect 231676 48628 231728 48680
rect 308036 48560 308088 48612
rect 309048 48560 309100 48612
rect 368848 48560 368900 48612
rect 369768 48560 369820 48612
rect 375932 48560 375984 48612
rect 376668 48560 376720 48612
rect 195980 48492 196032 48544
rect 197268 48492 197320 48544
rect 405740 48492 405792 48544
rect 406936 48492 406988 48544
rect 510620 48492 510672 48544
rect 511908 48492 511960 48544
rect 82820 48424 82872 48476
rect 84016 48424 84068 48476
rect 176936 48424 176988 48476
rect 177948 48424 178000 48476
rect 290188 48424 290240 48476
rect 291108 48424 291160 48476
rect 298468 48424 298520 48476
rect 299388 48424 299440 48476
rect 317604 48288 317656 48340
rect 318708 48288 318760 48340
rect 422392 48288 422444 48340
rect 423588 48288 423640 48340
rect 151912 47608 151964 47660
rect 212540 47608 212592 47660
rect 262772 47608 262824 47660
rect 322940 47608 322992 47660
rect 84108 47540 84160 47592
rect 144920 47540 144972 47592
rect 205548 47540 205600 47592
rect 266360 47540 266412 47592
rect 316408 47540 316460 47592
rect 376760 47540 376812 47592
rect 433248 47540 433300 47592
rect 494060 47540 494112 47592
rect 501052 47540 501104 47592
rect 561680 47540 561732 47592
rect 407212 46903 407264 46912
rect 407212 46869 407221 46903
rect 407221 46869 407255 46903
rect 407255 46869 407264 46903
rect 407212 46860 407264 46869
rect 443184 46903 443236 46912
rect 443184 46869 443193 46903
rect 443193 46869 443227 46903
rect 443227 46869 443236 46903
rect 443184 46860 443236 46869
rect 449992 46903 450044 46912
rect 449992 46869 450001 46903
rect 450001 46869 450035 46903
rect 450035 46869 450044 46903
rect 449992 46860 450044 46869
rect 535460 46903 535512 46912
rect 535460 46869 535469 46903
rect 535469 46869 535503 46903
rect 535503 46869 535512 46903
rect 535460 46860 535512 46869
rect 201960 46248 202012 46300
rect 262220 46248 262272 46300
rect 312820 46248 312872 46300
rect 374092 46248 374144 46300
rect 80428 46180 80480 46232
rect 140780 46180 140832 46232
rect 148324 46180 148376 46232
rect 209872 46180 209924 46232
rect 259184 46180 259236 46232
rect 320180 46180 320232 46232
rect 369952 46180 370004 46232
rect 430580 46180 430632 46232
rect 451004 46180 451056 46232
rect 512000 46180 512052 46232
rect 515404 46180 515456 46232
rect 575480 46180 575532 46232
rect 256608 44956 256660 45008
rect 316040 44956 316092 45008
rect 198648 44888 198700 44940
rect 259460 44888 259512 44940
rect 77208 44820 77260 44872
rect 138020 44820 138072 44872
rect 144736 44820 144788 44872
rect 205640 44820 205692 44872
rect 310336 44820 310388 44872
rect 369860 44820 369912 44872
rect 415216 44820 415268 44872
rect 476120 44820 476172 44872
rect 493876 44820 493928 44872
rect 554780 44820 554832 44872
rect 195888 43460 195940 43512
rect 255320 43460 255372 43512
rect 302056 43460 302108 43512
rect 362960 43460 363012 43512
rect 409788 43460 409840 43512
rect 469220 43460 469272 43512
rect 74356 43392 74408 43444
rect 133880 43392 133932 43444
rect 142068 43392 142120 43444
rect 201500 43392 201552 43444
rect 249616 43392 249668 43444
rect 309140 43392 309192 43444
rect 362776 43392 362828 43444
rect 423680 43392 423732 43444
rect 511816 43392 511868 43444
rect 571432 43392 571484 43444
rect 135168 42100 135220 42152
rect 194600 42100 194652 42152
rect 245568 42100 245620 42152
rect 305000 42100 305052 42152
rect 360108 42100 360160 42152
rect 419540 42100 419592 42152
rect 70308 42032 70360 42084
rect 131120 42032 131172 42084
rect 191748 42032 191800 42084
rect 252652 42032 252704 42084
rect 299388 42032 299440 42084
rect 358820 42032 358872 42084
rect 406936 42032 406988 42084
rect 466460 42032 466512 42084
rect 520096 42032 520148 42084
rect 579620 42032 579672 42084
rect 523684 41352 523736 41404
rect 580172 41352 580224 41404
rect 188988 40740 189040 40792
rect 248420 40740 248472 40792
rect 292488 40740 292540 40792
rect 351920 40740 351972 40792
rect 402888 40740 402940 40792
rect 462320 40740 462372 40792
rect 131028 40672 131080 40724
rect 191840 40672 191892 40724
rect 241336 40672 241388 40724
rect 302240 40672 302292 40724
rect 349068 40672 349120 40724
rect 408500 40672 408552 40724
rect 424968 40672 425020 40724
rect 485780 40672 485832 40724
rect 288348 39448 288400 39500
rect 347780 39448 347832 39500
rect 184848 39380 184900 39432
rect 244280 39380 244332 39432
rect 342168 39380 342220 39432
rect 401600 39380 401652 39432
rect 126796 39312 126848 39364
rect 187700 39312 187752 39364
rect 238668 39312 238720 39364
rect 298100 39312 298152 39364
rect 398748 39312 398800 39364
rect 459652 39312 459704 39364
rect 477408 39312 477460 39364
rect 536840 39312 536892 39364
rect 369860 38564 369912 38616
rect 369952 38564 370004 38616
rect 124128 37952 124180 38004
rect 183560 37952 183612 38004
rect 234528 37952 234580 38004
rect 295340 37952 295392 38004
rect 338028 37952 338080 38004
rect 420828 37952 420880 38004
rect 480260 37952 480312 38004
rect 180708 37884 180760 37936
rect 241520 37884 241572 37936
rect 284116 37884 284168 37936
rect 345020 37884 345072 37936
rect 395988 37884 396040 37936
rect 455420 37884 455472 37936
rect 485596 37884 485648 37936
rect 545120 37884 545172 37936
rect 398840 37315 398892 37324
rect 398840 37281 398849 37315
rect 398849 37281 398883 37315
rect 398883 37281 398892 37315
rect 398840 37272 398892 37281
rect 407212 37315 407264 37324
rect 407212 37281 407221 37315
rect 407221 37281 407255 37315
rect 407255 37281 407264 37315
rect 407212 37272 407264 37281
rect 443184 37315 443236 37324
rect 443184 37281 443193 37315
rect 443193 37281 443227 37315
rect 443227 37281 443236 37315
rect 443184 37272 443236 37281
rect 449992 37315 450044 37324
rect 449992 37281 450001 37315
rect 450001 37281 450035 37315
rect 450035 37281 450044 37315
rect 449992 37272 450044 37281
rect 535460 37315 535512 37324
rect 535460 37281 535469 37315
rect 535469 37281 535503 37315
rect 535503 37281 535512 37315
rect 535460 37272 535512 37281
rect 177948 36592 178000 36644
rect 237380 36592 237432 36644
rect 281448 36592 281500 36644
rect 340880 36592 340932 36644
rect 391848 36592 391900 36644
rect 451280 36592 451332 36644
rect 119988 36524 120040 36576
rect 180800 36524 180852 36576
rect 231676 36524 231728 36576
rect 291200 36524 291252 36576
rect 335268 36524 335320 36576
rect 394700 36524 394752 36576
rect 459376 36524 459428 36576
rect 520372 36524 520424 36576
rect 3332 35844 3384 35896
rect 60004 35844 60056 35896
rect 117228 35232 117280 35284
rect 176660 35232 176712 35284
rect 227628 35232 227680 35284
rect 287060 35232 287112 35284
rect 331128 35232 331180 35284
rect 390560 35232 390612 35284
rect 170956 35164 171008 35216
rect 230480 35164 230532 35216
rect 277308 35164 277360 35216
rect 338120 35164 338172 35216
rect 389088 35164 389140 35216
rect 448520 35164 448572 35216
rect 456708 35164 456760 35216
rect 274548 33872 274600 33924
rect 333980 33872 334032 33924
rect 113088 33804 113140 33856
rect 173900 33804 173952 33856
rect 223396 33804 223448 33856
rect 284300 33804 284352 33856
rect 166908 33736 166960 33788
rect 227812 33736 227864 33788
rect 328276 33736 328328 33788
rect 387800 33736 387852 33788
rect 441436 33736 441488 33788
rect 502432 33736 502484 33788
rect 110328 32444 110380 32496
rect 169760 32444 169812 32496
rect 220728 32444 220780 32496
rect 280160 32444 280212 32496
rect 324228 32444 324280 32496
rect 383660 32444 383712 32496
rect 162676 32376 162728 32428
rect 223580 32376 223632 32428
rect 270408 32376 270460 32428
rect 331220 32376 331272 32428
rect 384948 32376 385000 32428
rect 444380 32376 444432 32428
rect 449716 32376 449768 32428
rect 509240 32376 509292 32428
rect 510528 32376 510580 32428
rect 569960 32376 570012 32428
rect 160008 31084 160060 31136
rect 219440 31084 219492 31136
rect 267648 31084 267700 31136
rect 327080 31084 327132 31136
rect 378048 31084 378100 31136
rect 437480 31084 437532 31136
rect 106188 31016 106240 31068
rect 167092 31016 167144 31068
rect 216588 31016 216640 31068
rect 277400 31016 277452 31068
rect 320088 31016 320140 31068
rect 380900 31016 380952 31068
rect 445668 31016 445720 31068
rect 505100 31016 505152 31068
rect 506388 31016 506440 31068
rect 565820 31016 565872 31068
rect 523776 30268 523828 30320
rect 580172 30268 580224 30320
rect 213828 29724 213880 29776
rect 273260 29724 273312 29776
rect 155868 29656 155920 29708
rect 216680 29656 216732 29708
rect 306288 29656 306340 29708
rect 365720 29656 365772 29708
rect 102048 29588 102100 29640
rect 162860 29588 162912 29640
rect 252468 29588 252520 29640
rect 313372 29588 313424 29640
rect 367008 29588 367060 29640
rect 426440 29588 426492 29640
rect 438768 29588 438820 29640
rect 498200 29588 498252 29640
rect 407212 29112 407264 29164
rect 407212 28976 407264 29028
rect 516140 29019 516192 29028
rect 516140 28985 516149 29019
rect 516149 28985 516183 29019
rect 516183 28985 516192 29019
rect 516140 28976 516192 28985
rect 272524 28296 272576 28348
rect 331312 28296 331364 28348
rect 97908 28228 97960 28280
rect 158812 28228 158864 28280
rect 165528 28228 165580 28280
rect 226340 28228 226392 28280
rect 244188 28228 244240 28280
rect 305092 28228 305144 28280
rect 322848 28228 322900 28280
rect 382372 28228 382424 28280
rect 434628 28228 434680 28280
rect 494152 28228 494204 28280
rect 495348 28228 495400 28280
rect 554872 28228 554924 28280
rect 369860 27548 369912 27600
rect 370504 27548 370556 27600
rect 398840 27591 398892 27600
rect 398840 27557 398849 27591
rect 398849 27557 398883 27591
rect 398883 27557 398892 27591
rect 398840 27548 398892 27557
rect 407212 27591 407264 27600
rect 407212 27557 407221 27591
rect 407221 27557 407255 27591
rect 407255 27557 407264 27591
rect 407212 27548 407264 27557
rect 443184 27548 443236 27600
rect 449992 27548 450044 27600
rect 450360 27548 450412 27600
rect 535460 27591 535512 27600
rect 535460 27557 535469 27591
rect 535469 27557 535503 27591
rect 535503 27557 535512 27591
rect 535460 27548 535512 27557
rect 275836 26936 275888 26988
rect 335360 26936 335412 26988
rect 431868 26936 431920 26988
rect 491300 26936 491352 26988
rect 93768 26868 93820 26920
rect 154580 26868 154632 26920
rect 158628 26868 158680 26920
rect 218152 26868 218204 26920
rect 237288 26868 237340 26920
rect 296812 26868 296864 26920
rect 311808 26868 311860 26920
rect 372620 26868 372672 26920
rect 373908 26868 373960 26920
rect 433340 26868 433392 26920
rect 492588 26868 492640 26920
rect 552020 26868 552072 26920
rect 353208 25576 353260 25628
rect 412640 25576 412692 25628
rect 91008 25508 91060 25560
rect 150532 25508 150584 25560
rect 154488 25508 154540 25560
rect 215300 25508 215352 25560
rect 226248 25508 226300 25560
rect 287152 25508 287204 25560
rect 293776 25508 293828 25560
rect 354680 25508 354732 25560
rect 427728 25508 427780 25560
rect 487160 25508 487212 25560
rect 488448 25508 488500 25560
rect 547880 25508 547932 25560
rect 278688 24148 278740 24200
rect 339500 24148 339552 24200
rect 86868 24080 86920 24132
rect 147680 24080 147732 24132
rect 151728 24080 151780 24132
rect 211160 24080 211212 24132
rect 215116 24080 215168 24132
rect 276020 24080 276072 24132
rect 286968 24080 287020 24132
rect 347872 24080 347924 24132
rect 351828 24080 351880 24132
rect 411260 24080 411312 24132
rect 423496 24080 423548 24132
rect 484400 24080 484452 24132
rect 499488 24080 499540 24132
rect 558920 24080 558972 24132
rect 275928 22788 275980 22840
rect 336740 22788 336792 22840
rect 344928 22788 344980 22840
rect 404360 22788 404412 22840
rect 84016 22720 84068 22772
rect 143540 22720 143592 22772
rect 147588 22720 147640 22772
rect 208400 22720 208452 22772
rect 212448 22720 212500 22772
rect 271880 22720 271932 22772
rect 285588 22720 285640 22772
rect 346400 22720 346452 22772
rect 419448 22720 419500 22772
rect 478880 22720 478932 22772
rect 79968 21360 80020 21412
rect 140872 21360 140924 21412
rect 144828 21360 144880 21412
rect 204260 21360 204312 21412
rect 205456 21360 205508 21412
rect 264980 21360 265032 21412
rect 269028 21360 269080 21412
rect 329840 21360 329892 21412
rect 336556 21360 336608 21412
rect 397460 21360 397512 21412
rect 412548 21360 412600 21412
rect 471980 21360 472032 21412
rect 474648 21360 474700 21412
rect 534080 21360 534132 21412
rect 75828 19932 75880 19984
rect 136640 19932 136692 19984
rect 140688 19932 140740 19984
rect 201592 19932 201644 19984
rect 208308 19932 208360 19984
rect 269120 19932 269172 19984
rect 273168 19932 273220 19984
rect 332600 19932 332652 19984
rect 333888 19932 333940 19984
rect 393320 19932 393372 19984
rect 408408 19932 408460 19984
rect 467840 19932 467892 19984
rect 470508 19932 470560 19984
rect 529940 19932 529992 19984
rect 333980 19295 334032 19304
rect 333980 19261 333989 19295
rect 333989 19261 334023 19295
rect 334023 19261 334032 19295
rect 333980 19252 334032 19261
rect 345020 19295 345072 19304
rect 345020 19261 345029 19295
rect 345029 19261 345063 19295
rect 345063 19261 345072 19295
rect 345020 19252 345072 19261
rect 372620 19295 372672 19304
rect 372620 19261 372629 19295
rect 372629 19261 372663 19295
rect 372663 19261 372672 19295
rect 372620 19252 372672 19261
rect 394700 19295 394752 19304
rect 394700 19261 394709 19295
rect 394709 19261 394743 19295
rect 394743 19261 394752 19295
rect 394700 19252 394752 19261
rect 397460 19295 397512 19304
rect 397460 19261 397469 19295
rect 397469 19261 397503 19295
rect 397503 19261 397512 19295
rect 397460 19252 397512 19261
rect 515956 19252 516008 19304
rect 516140 19252 516192 19304
rect 73068 18572 73120 18624
rect 132592 18572 132644 18624
rect 136456 18572 136508 18624
rect 197360 18572 197412 18624
rect 201408 18572 201460 18624
rect 262312 18572 262364 18624
rect 266268 18572 266320 18624
rect 325700 18572 325752 18624
rect 329748 18572 329800 18624
rect 390652 18572 390704 18624
rect 405648 18572 405700 18624
rect 465080 18572 465132 18624
rect 467748 18572 467800 18624
rect 527272 18572 527324 18624
rect 523868 17892 523920 17944
rect 580080 17892 580132 17944
rect 401508 17280 401560 17332
rect 460940 17280 460992 17332
rect 129648 17212 129700 17264
rect 190460 17212 190512 17264
rect 197176 17212 197228 17264
rect 258080 17212 258132 17264
rect 262128 17212 262180 17264
rect 321652 17212 321704 17264
rect 326988 17212 327040 17264
rect 386420 17212 386472 17264
rect 452568 17212 452620 17264
rect 512092 17212 512144 17264
rect 126888 15920 126940 15972
rect 186320 15920 186372 15972
rect 315948 15920 316000 15972
rect 375380 15920 375432 15972
rect 66904 15852 66956 15904
rect 126980 15852 127032 15904
rect 194508 15852 194560 15904
rect 253940 15852 253992 15904
rect 257896 15852 257948 15904
rect 318800 15852 318852 15904
rect 397368 15852 397420 15904
rect 458180 15852 458232 15904
rect 469128 15852 469180 15904
rect 528652 15852 528704 15904
rect 248328 14492 248380 14544
rect 307760 14492 307812 14544
rect 355968 14492 356020 14544
rect 416872 14492 416924 14544
rect 448428 14492 448480 14544
rect 507860 14492 507912 14544
rect 122748 14424 122800 14476
rect 183652 14424 183704 14476
rect 187608 14424 187660 14476
rect 247040 14424 247092 14476
rect 304908 14424 304960 14476
rect 365812 14424 365864 14476
rect 413928 14424 413980 14476
rect 473360 14424 473412 14476
rect 509148 14424 509200 14476
rect 568580 14424 568632 14476
rect 309048 13132 309100 13184
rect 368480 13132 368532 13184
rect 118516 13064 118568 13116
rect 179420 13064 179472 13116
rect 183468 13064 183520 13116
rect 244372 13064 244424 13116
rect 251088 13064 251140 13116
rect 311900 13064 311952 13116
rect 381544 13064 381596 13116
rect 441620 13064 441672 13116
rect 444288 13064 444340 13116
rect 503720 13064 503772 13116
rect 505008 13064 505060 13116
rect 564440 13064 564492 13116
rect 336740 12452 336792 12504
rect 338120 12452 338172 12504
rect 346400 12452 346452 12504
rect 331312 12384 331364 12436
rect 332416 12384 332468 12436
rect 332600 12384 332652 12436
rect 333612 12384 333664 12436
rect 335360 12384 335412 12436
rect 335912 12384 335964 12436
rect 337108 12316 337160 12368
rect 340880 12384 340932 12436
rect 341892 12384 341944 12436
rect 338304 12316 338356 12368
rect 351920 12384 351972 12436
rect 352564 12384 352616 12436
rect 393320 12384 393372 12436
rect 394240 12384 394292 12436
rect 401600 12384 401652 12436
rect 402520 12384 402572 12436
rect 404360 12384 404412 12436
rect 404912 12384 404964 12436
rect 448520 12384 448572 12436
rect 448980 12384 449032 12436
rect 529940 12384 529992 12436
rect 531044 12384 531096 12436
rect 534080 12384 534132 12436
rect 534540 12384 534592 12436
rect 542360 12384 542412 12436
rect 542912 12384 542964 12436
rect 346676 12316 346728 12368
rect 407212 12291 407264 12300
rect 407212 12257 407221 12291
rect 407221 12257 407255 12291
rect 407255 12257 407264 12291
rect 407212 12248 407264 12257
rect 351184 11772 351236 11824
rect 406108 11772 406160 11824
rect 441528 11772 441580 11824
rect 500960 11772 501012 11824
rect 115848 11704 115900 11756
rect 175372 11704 175424 11756
rect 179236 11704 179288 11756
rect 240140 11704 240192 11756
rect 241428 11704 241480 11756
rect 300860 11704 300912 11756
rect 302148 11704 302200 11756
rect 361580 11704 361632 11756
rect 416688 11704 416740 11756
rect 477592 11704 477644 11756
rect 502156 11704 502208 11756
rect 563152 11704 563204 11756
rect 176568 10344 176620 10396
rect 236092 10344 236144 10396
rect 298008 10344 298060 10396
rect 357440 10344 357492 10396
rect 111708 10276 111760 10328
rect 172520 10276 172572 10328
rect 233148 10276 233200 10328
rect 293960 10276 294012 10328
rect 303528 10276 303580 10328
rect 364524 10276 364576 10328
rect 367744 10276 367796 10328
rect 415400 10276 415452 10328
rect 437388 10276 437440 10328
rect 496820 10276 496872 10328
rect 498108 10276 498160 10328
rect 557540 10276 557592 10328
rect 334716 9664 334768 9716
rect 345480 9664 345532 9716
rect 372896 9664 372948 9716
rect 395436 9664 395488 9716
rect 397828 9664 397880 9716
rect 399024 9664 399076 9716
rect 443000 9707 443052 9716
rect 443000 9673 443009 9707
rect 443009 9673 443043 9707
rect 443043 9673 443052 9707
rect 443000 9664 443052 9673
rect 535736 9664 535788 9716
rect 411260 9596 411312 9648
rect 419540 9596 419592 9648
rect 516140 9596 516192 9648
rect 520372 9596 520424 9648
rect 230388 8984 230440 9036
rect 290740 8984 290792 9036
rect 291108 8984 291160 9036
rect 351368 8984 351420 9036
rect 108948 8916 109000 8968
rect 169392 8916 169444 8968
rect 172428 8916 172480 8968
rect 233700 8916 233752 8968
rect 347688 8916 347740 8968
rect 408684 8916 408736 8968
rect 430488 8916 430540 8968
rect 490564 8916 490616 8968
rect 491208 8916 491260 8968
rect 551192 8916 551244 8968
rect 104808 7624 104860 7676
rect 165896 7624 165948 7676
rect 169668 7624 169720 7676
rect 230112 7624 230164 7676
rect 340788 7624 340840 7676
rect 401324 7624 401376 7676
rect 433340 7624 433392 7676
rect 434628 7624 434680 7676
rect 451280 7624 451332 7676
rect 452476 7624 452528 7676
rect 481548 7624 481600 7676
rect 541716 7624 541768 7676
rect 137928 7556 137980 7608
rect 199200 7556 199252 7608
rect 223488 7556 223540 7608
rect 283656 7556 283708 7608
rect 284208 7556 284260 7608
rect 344284 7556 344336 7608
rect 347780 7556 347832 7608
rect 349068 7556 349120 7608
rect 365720 7556 365772 7608
rect 366916 7556 366968 7608
rect 390560 7556 390612 7608
rect 391848 7556 391900 7608
rect 408500 7556 408552 7608
rect 409696 7556 409748 7608
rect 423588 7556 423640 7608
rect 483480 7556 483532 7608
rect 528652 7556 528704 7608
rect 529848 7556 529900 7608
rect 536840 7556 536892 7608
rect 538128 7556 538180 7608
rect 328368 7012 328420 7064
rect 162768 6264 162820 6316
rect 222936 6264 222988 6316
rect 219348 6196 219400 6248
rect 279976 6196 280028 6248
rect 282828 6196 282880 6248
rect 343088 6196 343140 6248
rect 100576 6128 100628 6180
rect 162308 6128 162360 6180
rect 209688 6128 209740 6180
rect 270592 6128 270644 6180
rect 280068 6128 280120 6180
rect 340696 6128 340748 6180
rect 345664 6128 345716 6180
rect 379980 6128 380032 6180
rect 426348 6128 426400 6180
rect 486976 6128 487028 6180
rect 369768 5448 369820 5500
rect 429936 5448 429988 5500
rect 358728 5380 358780 5432
rect 419172 5380 419224 5432
rect 473268 5380 473320 5432
rect 533436 5380 533488 5432
rect 387708 5312 387760 5364
rect 380808 5244 380860 5296
rect 394608 5312 394660 5364
rect 454868 5312 454920 5364
rect 463608 5312 463660 5364
rect 523868 5312 523920 5364
rect 440608 5244 440660 5296
rect 459468 5244 459520 5296
rect 519084 5244 519136 5296
rect 383568 5176 383620 5228
rect 447784 5176 447836 5228
rect 462228 5176 462280 5228
rect 522672 5176 522724 5228
rect 365628 5108 365680 5160
rect 426348 5108 426400 5160
rect 484308 5108 484360 5160
rect 544108 5108 544160 5160
rect 376668 5040 376720 5092
rect 437020 5040 437072 5092
rect 466368 5040 466420 5092
rect 526260 5040 526312 5092
rect 362868 4972 362920 5024
rect 422760 4972 422812 5024
rect 455328 4972 455380 5024
rect 515588 4972 515640 5024
rect 133788 4904 133840 4956
rect 194416 4904 194468 4956
rect 382372 4904 382424 4956
rect 383568 4904 383620 4956
rect 444196 4904 444248 4956
rect 480168 4904 480220 4956
rect 540520 4904 540572 4956
rect 66168 4836 66220 4888
rect 126612 4836 126664 4888
rect 190368 4836 190420 4888
rect 251456 4836 251508 4888
rect 255228 4836 255280 4888
rect 315764 4836 315816 4888
rect 372528 4836 372580 4888
rect 433524 4836 433576 4888
rect 68928 4768 68980 4820
rect 130200 4768 130252 4820
rect 173808 4768 173860 4820
rect 234804 4768 234856 4820
rect 295248 4768 295300 4820
rect 356152 4768 356204 4820
rect 390468 4700 390520 4752
rect 487068 4836 487120 4888
rect 547696 4836 547748 4888
rect 476028 4768 476080 4820
rect 536932 4768 536984 4820
rect 451280 4632 451332 4684
rect 143448 4088 143500 4140
rect 203892 4088 203944 4140
rect 246948 4088 247000 4140
rect 307392 4088 307444 4140
rect 307668 4088 307720 4140
rect 368020 4088 368072 4140
rect 379428 4088 379480 4140
rect 439412 4088 439464 4140
rect 460848 4088 460900 4140
rect 521476 4088 521528 4140
rect 521568 4088 521620 4140
rect 582196 4088 582248 4140
rect 132592 4020 132644 4072
rect 133788 4020 133840 4072
rect 150348 4020 150400 4072
rect 211068 4020 211120 4072
rect 257988 4020 258040 4072
rect 318064 4020 318116 4072
rect 336648 4020 336700 4072
rect 396632 4020 396684 4072
rect 440148 4020 440200 4072
rect 500132 4020 500184 4072
rect 518808 4020 518860 4072
rect 578608 4020 578660 4072
rect 92296 3952 92348 4004
rect 152740 3952 152792 4004
rect 161388 3952 161440 4004
rect 221740 3952 221792 4004
rect 264888 3952 264940 4004
rect 325240 3952 325292 4004
rect 343548 3952 343600 4004
rect 403716 3952 403768 4004
rect 415308 3952 415360 4004
rect 475108 3952 475160 4004
rect 496728 3952 496780 4004
rect 557172 3952 557224 4004
rect 114468 3884 114520 3936
rect 175280 3884 175332 3936
rect 215208 3884 215260 3936
rect 275284 3884 275336 3936
rect 293868 3884 293920 3936
rect 353760 3884 353812 3936
rect 393228 3884 393280 3936
rect 453672 3884 453724 3936
rect 453948 3884 454000 3936
rect 514392 3884 514444 3936
rect 514668 3884 514720 3936
rect 575020 3884 575072 3936
rect 95148 3816 95200 3868
rect 156328 3816 156380 3868
rect 201500 3816 201552 3868
rect 202696 3816 202748 3868
rect 206928 3816 206980 3868
rect 268108 3816 268160 3868
rect 289728 3816 289780 3868
rect 350264 3816 350316 3868
rect 386328 3816 386380 3868
rect 446588 3816 446640 3868
rect 447048 3816 447100 3868
rect 507216 3816 507268 3868
rect 511908 3816 511960 3868
rect 571340 3816 571392 3868
rect 121368 3748 121420 3800
rect 182548 3748 182600 3800
rect 200028 3748 200080 3800
rect 261024 3748 261076 3800
rect 262220 3748 262272 3800
rect 263416 3748 263468 3800
rect 296628 3748 296680 3800
rect 357348 3748 357400 3800
rect 400128 3748 400180 3800
rect 460848 3748 460900 3800
rect 507768 3748 507820 3800
rect 567844 3748 567896 3800
rect 88248 3680 88300 3732
rect 149244 3680 149296 3732
rect 153016 3680 153068 3732
rect 214656 3680 214708 3732
rect 222108 3680 222160 3732
rect 282460 3680 282512 3732
rect 300768 3680 300820 3732
rect 360936 3680 360988 3732
rect 371608 3680 371660 3732
rect 411168 3680 411220 3732
rect 471520 3680 471572 3732
rect 503628 3680 503680 3732
rect 564348 3680 564400 3732
rect 78588 3612 78640 3664
rect 139676 3612 139728 3664
rect 157248 3612 157300 3664
rect 218060 3612 218112 3664
rect 242808 3612 242860 3664
rect 71688 3544 71740 3596
rect 132500 3544 132552 3596
rect 1676 3476 1728 3528
rect 63500 3476 63552 3528
rect 74448 3476 74500 3528
rect 136088 3544 136140 3596
rect 150532 3544 150584 3596
rect 151544 3544 151596 3596
rect 164148 3544 164200 3596
rect 225328 3544 225380 3596
rect 236092 3544 236144 3596
rect 237196 3544 237248 3596
rect 244280 3544 244332 3596
rect 245568 3544 245620 3596
rect 249708 3612 249760 3664
rect 310980 3612 311032 3664
rect 303804 3544 303856 3596
rect 310428 3544 310480 3596
rect 314568 3544 314620 3596
rect 140780 3476 140832 3528
rect 142068 3476 142120 3528
rect 171048 3476 171100 3528
rect 232504 3476 232556 3528
rect 235908 3476 235960 3528
rect 296720 3476 296772 3528
rect 305000 3476 305052 3528
rect 306196 3476 306248 3528
rect 572 3408 624 3460
rect 62120 3408 62172 3460
rect 128268 3408 128320 3460
rect 183560 3408 183612 3460
rect 184848 3408 184900 3460
rect 218152 3408 218204 3460
rect 219348 3408 219400 3460
rect 231768 3408 231820 3460
rect 293132 3408 293184 3460
rect 136548 3340 136600 3392
rect 196808 3340 196860 3392
rect 229008 3340 229060 3392
rect 289544 3340 289596 3392
rect 125508 3272 125560 3324
rect 186044 3272 186096 3324
rect 193128 3272 193180 3324
rect 253848 3272 253900 3324
rect 270500 3272 270552 3324
rect 271696 3272 271748 3324
rect 321652 3544 321704 3596
rect 322848 3544 322900 3596
rect 371148 3612 371200 3664
rect 432328 3612 432380 3664
rect 436008 3612 436060 3664
rect 496544 3612 496596 3664
rect 500868 3612 500920 3664
rect 560760 3612 560812 3664
rect 422208 3544 422260 3596
rect 482284 3544 482336 3596
rect 494152 3544 494204 3596
rect 495348 3544 495400 3596
rect 517428 3544 517480 3596
rect 577412 3544 577464 3596
rect 418068 3476 418120 3528
rect 478696 3476 478748 3528
rect 493968 3476 494020 3528
rect 553584 3476 553636 3528
rect 571432 3476 571484 3528
rect 572628 3476 572680 3528
rect 321468 3408 321520 3460
rect 382280 3408 382332 3460
rect 429108 3408 429160 3460
rect 489368 3408 489420 3460
rect 513288 3408 513340 3460
rect 573824 3408 573876 3460
rect 332508 3340 332560 3392
rect 393044 3340 393096 3392
rect 467840 3340 467892 3392
rect 469128 3340 469180 3392
rect 478788 3340 478840 3392
rect 539324 3340 539376 3392
rect 375196 3272 375248 3324
rect 389456 3272 389508 3324
rect 464988 3272 465040 3324
rect 525064 3272 525116 3324
rect 118608 3204 118660 3256
rect 100668 3136 100720 3188
rect 161112 3136 161164 3188
rect 175372 3204 175424 3256
rect 176568 3204 176620 3256
rect 189632 3204 189684 3256
rect 197268 3204 197320 3256
rect 257436 3204 257488 3256
rect 318708 3204 318760 3256
rect 378784 3204 378836 3256
rect 442908 3204 442960 3256
rect 503628 3204 503680 3256
rect 178960 3136 179012 3188
rect 179328 3136 179380 3188
rect 239588 3136 239640 3188
rect 240048 3136 240100 3188
rect 300308 3136 300360 3188
rect 350448 3136 350500 3188
rect 410892 3136 410944 3188
rect 458088 3136 458140 3188
rect 517888 3136 517940 3188
rect 99288 3068 99340 3120
rect 159916 3068 159968 3120
rect 186228 3068 186280 3120
rect 246764 3068 246816 3120
rect 354588 3068 354640 3120
rect 414480 3068 414532 3120
rect 471888 3068 471940 3120
rect 532240 3068 532292 3120
rect 107568 3000 107620 3052
rect 168196 3000 168248 3052
rect 204168 3000 204220 3052
rect 264612 3000 264664 3052
rect 361488 3000 361540 3052
rect 421564 3000 421616 3052
rect 433156 3000 433208 3052
rect 492956 3000 493008 3052
rect 357164 2932 357216 2984
rect 417976 2932 418028 2984
rect 325608 2864 325660 2916
rect 385868 2864 385920 2916
rect 368480 2796 368532 2848
rect 412640 2796 412692 2848
rect 423680 2796 423732 2848
rect 426440 2796 426492 2848
rect 427912 2796 427964 2848
rect 434812 2796 434864 2848
rect 437480 2796 437532 2848
rect 441620 2796 441672 2848
rect 444380 2796 444432 2848
rect 369216 2728 369268 2780
rect 413284 2728 413336 2780
rect 423956 2728 424008 2780
rect 427544 2728 427596 2780
rect 438216 2728 438268 2780
rect 441804 2728 441856 2780
rect 445392 2728 445444 2780
rect 287060 2456 287112 2508
rect 288348 2456 288400 2508
rect 354680 552 354732 604
rect 354956 552 355008 604
rect 357440 552 357492 604
rect 358544 552 358596 604
rect 358820 552 358872 604
rect 359740 552 359792 604
rect 361580 552 361632 604
rect 362132 552 362184 604
rect 370412 552 370464 604
rect 370504 552 370556 604
rect 372804 552 372856 604
rect 372896 552 372948 604
rect 375380 552 375432 604
rect 376392 552 376444 604
rect 376760 552 376812 604
rect 377588 552 377640 604
rect 383660 552 383712 604
rect 384672 552 384724 604
rect 386420 552 386472 604
rect 387064 552 387116 604
rect 387800 552 387852 604
rect 388260 552 388312 604
rect 397828 552 397880 604
rect 397920 552 397972 604
rect 412088 595 412140 604
rect 412088 561 412097 595
rect 412097 561 412131 595
rect 412131 561 412140 595
rect 412088 552 412140 561
rect 420368 595 420420 604
rect 420368 561 420377 595
rect 420377 561 420411 595
rect 420411 561 420420 595
rect 420368 552 420420 561
rect 428740 595 428792 604
rect 428740 561 428749 595
rect 428749 561 428783 595
rect 428783 561 428792 595
rect 428740 552 428792 561
rect 430488 552 430540 604
rect 431132 552 431184 604
rect 435824 595 435876 604
rect 435824 561 435833 595
rect 435833 561 435867 595
rect 435867 561 435876 595
rect 435824 552 435876 561
rect 450176 552 450228 604
rect 450360 552 450412 604
rect 455420 552 455472 604
rect 456064 552 456116 604
rect 456892 552 456944 604
rect 457260 552 457312 604
rect 471980 552 472032 604
rect 472716 552 472768 604
rect 473360 552 473412 604
rect 473912 552 473964 604
rect 478880 552 478932 604
rect 479892 552 479944 604
rect 516784 595 516836 604
rect 516784 561 516793 595
rect 516793 561 516827 595
rect 516827 561 516836 595
rect 516784 552 516836 561
rect 520280 595 520332 604
rect 520280 561 520289 595
rect 520289 561 520323 595
rect 520323 561 520332 595
rect 520280 552 520332 561
rect 527272 552 527324 604
rect 527456 552 527508 604
rect 579620 552 579672 604
rect 579804 552 579856 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3436 630630 3464 667927
rect 3528 645862 3556 682207
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654838 8064 663734
rect 24780 654906 24808 699654
rect 41340 654974 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 692782 72740 698278
rect 72700 692776 72752 692782
rect 72700 692718 72752 692724
rect 72516 683256 72568 683262
rect 72516 683198 72568 683204
rect 72528 683126 72556 683198
rect 72516 683120 72568 683126
rect 72516 683062 72568 683068
rect 72700 678904 72752 678910
rect 72700 678846 72752 678852
rect 72712 669322 72740 678846
rect 72700 669316 72752 669322
rect 72700 669258 72752 669264
rect 72884 669316 72936 669322
rect 72884 669258 72936 669264
rect 72896 666534 72924 669258
rect 72884 666528 72936 666534
rect 72884 666470 72936 666476
rect 72792 656940 72844 656946
rect 72792 656882 72844 656888
rect 72804 655042 72832 656882
rect 72792 655036 72844 655042
rect 72792 654978 72844 654984
rect 41328 654968 41380 654974
rect 41328 654910 41380 654916
rect 24768 654900 24820 654906
rect 24768 654842 24820 654848
rect 87512 654900 87564 654906
rect 87512 654842 87564 654848
rect 8024 654832 8076 654838
rect 8024 654774 8076 654780
rect 70492 654832 70544 654838
rect 70492 654774 70544 654780
rect 3606 653576 3662 653585
rect 3606 653511 3662 653520
rect 3516 645856 3568 645862
rect 3516 645798 3568 645804
rect 3424 630624 3476 630630
rect 3424 630566 3476 630572
rect 3514 624880 3570 624889
rect 3514 624815 3570 624824
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 587858 3464 610399
rect 3528 603090 3556 624815
rect 3620 616826 3648 653511
rect 70504 651916 70532 654774
rect 87524 651916 87552 654842
rect 89640 654838 89668 699654
rect 104532 654968 104584 654974
rect 104532 654910 104584 654916
rect 89628 654832 89680 654838
rect 89628 654774 89680 654780
rect 104544 651916 104572 654910
rect 106200 654906 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 655042 137784 663734
rect 121552 655036 121604 655042
rect 121552 654978 121604 654984
rect 137744 655036 137796 655042
rect 137744 654978 137796 654984
rect 106188 654900 106240 654906
rect 106188 654842 106240 654848
rect 121564 651916 121592 654978
rect 154316 654974 154344 663734
rect 154304 654968 154356 654974
rect 154304 654910 154356 654916
rect 155592 654900 155644 654906
rect 155592 654842 155644 654848
rect 138572 654832 138624 654838
rect 138572 654774 138624 654780
rect 138584 651916 138612 654774
rect 155604 651916 155632 654842
rect 171060 654838 171088 700198
rect 172704 655036 172756 655042
rect 172704 654978 172756 654984
rect 171048 654832 171100 654838
rect 171048 654774 171100 654780
rect 172716 651916 172744 654978
rect 189724 654968 189776 654974
rect 189724 654910 189776 654916
rect 189736 651916 189764 654910
rect 202800 654906 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 679046 219112 685850
rect 219072 679040 219124 679046
rect 219072 678982 219124 678988
rect 218980 678972 219032 678978
rect 218980 678914 219032 678920
rect 218992 669322 219020 678914
rect 218980 669316 219032 669322
rect 218980 669258 219032 669264
rect 219164 669316 219216 669322
rect 219164 669258 219216 669264
rect 219176 666534 219204 669258
rect 219164 666528 219216 666534
rect 219164 666470 219216 666476
rect 219072 656940 219124 656946
rect 219072 656882 219124 656888
rect 219084 654974 219112 656882
rect 219072 654968 219124 654974
rect 219072 654910 219124 654916
rect 202788 654900 202840 654906
rect 202788 654842 202840 654848
rect 223764 654900 223816 654906
rect 223764 654842 223816 654848
rect 206744 654832 206796 654838
rect 206744 654774 206796 654780
rect 206756 651916 206784 654774
rect 223776 651916 223804 654842
rect 235920 654838 235948 699654
rect 240784 654968 240836 654974
rect 240784 654910 240836 654916
rect 235908 654832 235960 654838
rect 235908 654774 235960 654780
rect 240796 651916 240824 654910
rect 267660 654838 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 343548 700324 343600 700330
rect 343548 700266 343600 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 326988 699712 327040 699718
rect 326988 699654 327040 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654838 284064 663734
rect 257896 654832 257948 654838
rect 257896 654774 257948 654780
rect 267648 654832 267700 654838
rect 267648 654774 267700 654780
rect 274916 654832 274968 654838
rect 274916 654774 274968 654780
rect 284024 654832 284076 654838
rect 284024 654774 284076 654780
rect 291936 654832 291988 654838
rect 291936 654774 291988 654780
rect 257908 651916 257936 654774
rect 274928 651916 274956 654774
rect 291948 651916 291976 654774
rect 300780 654158 300808 699654
rect 327000 655178 327028 699654
rect 325976 655172 326028 655178
rect 325976 655114 326028 655120
rect 326988 655172 327040 655178
rect 326988 655114 327040 655120
rect 300768 654152 300820 654158
rect 300768 654094 300820 654100
rect 308956 654152 309008 654158
rect 308956 654094 309008 654100
rect 308968 651916 308996 654094
rect 325988 651916 326016 655114
rect 343560 651794 343588 700266
rect 364996 699718 365024 703520
rect 394608 700392 394660 700398
rect 394608 700334 394660 700340
rect 378048 700324 378100 700330
rect 378048 700266 378100 700272
rect 360108 699712 360160 699718
rect 360108 699654 360160 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 360120 651916 360148 699654
rect 378060 655518 378088 700266
rect 377128 655512 377180 655518
rect 377128 655454 377180 655460
rect 378048 655512 378100 655518
rect 378048 655454 378100 655460
rect 377140 651916 377168 655454
rect 394620 651794 394648 700334
rect 397472 700330 397500 703520
rect 411168 700460 411220 700466
rect 411168 700402 411220 700408
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 411180 651916 411208 700402
rect 413664 700398 413692 703520
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 445668 700392 445720 700398
rect 445668 700334 445720 700340
rect 429108 700324 429160 700330
rect 429108 700266 429160 700272
rect 429120 655518 429148 700266
rect 428188 655512 428240 655518
rect 428188 655454 428240 655460
rect 429108 655512 429160 655518
rect 429108 655454 429160 655460
rect 428200 651916 428228 655454
rect 445680 651930 445708 700334
rect 462332 700330 462360 703520
rect 463608 700460 463660 700466
rect 463608 700402 463660 700408
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 463620 655518 463648 700402
rect 478524 700398 478552 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 514668 700460 514720 700466
rect 514668 700402 514720 700408
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 496728 700392 496780 700398
rect 496728 700334 496780 700340
rect 480168 700324 480220 700330
rect 480168 700266 480220 700272
rect 480180 655518 480208 700266
rect 462320 655512 462372 655518
rect 462320 655454 462372 655460
rect 463608 655512 463660 655518
rect 463608 655454 463660 655460
rect 479340 655512 479392 655518
rect 479340 655454 479392 655460
rect 480168 655512 480220 655518
rect 480168 655454 480220 655460
rect 445326 651902 445708 651930
rect 462332 651916 462360 655454
rect 479352 651916 479380 655454
rect 496740 651930 496768 700334
rect 514680 655314 514708 700402
rect 527192 700330 527220 703520
rect 543476 700398 543504 703520
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 523776 696992 523828 696998
rect 523776 696934 523828 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 523684 685908 523736 685914
rect 523684 685850 523736 685856
rect 513380 655308 513432 655314
rect 513380 655250 513432 655256
rect 514668 655308 514720 655314
rect 514668 655250 514720 655256
rect 496386 651902 496768 651930
rect 513392 651916 513420 655250
rect 343022 651766 343588 651794
rect 394174 651766 394648 651794
rect 59360 645856 59412 645862
rect 59360 645798 59412 645804
rect 59372 644745 59400 645798
rect 59358 644736 59414 644745
rect 59358 644671 59414 644680
rect 523696 631961 523724 685850
rect 523788 645289 523816 696934
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 523774 645280 523830 645289
rect 523774 645215 523830 645224
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 523776 638988 523828 638994
rect 523776 638930 523828 638936
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 523682 631952 523738 631961
rect 523682 631887 523738 631896
rect 59360 630624 59412 630630
rect 59360 630566 59412 630572
rect 59372 630465 59400 630566
rect 59358 630456 59414 630465
rect 59358 630391 59414 630400
rect 3608 616820 3660 616826
rect 3608 616762 3660 616768
rect 59360 616820 59412 616826
rect 59360 616762 59412 616768
rect 59372 616185 59400 616762
rect 59358 616176 59414 616185
rect 59358 616111 59414 616120
rect 523132 605804 523184 605810
rect 523132 605746 523184 605752
rect 523144 605305 523172 605746
rect 523130 605296 523186 605305
rect 523130 605231 523186 605240
rect 3516 603084 3568 603090
rect 3516 603026 3568 603032
rect 59360 603084 59412 603090
rect 59360 603026 59412 603032
rect 59372 601905 59400 603026
rect 59358 601896 59414 601905
rect 59358 601831 59414 601840
rect 3514 596048 3570 596057
rect 3514 595983 3570 595992
rect 3424 587852 3476 587858
rect 3424 587794 3476 587800
rect 3528 574054 3556 595983
rect 523684 592068 523736 592074
rect 523684 592010 523736 592016
rect 59360 587852 59412 587858
rect 59360 587794 59412 587800
rect 59372 587625 59400 587794
rect 59358 587616 59414 587625
rect 59358 587551 59414 587560
rect 3516 574048 3568 574054
rect 3516 573990 3568 573996
rect 59360 574048 59412 574054
rect 59360 573990 59412 573996
rect 59372 573345 59400 573990
rect 59358 573336 59414 573345
rect 59358 573271 59414 573280
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 560250 3464 567287
rect 523132 565820 523184 565826
rect 523132 565762 523184 565768
rect 523144 565321 523172 565762
rect 523130 565312 523186 565321
rect 523130 565247 523186 565256
rect 3424 560244 3476 560250
rect 3424 560186 3476 560192
rect 59360 560244 59412 560250
rect 59360 560186 59412 560192
rect 59372 559065 59400 560186
rect 59358 559056 59414 559065
rect 59358 558991 59414 559000
rect 3422 553072 3478 553081
rect 3422 553007 3478 553016
rect 3436 545086 3464 553007
rect 523696 551993 523724 592010
rect 523788 591977 523816 638930
rect 580276 619614 580304 674591
rect 580446 651128 580502 651137
rect 580446 651063 580502 651072
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 524328 619608 524380 619614
rect 524328 619550 524380 619556
rect 580264 619608 580316 619614
rect 580264 619550 580316 619556
rect 524340 618633 524368 619550
rect 524326 618624 524382 618633
rect 524326 618559 524382 618568
rect 579802 592512 579858 592521
rect 579802 592447 579858 592456
rect 579816 592074 579844 592447
rect 579804 592068 579856 592074
rect 579804 592010 579856 592016
rect 523774 591968 523830 591977
rect 523774 591903 523830 591912
rect 580262 580816 580318 580825
rect 580262 580751 580318 580760
rect 524328 579624 524380 579630
rect 524328 579566 524380 579572
rect 524340 578649 524368 579566
rect 524326 578640 524382 578649
rect 524326 578575 524382 578584
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 523776 556232 523828 556238
rect 523776 556174 523828 556180
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 523682 551984 523738 551993
rect 523682 551919 523738 551928
rect 523500 545148 523552 545154
rect 523500 545090 523552 545096
rect 3424 545080 3476 545086
rect 3424 545022 3476 545028
rect 59360 545080 59412 545086
rect 59360 545022 59412 545028
rect 59372 544785 59400 545022
rect 59358 544776 59414 544785
rect 59358 544711 59414 544720
rect 3422 538656 3478 538665
rect 3422 538591 3478 538600
rect 3436 531282 3464 538591
rect 523512 538234 523540 545090
rect 523684 539572 523736 539578
rect 523684 539514 523736 539520
rect 523696 538665 523724 539514
rect 523682 538656 523738 538665
rect 523682 538591 523738 538600
rect 523512 538206 523724 538234
rect 3424 531276 3476 531282
rect 3424 531218 3476 531224
rect 59360 531276 59412 531282
rect 59360 531218 59412 531224
rect 59372 530505 59400 531218
rect 59358 530496 59414 530505
rect 59358 530431 59414 530440
rect 59358 516216 59414 516225
rect 3424 516180 3476 516186
rect 59358 516151 59360 516160
rect 3424 516122 3476 516128
rect 59412 516151 59414 516160
rect 59360 516122 59412 516128
rect 3436 509969 3464 516122
rect 523696 512009 523724 538206
rect 523788 525337 523816 556174
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580276 539578 580304 580751
rect 580368 579630 580396 627671
rect 580460 605810 580488 651063
rect 580448 605804 580500 605810
rect 580448 605746 580500 605752
rect 580446 604208 580502 604217
rect 580446 604143 580502 604152
rect 580356 579624 580408 579630
rect 580356 579566 580408 579572
rect 580460 565826 580488 604143
rect 580448 565820 580500 565826
rect 580448 565762 580500 565768
rect 580264 539572 580316 539578
rect 580264 539514 580316 539520
rect 580262 533896 580318 533905
rect 580262 533831 580318 533840
rect 523774 525328 523830 525337
rect 523774 525263 523830 525272
rect 523682 512000 523738 512009
rect 523682 511935 523738 511944
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 3422 509960 3478 509969
rect 3422 509895 3478 509904
rect 580184 509318 580212 510303
rect 523776 509312 523828 509318
rect 523776 509254 523828 509260
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 59358 501936 59414 501945
rect 59358 501871 59414 501880
rect 59372 501022 59400 501871
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 59360 501016 59412 501022
rect 59360 500958 59412 500964
rect 3344 495553 3372 500958
rect 523684 499520 523736 499526
rect 523684 499462 523736 499468
rect 523696 498681 523724 499462
rect 523682 498672 523738 498681
rect 523682 498607 523738 498616
rect 523684 498228 523736 498234
rect 523684 498170 523736 498176
rect 3330 495544 3386 495553
rect 3330 495479 3386 495488
rect 59358 487656 59414 487665
rect 59358 487591 59414 487600
rect 59372 487218 59400 487591
rect 3424 487212 3476 487218
rect 3424 487154 3476 487160
rect 59360 487212 59412 487218
rect 59360 487154 59412 487160
rect 3436 481137 3464 487154
rect 3422 481128 3478 481137
rect 3422 481063 3478 481072
rect 3424 473408 3476 473414
rect 59360 473408 59412 473414
rect 3424 473350 3476 473356
rect 59358 473376 59360 473385
rect 59412 473376 59414 473385
rect 3436 452441 3464 473350
rect 59358 473311 59414 473320
rect 523696 472025 523724 498170
rect 523788 485353 523816 509254
rect 580276 499526 580304 533831
rect 580264 499520 580316 499526
rect 580264 499462 580316 499468
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580262 486840 580318 486849
rect 580262 486775 580318 486784
rect 523774 485344 523830 485353
rect 523774 485279 523830 485288
rect 523682 472016 523738 472025
rect 523682 471951 523738 471960
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 523684 462392 523736 462398
rect 523684 462334 523736 462340
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 59358 459096 59414 459105
rect 59358 459031 59414 459040
rect 59372 458250 59400 459031
rect 3516 458244 3568 458250
rect 3516 458186 3568 458192
rect 59360 458244 59412 458250
rect 59360 458186 59412 458192
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 3424 444440 3476 444446
rect 3424 444382 3476 444388
rect 3436 423745 3464 444382
rect 3528 438025 3556 458186
rect 523696 445369 523724 462334
rect 580276 459542 580304 486775
rect 524328 459536 524380 459542
rect 524328 459478 524380 459484
rect 580264 459536 580316 459542
rect 580264 459478 580316 459484
rect 524340 458697 524368 459478
rect 524326 458688 524382 458697
rect 524326 458623 524382 458632
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 523776 451308 523828 451314
rect 523776 451250 523828 451256
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 523682 445360 523738 445369
rect 523682 445295 523738 445304
rect 59358 444816 59414 444825
rect 59358 444751 59414 444760
rect 59372 444446 59400 444751
rect 59360 444440 59412 444446
rect 59360 444382 59412 444388
rect 523684 438932 523736 438938
rect 523684 438874 523736 438880
rect 3514 438016 3570 438025
rect 3514 437951 3570 437960
rect 59358 430536 59414 430545
rect 59358 430471 59414 430480
rect 59372 429214 59400 430471
rect 3608 429208 3660 429214
rect 3608 429150 3660 429156
rect 59360 429208 59412 429214
rect 59360 429150 59412 429156
rect 3422 423736 3478 423745
rect 3422 423671 3478 423680
rect 3424 415472 3476 415478
rect 3424 415414 3476 415420
rect 3436 380633 3464 415414
rect 3516 401668 3568 401674
rect 3516 401610 3568 401616
rect 3422 380624 3478 380633
rect 3422 380559 3478 380568
rect 3528 366217 3556 401610
rect 3620 395049 3648 429150
rect 523696 418713 523724 438874
rect 523788 432041 523816 451250
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 523774 432032 523830 432041
rect 523774 431967 523830 431976
rect 523682 418704 523738 418713
rect 523682 418639 523738 418648
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 59358 416256 59414 416265
rect 59358 416191 59414 416200
rect 59372 415478 59400 416191
rect 580184 415478 580212 416463
rect 59360 415472 59412 415478
rect 59360 415414 59412 415420
rect 523684 415472 523736 415478
rect 523684 415414 523736 415420
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 523696 405385 523724 415414
rect 523682 405376 523738 405385
rect 523682 405311 523738 405320
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 523776 404388 523828 404394
rect 523776 404330 523828 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 59358 401976 59414 401985
rect 59358 401911 59414 401920
rect 59372 401674 59400 401911
rect 59360 401668 59412 401674
rect 59360 401610 59412 401616
rect 3606 395040 3662 395049
rect 3606 394975 3662 394984
rect 523788 392057 523816 404330
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 523774 392048 523830 392057
rect 523684 392012 523736 392018
rect 580184 392018 580212 392935
rect 523774 391983 523830 391992
rect 580172 392012 580224 392018
rect 523684 391954 523736 391960
rect 580172 391954 580224 391960
rect 60094 387696 60150 387705
rect 60094 387631 60150 387640
rect 59358 373416 59414 373425
rect 59358 373351 59414 373360
rect 59372 372638 59400 373351
rect 3608 372632 3660 372638
rect 3608 372574 3660 372580
rect 59360 372632 59412 372638
rect 59360 372574 59412 372580
rect 3514 366208 3570 366217
rect 3514 366143 3570 366152
rect 3516 358828 3568 358834
rect 3516 358770 3568 358776
rect 3332 338088 3384 338094
rect 3332 338030 3384 338036
rect 3344 337521 3372 338030
rect 3330 337512 3386 337521
rect 3330 337447 3386 337456
rect 3424 329860 3476 329866
rect 3424 329802 3476 329808
rect 3056 295316 3108 295322
rect 3056 295258 3108 295264
rect 3068 294409 3096 295258
rect 3054 294400 3110 294409
rect 3054 294335 3110 294344
rect 3436 280129 3464 329802
rect 3528 308825 3556 358770
rect 3620 323105 3648 372574
rect 59358 359136 59414 359145
rect 59358 359071 59414 359080
rect 59372 358834 59400 359071
rect 59360 358828 59412 358834
rect 59360 358770 59412 358776
rect 60002 344720 60058 344729
rect 60002 344655 60058 344664
rect 59358 330440 59414 330449
rect 59358 330375 59414 330384
rect 59372 329866 59400 330375
rect 59360 329860 59412 329866
rect 59360 329802 59412 329808
rect 3606 323096 3662 323105
rect 3606 323031 3662 323040
rect 59358 316160 59414 316169
rect 59358 316095 59414 316104
rect 59372 316062 59400 316095
rect 3608 316056 3660 316062
rect 3608 315998 3660 316004
rect 59360 316056 59412 316062
rect 59360 315998 59412 316004
rect 3514 308816 3570 308825
rect 3514 308751 3570 308760
rect 3516 287088 3568 287094
rect 3516 287030 3568 287036
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 3424 273284 3476 273290
rect 3424 273226 3476 273232
rect 3148 252544 3200 252550
rect 3148 252486 3200 252492
rect 3160 251297 3188 252486
rect 3146 251288 3202 251297
rect 3146 251223 3202 251232
rect 3436 222601 3464 273226
rect 3528 237017 3556 287030
rect 3620 265713 3648 315998
rect 60016 295322 60044 344655
rect 60108 338094 60136 387631
rect 523696 378729 523724 391954
rect 523682 378720 523738 378729
rect 523682 378655 523738 378664
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 524236 368552 524288 368558
rect 524236 368494 524288 368500
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 524248 365401 524276 368494
rect 524234 365392 524290 365401
rect 524234 365327 524290 365336
rect 580170 357912 580226 357921
rect 580170 357847 580226 357856
rect 580184 357474 580212 357847
rect 523684 357468 523736 357474
rect 523684 357410 523736 357416
rect 580172 357468 580224 357474
rect 580172 357410 580224 357416
rect 523696 351937 523724 357410
rect 523682 351928 523738 351937
rect 523682 351863 523738 351872
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345098 580212 346015
rect 523776 345092 523828 345098
rect 523776 345034 523828 345040
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 523788 338609 523816 345034
rect 523774 338600 523830 338609
rect 523774 338535 523830 338544
rect 60096 338088 60148 338094
rect 60096 338030 60148 338036
rect 524326 325272 524382 325281
rect 524326 325207 524382 325216
rect 524340 322930 524368 325207
rect 524328 322924 524380 322930
rect 524328 322866 524380 322872
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 524326 311944 524382 311953
rect 524326 311879 524382 311888
rect 524340 311846 524368 311879
rect 524328 311840 524380 311846
rect 524328 311782 524380 311788
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 60094 301880 60150 301889
rect 60094 301815 60150 301824
rect 60004 295316 60056 295322
rect 60004 295258 60056 295264
rect 59358 287600 59414 287609
rect 59358 287535 59414 287544
rect 59372 287094 59400 287535
rect 59360 287088 59412 287094
rect 59360 287030 59412 287036
rect 59358 273320 59414 273329
rect 59358 273255 59360 273264
rect 59412 273255 59414 273264
rect 59360 273226 59412 273232
rect 3606 265704 3662 265713
rect 3606 265639 3662 265648
rect 60002 259040 60058 259049
rect 60002 258975 60058 258984
rect 59358 244760 59414 244769
rect 59358 244695 59414 244704
rect 59372 244322 59400 244695
rect 3608 244316 3660 244322
rect 3608 244258 3660 244264
rect 59360 244316 59412 244322
rect 59360 244258 59412 244264
rect 3514 237008 3570 237017
rect 3514 236943 3570 236952
rect 3422 222592 3478 222601
rect 3422 222527 3478 222536
rect 3148 208344 3200 208350
rect 3148 208286 3200 208292
rect 3160 208185 3188 208286
rect 3146 208176 3202 208185
rect 3146 208111 3202 208120
rect 3516 201544 3568 201550
rect 3516 201486 3568 201492
rect 3424 165572 3476 165578
rect 3424 165514 3476 165520
rect 3436 165073 3464 165514
rect 3422 165064 3478 165073
rect 3422 164999 3478 165008
rect 3424 158772 3476 158778
rect 3424 158714 3476 158720
rect 2964 122800 3016 122806
rect 2964 122742 3016 122748
rect 2976 122097 3004 122742
rect 2962 122088 3018 122097
rect 2962 122023 3018 122032
rect 3436 107681 3464 158714
rect 3528 150793 3556 201486
rect 3620 193905 3648 244258
rect 59358 230480 59414 230489
rect 59358 230415 59414 230424
rect 59372 229158 59400 230415
rect 3700 229152 3752 229158
rect 3700 229094 3752 229100
rect 59360 229152 59412 229158
rect 59360 229094 59412 229100
rect 3606 193896 3662 193905
rect 3606 193831 3662 193840
rect 3608 186380 3660 186386
rect 3608 186322 3660 186328
rect 3514 150784 3570 150793
rect 3514 150719 3570 150728
rect 3620 136377 3648 186322
rect 3712 179489 3740 229094
rect 60016 208350 60044 258975
rect 60108 252550 60136 301815
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580184 298790 580212 299095
rect 524328 298784 524380 298790
rect 524328 298726 524380 298732
rect 580172 298784 580224 298790
rect 580172 298726 580224 298732
rect 524340 298625 524368 298726
rect 524326 298616 524382 298625
rect 524326 298551 524382 298560
rect 523682 285288 523738 285297
rect 523682 285223 523738 285232
rect 523696 276010 523724 285223
rect 523684 276004 523736 276010
rect 523684 275946 523736 275952
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 523682 271960 523738 271969
rect 523682 271895 523738 271904
rect 523696 264926 523724 271895
rect 523684 264920 523736 264926
rect 523684 264862 523736 264868
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 523682 258632 523738 258641
rect 523682 258567 523738 258576
rect 523696 252550 523724 258567
rect 60096 252544 60148 252550
rect 60096 252486 60148 252492
rect 523684 252544 523736 252550
rect 523684 252486 523736 252492
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 523682 245304 523738 245313
rect 523682 245239 523738 245248
rect 523696 229090 523724 245239
rect 523774 231976 523830 231985
rect 523774 231911 523830 231920
rect 523684 229084 523736 229090
rect 523684 229026 523736 229032
rect 523788 218006 523816 231911
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 523866 218648 523922 218657
rect 523866 218583 523922 218592
rect 523776 218000 523828 218006
rect 523776 217942 523828 217948
rect 60094 216200 60150 216209
rect 60094 216135 60150 216144
rect 60004 208344 60056 208350
rect 60004 208286 60056 208292
rect 59358 201920 59414 201929
rect 59358 201855 59414 201864
rect 59372 201550 59400 201855
rect 59360 201544 59412 201550
rect 59360 201486 59412 201492
rect 59358 187640 59414 187649
rect 59358 187575 59414 187584
rect 59372 186386 59400 187575
rect 59360 186380 59412 186386
rect 59360 186322 59412 186328
rect 3698 179480 3754 179489
rect 3698 179415 3754 179424
rect 60002 173360 60058 173369
rect 60002 173295 60058 173304
rect 59358 159080 59414 159089
rect 59358 159015 59414 159024
rect 59372 158778 59400 159015
rect 59360 158772 59412 158778
rect 59360 158714 59412 158720
rect 59358 144800 59414 144809
rect 59358 144735 59414 144744
rect 59372 143614 59400 144735
rect 3700 143608 3752 143614
rect 3700 143550 3752 143556
rect 59360 143608 59412 143614
rect 59360 143550 59412 143556
rect 3606 136368 3662 136377
rect 3606 136303 3662 136312
rect 3516 116000 3568 116006
rect 3516 115942 3568 115948
rect 3422 107672 3478 107681
rect 3422 107607 3478 107616
rect 3056 80028 3108 80034
rect 3056 79970 3108 79976
rect 3068 78985 3096 79970
rect 3054 78976 3110 78985
rect 3054 78911 3110 78920
rect 3424 73228 3476 73234
rect 3424 73170 3476 73176
rect 3332 35896 3384 35902
rect 3330 35864 3332 35873
rect 3384 35864 3386 35873
rect 3330 35799 3386 35808
rect 3436 21457 3464 73170
rect 3528 64569 3556 115942
rect 3608 100768 3660 100774
rect 3608 100710 3660 100716
rect 3514 64560 3570 64569
rect 3514 64495 3570 64504
rect 3516 57996 3568 58002
rect 3516 57938 3568 57944
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3528 7177 3556 57938
rect 3620 50153 3648 100710
rect 3712 93265 3740 143550
rect 60016 122806 60044 173295
rect 60108 165578 60136 216135
rect 523880 205630 523908 218583
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 523868 205624 523920 205630
rect 523868 205566 523920 205572
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 523682 205320 523738 205329
rect 523682 205255 523738 205264
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 523696 182170 523724 205255
rect 523774 191992 523830 192001
rect 523774 191927 523830 191936
rect 523684 182164 523736 182170
rect 523684 182106 523736 182112
rect 523788 171086 523816 191927
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 523866 178664 523922 178673
rect 523866 178599 523922 178608
rect 523776 171080 523828 171086
rect 523776 171022 523828 171028
rect 60096 165572 60148 165578
rect 60096 165514 60148 165520
rect 523682 165336 523738 165345
rect 523682 165271 523738 165280
rect 523696 135250 523724 165271
rect 523880 158710 523908 178599
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 523868 158704 523920 158710
rect 523868 158646 523920 158652
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 523774 152008 523830 152017
rect 523774 151943 523830 151952
rect 523684 135244 523736 135250
rect 523684 135186 523736 135192
rect 60094 130520 60150 130529
rect 60094 130455 60150 130464
rect 60004 122800 60056 122806
rect 60004 122742 60056 122748
rect 59358 116240 59414 116249
rect 59358 116175 59414 116184
rect 59372 116006 59400 116175
rect 59360 116000 59412 116006
rect 59360 115942 59412 115948
rect 59358 101960 59414 101969
rect 59358 101895 59414 101904
rect 59372 100774 59400 101895
rect 59360 100768 59412 100774
rect 59360 100710 59412 100716
rect 3698 93256 3754 93265
rect 3698 93191 3754 93200
rect 60002 87680 60058 87689
rect 60002 87615 60058 87624
rect 59358 73400 59414 73409
rect 59358 73335 59414 73344
rect 59372 73234 59400 73335
rect 59360 73228 59412 73234
rect 59360 73170 59412 73176
rect 59358 59120 59414 59129
rect 59358 59055 59414 59064
rect 59372 58002 59400 59055
rect 59360 57996 59412 58002
rect 59360 57938 59412 57944
rect 3606 50144 3662 50153
rect 3606 50079 3662 50088
rect 60016 35902 60044 87615
rect 60108 80034 60136 130455
rect 523682 125352 523738 125361
rect 523682 125287 523738 125296
rect 523696 88330 523724 125287
rect 523788 124166 523816 151943
rect 523866 138680 523922 138689
rect 523866 138615 523922 138624
rect 523776 124160 523828 124166
rect 523776 124102 523828 124108
rect 523774 112024 523830 112033
rect 523774 111959 523830 111968
rect 523684 88324 523736 88330
rect 523684 88266 523736 88272
rect 523682 85368 523738 85377
rect 523682 85303 523738 85312
rect 60096 80028 60148 80034
rect 60096 79970 60148 79976
rect 62132 52006 62606 52034
rect 63512 52006 63710 52034
rect 60004 35896 60056 35902
rect 60004 35838 60056 35844
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 62132 3466 62160 52006
rect 63512 3534 63540 52006
rect 64892 48754 64920 52020
rect 66088 48822 66116 52020
rect 67284 49026 67312 52020
rect 68494 52006 68968 52034
rect 69690 52006 70348 52034
rect 67272 49020 67324 49026
rect 67272 48962 67324 48968
rect 66076 48816 66128 48822
rect 66076 48758 66128 48764
rect 66904 48816 66956 48822
rect 66904 48758 66956 48764
rect 64880 48748 64932 48754
rect 64880 48690 64932 48696
rect 66168 48748 66220 48754
rect 66168 48690 66220 48696
rect 66180 4894 66208 48690
rect 66916 15910 66944 48758
rect 66904 15904 66956 15910
rect 66904 15846 66956 15852
rect 66168 4888 66220 4894
rect 66168 4830 66220 4836
rect 68940 4826 68968 52006
rect 70320 42090 70348 52006
rect 70872 48822 70900 52020
rect 72068 48822 72096 52020
rect 73264 48822 73292 52020
rect 70860 48816 70912 48822
rect 70860 48758 70912 48764
rect 71688 48816 71740 48822
rect 71688 48758 71740 48764
rect 72056 48816 72108 48822
rect 72056 48758 72108 48764
rect 73068 48816 73120 48822
rect 73068 48758 73120 48764
rect 73252 48816 73304 48822
rect 73252 48758 73304 48764
rect 74356 48816 74408 48822
rect 74356 48758 74408 48764
rect 70308 42084 70360 42090
rect 70308 42026 70360 42032
rect 68928 4820 68980 4826
rect 68928 4762 68980 4768
rect 71700 3602 71728 48758
rect 73080 18630 73108 48758
rect 74368 43450 74396 48758
rect 74356 43444 74408 43450
rect 74356 43386 74408 43392
rect 73068 18624 73120 18630
rect 73068 18566 73120 18572
rect 71688 3596 71740 3602
rect 71688 3538 71740 3544
rect 74460 3534 74488 52020
rect 75670 52006 75868 52034
rect 76866 52006 77248 52034
rect 78062 52006 78628 52034
rect 79258 52006 80008 52034
rect 75840 19990 75868 52006
rect 77220 44878 77248 52006
rect 77208 44872 77260 44878
rect 77208 44814 77260 44820
rect 75828 19984 75880 19990
rect 75828 19926 75880 19932
rect 78600 3670 78628 52006
rect 79980 21418 80008 52006
rect 80440 46238 80468 52020
rect 81636 49502 81664 52020
rect 81624 49496 81676 49502
rect 81624 49438 81676 49444
rect 82832 48482 82860 52020
rect 84042 52006 84148 52034
rect 85238 52006 85528 52034
rect 86434 52006 86908 52034
rect 87630 52006 88288 52034
rect 82820 48476 82872 48482
rect 82820 48418 82872 48424
rect 84016 48476 84068 48482
rect 84016 48418 84068 48424
rect 80428 46232 80480 46238
rect 80428 46174 80480 46180
rect 84028 22778 84056 48418
rect 84120 47598 84148 52006
rect 84108 47592 84160 47598
rect 84108 47534 84160 47540
rect 84016 22772 84068 22778
rect 84016 22714 84068 22720
rect 79968 21412 80020 21418
rect 79968 21354 80020 21360
rect 78588 3664 78640 3670
rect 78588 3606 78640 3612
rect 63500 3528 63552 3534
rect 63500 3470 63552 3476
rect 74448 3528 74500 3534
rect 85500 3505 85528 52006
rect 86880 24138 86908 52006
rect 86868 24132 86920 24138
rect 86868 24074 86920 24080
rect 88260 3738 88288 52006
rect 88720 49094 88748 52020
rect 88708 49088 88760 49094
rect 88708 49030 88760 49036
rect 89916 48822 89944 52020
rect 91112 48822 91140 52020
rect 92322 52006 92428 52034
rect 93518 52006 93808 52034
rect 94714 52006 95188 52034
rect 89904 48816 89956 48822
rect 89904 48758 89956 48764
rect 91008 48816 91060 48822
rect 91008 48758 91060 48764
rect 91100 48816 91152 48822
rect 91100 48758 91152 48764
rect 92296 48816 92348 48822
rect 92296 48758 92348 48764
rect 91020 25566 91048 48758
rect 91008 25560 91060 25566
rect 91008 25502 91060 25508
rect 92308 4010 92336 48758
rect 92296 4004 92348 4010
rect 92296 3946 92348 3952
rect 88248 3732 88300 3738
rect 88248 3674 88300 3680
rect 74448 3470 74500 3476
rect 85486 3496 85542 3505
rect 62120 3460 62172 3466
rect 85486 3431 85542 3440
rect 62120 3402 62172 3408
rect 92400 3369 92428 52006
rect 93780 26926 93808 52006
rect 93768 26920 93820 26926
rect 93768 26862 93820 26868
rect 95160 3874 95188 52006
rect 95896 49298 95924 52020
rect 95884 49292 95936 49298
rect 95884 49234 95936 49240
rect 97092 48822 97120 52020
rect 98288 48822 98316 52020
rect 99484 48822 99512 52020
rect 100588 52006 100694 52034
rect 101890 52006 102088 52034
rect 97080 48816 97132 48822
rect 97080 48758 97132 48764
rect 97908 48816 97960 48822
rect 97908 48758 97960 48764
rect 98276 48816 98328 48822
rect 98276 48758 98328 48764
rect 99288 48816 99340 48822
rect 99288 48758 99340 48764
rect 99472 48816 99524 48822
rect 99472 48758 99524 48764
rect 97920 28286 97948 48758
rect 97908 28280 97960 28286
rect 97908 28222 97960 28228
rect 95148 3868 95200 3874
rect 95148 3810 95200 3816
rect 92386 3360 92442 3369
rect 92386 3295 92442 3304
rect 99300 3126 99328 48758
rect 100588 6186 100616 52006
rect 100668 48816 100720 48822
rect 100668 48758 100720 48764
rect 100576 6180 100628 6186
rect 100576 6122 100628 6128
rect 100680 3194 100708 48758
rect 102060 29646 102088 52006
rect 103072 49162 103100 52020
rect 104282 52006 104848 52034
rect 103060 49156 103112 49162
rect 103060 49098 103112 49104
rect 102048 29640 102100 29646
rect 102048 29582 102100 29588
rect 104820 7682 104848 52006
rect 105464 48822 105492 52020
rect 106660 48822 106688 52020
rect 107856 48822 107884 52020
rect 109052 48822 109080 52020
rect 110248 49434 110276 52020
rect 111458 52006 111748 52034
rect 112654 52006 113128 52034
rect 110236 49428 110288 49434
rect 110236 49370 110288 49376
rect 105452 48816 105504 48822
rect 105452 48758 105504 48764
rect 106188 48816 106240 48822
rect 106188 48758 106240 48764
rect 106648 48816 106700 48822
rect 106648 48758 106700 48764
rect 107568 48816 107620 48822
rect 107568 48758 107620 48764
rect 107844 48816 107896 48822
rect 107844 48758 107896 48764
rect 108948 48816 109000 48822
rect 108948 48758 109000 48764
rect 109040 48816 109092 48822
rect 109040 48758 109092 48764
rect 110328 48816 110380 48822
rect 110328 48758 110380 48764
rect 106200 31074 106228 48758
rect 106188 31068 106240 31074
rect 106188 31010 106240 31016
rect 104808 7676 104860 7682
rect 104808 7618 104860 7624
rect 100668 3188 100720 3194
rect 100668 3130 100720 3136
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 107580 3058 107608 48758
rect 108960 8974 108988 48758
rect 110340 32502 110368 48758
rect 110328 32496 110380 32502
rect 110328 32438 110380 32444
rect 111720 10334 111748 52006
rect 113100 33862 113128 52006
rect 113744 48822 113772 52020
rect 114940 48822 114968 52020
rect 116136 48822 116164 52020
rect 117332 48822 117360 52020
rect 113732 48816 113784 48822
rect 113732 48758 113784 48764
rect 114468 48816 114520 48822
rect 114468 48758 114520 48764
rect 114928 48816 114980 48822
rect 114928 48758 114980 48764
rect 115848 48816 115900 48822
rect 115848 48758 115900 48764
rect 116124 48816 116176 48822
rect 116124 48758 116176 48764
rect 117228 48816 117280 48822
rect 117228 48758 117280 48764
rect 117320 48816 117372 48822
rect 117320 48758 117372 48764
rect 113088 33856 113140 33862
rect 113088 33798 113140 33804
rect 111708 10328 111760 10334
rect 111708 10270 111760 10276
rect 108948 8968 109000 8974
rect 108948 8910 109000 8916
rect 114480 3942 114508 48758
rect 115860 11762 115888 48758
rect 117240 35290 117268 48758
rect 117228 35284 117280 35290
rect 117228 35226 117280 35232
rect 118528 13122 118556 52020
rect 119738 52006 120028 52034
rect 120934 52006 121408 52034
rect 122130 52006 122788 52034
rect 118608 48816 118660 48822
rect 118608 48758 118660 48764
rect 118516 13116 118568 13122
rect 118516 13058 118568 13064
rect 115848 11756 115900 11762
rect 115848 11698 115900 11704
rect 114468 3936 114520 3942
rect 114468 3878 114520 3884
rect 118620 3262 118648 48758
rect 120000 36582 120028 52006
rect 119988 36576 120040 36582
rect 119988 36518 120040 36524
rect 121380 3806 121408 52006
rect 122760 14482 122788 52006
rect 123312 48754 123340 52020
rect 124508 48822 124536 52020
rect 124496 48816 124548 48822
rect 124496 48758 124548 48764
rect 125508 48816 125560 48822
rect 125508 48758 125560 48764
rect 123300 48748 123352 48754
rect 123300 48690 123352 48696
rect 124128 48748 124180 48754
rect 124128 48690 124180 48696
rect 124140 38010 124168 48690
rect 124128 38004 124180 38010
rect 124128 37946 124180 37952
rect 122748 14476 122800 14482
rect 122748 14418 122800 14424
rect 121368 3800 121420 3806
rect 121368 3742 121420 3748
rect 125520 3330 125548 48758
rect 125704 48686 125732 52020
rect 126808 52006 126914 52034
rect 128110 52006 128308 52034
rect 129306 52006 129688 52034
rect 130502 52006 131068 52034
rect 125692 48680 125744 48686
rect 125692 48622 125744 48628
rect 126808 39370 126836 52006
rect 126888 48680 126940 48686
rect 126888 48622 126940 48628
rect 126796 39364 126848 39370
rect 126796 39306 126848 39312
rect 126900 15978 126928 48622
rect 126888 15972 126940 15978
rect 126888 15914 126940 15920
rect 126980 15904 127032 15910
rect 126980 15846 127032 15852
rect 126612 4888 126664 4894
rect 126612 4830 126664 4836
rect 125508 3324 125560 3330
rect 125508 3266 125560 3272
rect 118608 3256 118660 3262
rect 118608 3198 118660 3204
rect 107568 3052 107620 3058
rect 107568 2994 107620 3000
rect 126624 480 126652 4830
rect 126992 3482 127020 15846
rect 126992 3454 127848 3482
rect 128280 3466 128308 52006
rect 128452 49020 128504 49026
rect 128452 48962 128504 48968
rect 128464 3482 128492 48962
rect 129660 17270 129688 52006
rect 131040 40730 131068 52006
rect 131684 49230 131712 52020
rect 131672 49224 131724 49230
rect 131672 49166 131724 49172
rect 132880 48822 132908 52020
rect 134076 48822 134104 52020
rect 135272 48822 135300 52020
rect 132868 48816 132920 48822
rect 132868 48758 132920 48764
rect 133788 48816 133840 48822
rect 133788 48758 133840 48764
rect 134064 48816 134116 48822
rect 134064 48758 134116 48764
rect 135168 48816 135220 48822
rect 135168 48758 135220 48764
rect 135260 48816 135312 48822
rect 135260 48758 135312 48764
rect 131120 42084 131172 42090
rect 131120 42026 131172 42032
rect 131028 40724 131080 40730
rect 131028 40666 131080 40672
rect 129648 17264 129700 17270
rect 129648 17206 129700 17212
rect 130200 4820 130252 4826
rect 130200 4762 130252 4768
rect 127820 480 127848 3454
rect 128268 3460 128320 3466
rect 128464 3454 129044 3482
rect 128268 3402 128320 3408
rect 129016 480 129044 3454
rect 130212 480 130240 4762
rect 131132 3482 131160 42026
rect 132592 18624 132644 18630
rect 132592 18566 132644 18572
rect 132604 4078 132632 18566
rect 133800 4962 133828 48758
rect 133880 43444 133932 43450
rect 133880 43386 133932 43392
rect 133788 4956 133840 4962
rect 133788 4898 133840 4904
rect 132592 4072 132644 4078
rect 132592 4014 132644 4020
rect 133788 4072 133840 4078
rect 133788 4014 133840 4020
rect 132500 3596 132552 3602
rect 132500 3538 132552 3544
rect 131132 3454 131436 3482
rect 131408 480 131436 3454
rect 132512 3346 132540 3538
rect 132512 3318 132632 3346
rect 132604 480 132632 3318
rect 133800 480 133828 4014
rect 133892 3346 133920 43386
rect 135180 42158 135208 48758
rect 135168 42152 135220 42158
rect 135168 42094 135220 42100
rect 136468 18630 136496 52020
rect 137678 52006 137968 52034
rect 136548 48816 136600 48822
rect 136548 48758 136600 48764
rect 136456 18624 136508 18630
rect 136456 18566 136508 18572
rect 136088 3596 136140 3602
rect 136088 3538 136140 3544
rect 133892 3318 134932 3346
rect 134904 480 134932 3318
rect 136100 480 136128 3538
rect 136560 3398 136588 48758
rect 136640 19984 136692 19990
rect 136640 19926 136692 19932
rect 136548 3392 136600 3398
rect 136548 3334 136600 3340
rect 136652 3346 136680 19926
rect 137940 7614 137968 52006
rect 138860 49366 138888 52020
rect 139978 52006 140728 52034
rect 138848 49360 138900 49366
rect 138848 49302 138900 49308
rect 138020 44872 138072 44878
rect 138020 44814 138072 44820
rect 137928 7608 137980 7614
rect 137928 7550 137980 7556
rect 138032 3346 138060 44814
rect 140700 19990 140728 52006
rect 141160 48822 141188 52020
rect 142252 49496 142304 49502
rect 142252 49438 142304 49444
rect 141148 48816 141200 48822
rect 141148 48758 141200 48764
rect 142068 48816 142120 48822
rect 142068 48758 142120 48764
rect 140780 46232 140832 46238
rect 140780 46174 140832 46180
rect 140688 19984 140740 19990
rect 140688 19926 140740 19932
rect 139676 3664 139728 3670
rect 139676 3606 139728 3612
rect 136652 3318 137324 3346
rect 138032 3318 138520 3346
rect 137296 480 137324 3318
rect 138492 480 138520 3318
rect 139688 480 139716 3606
rect 140792 3534 140820 46174
rect 142080 43450 142108 48758
rect 142068 43444 142120 43450
rect 142068 43386 142120 43392
rect 140872 21412 140924 21418
rect 140872 21354 140924 21360
rect 140780 3528 140832 3534
rect 140780 3470 140832 3476
rect 140884 480 140912 21354
rect 142068 3528 142120 3534
rect 142068 3470 142120 3476
rect 142080 480 142108 3470
rect 142264 3346 142292 49438
rect 142356 48822 142384 52020
rect 143552 48822 143580 52020
rect 142344 48816 142396 48822
rect 142344 48758 142396 48764
rect 143448 48816 143500 48822
rect 143448 48758 143500 48764
rect 143540 48816 143592 48822
rect 143540 48758 143592 48764
rect 143460 4146 143488 48758
rect 144748 44878 144776 52020
rect 145944 49026 145972 52020
rect 147154 52006 147628 52034
rect 145932 49020 145984 49026
rect 145932 48962 145984 48968
rect 144828 48816 144880 48822
rect 144828 48758 144880 48764
rect 144736 44872 144788 44878
rect 144736 44814 144788 44820
rect 143540 22772 143592 22778
rect 143540 22714 143592 22720
rect 143448 4140 143500 4146
rect 143448 4082 143500 4088
rect 143552 3346 143580 22714
rect 144840 21418 144868 48758
rect 144920 47592 144972 47598
rect 144920 47534 144972 47540
rect 144828 21412 144880 21418
rect 144828 21354 144880 21360
rect 144932 3346 144960 47534
rect 147600 22778 147628 52006
rect 148336 46238 148364 52020
rect 149532 48822 149560 52020
rect 150624 49088 150676 49094
rect 150624 49030 150676 49036
rect 149520 48816 149572 48822
rect 149520 48758 149572 48764
rect 150348 48816 150400 48822
rect 150348 48758 150400 48764
rect 148324 46232 148376 46238
rect 148324 46174 148376 46180
rect 147680 24132 147732 24138
rect 147680 24074 147732 24080
rect 147588 22772 147640 22778
rect 147588 22714 147640 22720
rect 146850 3496 146906 3505
rect 146850 3431 146906 3440
rect 142264 3318 143304 3346
rect 143552 3318 144500 3346
rect 144932 3318 145696 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3318
rect 146864 480 146892 3431
rect 147692 3346 147720 24074
rect 150360 4078 150388 48758
rect 150532 25560 150584 25566
rect 150532 25502 150584 25508
rect 150348 4072 150400 4078
rect 150348 4014 150400 4020
rect 149244 3732 149296 3738
rect 149244 3674 149296 3680
rect 147692 3318 148088 3346
rect 148060 480 148088 3318
rect 149256 480 149284 3674
rect 150544 3602 150572 25502
rect 150532 3596 150584 3602
rect 150532 3538 150584 3544
rect 150636 3482 150664 49030
rect 150728 48822 150756 52020
rect 150716 48816 150768 48822
rect 150716 48758 150768 48764
rect 151728 48816 151780 48822
rect 151728 48758 151780 48764
rect 151740 24138 151768 48758
rect 151924 47666 151952 52020
rect 153028 52006 153134 52034
rect 154330 52006 154528 52034
rect 155526 52006 155908 52034
rect 156722 52006 157288 52034
rect 151912 47660 151964 47666
rect 151912 47602 151964 47608
rect 151728 24132 151780 24138
rect 151728 24074 151780 24080
rect 152740 4004 152792 4010
rect 152740 3946 152792 3952
rect 151544 3596 151596 3602
rect 151544 3538 151596 3544
rect 150452 3454 150664 3482
rect 150452 480 150480 3454
rect 151556 480 151584 3538
rect 152752 480 152780 3946
rect 153028 3738 153056 52006
rect 154500 25566 154528 52006
rect 155880 29714 155908 52006
rect 155868 29708 155920 29714
rect 155868 29650 155920 29656
rect 154580 26920 154632 26926
rect 154580 26862 154632 26868
rect 154488 25560 154540 25566
rect 154488 25502 154540 25508
rect 153016 3732 153068 3738
rect 153016 3674 153068 3680
rect 153934 3360 153990 3369
rect 154592 3346 154620 26862
rect 156328 3868 156380 3874
rect 156328 3810 156380 3816
rect 154592 3318 155172 3346
rect 153934 3295 153990 3304
rect 153948 480 153976 3295
rect 155144 480 155172 3318
rect 156340 480 156368 3810
rect 157260 3670 157288 52006
rect 157432 49292 157484 49298
rect 157432 49234 157484 49240
rect 157248 3664 157300 3670
rect 157248 3606 157300 3612
rect 157444 1578 157472 49234
rect 157904 48754 157932 52020
rect 159100 48822 159128 52020
rect 160296 48822 160324 52020
rect 161492 48822 161520 52020
rect 159088 48816 159140 48822
rect 159088 48758 159140 48764
rect 160008 48816 160060 48822
rect 160008 48758 160060 48764
rect 160284 48816 160336 48822
rect 160284 48758 160336 48764
rect 161388 48816 161440 48822
rect 161388 48758 161440 48764
rect 161480 48816 161532 48822
rect 161480 48758 161532 48764
rect 157892 48748 157944 48754
rect 157892 48690 157944 48696
rect 158628 48748 158680 48754
rect 158628 48690 158680 48696
rect 158640 26926 158668 48690
rect 160020 31142 160048 48758
rect 160008 31136 160060 31142
rect 160008 31078 160060 31084
rect 158812 28280 158864 28286
rect 158812 28222 158864 28228
rect 158628 26920 158680 26926
rect 158628 26862 158680 26868
rect 158824 1578 158852 28222
rect 161400 4010 161428 48758
rect 162688 32434 162716 52020
rect 163898 52006 164188 52034
rect 165002 52006 165568 52034
rect 162768 48816 162820 48822
rect 162768 48758 162820 48764
rect 162676 32428 162728 32434
rect 162676 32370 162728 32376
rect 162780 6322 162808 48758
rect 162860 29640 162912 29646
rect 162860 29582 162912 29588
rect 162768 6316 162820 6322
rect 162768 6258 162820 6264
rect 162308 6180 162360 6186
rect 162308 6122 162360 6128
rect 161388 4004 161440 4010
rect 161388 3946 161440 3952
rect 161112 3188 161164 3194
rect 161112 3130 161164 3136
rect 159916 3120 159968 3126
rect 159916 3062 159968 3068
rect 157444 1550 157564 1578
rect 157536 480 157564 1550
rect 158732 1550 158852 1578
rect 158732 480 158760 1550
rect 159928 480 159956 3062
rect 161124 480 161152 3130
rect 162320 480 162348 6122
rect 162872 3482 162900 29582
rect 164160 3602 164188 52006
rect 164332 49156 164384 49162
rect 164332 49098 164384 49104
rect 164148 3596 164200 3602
rect 164148 3538 164200 3544
rect 164344 3482 164372 49098
rect 165540 28286 165568 52006
rect 166184 48822 166212 52020
rect 167380 49502 167408 52020
rect 167368 49496 167420 49502
rect 167368 49438 167420 49444
rect 168576 48822 168604 52020
rect 169772 48822 169800 52020
rect 170982 52006 171088 52034
rect 172178 52006 172468 52034
rect 173374 52006 173848 52034
rect 166172 48816 166224 48822
rect 166172 48758 166224 48764
rect 166908 48816 166960 48822
rect 166908 48758 166960 48764
rect 168564 48816 168616 48822
rect 168564 48758 168616 48764
rect 169668 48816 169720 48822
rect 169668 48758 169720 48764
rect 169760 48816 169812 48822
rect 169760 48758 169812 48764
rect 170956 48816 171008 48822
rect 170956 48758 171008 48764
rect 166920 33794 166948 48758
rect 166908 33788 166960 33794
rect 166908 33730 166960 33736
rect 167092 31068 167144 31074
rect 167092 31010 167144 31016
rect 165528 28280 165580 28286
rect 165528 28222 165580 28228
rect 165896 7676 165948 7682
rect 165896 7618 165948 7624
rect 162872 3454 163544 3482
rect 164344 3454 164740 3482
rect 163516 480 163544 3454
rect 164712 480 164740 3454
rect 165908 480 165936 7618
rect 167104 480 167132 31010
rect 169392 8968 169444 8974
rect 169392 8910 169444 8916
rect 168196 3052 168248 3058
rect 168196 2994 168248 3000
rect 168208 480 168236 2994
rect 169404 480 169432 8910
rect 169680 7682 169708 48758
rect 170968 35222 170996 48758
rect 170956 35216 171008 35222
rect 170956 35158 171008 35164
rect 169760 32496 169812 32502
rect 169760 32438 169812 32444
rect 169668 7676 169720 7682
rect 169668 7618 169720 7624
rect 169772 3482 169800 32438
rect 171060 3534 171088 52006
rect 171232 49428 171284 49434
rect 171232 49370 171284 49376
rect 171048 3528 171100 3534
rect 169772 3454 170628 3482
rect 171048 3470 171100 3476
rect 170600 480 170628 3454
rect 171244 3346 171272 49370
rect 172440 8974 172468 52006
rect 172520 10328 172572 10334
rect 172520 10270 172572 10276
rect 172428 8968 172480 8974
rect 172428 8910 172480 8916
rect 172532 3346 172560 10270
rect 173820 4826 173848 52006
rect 174556 49298 174584 52020
rect 174544 49292 174596 49298
rect 174544 49234 174596 49240
rect 175752 48822 175780 52020
rect 175740 48816 175792 48822
rect 175740 48758 175792 48764
rect 176568 48816 176620 48822
rect 176568 48758 176620 48764
rect 173900 33856 173952 33862
rect 173900 33798 173952 33804
rect 173808 4820 173860 4826
rect 173808 4762 173860 4768
rect 173912 3346 173940 33798
rect 175372 11756 175424 11762
rect 175372 11698 175424 11704
rect 175280 3936 175332 3942
rect 175280 3878 175332 3884
rect 171244 3318 171824 3346
rect 172532 3318 173020 3346
rect 173912 3318 174216 3346
rect 171796 480 171824 3318
rect 172992 480 173020 3318
rect 174188 480 174216 3318
rect 175292 2258 175320 3878
rect 175384 3262 175412 11698
rect 176580 10402 176608 48758
rect 176948 48482 176976 52020
rect 178144 48822 178172 52020
rect 179248 52006 179354 52034
rect 180550 52006 180748 52034
rect 178132 48816 178184 48822
rect 178132 48758 178184 48764
rect 176936 48476 176988 48482
rect 176936 48418 176988 48424
rect 177948 48476 178000 48482
rect 177948 48418 178000 48424
rect 177960 36650 177988 48418
rect 177948 36644 178000 36650
rect 177948 36586 178000 36592
rect 176660 35284 176712 35290
rect 176660 35226 176712 35232
rect 176568 10396 176620 10402
rect 176568 10338 176620 10344
rect 176672 3346 176700 35226
rect 179248 11762 179276 52006
rect 179328 48816 179380 48822
rect 179328 48758 179380 48764
rect 179236 11756 179288 11762
rect 179236 11698 179288 11704
rect 176672 3318 177804 3346
rect 175372 3256 175424 3262
rect 175372 3198 175424 3204
rect 176568 3256 176620 3262
rect 176568 3198 176620 3204
rect 175292 2230 175412 2258
rect 175384 480 175412 2230
rect 176580 480 176608 3198
rect 177776 480 177804 3318
rect 179340 3194 179368 48758
rect 180720 37942 180748 52006
rect 181732 49162 181760 52020
rect 182942 52006 183508 52034
rect 184138 52006 184888 52034
rect 181720 49156 181772 49162
rect 181720 49098 181772 49104
rect 180708 37936 180760 37942
rect 180708 37878 180760 37884
rect 180800 36576 180852 36582
rect 180800 36518 180852 36524
rect 179420 13116 179472 13122
rect 179420 13058 179472 13064
rect 179432 3346 179460 13058
rect 180812 3346 180840 36518
rect 183480 13122 183508 52006
rect 184860 39438 184888 52006
rect 185320 48822 185348 52020
rect 185308 48816 185360 48822
rect 185308 48758 185360 48764
rect 186228 48816 186280 48822
rect 186228 48758 186280 48764
rect 184848 39432 184900 39438
rect 184848 39374 184900 39380
rect 183560 38004 183612 38010
rect 183560 37946 183612 37952
rect 183468 13116 183520 13122
rect 183468 13058 183520 13064
rect 182548 3800 182600 3806
rect 182548 3742 182600 3748
rect 179432 3318 180196 3346
rect 180812 3318 181392 3346
rect 178960 3188 179012 3194
rect 178960 3130 179012 3136
rect 179328 3188 179380 3194
rect 179328 3130 179380 3136
rect 178972 480 179000 3130
rect 180168 480 180196 3318
rect 181364 480 181392 3318
rect 182560 480 182588 3742
rect 183572 3466 183600 37946
rect 183652 14476 183704 14482
rect 183652 14418 183704 14424
rect 183664 3482 183692 14418
rect 183560 3460 183612 3466
rect 183664 3454 183784 3482
rect 183560 3402 183612 3408
rect 183756 480 183784 3454
rect 184848 3460 184900 3466
rect 184848 3402 184900 3408
rect 184860 480 184888 3402
rect 186044 3324 186096 3330
rect 186044 3266 186096 3272
rect 186056 480 186084 3266
rect 186240 3126 186268 48758
rect 186516 48686 186544 52020
rect 187712 48822 187740 52020
rect 188908 49094 188936 52020
rect 190118 52006 190408 52034
rect 191222 52006 191788 52034
rect 192418 52006 193168 52034
rect 188896 49088 188948 49094
rect 188896 49030 188948 49036
rect 187700 48816 187752 48822
rect 187700 48758 187752 48764
rect 188988 48816 189040 48822
rect 188988 48758 189040 48764
rect 186504 48680 186556 48686
rect 186504 48622 186556 48628
rect 187608 48680 187660 48686
rect 187608 48622 187660 48628
rect 186320 15972 186372 15978
rect 186320 15914 186372 15920
rect 186332 3346 186360 15914
rect 187620 14482 187648 48622
rect 189000 40798 189028 48758
rect 188988 40792 189040 40798
rect 188988 40734 189040 40740
rect 187700 39364 187752 39370
rect 187700 39306 187752 39312
rect 187608 14476 187660 14482
rect 187608 14418 187660 14424
rect 187712 3346 187740 39306
rect 190380 4894 190408 52006
rect 191760 42090 191788 52006
rect 191748 42084 191800 42090
rect 191748 42026 191800 42032
rect 191840 40724 191892 40730
rect 191840 40666 191892 40672
rect 190460 17264 190512 17270
rect 190460 17206 190512 17212
rect 190368 4888 190420 4894
rect 190368 4830 190420 4836
rect 190472 3346 190500 17206
rect 191852 3346 191880 40666
rect 186332 3318 187280 3346
rect 187712 3318 188476 3346
rect 190472 3318 190868 3346
rect 191852 3318 192064 3346
rect 193140 3330 193168 52006
rect 193404 49224 193456 49230
rect 193404 49166 193456 49172
rect 193416 3346 193444 49166
rect 193600 48822 193628 52020
rect 194796 48822 194824 52020
rect 193588 48816 193640 48822
rect 193588 48758 193640 48764
rect 194508 48816 194560 48822
rect 194508 48758 194560 48764
rect 194784 48816 194836 48822
rect 194784 48758 194836 48764
rect 195888 48816 195940 48822
rect 195888 48758 195940 48764
rect 194520 15910 194548 48758
rect 195900 43518 195928 48758
rect 195992 48550 196020 52020
rect 195980 48544 196032 48550
rect 195980 48486 196032 48492
rect 195888 43512 195940 43518
rect 195888 43454 195940 43460
rect 194600 42152 194652 42158
rect 194600 42094 194652 42100
rect 194508 15904 194560 15910
rect 194508 15846 194560 15852
rect 194416 4956 194468 4962
rect 194416 4898 194468 4904
rect 186228 3120 186280 3126
rect 186228 3062 186280 3068
rect 187252 480 187280 3318
rect 188448 480 188476 3318
rect 189632 3256 189684 3262
rect 189632 3198 189684 3204
rect 189644 480 189672 3198
rect 190840 480 190868 3318
rect 192036 480 192064 3318
rect 193128 3324 193180 3330
rect 193128 3266 193180 3272
rect 193232 3318 193444 3346
rect 193232 480 193260 3318
rect 194428 480 194456 4898
rect 194612 3346 194640 42094
rect 197188 17270 197216 52020
rect 198398 52006 198688 52034
rect 199594 52006 200068 52034
rect 200790 52006 201448 52034
rect 197268 48544 197320 48550
rect 197268 48486 197320 48492
rect 197176 17264 197228 17270
rect 197176 17206 197228 17212
rect 196808 3392 196860 3398
rect 194612 3318 195652 3346
rect 196808 3334 196860 3340
rect 195624 480 195652 3318
rect 196820 480 196848 3334
rect 197280 3262 197308 48486
rect 198660 44946 198688 52006
rect 198648 44940 198700 44946
rect 198648 44882 198700 44888
rect 197360 18624 197412 18630
rect 197360 18566 197412 18572
rect 197372 3346 197400 18566
rect 199200 7608 199252 7614
rect 199200 7550 199252 7556
rect 197372 3318 198044 3346
rect 197268 3256 197320 3262
rect 197268 3198 197320 3204
rect 198016 480 198044 3318
rect 199212 480 199240 7550
rect 200040 3806 200068 52006
rect 200212 49360 200264 49366
rect 200212 49302 200264 49308
rect 200028 3800 200080 3806
rect 200028 3742 200080 3748
rect 200224 3346 200252 49302
rect 201420 18630 201448 52006
rect 201972 46306 202000 52020
rect 203168 48822 203196 52020
rect 204364 48822 204392 52020
rect 203156 48816 203208 48822
rect 203156 48758 203208 48764
rect 204168 48816 204220 48822
rect 204168 48758 204220 48764
rect 204352 48816 204404 48822
rect 204352 48758 204404 48764
rect 205456 48816 205508 48822
rect 205456 48758 205508 48764
rect 201960 46300 202012 46306
rect 201960 46242 202012 46248
rect 201500 43444 201552 43450
rect 201500 43386 201552 43392
rect 201408 18624 201460 18630
rect 201408 18566 201460 18572
rect 201512 3874 201540 43386
rect 201592 19984 201644 19990
rect 201592 19926 201644 19932
rect 201500 3868 201552 3874
rect 201500 3810 201552 3816
rect 201604 3482 201632 19926
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 202696 3868 202748 3874
rect 202696 3810 202748 3816
rect 201512 3454 201632 3482
rect 200224 3318 200436 3346
rect 200408 480 200436 3318
rect 201512 480 201540 3454
rect 202708 480 202736 3810
rect 203904 480 203932 4082
rect 204180 3058 204208 48758
rect 205468 21418 205496 48758
rect 205560 47598 205588 52020
rect 206770 52006 206968 52034
rect 207966 52006 208348 52034
rect 209162 52006 209728 52034
rect 205548 47592 205600 47598
rect 205548 47534 205600 47540
rect 205640 44872 205692 44878
rect 205640 44814 205692 44820
rect 204260 21412 204312 21418
rect 204260 21354 204312 21360
rect 205456 21412 205508 21418
rect 205456 21354 205508 21360
rect 204272 3346 204300 21354
rect 205652 3346 205680 44814
rect 206940 3874 206968 52006
rect 207112 49020 207164 49026
rect 207112 48962 207164 48968
rect 206928 3868 206980 3874
rect 206928 3810 206980 3816
rect 207124 3346 207152 48962
rect 208320 19990 208348 52006
rect 208400 22772 208452 22778
rect 208400 22714 208452 22720
rect 208308 19984 208360 19990
rect 208308 19926 208360 19932
rect 208412 3346 208440 22714
rect 209700 6186 209728 52006
rect 210344 49366 210372 52020
rect 210332 49360 210384 49366
rect 210332 49302 210384 49308
rect 211540 48822 211568 52020
rect 212736 48822 212764 52020
rect 213932 48822 213960 52020
rect 211528 48816 211580 48822
rect 211528 48758 211580 48764
rect 212448 48816 212500 48822
rect 212448 48758 212500 48764
rect 212724 48816 212776 48822
rect 212724 48758 212776 48764
rect 213828 48816 213880 48822
rect 213828 48758 213880 48764
rect 213920 48816 213972 48822
rect 213920 48758 213972 48764
rect 209872 46232 209924 46238
rect 209872 46174 209924 46180
rect 209688 6180 209740 6186
rect 209688 6122 209740 6128
rect 204272 3318 205128 3346
rect 205652 3318 206324 3346
rect 207124 3318 207520 3346
rect 208412 3318 208716 3346
rect 204168 3052 204220 3058
rect 204168 2994 204220 3000
rect 205100 480 205128 3318
rect 206296 480 206324 3318
rect 207492 480 207520 3318
rect 208688 480 208716 3318
rect 209884 480 209912 46174
rect 211160 24132 211212 24138
rect 211160 24074 211212 24080
rect 211068 4072 211120 4078
rect 211068 4014 211120 4020
rect 211080 480 211108 4014
rect 211172 3346 211200 24074
rect 212460 22778 212488 48758
rect 212540 47660 212592 47666
rect 212540 47602 212592 47608
rect 212448 22772 212500 22778
rect 212448 22714 212500 22720
rect 212552 3346 212580 47602
rect 213840 29782 213868 48758
rect 213828 29776 213880 29782
rect 213828 29718 213880 29724
rect 215128 24138 215156 52020
rect 216246 52006 216628 52034
rect 215208 48816 215260 48822
rect 215208 48758 215260 48764
rect 215116 24132 215168 24138
rect 215116 24074 215168 24080
rect 215220 3942 215248 48758
rect 216600 31074 216628 52006
rect 217428 49230 217456 52020
rect 217416 49224 217468 49230
rect 217416 49166 217468 49172
rect 218624 48822 218652 52020
rect 219820 48822 219848 52020
rect 221016 48822 221044 52020
rect 222212 48822 222240 52020
rect 218612 48816 218664 48822
rect 218612 48758 218664 48764
rect 219348 48816 219400 48822
rect 219348 48758 219400 48764
rect 219808 48816 219860 48822
rect 219808 48758 219860 48764
rect 220728 48816 220780 48822
rect 220728 48758 220780 48764
rect 221004 48816 221056 48822
rect 221004 48758 221056 48764
rect 222108 48816 222160 48822
rect 222108 48758 222160 48764
rect 222200 48816 222252 48822
rect 222200 48758 222252 48764
rect 216588 31068 216640 31074
rect 216588 31010 216640 31016
rect 216680 29708 216732 29714
rect 216680 29650 216732 29656
rect 215300 25560 215352 25566
rect 215300 25502 215352 25508
rect 215208 3936 215260 3942
rect 215208 3878 215260 3884
rect 214656 3732 214708 3738
rect 214656 3674 214708 3680
rect 211172 3318 212304 3346
rect 212552 3318 213500 3346
rect 212276 480 212304 3318
rect 213472 480 213500 3318
rect 214668 480 214696 3674
rect 215312 3346 215340 25502
rect 216692 3346 216720 29650
rect 218152 26920 218204 26926
rect 218152 26862 218204 26868
rect 218060 3664 218112 3670
rect 218060 3606 218112 3612
rect 218072 3346 218100 3606
rect 218164 3466 218192 26862
rect 219360 6254 219388 48758
rect 220740 32502 220768 48758
rect 220728 32496 220780 32502
rect 220728 32438 220780 32444
rect 219440 31136 219492 31142
rect 219440 31078 219492 31084
rect 219348 6248 219400 6254
rect 219348 6190 219400 6196
rect 218152 3460 218204 3466
rect 218152 3402 218204 3408
rect 219348 3460 219400 3466
rect 219348 3402 219400 3408
rect 215312 3318 215892 3346
rect 216692 3318 217088 3346
rect 218072 3318 218192 3346
rect 215864 480 215892 3318
rect 217060 480 217088 3318
rect 218164 480 218192 3318
rect 219360 480 219388 3402
rect 219452 3346 219480 31078
rect 221740 4004 221792 4010
rect 221740 3946 221792 3952
rect 219452 3318 220584 3346
rect 220556 480 220584 3318
rect 221752 480 221780 3946
rect 222120 3738 222148 48758
rect 223408 33862 223436 52020
rect 224604 49026 224632 52020
rect 225814 52006 226288 52034
rect 227010 52006 227668 52034
rect 224592 49020 224644 49026
rect 224592 48962 224644 48968
rect 223488 48816 223540 48822
rect 223488 48758 223540 48764
rect 223396 33856 223448 33862
rect 223396 33798 223448 33804
rect 223500 7614 223528 48758
rect 223580 32428 223632 32434
rect 223580 32370 223632 32376
rect 223488 7608 223540 7614
rect 223488 7550 223540 7556
rect 222936 6316 222988 6322
rect 222936 6258 222988 6264
rect 222108 3732 222160 3738
rect 222108 3674 222160 3680
rect 222948 480 222976 6258
rect 223592 3346 223620 32370
rect 226260 25566 226288 52006
rect 227640 35290 227668 52006
rect 227904 49496 227956 49502
rect 227904 49438 227956 49444
rect 227628 35284 227680 35290
rect 227628 35226 227680 35232
rect 227812 33788 227864 33794
rect 227812 33730 227864 33736
rect 226340 28280 226392 28286
rect 226340 28222 226392 28228
rect 226248 25560 226300 25566
rect 226248 25502 226300 25508
rect 225328 3596 225380 3602
rect 225328 3538 225380 3544
rect 223592 3318 224172 3346
rect 224144 480 224172 3318
rect 225340 480 225368 3538
rect 226352 3448 226380 28222
rect 227824 3482 227852 33730
rect 227732 3454 227852 3482
rect 226352 3420 226564 3448
rect 226536 480 226564 3420
rect 227732 480 227760 3454
rect 227916 3346 227944 49438
rect 228192 48822 228220 52020
rect 229388 48822 229416 52020
rect 228180 48816 228232 48822
rect 228180 48758 228232 48764
rect 229008 48816 229060 48822
rect 229008 48758 229060 48764
rect 229376 48816 229428 48822
rect 229376 48758 229428 48764
rect 230388 48816 230440 48822
rect 230388 48758 230440 48764
rect 229020 3398 229048 48758
rect 230400 9042 230428 48758
rect 230584 48686 230612 52020
rect 230572 48680 230624 48686
rect 230572 48622 230624 48628
rect 231676 48680 231728 48686
rect 231676 48622 231728 48628
rect 231688 36582 231716 48622
rect 231676 36576 231728 36582
rect 231676 36518 231728 36524
rect 230480 35216 230532 35222
rect 230480 35158 230532 35164
rect 230388 9036 230440 9042
rect 230388 8978 230440 8984
rect 230112 7676 230164 7682
rect 230112 7618 230164 7624
rect 229008 3392 229060 3398
rect 227916 3318 228956 3346
rect 229008 3334 229060 3340
rect 228928 480 228956 3318
rect 230124 480 230152 7618
rect 230492 3482 230520 35158
rect 230492 3454 231348 3482
rect 231780 3466 231808 52020
rect 232990 52006 233188 52034
rect 234186 52006 234568 52034
rect 235382 52006 235948 52034
rect 236578 52006 237328 52034
rect 233160 10334 233188 52006
rect 234540 38010 234568 52006
rect 234528 38004 234580 38010
rect 234528 37946 234580 37952
rect 233148 10328 233200 10334
rect 233148 10270 233200 10276
rect 233700 8968 233752 8974
rect 233700 8910 233752 8916
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 231320 480 231348 3454
rect 231768 3460 231820 3466
rect 231768 3402 231820 3408
rect 232516 480 232544 3470
rect 233712 480 233740 8910
rect 234804 4820 234856 4826
rect 234804 4762 234856 4768
rect 234816 480 234844 4762
rect 235920 3534 235948 52006
rect 236184 49292 236236 49298
rect 236184 49234 236236 49240
rect 236092 10396 236144 10402
rect 236092 10338 236144 10344
rect 236104 3602 236132 10338
rect 236092 3596 236144 3602
rect 236092 3538 236144 3544
rect 235908 3528 235960 3534
rect 236196 3482 236224 49234
rect 237300 26926 237328 52006
rect 237760 48822 237788 52020
rect 238956 48822 238984 52020
rect 240152 48822 240180 52020
rect 237748 48816 237800 48822
rect 237748 48758 237800 48764
rect 238668 48816 238720 48822
rect 238668 48758 238720 48764
rect 238944 48816 238996 48822
rect 238944 48758 238996 48764
rect 240048 48816 240100 48822
rect 240048 48758 240100 48764
rect 240140 48816 240192 48822
rect 240140 48758 240192 48764
rect 238680 39370 238708 48758
rect 238668 39364 238720 39370
rect 238668 39306 238720 39312
rect 237380 36644 237432 36650
rect 237380 36586 237432 36592
rect 237288 26920 237340 26926
rect 237288 26862 237340 26868
rect 237196 3596 237248 3602
rect 237196 3538 237248 3544
rect 235908 3470 235960 3476
rect 236012 3454 236224 3482
rect 236012 480 236040 3454
rect 237208 480 237236 3538
rect 237392 3482 237420 36586
rect 237392 3454 238432 3482
rect 238404 480 238432 3454
rect 240060 3194 240088 48758
rect 241348 40730 241376 52020
rect 242466 52006 242848 52034
rect 243662 52006 244228 52034
rect 244858 52006 245608 52034
rect 241428 48816 241480 48822
rect 241428 48758 241480 48764
rect 241336 40724 241388 40730
rect 241336 40666 241388 40672
rect 241440 11762 241468 48758
rect 241520 37936 241572 37942
rect 241520 37878 241572 37884
rect 240140 11756 240192 11762
rect 240140 11698 240192 11704
rect 241428 11756 241480 11762
rect 241428 11698 241480 11704
rect 240152 3346 240180 11698
rect 241532 3346 241560 37878
rect 242820 3670 242848 52006
rect 242992 49156 243044 49162
rect 242992 49098 243044 49104
rect 242808 3664 242860 3670
rect 242808 3606 242860 3612
rect 243004 3346 243032 49098
rect 244200 28286 244228 52006
rect 245580 42158 245608 52006
rect 246040 48822 246068 52020
rect 247236 48822 247264 52020
rect 248432 48822 248460 52020
rect 249642 52006 249748 52034
rect 250838 52006 251128 52034
rect 252034 52006 252508 52034
rect 246028 48816 246080 48822
rect 246028 48758 246080 48764
rect 246948 48816 247000 48822
rect 246948 48758 247000 48764
rect 247224 48816 247276 48822
rect 247224 48758 247276 48764
rect 248328 48816 248380 48822
rect 248328 48758 248380 48764
rect 248420 48816 248472 48822
rect 248420 48758 248472 48764
rect 249616 48816 249668 48822
rect 249616 48758 249668 48764
rect 245568 42152 245620 42158
rect 245568 42094 245620 42100
rect 244280 39432 244332 39438
rect 244280 39374 244332 39380
rect 244188 28280 244240 28286
rect 244188 28222 244240 28228
rect 244292 3602 244320 39374
rect 244372 13116 244424 13122
rect 244372 13058 244424 13064
rect 244280 3596 244332 3602
rect 244280 3538 244332 3544
rect 240152 3318 240824 3346
rect 241532 3318 242020 3346
rect 243004 3318 243216 3346
rect 239588 3188 239640 3194
rect 239588 3130 239640 3136
rect 240048 3188 240100 3194
rect 240048 3130 240100 3136
rect 239600 480 239628 3130
rect 240796 480 240824 3318
rect 241992 480 242020 3318
rect 243188 480 243216 3318
rect 244384 480 244412 13058
rect 246960 4146 246988 48758
rect 248340 14550 248368 48758
rect 249628 43450 249656 48758
rect 249616 43444 249668 43450
rect 249616 43386 249668 43392
rect 248420 40792 248472 40798
rect 248420 40734 248472 40740
rect 248328 14544 248380 14550
rect 248328 14486 248380 14492
rect 247040 14476 247092 14482
rect 247040 14418 247092 14424
rect 246948 4140 247000 4146
rect 246948 4082 247000 4088
rect 245568 3596 245620 3602
rect 245568 3538 245620 3544
rect 245580 480 245608 3538
rect 247052 3346 247080 14418
rect 248432 3346 248460 40734
rect 249720 3670 249748 52006
rect 249892 49088 249944 49094
rect 249892 49030 249944 49036
rect 249708 3664 249760 3670
rect 249708 3606 249760 3612
rect 249904 3346 249932 49030
rect 251100 13122 251128 52006
rect 252480 29646 252508 52006
rect 253216 49298 253244 52020
rect 253204 49292 253256 49298
rect 253204 49234 253256 49240
rect 254412 48822 254440 52020
rect 255608 48822 255636 52020
rect 256804 48822 256832 52020
rect 257908 52006 258014 52034
rect 254400 48816 254452 48822
rect 254400 48758 254452 48764
rect 255228 48816 255280 48822
rect 255228 48758 255280 48764
rect 255596 48816 255648 48822
rect 255596 48758 255648 48764
rect 256608 48816 256660 48822
rect 256608 48758 256660 48764
rect 256792 48816 256844 48822
rect 256792 48758 256844 48764
rect 252652 42084 252704 42090
rect 252652 42026 252704 42032
rect 252468 29640 252520 29646
rect 252468 29582 252520 29588
rect 251088 13116 251140 13122
rect 251088 13058 251140 13064
rect 251456 4888 251508 4894
rect 251456 4830 251508 4836
rect 247052 3318 248000 3346
rect 248432 3318 249196 3346
rect 249904 3318 250392 3346
rect 246764 3120 246816 3126
rect 246764 3062 246816 3068
rect 246776 480 246804 3062
rect 247972 480 248000 3318
rect 249168 480 249196 3318
rect 250364 480 250392 3318
rect 251468 480 251496 4830
rect 252664 480 252692 42026
rect 253940 15904 253992 15910
rect 253940 15846 253992 15852
rect 253952 3346 253980 15846
rect 255240 4894 255268 48758
rect 256620 45014 256648 48758
rect 256608 45008 256660 45014
rect 256608 44950 256660 44956
rect 255320 43512 255372 43518
rect 255320 43454 255372 43460
rect 255228 4888 255280 4894
rect 255228 4830 255280 4836
rect 255332 3346 255360 43454
rect 257908 15910 257936 52006
rect 257988 48816 258040 48822
rect 257988 48758 258040 48764
rect 257896 15904 257948 15910
rect 257896 15846 257948 15852
rect 258000 4078 258028 48758
rect 259196 46238 259224 52020
rect 260392 49162 260420 52020
rect 261602 52006 262168 52034
rect 260380 49156 260432 49162
rect 260380 49098 260432 49104
rect 259184 46232 259236 46238
rect 259184 46174 259236 46180
rect 259460 44940 259512 44946
rect 259460 44882 259512 44888
rect 258080 17264 258132 17270
rect 258080 17206 258132 17212
rect 257988 4072 258040 4078
rect 257988 4014 258040 4020
rect 258092 3482 258120 17206
rect 259472 3482 259500 44882
rect 262140 17270 262168 52006
rect 262784 47666 262812 52020
rect 263980 48822 264008 52020
rect 265176 48822 265204 52020
rect 266372 48822 266400 52020
rect 267476 49094 267504 52020
rect 268686 52006 269068 52034
rect 269882 52006 270448 52034
rect 267464 49088 267516 49094
rect 267464 49030 267516 49036
rect 263968 48816 264020 48822
rect 263968 48758 264020 48764
rect 264888 48816 264940 48822
rect 264888 48758 264940 48764
rect 265164 48816 265216 48822
rect 265164 48758 265216 48764
rect 266268 48816 266320 48822
rect 266268 48758 266320 48764
rect 266360 48816 266412 48822
rect 266360 48758 266412 48764
rect 267648 48816 267700 48822
rect 267648 48758 267700 48764
rect 262772 47660 262824 47666
rect 262772 47602 262824 47608
rect 262220 46300 262272 46306
rect 262220 46242 262272 46248
rect 262128 17264 262180 17270
rect 262128 17206 262180 17212
rect 262232 3806 262260 46242
rect 262312 18624 262364 18630
rect 262312 18566 262364 18572
rect 261024 3800 261076 3806
rect 261024 3742 261076 3748
rect 262220 3800 262272 3806
rect 262220 3742 262272 3748
rect 258092 3454 258672 3482
rect 259472 3454 259868 3482
rect 253848 3324 253900 3330
rect 253952 3318 255084 3346
rect 255332 3318 256280 3346
rect 253848 3266 253900 3272
rect 253860 480 253888 3266
rect 255056 480 255084 3318
rect 256252 480 256280 3318
rect 257436 3256 257488 3262
rect 257436 3198 257488 3204
rect 257448 480 257476 3198
rect 258644 480 258672 3454
rect 259840 480 259868 3454
rect 261036 480 261064 3742
rect 262324 3482 262352 18566
rect 264900 4010 264928 48758
rect 264980 21412 265032 21418
rect 264980 21354 265032 21360
rect 264888 4004 264940 4010
rect 264888 3946 264940 3952
rect 263416 3800 263468 3806
rect 263416 3742 263468 3748
rect 262232 3454 262352 3482
rect 262232 480 262260 3454
rect 263428 480 263456 3742
rect 264992 3482 265020 21354
rect 266280 18630 266308 48758
rect 266360 47592 266412 47598
rect 266360 47534 266412 47540
rect 266268 18624 266320 18630
rect 266268 18566 266320 18572
rect 266372 3482 266400 47534
rect 267660 31142 267688 48758
rect 267648 31136 267700 31142
rect 267648 31078 267700 31084
rect 269040 21418 269068 52006
rect 270420 32434 270448 52006
rect 270500 49360 270552 49366
rect 270500 49302 270552 49308
rect 270408 32428 270460 32434
rect 270408 32370 270460 32376
rect 269028 21412 269080 21418
rect 269028 21354 269080 21360
rect 269120 19984 269172 19990
rect 269120 19926 269172 19932
rect 268108 3868 268160 3874
rect 268108 3810 268160 3816
rect 264992 3454 265848 3482
rect 266372 3454 267044 3482
rect 264612 3052 264664 3058
rect 264612 2994 264664 3000
rect 264624 480 264652 2994
rect 265820 480 265848 3454
rect 267016 480 267044 3454
rect 268120 480 268148 3810
rect 269132 3482 269160 19926
rect 269132 3454 269344 3482
rect 269316 480 269344 3454
rect 270512 3330 270540 49302
rect 271064 48754 271092 52020
rect 272260 48822 272288 52020
rect 273456 48822 273484 52020
rect 274652 48822 274680 52020
rect 275862 52006 275968 52034
rect 277058 52006 277348 52034
rect 278254 52006 278728 52034
rect 279450 52006 280108 52034
rect 272248 48816 272300 48822
rect 272248 48758 272300 48764
rect 273168 48816 273220 48822
rect 273168 48758 273220 48764
rect 273444 48816 273496 48822
rect 273444 48758 273496 48764
rect 274548 48816 274600 48822
rect 274548 48758 274600 48764
rect 274640 48816 274692 48822
rect 274640 48758 274692 48764
rect 275836 48816 275888 48822
rect 275836 48758 275888 48764
rect 271052 48748 271104 48754
rect 271052 48690 271104 48696
rect 272524 48748 272576 48754
rect 272524 48690 272576 48696
rect 272536 28354 272564 48690
rect 272524 28348 272576 28354
rect 272524 28290 272576 28296
rect 271880 22772 271932 22778
rect 271880 22714 271932 22720
rect 270592 6180 270644 6186
rect 270592 6122 270644 6128
rect 270500 3324 270552 3330
rect 270500 3266 270552 3272
rect 270604 3210 270632 6122
rect 271892 3482 271920 22714
rect 273180 19990 273208 48758
rect 274560 33930 274588 48758
rect 274548 33924 274600 33930
rect 274548 33866 274600 33872
rect 273260 29776 273312 29782
rect 273260 29718 273312 29724
rect 273168 19984 273220 19990
rect 273168 19926 273220 19932
rect 273272 3482 273300 29718
rect 275848 26994 275876 48758
rect 275836 26988 275888 26994
rect 275836 26930 275888 26936
rect 275940 22846 275968 52006
rect 277320 35222 277348 52006
rect 277308 35216 277360 35222
rect 277308 35158 277360 35164
rect 277400 31068 277452 31074
rect 277400 31010 277452 31016
rect 276020 24132 276072 24138
rect 276020 24074 276072 24080
rect 275928 22840 275980 22846
rect 275928 22782 275980 22788
rect 275284 3936 275336 3942
rect 275284 3878 275336 3884
rect 271892 3454 272932 3482
rect 273272 3454 274128 3482
rect 271696 3324 271748 3330
rect 271696 3266 271748 3272
rect 270512 3182 270632 3210
rect 270512 480 270540 3182
rect 271708 480 271736 3266
rect 272904 480 272932 3454
rect 274100 480 274128 3454
rect 275296 480 275324 3878
rect 276032 3482 276060 24074
rect 276032 3454 276520 3482
rect 276492 480 276520 3454
rect 277412 3346 277440 31010
rect 278700 24206 278728 52006
rect 278964 49224 279016 49230
rect 278964 49166 279016 49172
rect 278688 24200 278740 24206
rect 278688 24142 278740 24148
rect 277412 3318 277716 3346
rect 277688 480 277716 3318
rect 278976 2496 279004 49166
rect 279976 6248 280028 6254
rect 279976 6190 280028 6196
rect 279988 6066 280016 6190
rect 280080 6186 280108 52006
rect 280632 48822 280660 52020
rect 281828 48822 281856 52020
rect 283024 48822 283052 52020
rect 284128 52006 284234 52034
rect 285430 52006 285628 52034
rect 286626 52006 287008 52034
rect 287822 52006 288388 52034
rect 289018 52006 289768 52034
rect 280620 48816 280672 48822
rect 280620 48758 280672 48764
rect 281448 48816 281500 48822
rect 281448 48758 281500 48764
rect 281816 48816 281868 48822
rect 281816 48758 281868 48764
rect 282828 48816 282880 48822
rect 282828 48758 282880 48764
rect 283012 48816 283064 48822
rect 283012 48758 283064 48764
rect 281460 36650 281488 48758
rect 281448 36644 281500 36650
rect 281448 36586 281500 36592
rect 280160 32496 280212 32502
rect 280160 32438 280212 32444
rect 280068 6180 280120 6186
rect 280068 6122 280120 6128
rect 279988 6038 280108 6066
rect 278884 2468 279004 2496
rect 278884 480 278912 2468
rect 280080 480 280108 6038
rect 280172 3346 280200 32438
rect 282840 6254 282868 48758
rect 284128 37942 284156 52006
rect 284208 48816 284260 48822
rect 284208 48758 284260 48764
rect 284116 37936 284168 37942
rect 284116 37878 284168 37884
rect 284220 7614 284248 48758
rect 284300 33856 284352 33862
rect 284300 33798 284352 33804
rect 283656 7608 283708 7614
rect 283656 7550 283708 7556
rect 284208 7608 284260 7614
rect 284208 7550 284260 7556
rect 282828 6248 282880 6254
rect 282828 6190 282880 6196
rect 282460 3732 282512 3738
rect 282460 3674 282512 3680
rect 280172 3318 281304 3346
rect 281276 480 281304 3318
rect 282472 480 282500 3674
rect 283668 480 283696 7550
rect 284312 3346 284340 33798
rect 285600 22778 285628 52006
rect 285772 49020 285824 49026
rect 285772 48962 285824 48968
rect 285588 22772 285640 22778
rect 285588 22714 285640 22720
rect 285784 3346 285812 48962
rect 286980 24138 287008 52006
rect 288360 39506 288388 52006
rect 288348 39500 288400 39506
rect 288348 39442 288400 39448
rect 287060 35284 287112 35290
rect 287060 35226 287112 35232
rect 286968 24132 287020 24138
rect 286968 24074 287020 24080
rect 284312 3318 284800 3346
rect 285784 3318 285996 3346
rect 284772 480 284800 3318
rect 285968 480 285996 3318
rect 287072 2514 287100 35226
rect 287152 25560 287204 25566
rect 287152 25502 287204 25508
rect 287060 2508 287112 2514
rect 287060 2450 287112 2456
rect 287164 480 287192 25502
rect 289740 3874 289768 52006
rect 290200 48482 290228 52020
rect 291396 48822 291424 52020
rect 292592 48822 292620 52020
rect 293710 52006 293816 52034
rect 294906 52006 295288 52034
rect 296102 52006 296668 52034
rect 297298 52006 298048 52034
rect 291384 48816 291436 48822
rect 291384 48758 291436 48764
rect 292488 48816 292540 48822
rect 292488 48758 292540 48764
rect 292580 48816 292632 48822
rect 292580 48758 292632 48764
rect 290188 48476 290240 48482
rect 290188 48418 290240 48424
rect 291108 48476 291160 48482
rect 291108 48418 291160 48424
rect 291120 9042 291148 48418
rect 292500 40798 292528 48758
rect 292488 40792 292540 40798
rect 292488 40734 292540 40740
rect 291200 36576 291252 36582
rect 291200 36518 291252 36524
rect 290740 9036 290792 9042
rect 290740 8978 290792 8984
rect 291108 9036 291160 9042
rect 291108 8978 291160 8984
rect 289728 3868 289780 3874
rect 289728 3810 289780 3816
rect 289544 3392 289596 3398
rect 289544 3334 289596 3340
rect 288348 2508 288400 2514
rect 288348 2450 288400 2456
rect 288360 480 288388 2450
rect 289556 480 289584 3334
rect 290752 480 290780 8978
rect 291212 3346 291240 36518
rect 293788 25566 293816 52006
rect 293868 48816 293920 48822
rect 293868 48758 293920 48764
rect 293776 25560 293828 25566
rect 293776 25502 293828 25508
rect 293880 3942 293908 48758
rect 293960 10328 294012 10334
rect 293960 10270 294012 10276
rect 293868 3936 293920 3942
rect 293868 3878 293920 3884
rect 293132 3460 293184 3466
rect 293132 3402 293184 3408
rect 291212 3318 291976 3346
rect 291948 480 291976 3318
rect 293144 480 293172 3402
rect 293972 3346 294000 10270
rect 295260 4826 295288 52006
rect 295340 38004 295392 38010
rect 295340 37946 295392 37952
rect 295248 4820 295300 4826
rect 295248 4762 295300 4768
rect 295352 3346 295380 37946
rect 296640 3806 296668 52006
rect 296812 26920 296864 26926
rect 296812 26862 296864 26868
rect 296628 3800 296680 3806
rect 296628 3742 296680 3748
rect 296720 3528 296772 3534
rect 296720 3470 296772 3476
rect 296824 3482 296852 26862
rect 298020 10402 298048 52006
rect 298480 48482 298508 52020
rect 299676 48822 299704 52020
rect 300872 48822 300900 52020
rect 299664 48816 299716 48822
rect 299664 48758 299716 48764
rect 300768 48816 300820 48822
rect 300768 48758 300820 48764
rect 300860 48816 300912 48822
rect 300860 48758 300912 48764
rect 298468 48476 298520 48482
rect 298468 48418 298520 48424
rect 299388 48476 299440 48482
rect 299388 48418 299440 48424
rect 299400 42090 299428 48418
rect 299388 42084 299440 42090
rect 299388 42026 299440 42032
rect 298100 39364 298152 39370
rect 298100 39306 298152 39312
rect 298008 10396 298060 10402
rect 298008 10338 298060 10344
rect 298112 3482 298140 39306
rect 300780 3738 300808 48758
rect 302068 43518 302096 52020
rect 303278 52006 303568 52034
rect 304474 52006 304948 52034
rect 305670 52006 306328 52034
rect 302148 48816 302200 48822
rect 302148 48758 302200 48764
rect 302056 43512 302108 43518
rect 302056 43454 302108 43460
rect 302160 11762 302188 48758
rect 302240 40724 302292 40730
rect 302240 40666 302292 40672
rect 300860 11756 300912 11762
rect 300860 11698 300912 11704
rect 302148 11756 302200 11762
rect 302148 11698 302200 11704
rect 300768 3732 300820 3738
rect 300768 3674 300820 3680
rect 300872 3482 300900 11698
rect 302252 3482 302280 40666
rect 303540 10334 303568 52006
rect 304920 14482 304948 52006
rect 305000 42152 305052 42158
rect 305000 42094 305052 42100
rect 304908 14476 304960 14482
rect 304908 14418 304960 14424
rect 303528 10328 303580 10334
rect 303528 10270 303580 10276
rect 303804 3596 303856 3602
rect 303804 3538 303856 3544
rect 293972 3318 294368 3346
rect 295352 3318 295564 3346
rect 294340 480 294368 3318
rect 295536 480 295564 3318
rect 296732 480 296760 3470
rect 296824 3454 297956 3482
rect 298112 3454 299152 3482
rect 300872 3454 301452 3482
rect 302252 3454 302648 3482
rect 297928 480 297956 3454
rect 299124 480 299152 3454
rect 300308 3188 300360 3194
rect 300308 3130 300360 3136
rect 300320 480 300348 3130
rect 301424 480 301452 3454
rect 302620 480 302648 3454
rect 303816 480 303844 3538
rect 305012 3534 305040 42094
rect 306300 29714 306328 52006
rect 306852 48822 306880 52020
rect 306840 48816 306892 48822
rect 306840 48758 306892 48764
rect 307668 48816 307720 48822
rect 307668 48758 307720 48764
rect 306288 29708 306340 29714
rect 306288 29650 306340 29656
rect 305092 28280 305144 28286
rect 305092 28222 305144 28228
rect 305000 3528 305052 3534
rect 305000 3470 305052 3476
rect 305104 1578 305132 28222
rect 307680 4146 307708 48758
rect 308048 48618 308076 52020
rect 309244 48822 309272 52020
rect 309232 48816 309284 48822
rect 309232 48758 309284 48764
rect 310336 48816 310388 48822
rect 310336 48758 310388 48764
rect 308036 48612 308088 48618
rect 308036 48554 308088 48560
rect 309048 48612 309100 48618
rect 309048 48554 309100 48560
rect 307760 14544 307812 14550
rect 307760 14486 307812 14492
rect 307392 4140 307444 4146
rect 307392 4082 307444 4088
rect 307668 4140 307720 4146
rect 307668 4082 307720 4088
rect 306196 3528 306248 3534
rect 306196 3470 306248 3476
rect 305012 1550 305132 1578
rect 305012 480 305040 1550
rect 306208 480 306236 3470
rect 307404 480 307432 4082
rect 307772 3346 307800 14486
rect 309060 13190 309088 48554
rect 310348 44878 310376 48758
rect 310336 44872 310388 44878
rect 310336 44814 310388 44820
rect 309140 43444 309192 43450
rect 309140 43386 309192 43392
rect 309048 13184 309100 13190
rect 309048 13126 309100 13132
rect 309152 3346 309180 43386
rect 310440 3602 310468 52020
rect 311650 52006 311848 52034
rect 311820 26926 311848 52006
rect 312832 46306 312860 52020
rect 314042 52006 314608 52034
rect 313464 49292 313516 49298
rect 313464 49234 313516 49240
rect 312820 46300 312872 46306
rect 312820 46242 312872 46248
rect 313372 29640 313424 29646
rect 313372 29582 313424 29588
rect 311808 26920 311860 26926
rect 311808 26862 311860 26868
rect 311900 13116 311952 13122
rect 311900 13058 311952 13064
rect 310980 3664 311032 3670
rect 310980 3606 311032 3612
rect 310428 3596 310480 3602
rect 310428 3538 310480 3544
rect 307772 3318 308628 3346
rect 309152 3318 309824 3346
rect 308600 480 308628 3318
rect 309796 480 309824 3318
rect 310992 480 311020 3606
rect 311912 3346 311940 13058
rect 311912 3318 312216 3346
rect 312188 480 312216 3318
rect 313384 480 313412 29582
rect 313476 3346 313504 49234
rect 314580 3602 314608 52006
rect 315224 48754 315252 52020
rect 315212 48748 315264 48754
rect 315212 48690 315264 48696
rect 315948 48748 316000 48754
rect 315948 48690 316000 48696
rect 315960 15978 315988 48690
rect 316420 47598 316448 52020
rect 317616 48346 317644 52020
rect 318720 49026 318748 52020
rect 319930 52006 320128 52034
rect 321126 52006 321508 52034
rect 322322 52006 322888 52034
rect 318708 49020 318760 49026
rect 318708 48962 318760 48968
rect 317604 48340 317656 48346
rect 317604 48282 317656 48288
rect 318708 48340 318760 48346
rect 318708 48282 318760 48288
rect 316408 47592 316460 47598
rect 316408 47534 316460 47540
rect 316040 45008 316092 45014
rect 316040 44950 316092 44956
rect 315948 15972 316000 15978
rect 315948 15914 316000 15920
rect 315764 4888 315816 4894
rect 315764 4830 315816 4836
rect 314568 3596 314620 3602
rect 314568 3538 314620 3544
rect 313476 3318 314608 3346
rect 314580 480 314608 3318
rect 315776 480 315804 4830
rect 316052 3346 316080 44950
rect 318064 4072 318116 4078
rect 318064 4014 318116 4020
rect 316052 3318 317000 3346
rect 316972 480 317000 3318
rect 318076 480 318104 4014
rect 318720 3262 318748 48282
rect 320100 31074 320128 52006
rect 320180 46232 320232 46238
rect 320180 46174 320232 46180
rect 320088 31068 320140 31074
rect 320088 31010 320140 31016
rect 318800 15904 318852 15910
rect 318800 15846 318852 15852
rect 318812 3346 318840 15846
rect 320192 3346 320220 46174
rect 321480 3466 321508 52006
rect 321744 49156 321796 49162
rect 321744 49098 321796 49104
rect 321652 17264 321704 17270
rect 321652 17206 321704 17212
rect 321664 3602 321692 17206
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 321756 3482 321784 49098
rect 322860 28286 322888 52006
rect 323504 48822 323532 52020
rect 324700 48822 324728 52020
rect 325896 48822 325924 52020
rect 327092 48822 327120 52020
rect 328302 52006 328408 52034
rect 329498 52006 329788 52034
rect 330694 52006 331168 52034
rect 331890 52006 332548 52034
rect 323492 48816 323544 48822
rect 323492 48758 323544 48764
rect 324228 48816 324280 48822
rect 324228 48758 324280 48764
rect 324688 48816 324740 48822
rect 324688 48758 324740 48764
rect 325608 48816 325660 48822
rect 325608 48758 325660 48764
rect 325884 48816 325936 48822
rect 325884 48758 325936 48764
rect 326988 48816 327040 48822
rect 326988 48758 327040 48764
rect 327080 48816 327132 48822
rect 327080 48758 327132 48764
rect 328276 48816 328328 48822
rect 328276 48758 328328 48764
rect 322940 47660 322992 47666
rect 322940 47602 322992 47608
rect 322848 28280 322900 28286
rect 322848 28222 322900 28228
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 321468 3460 321520 3466
rect 321468 3402 321520 3408
rect 321664 3454 321784 3482
rect 318812 3318 319300 3346
rect 320192 3318 320496 3346
rect 318708 3256 318760 3262
rect 318708 3198 318760 3204
rect 319272 480 319300 3318
rect 320468 480 320496 3318
rect 321664 480 321692 3454
rect 322860 480 322888 3538
rect 322952 3346 322980 47602
rect 324240 32502 324268 48758
rect 324228 32496 324280 32502
rect 324228 32438 324280 32444
rect 325240 4004 325292 4010
rect 325240 3946 325292 3952
rect 322952 3318 324084 3346
rect 324056 480 324084 3318
rect 325252 480 325280 3946
rect 325620 2922 325648 48758
rect 325700 18624 325752 18630
rect 325700 18566 325752 18572
rect 325712 3346 325740 18566
rect 327000 17270 327028 48758
rect 328288 33794 328316 48758
rect 328276 33788 328328 33794
rect 328276 33730 328328 33736
rect 327080 31136 327132 31142
rect 327080 31078 327132 31084
rect 326988 17264 327040 17270
rect 326988 17206 327040 17212
rect 327092 3346 327120 31078
rect 328380 7070 328408 52006
rect 328552 49088 328604 49094
rect 328552 49030 328604 49036
rect 328368 7064 328420 7070
rect 328368 7006 328420 7012
rect 328564 3346 328592 49030
rect 329760 18630 329788 52006
rect 331140 35290 331168 52006
rect 331128 35284 331180 35290
rect 331128 35226 331180 35232
rect 331220 32428 331272 32434
rect 331220 32370 331272 32376
rect 329840 21412 329892 21418
rect 329840 21354 329892 21360
rect 329748 18624 329800 18630
rect 329748 18566 329800 18572
rect 329852 3346 329880 21354
rect 325712 3318 326476 3346
rect 327092 3318 327672 3346
rect 328564 3318 328868 3346
rect 329852 3318 330064 3346
rect 325608 2916 325660 2922
rect 325608 2858 325660 2864
rect 326448 480 326476 3318
rect 327644 480 327672 3318
rect 328840 480 328868 3318
rect 330036 480 330064 3318
rect 331232 480 331260 32370
rect 331312 28348 331364 28354
rect 331312 28290 331364 28296
rect 331324 12442 331352 28290
rect 331312 12436 331364 12442
rect 331312 12378 331364 12384
rect 332416 12436 332468 12442
rect 332416 12378 332468 12384
rect 332428 480 332456 12378
rect 332520 3398 332548 52006
rect 333072 48822 333100 52020
rect 334268 48822 334296 52020
rect 335464 48822 335492 52020
rect 336568 52006 336674 52034
rect 337870 52006 338068 52034
rect 339066 52006 339448 52034
rect 340262 52006 340828 52034
rect 341458 52006 342208 52034
rect 333060 48816 333112 48822
rect 333060 48758 333112 48764
rect 333888 48816 333940 48822
rect 333888 48758 333940 48764
rect 334256 48816 334308 48822
rect 334256 48758 334308 48764
rect 335268 48816 335320 48822
rect 335268 48758 335320 48764
rect 335452 48816 335504 48822
rect 335452 48758 335504 48764
rect 333900 19990 333928 48758
rect 335280 36582 335308 48758
rect 335268 36576 335320 36582
rect 335268 36518 335320 36524
rect 333980 33924 334032 33930
rect 333980 33866 334032 33872
rect 332600 19984 332652 19990
rect 332600 19926 332652 19932
rect 333888 19984 333940 19990
rect 333888 19926 333940 19932
rect 332612 12442 332640 19926
rect 333992 19310 334020 33866
rect 335360 26988 335412 26994
rect 335360 26930 335412 26936
rect 333980 19304 334032 19310
rect 333980 19246 334032 19252
rect 335372 12442 335400 26930
rect 336568 21418 336596 52006
rect 336648 48816 336700 48822
rect 336648 48758 336700 48764
rect 336556 21412 336608 21418
rect 336556 21354 336608 21360
rect 332600 12436 332652 12442
rect 332600 12378 332652 12384
rect 333612 12436 333664 12442
rect 333612 12378 333664 12384
rect 335360 12436 335412 12442
rect 335360 12378 335412 12384
rect 335912 12436 335964 12442
rect 335912 12378 335964 12384
rect 332508 3392 332560 3398
rect 332508 3334 332560 3340
rect 333624 480 333652 12378
rect 334716 9716 334768 9722
rect 334716 9658 334768 9664
rect 334728 480 334756 9658
rect 335924 480 335952 12378
rect 336660 4078 336688 48758
rect 338040 38010 338068 52006
rect 338028 38004 338080 38010
rect 338028 37946 338080 37952
rect 338120 35216 338172 35222
rect 338120 35158 338172 35164
rect 336740 22840 336792 22846
rect 336740 22782 336792 22788
rect 336752 12510 336780 22782
rect 338132 12510 338160 35158
rect 336740 12504 336792 12510
rect 336740 12446 336792 12452
rect 338120 12504 338172 12510
rect 338120 12446 338172 12452
rect 337108 12368 337160 12374
rect 337108 12310 337160 12316
rect 338304 12368 338356 12374
rect 338304 12310 338356 12316
rect 336648 4072 336700 4078
rect 336648 4014 336700 4020
rect 337120 480 337148 12310
rect 338316 480 338344 12310
rect 339420 3369 339448 52006
rect 339500 24200 339552 24206
rect 339500 24142 339552 24148
rect 339406 3360 339462 3369
rect 339406 3295 339462 3304
rect 339512 480 339540 24142
rect 340800 7682 340828 52006
rect 342180 39438 342208 52006
rect 342640 48822 342668 52020
rect 343744 48822 343772 52020
rect 344940 49094 344968 52020
rect 346136 49162 346164 52020
rect 347346 52006 347728 52034
rect 348542 52006 349108 52034
rect 349738 52006 350488 52034
rect 346124 49156 346176 49162
rect 346124 49098 346176 49104
rect 344928 49088 344980 49094
rect 344928 49030 344980 49036
rect 345664 49020 345716 49026
rect 345664 48962 345716 48968
rect 342628 48816 342680 48822
rect 342628 48758 342680 48764
rect 343548 48816 343600 48822
rect 343548 48758 343600 48764
rect 343732 48816 343784 48822
rect 343732 48758 343784 48764
rect 344928 48816 344980 48822
rect 344928 48758 344980 48764
rect 342168 39432 342220 39438
rect 342168 39374 342220 39380
rect 340880 36644 340932 36650
rect 340880 36586 340932 36592
rect 340892 12442 340920 36586
rect 340880 12436 340932 12442
rect 340880 12378 340932 12384
rect 341892 12436 341944 12442
rect 341892 12378 341944 12384
rect 340788 7676 340840 7682
rect 340788 7618 340840 7624
rect 340696 6180 340748 6186
rect 340696 6122 340748 6128
rect 340708 480 340736 6122
rect 341904 480 341932 12378
rect 343088 6248 343140 6254
rect 343088 6190 343140 6196
rect 343100 480 343128 6190
rect 343560 4010 343588 48758
rect 344940 22846 344968 48758
rect 345020 37936 345072 37942
rect 345020 37878 345072 37884
rect 344928 22840 344980 22846
rect 344928 22782 344980 22788
rect 345032 19310 345060 37878
rect 345020 19304 345072 19310
rect 345020 19246 345072 19252
rect 345480 9716 345532 9722
rect 345480 9658 345532 9664
rect 344284 7608 344336 7614
rect 344284 7550 344336 7556
rect 343548 4004 343600 4010
rect 343548 3946 343600 3952
rect 344296 480 344324 7550
rect 345492 480 345520 9658
rect 345676 6186 345704 48962
rect 346400 22772 346452 22778
rect 346400 22714 346452 22720
rect 346412 12510 346440 22714
rect 346400 12504 346452 12510
rect 346400 12446 346452 12452
rect 346676 12368 346728 12374
rect 346676 12310 346728 12316
rect 345664 6180 345716 6186
rect 345664 6122 345716 6128
rect 346688 480 346716 12310
rect 347700 8974 347728 52006
rect 349080 40730 349108 52006
rect 349068 40724 349120 40730
rect 349068 40666 349120 40672
rect 347780 39500 347832 39506
rect 347780 39442 347832 39448
rect 347688 8968 347740 8974
rect 347688 8910 347740 8916
rect 347792 7614 347820 39442
rect 347872 24132 347924 24138
rect 347872 24074 347924 24080
rect 347780 7608 347832 7614
rect 347780 7550 347832 7556
rect 347884 480 347912 24074
rect 349068 7608 349120 7614
rect 349068 7550 349120 7556
rect 349080 480 349108 7550
rect 350264 3868 350316 3874
rect 350264 3810 350316 3816
rect 350276 480 350304 3810
rect 350460 3194 350488 52006
rect 350920 48822 350948 52020
rect 351184 49088 351236 49094
rect 351184 49030 351236 49036
rect 350908 48816 350960 48822
rect 350908 48758 350960 48764
rect 351196 11830 351224 49030
rect 352116 48822 352144 52020
rect 353312 48822 353340 52020
rect 354508 49026 354536 52020
rect 355718 52006 356008 52034
rect 356914 52006 357388 52034
rect 358110 52006 358768 52034
rect 354496 49020 354548 49026
rect 354496 48962 354548 48968
rect 351828 48816 351880 48822
rect 351828 48758 351880 48764
rect 352104 48816 352156 48822
rect 352104 48758 352156 48764
rect 353208 48816 353260 48822
rect 353208 48758 353260 48764
rect 353300 48816 353352 48822
rect 353300 48758 353352 48764
rect 354588 48816 354640 48822
rect 354588 48758 354640 48764
rect 351840 24138 351868 48758
rect 351920 40792 351972 40798
rect 351920 40734 351972 40740
rect 351828 24132 351880 24138
rect 351828 24074 351880 24080
rect 351932 12442 351960 40734
rect 353220 25634 353248 48758
rect 353208 25628 353260 25634
rect 353208 25570 353260 25576
rect 351920 12436 351972 12442
rect 351920 12378 351972 12384
rect 352564 12436 352616 12442
rect 352564 12378 352616 12384
rect 351184 11824 351236 11830
rect 351184 11766 351236 11772
rect 351368 9036 351420 9042
rect 351368 8978 351420 8984
rect 350448 3188 350500 3194
rect 350448 3130 350500 3136
rect 351380 480 351408 8978
rect 352576 480 352604 12378
rect 353760 3936 353812 3942
rect 353760 3878 353812 3884
rect 353772 480 353800 3878
rect 354600 3126 354628 48758
rect 354680 25560 354732 25566
rect 354680 25502 354732 25508
rect 354588 3120 354640 3126
rect 354588 3062 354640 3068
rect 354692 610 354720 25502
rect 355980 14550 356008 52006
rect 355968 14544 356020 14550
rect 355968 14486 356020 14492
rect 357360 7698 357388 52006
rect 357440 10396 357492 10402
rect 357440 10338 357492 10344
rect 357176 7670 357388 7698
rect 356152 4820 356204 4826
rect 356152 4762 356204 4768
rect 354680 604 354732 610
rect 354680 546 354732 552
rect 354956 604 355008 610
rect 354956 546 355008 552
rect 354968 480 354996 546
rect 356164 480 356192 4762
rect 357176 2990 357204 7670
rect 357348 3800 357400 3806
rect 357348 3742 357400 3748
rect 357164 2984 357216 2990
rect 357164 2926 357216 2932
rect 357360 480 357388 3742
rect 357452 610 357480 10338
rect 358740 5438 358768 52006
rect 359292 48822 359320 52020
rect 360488 48822 360516 52020
rect 361684 48822 361712 52020
rect 362788 52006 362894 52034
rect 364090 52006 364288 52034
rect 365286 52006 365668 52034
rect 366482 52006 367048 52034
rect 359280 48816 359332 48822
rect 359280 48758 359332 48764
rect 360108 48816 360160 48822
rect 360108 48758 360160 48764
rect 360476 48816 360528 48822
rect 360476 48758 360528 48764
rect 361488 48816 361540 48822
rect 361488 48758 361540 48764
rect 361672 48816 361724 48822
rect 361672 48758 361724 48764
rect 360120 42158 360148 48758
rect 360108 42152 360160 42158
rect 360108 42094 360160 42100
rect 358820 42084 358872 42090
rect 358820 42026 358872 42032
rect 358728 5432 358780 5438
rect 358728 5374 358780 5380
rect 358832 610 358860 42026
rect 360936 3732 360988 3738
rect 360936 3674 360988 3680
rect 357440 604 357492 610
rect 357440 546 357492 552
rect 358544 604 358596 610
rect 358544 546 358596 552
rect 358820 604 358872 610
rect 358820 546 358872 552
rect 359740 604 359792 610
rect 359740 546 359792 552
rect 358556 480 358584 546
rect 359752 480 359780 546
rect 360948 480 360976 3674
rect 361500 3058 361528 48758
rect 362788 43450 362816 52006
rect 362868 48816 362920 48822
rect 362868 48758 362920 48764
rect 362776 43444 362828 43450
rect 362776 43386 362828 43392
rect 361580 11756 361632 11762
rect 361580 11698 361632 11704
rect 361488 3052 361540 3058
rect 361488 2994 361540 3000
rect 361592 610 361620 11698
rect 362880 5030 362908 48758
rect 362960 43512 363012 43518
rect 362960 43454 363012 43460
rect 362868 5024 362920 5030
rect 362868 4966 362920 4972
rect 362972 626 363000 43454
rect 364260 3505 364288 52006
rect 364524 10328 364576 10334
rect 364524 10270 364576 10276
rect 364246 3496 364302 3505
rect 364246 3431 364302 3440
rect 361580 604 361632 610
rect 361580 546 361632 552
rect 362132 604 362184 610
rect 362972 598 363368 626
rect 362132 546 362184 552
rect 362144 480 362172 546
rect 363340 480 363368 598
rect 364536 480 364564 10270
rect 365640 5166 365668 52006
rect 365720 29708 365772 29714
rect 365720 29650 365772 29656
rect 365732 7614 365760 29650
rect 367020 29646 367048 52006
rect 367664 49298 367692 52020
rect 367652 49292 367704 49298
rect 367652 49234 367704 49240
rect 367744 49020 367796 49026
rect 367744 48962 367796 48968
rect 367008 29640 367060 29646
rect 367008 29582 367060 29588
rect 365812 14476 365864 14482
rect 365812 14418 365864 14424
rect 365720 7608 365772 7614
rect 365720 7550 365772 7556
rect 365628 5160 365680 5166
rect 365628 5102 365680 5108
rect 365824 1442 365852 14418
rect 367756 10334 367784 48962
rect 368860 48618 368888 52020
rect 368848 48612 368900 48618
rect 368848 48554 368900 48560
rect 369768 48612 369820 48618
rect 369768 48554 369820 48560
rect 368480 13184 368532 13190
rect 368480 13126 368532 13132
rect 367744 10328 367796 10334
rect 367744 10270 367796 10276
rect 366916 7608 366968 7614
rect 366916 7550 366968 7556
rect 365732 1414 365852 1442
rect 365732 480 365760 1414
rect 366928 480 366956 7550
rect 368020 4140 368072 4146
rect 368020 4082 368072 4088
rect 368032 480 368060 4082
rect 368492 2854 368520 13126
rect 369780 5506 369808 48554
rect 369964 46238 369992 52020
rect 369952 46232 370004 46238
rect 369952 46174 370004 46180
rect 369860 44872 369912 44878
rect 369860 44814 369912 44820
rect 369872 38622 369900 44814
rect 369860 38616 369912 38622
rect 369860 38558 369912 38564
rect 369952 38616 370004 38622
rect 369952 38558 370004 38564
rect 369964 29050 369992 38558
rect 369872 29022 369992 29050
rect 369872 27606 369900 29022
rect 369860 27600 369912 27606
rect 369860 27542 369912 27548
rect 370504 27600 370556 27606
rect 370504 27542 370556 27548
rect 369768 5500 369820 5506
rect 369768 5442 369820 5448
rect 368480 2848 368532 2854
rect 368480 2790 368532 2796
rect 369216 2780 369268 2786
rect 369216 2722 369268 2728
rect 369228 480 369256 2722
rect 370516 610 370544 27542
rect 371160 3670 371188 52020
rect 372370 52006 372568 52034
rect 373566 52006 373948 52034
rect 372540 4894 372568 52006
rect 373920 26926 373948 52006
rect 374748 49230 374776 52020
rect 374736 49224 374788 49230
rect 374736 49166 374788 49172
rect 375944 48618 375972 52020
rect 377140 48822 377168 52020
rect 378336 48822 378364 52020
rect 379532 48890 379560 52020
rect 379520 48884 379572 48890
rect 379520 48826 379572 48832
rect 380728 48822 380756 52020
rect 381924 49026 381952 52020
rect 383134 52006 383608 52034
rect 384330 52006 384988 52034
rect 381912 49020 381964 49026
rect 381912 48962 381964 48968
rect 380808 48884 380860 48890
rect 380808 48826 380860 48832
rect 377128 48816 377180 48822
rect 377128 48758 377180 48764
rect 378048 48816 378100 48822
rect 378048 48758 378100 48764
rect 378324 48816 378376 48822
rect 378324 48758 378376 48764
rect 379428 48816 379480 48822
rect 379428 48758 379480 48764
rect 380716 48816 380768 48822
rect 380716 48758 380768 48764
rect 375932 48612 375984 48618
rect 375932 48554 375984 48560
rect 376668 48612 376720 48618
rect 376668 48554 376720 48560
rect 374092 46300 374144 46306
rect 374092 46242 374144 46248
rect 372620 26920 372672 26926
rect 372620 26862 372672 26868
rect 373908 26920 373960 26926
rect 373908 26862 373960 26868
rect 372632 19310 372660 26862
rect 372620 19304 372672 19310
rect 372620 19246 372672 19252
rect 372896 9716 372948 9722
rect 372896 9658 372948 9664
rect 372528 4888 372580 4894
rect 372528 4830 372580 4836
rect 371608 3732 371660 3738
rect 371608 3674 371660 3680
rect 371148 3664 371200 3670
rect 371148 3606 371200 3612
rect 370412 604 370464 610
rect 370412 546 370464 552
rect 370504 604 370556 610
rect 370504 546 370556 552
rect 370424 480 370452 546
rect 371620 480 371648 3674
rect 372908 610 372936 9658
rect 374104 4842 374132 46242
rect 375380 15972 375432 15978
rect 375380 15914 375432 15920
rect 374012 4814 374132 4842
rect 372804 604 372856 610
rect 372804 546 372856 552
rect 372896 604 372948 610
rect 372896 546 372948 552
rect 372816 480 372844 546
rect 374012 480 374040 4814
rect 375196 3324 375248 3330
rect 375196 3266 375248 3272
rect 375208 480 375236 3266
rect 375392 610 375420 15914
rect 376680 5098 376708 48554
rect 376760 47592 376812 47598
rect 376760 47534 376812 47540
rect 376668 5092 376720 5098
rect 376668 5034 376720 5040
rect 376772 610 376800 47534
rect 378060 31142 378088 48758
rect 378048 31136 378100 31142
rect 378048 31078 378100 31084
rect 379440 4146 379468 48758
rect 379980 6180 380032 6186
rect 379980 6122 380032 6128
rect 379428 4140 379480 4146
rect 379428 4082 379480 4088
rect 378784 3256 378836 3262
rect 378784 3198 378836 3204
rect 375380 604 375432 610
rect 375380 546 375432 552
rect 376392 604 376444 610
rect 376392 546 376444 552
rect 376760 604 376812 610
rect 376760 546 376812 552
rect 377588 604 377640 610
rect 377588 546 377640 552
rect 376404 480 376432 546
rect 377600 480 377628 546
rect 378796 480 378824 3198
rect 379992 480 380020 6122
rect 380820 5302 380848 48826
rect 381544 48816 381596 48822
rect 381544 48758 381596 48764
rect 380900 31068 380952 31074
rect 380900 31010 380952 31016
rect 380808 5296 380860 5302
rect 380808 5238 380860 5244
rect 380912 626 380940 31010
rect 381556 13122 381584 48758
rect 382372 28280 382424 28286
rect 382372 28222 382424 28228
rect 381544 13116 381596 13122
rect 381544 13058 381596 13064
rect 382384 4962 382412 28222
rect 383580 5234 383608 52006
rect 383660 32496 383712 32502
rect 383660 32438 383712 32444
rect 383568 5228 383620 5234
rect 383568 5170 383620 5176
rect 382372 4956 382424 4962
rect 382372 4898 382424 4904
rect 383568 4956 383620 4962
rect 383568 4898 383620 4904
rect 382280 3460 382332 3466
rect 382280 3402 382332 3408
rect 382292 3346 382320 3402
rect 382292 3318 382412 3346
rect 380912 598 381124 626
rect 381096 592 381124 598
rect 381096 564 381216 592
rect 381188 480 381216 564
rect 382384 480 382412 3318
rect 383580 480 383608 4898
rect 383672 610 383700 32438
rect 384960 32434 384988 52006
rect 385512 48754 385540 52020
rect 386708 48822 386736 52020
rect 387904 48822 387932 52020
rect 389100 49094 389128 52020
rect 390310 52006 390508 52034
rect 391506 52006 391888 52034
rect 392702 52006 393268 52034
rect 393898 52006 394648 52034
rect 389088 49088 389140 49094
rect 389088 49030 389140 49036
rect 386696 48816 386748 48822
rect 386696 48758 386748 48764
rect 387708 48816 387760 48822
rect 387708 48758 387760 48764
rect 387892 48816 387944 48822
rect 387892 48758 387944 48764
rect 389088 48816 389140 48822
rect 389088 48758 389140 48764
rect 385500 48748 385552 48754
rect 385500 48690 385552 48696
rect 386328 48748 386380 48754
rect 386328 48690 386380 48696
rect 384948 32428 385000 32434
rect 384948 32370 385000 32376
rect 386340 3874 386368 48690
rect 386420 17264 386472 17270
rect 386420 17206 386472 17212
rect 386328 3868 386380 3874
rect 386328 3810 386380 3816
rect 385868 2916 385920 2922
rect 385868 2858 385920 2864
rect 383660 604 383712 610
rect 383660 546 383712 552
rect 384672 604 384724 610
rect 384672 546 384724 552
rect 384684 480 384712 546
rect 385880 480 385908 2858
rect 386432 610 386460 17206
rect 387720 5370 387748 48758
rect 389100 35222 389128 48758
rect 389088 35216 389140 35222
rect 389088 35158 389140 35164
rect 387800 33788 387852 33794
rect 387800 33730 387852 33736
rect 387708 5364 387760 5370
rect 387708 5306 387760 5312
rect 387812 610 387840 33730
rect 390480 4758 390508 52006
rect 391860 36650 391888 52006
rect 391848 36644 391900 36650
rect 391848 36586 391900 36592
rect 390560 35284 390612 35290
rect 390560 35226 390612 35232
rect 390572 7614 390600 35226
rect 390652 18624 390704 18630
rect 390652 18566 390704 18572
rect 390560 7608 390612 7614
rect 390560 7550 390612 7556
rect 390468 4752 390520 4758
rect 390468 4694 390520 4700
rect 389456 3324 389508 3330
rect 389456 3266 389508 3272
rect 386420 604 386472 610
rect 386420 546 386472 552
rect 387064 604 387116 610
rect 387064 546 387116 552
rect 387800 604 387852 610
rect 387800 546 387852 552
rect 388260 604 388312 610
rect 388260 546 388312 552
rect 387076 480 387104 546
rect 388272 480 388300 546
rect 389468 480 389496 3266
rect 390664 480 390692 18566
rect 391848 7608 391900 7614
rect 391848 7550 391900 7556
rect 391860 480 391888 7550
rect 393240 3942 393268 52006
rect 393320 19984 393372 19990
rect 393320 19926 393372 19932
rect 393332 12442 393360 19926
rect 393320 12436 393372 12442
rect 393320 12378 393372 12384
rect 394240 12436 394292 12442
rect 394240 12378 394292 12384
rect 393228 3936 393280 3942
rect 393228 3878 393280 3884
rect 393044 3392 393096 3398
rect 393044 3334 393096 3340
rect 393056 480 393084 3334
rect 394252 480 394280 12378
rect 394620 5370 394648 52006
rect 394988 48822 395016 52020
rect 396184 49366 396212 52020
rect 396172 49360 396224 49366
rect 396172 49302 396224 49308
rect 394976 48816 395028 48822
rect 394976 48758 395028 48764
rect 395988 48816 396040 48822
rect 395988 48758 396040 48764
rect 396000 37942 396028 48758
rect 395988 37936 396040 37942
rect 395988 37878 396040 37884
rect 394700 36576 394752 36582
rect 394700 36518 394752 36524
rect 394712 19310 394740 36518
rect 394700 19304 394752 19310
rect 394700 19246 394752 19252
rect 397380 15910 397408 52020
rect 398590 52006 398788 52034
rect 399786 52006 400168 52034
rect 400982 52006 401548 52034
rect 402178 52006 402928 52034
rect 398760 39370 398788 52006
rect 398748 39364 398800 39370
rect 398748 39306 398800 39312
rect 398840 37324 398892 37330
rect 398840 37266 398892 37272
rect 398852 27606 398880 37266
rect 398840 27600 398892 27606
rect 398840 27542 398892 27548
rect 397460 21412 397512 21418
rect 397460 21354 397512 21360
rect 397472 19310 397500 21354
rect 397460 19304 397512 19310
rect 397460 19246 397512 19252
rect 397368 15904 397420 15910
rect 397368 15846 397420 15852
rect 395436 9716 395488 9722
rect 395436 9658 395488 9664
rect 397828 9716 397880 9722
rect 397828 9658 397880 9664
rect 399024 9716 399076 9722
rect 399024 9658 399076 9664
rect 394608 5364 394660 5370
rect 394608 5306 394660 5312
rect 395448 480 395476 9658
rect 397840 9602 397868 9658
rect 397840 9574 397960 9602
rect 396632 4072 396684 4078
rect 396632 4014 396684 4020
rect 396644 480 396672 4014
rect 397932 610 397960 9574
rect 397828 604 397880 610
rect 397828 546 397880 552
rect 397920 604 397972 610
rect 397920 546 397972 552
rect 397840 480 397868 546
rect 399036 480 399064 9658
rect 400140 3806 400168 52006
rect 401520 17338 401548 52006
rect 402900 40798 402928 52006
rect 403360 49434 403388 52020
rect 403348 49428 403400 49434
rect 403348 49370 403400 49376
rect 404556 48822 404584 52020
rect 404544 48816 404596 48822
rect 404544 48758 404596 48764
rect 405648 48816 405700 48822
rect 405648 48758 405700 48764
rect 402888 40792 402940 40798
rect 402888 40734 402940 40740
rect 401600 39432 401652 39438
rect 401600 39374 401652 39380
rect 401508 17332 401560 17338
rect 401508 17274 401560 17280
rect 401612 12442 401640 39374
rect 404360 22840 404412 22846
rect 404360 22782 404412 22788
rect 404372 12442 404400 22782
rect 405660 18630 405688 48758
rect 405752 48550 405780 52020
rect 406962 52006 407068 52034
rect 408158 52006 408448 52034
rect 409354 52006 409828 52034
rect 410550 52006 411208 52034
rect 405740 48544 405792 48550
rect 405740 48486 405792 48492
rect 406936 48544 406988 48550
rect 406936 48486 406988 48492
rect 406948 42090 406976 48486
rect 406936 42084 406988 42090
rect 406936 42026 406988 42032
rect 405648 18624 405700 18630
rect 405648 18566 405700 18572
rect 401600 12436 401652 12442
rect 401600 12378 401652 12384
rect 402520 12436 402572 12442
rect 402520 12378 402572 12384
rect 404360 12436 404412 12442
rect 404360 12378 404412 12384
rect 404912 12436 404964 12442
rect 404912 12378 404964 12384
rect 401324 7676 401376 7682
rect 401324 7618 401376 7624
rect 400128 3800 400180 3806
rect 400128 3742 400180 3748
rect 400218 3360 400274 3369
rect 400218 3295 400274 3304
rect 400232 480 400260 3295
rect 401336 480 401364 7618
rect 402532 480 402560 12378
rect 403716 4004 403768 4010
rect 403716 3946 403768 3952
rect 403728 480 403756 3946
rect 404924 480 404952 12378
rect 406108 11824 406160 11830
rect 406108 11766 406160 11772
rect 406120 480 406148 11766
rect 407040 3369 407068 52006
rect 407212 49156 407264 49162
rect 407212 49098 407264 49104
rect 407224 46918 407252 49098
rect 407212 46912 407264 46918
rect 407212 46854 407264 46860
rect 407212 37324 407264 37330
rect 407212 37266 407264 37272
rect 407224 29170 407252 37266
rect 407212 29164 407264 29170
rect 407212 29106 407264 29112
rect 407212 29028 407264 29034
rect 407212 28970 407264 28976
rect 407224 27606 407252 28970
rect 407212 27600 407264 27606
rect 407212 27542 407264 27548
rect 408420 19990 408448 52006
rect 409800 43518 409828 52006
rect 409788 43512 409840 43518
rect 409788 43454 409840 43460
rect 408500 40724 408552 40730
rect 408500 40666 408552 40672
rect 408408 19984 408460 19990
rect 408408 19926 408460 19932
rect 407212 12300 407264 12306
rect 407212 12242 407264 12248
rect 407026 3360 407082 3369
rect 407026 3295 407082 3304
rect 407224 3176 407252 12242
rect 408512 7614 408540 40666
rect 408684 8968 408736 8974
rect 408684 8910 408736 8916
rect 408500 7608 408552 7614
rect 408500 7550 408552 7556
rect 408696 7426 408724 8910
rect 409696 7608 409748 7614
rect 409696 7550 409748 7556
rect 408512 7398 408724 7426
rect 407224 3148 407344 3176
rect 407316 480 407344 3148
rect 408512 480 408540 7398
rect 409708 480 409736 7550
rect 411180 3738 411208 52006
rect 411732 48822 411760 52020
rect 412928 48822 412956 52020
rect 414124 48822 414152 52020
rect 415228 52006 415334 52034
rect 416530 52006 416728 52034
rect 417726 52006 418108 52034
rect 418922 52006 419488 52034
rect 411720 48816 411772 48822
rect 411720 48758 411772 48764
rect 412548 48816 412600 48822
rect 412548 48758 412600 48764
rect 412916 48816 412968 48822
rect 412916 48758 412968 48764
rect 413928 48816 413980 48822
rect 413928 48758 413980 48764
rect 414112 48816 414164 48822
rect 414112 48758 414164 48764
rect 411260 24132 411312 24138
rect 411260 24074 411312 24080
rect 411272 9654 411300 24074
rect 412560 21418 412588 48758
rect 412640 25628 412692 25634
rect 412640 25570 412692 25576
rect 412548 21412 412600 21418
rect 412548 21354 412600 21360
rect 411260 9648 411312 9654
rect 411260 9590 411312 9596
rect 411168 3732 411220 3738
rect 411168 3674 411220 3680
rect 410892 3188 410944 3194
rect 410892 3130 410944 3136
rect 410904 480 410932 3130
rect 412652 2854 412680 25570
rect 413940 14482 413968 48758
rect 415228 44878 415256 52006
rect 415308 48816 415360 48822
rect 415308 48758 415360 48764
rect 415216 44872 415268 44878
rect 415216 44814 415268 44820
rect 413928 14476 413980 14482
rect 413928 14418 413980 14424
rect 415320 4010 415348 48758
rect 416700 11762 416728 52006
rect 416872 14544 416924 14550
rect 416872 14486 416924 14492
rect 416688 11756 416740 11762
rect 416688 11698 416740 11704
rect 415400 10328 415452 10334
rect 415400 10270 415452 10276
rect 415308 4004 415360 4010
rect 415308 3946 415360 3952
rect 414480 3120 414532 3126
rect 414480 3062 414532 3068
rect 412640 2848 412692 2854
rect 412640 2790 412692 2796
rect 413284 2780 413336 2786
rect 413284 2722 413336 2728
rect 412088 604 412140 610
rect 412088 546 412140 552
rect 412100 480 412128 546
rect 413296 480 413324 2722
rect 414492 480 414520 3062
rect 415412 1034 415440 10270
rect 415412 1006 415716 1034
rect 415688 480 415716 1006
rect 416884 480 416912 14486
rect 418080 3534 418108 52006
rect 419460 22778 419488 52006
rect 420104 48822 420132 52020
rect 421208 48822 421236 52020
rect 420092 48816 420144 48822
rect 420092 48758 420144 48764
rect 420828 48816 420880 48822
rect 420828 48758 420880 48764
rect 421196 48816 421248 48822
rect 421196 48758 421248 48764
rect 422208 48816 422260 48822
rect 422208 48758 422260 48764
rect 419540 42152 419592 42158
rect 419540 42094 419592 42100
rect 419448 22772 419500 22778
rect 419448 22714 419500 22720
rect 419552 9654 419580 42094
rect 420840 38010 420868 48758
rect 420828 38004 420880 38010
rect 420828 37946 420880 37952
rect 419540 9648 419592 9654
rect 419540 9590 419592 9596
rect 419172 5432 419224 5438
rect 419172 5374 419224 5380
rect 418068 3528 418120 3534
rect 418068 3470 418120 3476
rect 417976 2984 418028 2990
rect 417976 2926 418028 2932
rect 417988 480 418016 2926
rect 419184 480 419212 5374
rect 422220 3602 422248 48758
rect 422404 48346 422432 52020
rect 423508 52006 423614 52034
rect 424810 52006 425008 52034
rect 426006 52006 426388 52034
rect 427202 52006 427768 52034
rect 422392 48340 422444 48346
rect 422392 48282 422444 48288
rect 423508 24138 423536 52006
rect 423588 48340 423640 48346
rect 423588 48282 423640 48288
rect 423496 24132 423548 24138
rect 423496 24074 423548 24080
rect 423600 7614 423628 48282
rect 423680 43444 423732 43450
rect 423680 43386 423732 43392
rect 423588 7608 423640 7614
rect 423588 7550 423640 7556
rect 422760 5024 422812 5030
rect 422760 4966 422812 4972
rect 422208 3596 422260 3602
rect 422208 3538 422260 3544
rect 421564 3052 421616 3058
rect 421564 2994 421616 3000
rect 420368 604 420420 610
rect 420368 546 420420 552
rect 420380 480 420408 546
rect 421576 480 421604 2994
rect 422772 480 422800 4966
rect 423692 2854 423720 43386
rect 424980 40730 425008 52006
rect 424968 40724 425020 40730
rect 424968 40666 425020 40672
rect 426360 6186 426388 52006
rect 426440 29640 426492 29646
rect 426440 29582 426492 29588
rect 426348 6180 426400 6186
rect 426348 6122 426400 6128
rect 426348 5160 426400 5166
rect 426348 5102 426400 5108
rect 425150 3496 425206 3505
rect 425150 3431 425206 3440
rect 423680 2848 423732 2854
rect 423680 2790 423732 2796
rect 423956 2780 424008 2786
rect 423956 2722 424008 2728
rect 423968 480 423996 2722
rect 425164 480 425192 3431
rect 426360 480 426388 5102
rect 426452 2854 426480 29582
rect 427740 25566 427768 52006
rect 427912 49292 427964 49298
rect 427912 49234 427964 49240
rect 427728 25560 427780 25566
rect 427728 25502 427780 25508
rect 427924 2854 427952 49234
rect 428384 48822 428412 52020
rect 429580 48822 429608 52020
rect 430776 48822 430804 52020
rect 431972 48822 432000 52020
rect 433182 52006 433288 52034
rect 434378 52006 434668 52034
rect 435574 52006 436048 52034
rect 436770 52006 437428 52034
rect 428372 48816 428424 48822
rect 428372 48758 428424 48764
rect 429108 48816 429160 48822
rect 429108 48758 429160 48764
rect 429568 48816 429620 48822
rect 429568 48758 429620 48764
rect 430488 48816 430540 48822
rect 430488 48758 430540 48764
rect 430764 48816 430816 48822
rect 430764 48758 430816 48764
rect 431868 48816 431920 48822
rect 431868 48758 431920 48764
rect 431960 48816 432012 48822
rect 431960 48758 432012 48764
rect 433156 48816 433208 48822
rect 433156 48758 433208 48764
rect 429120 3466 429148 48758
rect 430500 8974 430528 48758
rect 430580 46232 430632 46238
rect 430580 46174 430632 46180
rect 430488 8968 430540 8974
rect 430488 8910 430540 8916
rect 429936 5500 429988 5506
rect 429936 5442 429988 5448
rect 429108 3460 429160 3466
rect 429108 3402 429160 3408
rect 426440 2848 426492 2854
rect 426440 2790 426492 2796
rect 427912 2848 427964 2854
rect 427912 2790 427964 2796
rect 427544 2780 427596 2786
rect 427544 2722 427596 2728
rect 427556 480 427584 2722
rect 428740 604 428792 610
rect 428740 546 428792 552
rect 428752 480 428780 546
rect 429948 480 429976 5442
rect 430592 4876 430620 46174
rect 431880 26994 431908 48758
rect 431868 26988 431920 26994
rect 431868 26930 431920 26936
rect 430500 4848 430620 4876
rect 430500 610 430528 4848
rect 432328 3664 432380 3670
rect 432328 3606 432380 3612
rect 430488 604 430540 610
rect 430488 546 430540 552
rect 431132 604 431184 610
rect 431132 546 431184 552
rect 431144 480 431172 546
rect 432340 480 432368 3606
rect 433168 3058 433196 48758
rect 433260 47598 433288 52006
rect 433248 47592 433300 47598
rect 433248 47534 433300 47540
rect 434640 28286 434668 52006
rect 434812 49224 434864 49230
rect 434812 49166 434864 49172
rect 434628 28280 434680 28286
rect 434628 28222 434680 28228
rect 433340 26920 433392 26926
rect 433340 26862 433392 26868
rect 433352 7682 433380 26862
rect 433340 7676 433392 7682
rect 433340 7618 433392 7624
rect 434628 7676 434680 7682
rect 434628 7618 434680 7624
rect 433524 4888 433576 4894
rect 433524 4830 433576 4836
rect 433156 3052 433208 3058
rect 433156 2994 433208 3000
rect 433536 480 433564 4830
rect 434640 480 434668 7618
rect 434824 2854 434852 49166
rect 436020 3670 436048 52006
rect 437400 10334 437428 52006
rect 437952 48822 437980 52020
rect 439148 48822 439176 52020
rect 440344 48822 440372 52020
rect 441448 52006 441554 52034
rect 442750 52006 442948 52034
rect 443946 52006 444328 52034
rect 445142 52006 445708 52034
rect 437940 48816 437992 48822
rect 437940 48758 437992 48764
rect 438768 48816 438820 48822
rect 438768 48758 438820 48764
rect 439136 48816 439188 48822
rect 439136 48758 439188 48764
rect 440148 48816 440200 48822
rect 440148 48758 440200 48764
rect 440332 48816 440384 48822
rect 440332 48758 440384 48764
rect 437480 31136 437532 31142
rect 437480 31078 437532 31084
rect 437388 10328 437440 10334
rect 437388 10270 437440 10276
rect 437020 5092 437072 5098
rect 437020 5034 437072 5040
rect 436008 3664 436060 3670
rect 436008 3606 436060 3612
rect 434812 2848 434864 2854
rect 434812 2790 434864 2796
rect 435824 604 435876 610
rect 435824 546 435876 552
rect 435836 480 435864 546
rect 437032 480 437060 5034
rect 437492 2854 437520 31078
rect 438780 29646 438808 48758
rect 438768 29640 438820 29646
rect 438768 29582 438820 29588
rect 439412 4140 439464 4146
rect 439412 4082 439464 4088
rect 437480 2848 437532 2854
rect 437480 2790 437532 2796
rect 438216 2780 438268 2786
rect 438216 2722 438268 2728
rect 438228 480 438256 2722
rect 439424 480 439452 4082
rect 440160 4078 440188 48758
rect 441448 33794 441476 52006
rect 441528 48816 441580 48822
rect 441528 48758 441580 48764
rect 441436 33788 441488 33794
rect 441436 33730 441488 33736
rect 441540 11830 441568 48758
rect 441620 13116 441672 13122
rect 441620 13058 441672 13064
rect 441528 11824 441580 11830
rect 441528 11766 441580 11772
rect 440608 5296 440660 5302
rect 440608 5238 440660 5244
rect 440148 4072 440200 4078
rect 440148 4014 440200 4020
rect 440620 480 440648 5238
rect 441632 2854 441660 13058
rect 442920 3262 442948 52006
rect 443184 49020 443236 49026
rect 443184 48962 443236 48968
rect 443196 46918 443224 48962
rect 443184 46912 443236 46918
rect 443184 46854 443236 46860
rect 443184 37324 443236 37330
rect 443184 37266 443236 37272
rect 443196 27606 443224 37266
rect 443184 27600 443236 27606
rect 443184 27542 443236 27548
rect 444300 13122 444328 52006
rect 444380 32428 444432 32434
rect 444380 32370 444432 32376
rect 444288 13116 444340 13122
rect 444288 13058 444340 13064
rect 443000 9716 443052 9722
rect 443000 9658 443052 9664
rect 442908 3256 442960 3262
rect 442908 3198 442960 3204
rect 441620 2848 441672 2854
rect 441620 2790 441672 2796
rect 441804 2780 441856 2786
rect 441804 2722 441856 2728
rect 441816 480 441844 2722
rect 443012 480 443040 9658
rect 444196 4956 444248 4962
rect 444196 4898 444248 4904
rect 444208 480 444236 4898
rect 444392 2854 444420 32370
rect 445680 31074 445708 52006
rect 446232 48822 446260 52020
rect 447428 48822 447456 52020
rect 448624 48822 448652 52020
rect 446220 48816 446272 48822
rect 446220 48758 446272 48764
rect 447048 48816 447100 48822
rect 447048 48758 447100 48764
rect 447416 48816 447468 48822
rect 447416 48758 447468 48764
rect 448428 48816 448480 48822
rect 448428 48758 448480 48764
rect 448612 48816 448664 48822
rect 448612 48758 448664 48764
rect 449716 48816 449768 48822
rect 449716 48758 449768 48764
rect 445668 31068 445720 31074
rect 445668 31010 445720 31016
rect 447060 3874 447088 48758
rect 448440 14550 448468 48758
rect 448520 35216 448572 35222
rect 448520 35158 448572 35164
rect 448428 14544 448480 14550
rect 448428 14486 448480 14492
rect 448532 12442 448560 35158
rect 449728 32434 449756 48758
rect 449716 32428 449768 32434
rect 449716 32370 449768 32376
rect 448520 12436 448572 12442
rect 448520 12378 448572 12384
rect 448980 12436 449032 12442
rect 448980 12378 449032 12384
rect 447784 5228 447836 5234
rect 447784 5170 447836 5176
rect 446588 3868 446640 3874
rect 446588 3810 446640 3816
rect 447048 3868 447100 3874
rect 447048 3810 447100 3816
rect 444380 2848 444432 2854
rect 444380 2790 444432 2796
rect 445392 2780 445444 2786
rect 445392 2722 445444 2728
rect 445404 480 445432 2722
rect 446600 480 446628 3810
rect 447796 480 447824 5170
rect 448992 480 449020 12378
rect 449820 3505 449848 52020
rect 449992 49088 450044 49094
rect 449992 49030 450044 49036
rect 450004 46918 450032 49030
rect 449992 46912 450044 46918
rect 449992 46854 450044 46860
rect 451016 46238 451044 52020
rect 452226 52006 452608 52034
rect 453422 52006 453988 52034
rect 454618 52006 455368 52034
rect 451004 46232 451056 46238
rect 451004 46174 451056 46180
rect 449992 37324 450044 37330
rect 449992 37266 450044 37272
rect 450004 27606 450032 37266
rect 451280 36644 451332 36650
rect 451280 36586 451332 36592
rect 449992 27600 450044 27606
rect 449992 27542 450044 27548
rect 450360 27600 450412 27606
rect 450360 27542 450412 27548
rect 449806 3496 449862 3505
rect 449806 3431 449862 3440
rect 450372 610 450400 27542
rect 451292 7682 451320 36586
rect 452580 17270 452608 52006
rect 452568 17264 452620 17270
rect 452568 17206 452620 17212
rect 451280 7676 451332 7682
rect 451280 7618 451332 7624
rect 452476 7676 452528 7682
rect 452476 7618 452528 7624
rect 451280 4684 451332 4690
rect 451280 4626 451332 4632
rect 450176 604 450228 610
rect 450176 546 450228 552
rect 450360 604 450412 610
rect 450360 546 450412 552
rect 450188 480 450216 546
rect 451292 480 451320 4626
rect 452488 480 452516 7618
rect 453960 3942 453988 52006
rect 454868 5364 454920 5370
rect 454868 5306 454920 5312
rect 453672 3936 453724 3942
rect 453672 3878 453724 3884
rect 453948 3936 454000 3942
rect 453948 3878 454000 3884
rect 453684 480 453712 3878
rect 454880 480 454908 5306
rect 455340 5030 455368 52006
rect 455800 48822 455828 52020
rect 456892 49360 456944 49366
rect 456892 49302 456944 49308
rect 455788 48816 455840 48822
rect 455788 48758 455840 48764
rect 456708 48816 456760 48822
rect 456708 48758 456760 48764
rect 455420 37936 455472 37942
rect 455420 37878 455472 37884
rect 455328 5024 455380 5030
rect 455328 4966 455380 4972
rect 455432 610 455460 37878
rect 456720 35222 456748 48758
rect 456708 35216 456760 35222
rect 456708 35158 456760 35164
rect 456904 610 456932 49302
rect 456996 48822 457024 52020
rect 458192 48822 458220 52020
rect 456984 48816 457036 48822
rect 456984 48758 457036 48764
rect 458088 48816 458140 48822
rect 458088 48758 458140 48764
rect 458180 48816 458232 48822
rect 458180 48758 458232 48764
rect 458100 3194 458128 48758
rect 459388 36582 459416 52020
rect 460598 52006 460888 52034
rect 461794 52006 462268 52034
rect 462990 52006 463648 52034
rect 459468 48816 459520 48822
rect 459468 48758 459520 48764
rect 459376 36576 459428 36582
rect 459376 36518 459428 36524
rect 458180 15904 458232 15910
rect 458180 15846 458232 15852
rect 458088 3188 458140 3194
rect 458088 3130 458140 3136
rect 458192 626 458220 15846
rect 459480 5302 459508 48758
rect 459652 39364 459704 39370
rect 459652 39306 459704 39312
rect 459468 5296 459520 5302
rect 459468 5238 459520 5244
rect 455420 604 455472 610
rect 455420 546 455472 552
rect 456064 604 456116 610
rect 456064 546 456116 552
rect 456892 604 456944 610
rect 456892 546 456944 552
rect 457260 604 457312 610
rect 458192 598 458496 626
rect 457260 546 457312 552
rect 456076 480 456104 546
rect 457272 480 457300 546
rect 458468 480 458496 598
rect 459664 480 459692 39306
rect 460860 4146 460888 52006
rect 460940 17332 460992 17338
rect 460940 17274 460992 17280
rect 460848 4140 460900 4146
rect 460848 4082 460900 4088
rect 460848 3800 460900 3806
rect 460848 3742 460900 3748
rect 460860 480 460888 3742
rect 460952 3346 460980 17274
rect 462240 5234 462268 52006
rect 462320 40792 462372 40798
rect 462320 40734 462372 40740
rect 462228 5228 462280 5234
rect 462228 5170 462280 5176
rect 462332 3346 462360 40734
rect 463620 5370 463648 52006
rect 463792 49428 463844 49434
rect 463792 49370 463844 49376
rect 463608 5364 463660 5370
rect 463608 5306 463660 5312
rect 463804 3346 463832 49370
rect 464172 48822 464200 52020
rect 465368 48822 465396 52020
rect 466564 48822 466592 52020
rect 467760 49026 467788 52020
rect 468970 52006 469168 52034
rect 470166 52006 470548 52034
rect 471362 52006 471928 52034
rect 467748 49020 467800 49026
rect 467748 48962 467800 48968
rect 464160 48816 464212 48822
rect 464160 48758 464212 48764
rect 464988 48816 465040 48822
rect 464988 48758 465040 48764
rect 465356 48816 465408 48822
rect 465356 48758 465408 48764
rect 466368 48816 466420 48822
rect 466368 48758 466420 48764
rect 466552 48816 466604 48822
rect 466552 48758 466604 48764
rect 467748 48816 467800 48822
rect 467748 48758 467800 48764
rect 460952 3318 462084 3346
rect 462332 3318 463280 3346
rect 463804 3318 464476 3346
rect 465000 3330 465028 48758
rect 465080 18624 465132 18630
rect 465080 18566 465132 18572
rect 465092 3346 465120 18566
rect 466380 5098 466408 48758
rect 466460 42084 466512 42090
rect 466460 42026 466512 42032
rect 466368 5092 466420 5098
rect 466368 5034 466420 5040
rect 466472 3346 466500 42026
rect 467760 18630 467788 48758
rect 467840 19984 467892 19990
rect 467840 19926 467892 19932
rect 467748 18624 467800 18630
rect 467748 18566 467800 18572
rect 467852 3398 467880 19926
rect 469140 15910 469168 52006
rect 469220 43512 469272 43518
rect 469220 43454 469272 43460
rect 469128 15904 469180 15910
rect 469128 15846 469180 15852
rect 467840 3392 467892 3398
rect 462056 480 462084 3318
rect 463252 480 463280 3318
rect 464448 480 464476 3318
rect 464988 3324 465040 3330
rect 465092 3318 465672 3346
rect 466472 3318 466868 3346
rect 469128 3392 469180 3398
rect 467840 3334 467892 3340
rect 467930 3360 467986 3369
rect 464988 3266 465040 3272
rect 465644 480 465672 3318
rect 466840 480 466868 3318
rect 469128 3334 469180 3340
rect 469232 3346 469260 43454
rect 470520 19990 470548 52006
rect 470508 19984 470560 19990
rect 470508 19926 470560 19932
rect 471520 3732 471572 3738
rect 471520 3674 471572 3680
rect 467930 3295 467986 3304
rect 467944 480 467972 3295
rect 469140 480 469168 3334
rect 469232 3318 470364 3346
rect 470336 480 470364 3318
rect 471532 480 471560 3674
rect 471900 3126 471928 52006
rect 472452 48822 472480 52020
rect 473648 48822 473676 52020
rect 474844 49162 474872 52020
rect 474832 49156 474884 49162
rect 474832 49098 474884 49104
rect 472440 48816 472492 48822
rect 472440 48758 472492 48764
rect 473268 48816 473320 48822
rect 473268 48758 473320 48764
rect 473636 48816 473688 48822
rect 473636 48758 473688 48764
rect 474648 48816 474700 48822
rect 474648 48758 474700 48764
rect 471980 21412 472032 21418
rect 471980 21354 472032 21360
rect 471888 3120 471940 3126
rect 471888 3062 471940 3068
rect 471992 610 472020 21354
rect 473280 5438 473308 48758
rect 474660 21418 474688 48758
rect 474648 21412 474700 21418
rect 474648 21354 474700 21360
rect 473360 14476 473412 14482
rect 473360 14418 473412 14424
rect 473268 5432 473320 5438
rect 473268 5374 473320 5380
rect 473372 610 473400 14418
rect 476040 4826 476068 52020
rect 477250 52006 477448 52034
rect 478446 52006 478828 52034
rect 479642 52006 480208 52034
rect 476120 44872 476172 44878
rect 476120 44814 476172 44820
rect 476028 4820 476080 4826
rect 476028 4762 476080 4768
rect 475108 4004 475160 4010
rect 475108 3946 475160 3952
rect 471980 604 472032 610
rect 471980 546 472032 552
rect 472716 604 472768 610
rect 472716 546 472768 552
rect 473360 604 473412 610
rect 473360 546 473412 552
rect 473912 604 473964 610
rect 473912 546 473964 552
rect 472728 480 472756 546
rect 473924 480 473952 546
rect 475120 480 475148 3946
rect 476132 626 476160 44814
rect 477420 39370 477448 52006
rect 477408 39364 477460 39370
rect 477408 39306 477460 39312
rect 477592 11756 477644 11762
rect 477592 11698 477644 11704
rect 477604 626 477632 11698
rect 478696 3528 478748 3534
rect 478696 3470 478748 3476
rect 476132 598 476344 626
rect 476316 480 476344 598
rect 477512 598 477632 626
rect 477512 480 477540 598
rect 478708 480 478736 3470
rect 478800 3398 478828 52006
rect 478880 22772 478932 22778
rect 478880 22714 478932 22720
rect 478788 3392 478840 3398
rect 478788 3334 478840 3340
rect 478892 610 478920 22714
rect 480180 4962 480208 52006
rect 480824 48822 480852 52020
rect 482020 49230 482048 52020
rect 482008 49224 482060 49230
rect 482008 49166 482060 49172
rect 483216 48822 483244 52020
rect 484412 48822 484440 52020
rect 485622 52006 485728 52034
rect 486818 52006 487108 52034
rect 488014 52006 488488 52034
rect 480812 48816 480864 48822
rect 480812 48758 480864 48764
rect 481548 48816 481600 48822
rect 481548 48758 481600 48764
rect 483204 48816 483256 48822
rect 483204 48758 483256 48764
rect 484308 48816 484360 48822
rect 484308 48758 484360 48764
rect 484400 48816 484452 48822
rect 484400 48758 484452 48764
rect 485596 48816 485648 48822
rect 485596 48758 485648 48764
rect 480260 38004 480312 38010
rect 480260 37946 480312 37952
rect 480168 4956 480220 4962
rect 480168 4898 480220 4904
rect 480272 3346 480300 37946
rect 481560 7682 481588 48758
rect 481548 7676 481600 7682
rect 481548 7618 481600 7624
rect 483480 7608 483532 7614
rect 483480 7550 483532 7556
rect 482284 3596 482336 3602
rect 482284 3538 482336 3544
rect 480272 3318 481128 3346
rect 478880 604 478932 610
rect 478880 546 478932 552
rect 479892 604 479944 610
rect 479892 546 479944 552
rect 479904 480 479932 546
rect 481100 480 481128 3318
rect 482296 480 482324 3538
rect 483492 480 483520 7550
rect 484320 5166 484348 48758
rect 485608 37942 485636 48758
rect 485596 37936 485648 37942
rect 485596 37878 485648 37884
rect 484400 24132 484452 24138
rect 484400 24074 484452 24080
rect 484308 5160 484360 5166
rect 484308 5102 484360 5108
rect 484412 3346 484440 24074
rect 485700 3641 485728 52006
rect 485780 40724 485832 40730
rect 485780 40666 485832 40672
rect 485686 3632 485742 3641
rect 485686 3567 485742 3576
rect 484412 3318 484624 3346
rect 484596 480 484624 3318
rect 485792 480 485820 40666
rect 486976 6180 487028 6186
rect 486976 6122 487028 6128
rect 486988 480 487016 6122
rect 487080 4894 487108 52006
rect 488460 25566 488488 52006
rect 489196 49094 489224 52020
rect 489184 49088 489236 49094
rect 489184 49030 489236 49036
rect 490392 48822 490420 52020
rect 491588 48822 491616 52020
rect 492784 48822 492812 52020
rect 493888 52006 493994 52034
rect 495190 52006 495388 52034
rect 496386 52006 496768 52034
rect 497490 52006 498148 52034
rect 490380 48816 490432 48822
rect 490380 48758 490432 48764
rect 491208 48816 491260 48822
rect 491208 48758 491260 48764
rect 491576 48816 491628 48822
rect 491576 48758 491628 48764
rect 492588 48816 492640 48822
rect 492588 48758 492640 48764
rect 492772 48816 492824 48822
rect 492772 48758 492824 48764
rect 487160 25560 487212 25566
rect 487160 25502 487212 25508
rect 488448 25560 488500 25566
rect 488448 25502 488500 25508
rect 487068 4888 487120 4894
rect 487068 4830 487120 4836
rect 487172 3346 487200 25502
rect 491220 8974 491248 48758
rect 491300 26988 491352 26994
rect 491300 26930 491352 26936
rect 490564 8968 490616 8974
rect 490564 8910 490616 8916
rect 491208 8968 491260 8974
rect 491208 8910 491260 8916
rect 489368 3460 489420 3466
rect 489368 3402 489420 3408
rect 487172 3318 488212 3346
rect 488184 480 488212 3318
rect 489380 480 489408 3402
rect 490576 480 490604 8910
rect 491312 3482 491340 26930
rect 492600 26926 492628 48758
rect 493888 44878 493916 52006
rect 493968 48816 494020 48822
rect 493968 48758 494020 48764
rect 493876 44872 493928 44878
rect 493876 44814 493928 44820
rect 492588 26920 492640 26926
rect 492588 26862 492640 26868
rect 493980 3534 494008 48758
rect 494060 47592 494112 47598
rect 494060 47534 494112 47540
rect 493968 3528 494020 3534
rect 491312 3454 491800 3482
rect 493968 3470 494020 3476
rect 494072 3482 494100 47534
rect 495360 28286 495388 52006
rect 494152 28280 494204 28286
rect 494152 28222 494204 28228
rect 495348 28280 495400 28286
rect 495348 28222 495400 28228
rect 494164 3602 494192 28222
rect 496740 4010 496768 52006
rect 498120 10334 498148 52006
rect 498672 48822 498700 52020
rect 499868 48822 499896 52020
rect 498660 48816 498712 48822
rect 498660 48758 498712 48764
rect 499488 48816 499540 48822
rect 499488 48758 499540 48764
rect 499856 48816 499908 48822
rect 499856 48758 499908 48764
rect 500868 48816 500920 48822
rect 500868 48758 500920 48764
rect 498200 29640 498252 29646
rect 498200 29582 498252 29588
rect 496820 10328 496872 10334
rect 496820 10270 496872 10276
rect 498108 10328 498160 10334
rect 498108 10270 498160 10276
rect 496728 4004 496780 4010
rect 496728 3946 496780 3952
rect 496544 3664 496596 3670
rect 496544 3606 496596 3612
rect 494152 3596 494204 3602
rect 494152 3538 494204 3544
rect 495348 3596 495400 3602
rect 495348 3538 495400 3544
rect 494072 3454 494192 3482
rect 491772 480 491800 3454
rect 492956 3052 493008 3058
rect 492956 2994 493008 3000
rect 492968 480 492996 2994
rect 494164 480 494192 3454
rect 495360 480 495388 3538
rect 496556 480 496584 3606
rect 496832 3482 496860 10270
rect 498212 3482 498240 29582
rect 499500 24138 499528 48758
rect 499488 24132 499540 24138
rect 499488 24074 499540 24080
rect 500132 4072 500184 4078
rect 500132 4014 500184 4020
rect 496832 3454 497780 3482
rect 498212 3454 498976 3482
rect 497752 480 497780 3454
rect 498948 480 498976 3454
rect 500144 480 500172 4014
rect 500880 3670 500908 48758
rect 501064 47598 501092 52020
rect 502168 52006 502274 52034
rect 503470 52006 503668 52034
rect 504666 52006 505048 52034
rect 505862 52006 506428 52034
rect 507058 52006 507808 52034
rect 501052 47592 501104 47598
rect 501052 47534 501104 47540
rect 500960 11824 501012 11830
rect 500960 11766 501012 11772
rect 500868 3664 500920 3670
rect 500868 3606 500920 3612
rect 500972 762 501000 11766
rect 502168 11762 502196 52006
rect 502432 33788 502484 33794
rect 502432 33730 502484 33736
rect 502156 11756 502208 11762
rect 502156 11698 502208 11704
rect 500972 734 501276 762
rect 501248 480 501276 734
rect 502444 480 502472 33730
rect 503640 3738 503668 52006
rect 505020 13122 505048 52006
rect 506400 31074 506428 52006
rect 505100 31068 505152 31074
rect 505100 31010 505152 31016
rect 506388 31068 506440 31074
rect 506388 31010 506440 31016
rect 503720 13116 503772 13122
rect 503720 13058 503772 13064
rect 505008 13116 505060 13122
rect 505008 13058 505060 13064
rect 503628 3732 503680 3738
rect 503628 3674 503680 3680
rect 503732 3346 503760 13058
rect 505112 3346 505140 31010
rect 507216 3868 507268 3874
rect 507216 3810 507268 3816
rect 503732 3318 504864 3346
rect 505112 3318 506060 3346
rect 503628 3256 503680 3262
rect 503628 3198 503680 3204
rect 503640 480 503668 3198
rect 504836 480 504864 3318
rect 506032 480 506060 3318
rect 507228 480 507256 3810
rect 507780 3806 507808 52006
rect 508240 48822 508268 52020
rect 509436 48822 509464 52020
rect 508228 48816 508280 48822
rect 508228 48758 508280 48764
rect 509148 48816 509200 48822
rect 509148 48758 509200 48764
rect 509424 48816 509476 48822
rect 509424 48758 509476 48764
rect 510528 48816 510580 48822
rect 510528 48758 510580 48764
rect 507860 14544 507912 14550
rect 507860 14486 507912 14492
rect 507768 3800 507820 3806
rect 507768 3742 507820 3748
rect 507872 3346 507900 14486
rect 509160 14482 509188 48758
rect 510540 32434 510568 48758
rect 510632 48550 510660 52020
rect 510620 48544 510672 48550
rect 510620 48486 510672 48492
rect 511828 43450 511856 52020
rect 513038 52006 513328 52034
rect 514234 52006 514708 52034
rect 511908 48544 511960 48550
rect 511908 48486 511960 48492
rect 511816 43444 511868 43450
rect 511816 43386 511868 43392
rect 509240 32428 509292 32434
rect 509240 32370 509292 32376
rect 510528 32428 510580 32434
rect 510528 32370 510580 32376
rect 509148 14476 509200 14482
rect 509148 14418 509200 14424
rect 509252 3346 509280 32370
rect 511920 3874 511948 48486
rect 512000 46232 512052 46238
rect 512000 46174 512052 46180
rect 511908 3868 511960 3874
rect 511908 3810 511960 3816
rect 510802 3496 510858 3505
rect 510802 3431 510858 3440
rect 507872 3318 508452 3346
rect 509252 3318 509648 3346
rect 508424 480 508452 3318
rect 509620 480 509648 3318
rect 510816 480 510844 3431
rect 512012 480 512040 46174
rect 512092 17264 512144 17270
rect 512092 17206 512144 17212
rect 512104 3346 512132 17206
rect 513300 3466 513328 52006
rect 514680 3942 514708 52006
rect 515416 46238 515444 52020
rect 516612 48822 516640 52020
rect 517808 48822 517836 52020
rect 519004 48822 519032 52020
rect 516600 48816 516652 48822
rect 516600 48758 516652 48764
rect 517428 48816 517480 48822
rect 517428 48758 517480 48764
rect 517796 48816 517848 48822
rect 517796 48758 517848 48764
rect 518808 48816 518860 48822
rect 518808 48758 518860 48764
rect 518992 48816 519044 48822
rect 518992 48758 519044 48764
rect 520096 48816 520148 48822
rect 520096 48758 520148 48764
rect 515404 46232 515456 46238
rect 515404 46174 515456 46180
rect 516140 29028 516192 29034
rect 516140 28970 516192 28976
rect 516152 19310 516180 28970
rect 515956 19304 516008 19310
rect 515956 19246 516008 19252
rect 516140 19304 516192 19310
rect 516140 19246 516192 19252
rect 515968 9761 515996 19246
rect 515954 9752 516010 9761
rect 515954 9687 516010 9696
rect 516138 9752 516194 9761
rect 516138 9687 516194 9696
rect 516152 9654 516180 9687
rect 516140 9648 516192 9654
rect 516140 9590 516192 9596
rect 515588 5024 515640 5030
rect 515588 4966 515640 4972
rect 514392 3936 514444 3942
rect 514392 3878 514444 3884
rect 514668 3936 514720 3942
rect 514668 3878 514720 3884
rect 513288 3460 513340 3466
rect 513288 3402 513340 3408
rect 512104 3318 513236 3346
rect 513208 480 513236 3318
rect 514404 480 514432 3878
rect 515600 480 515628 4966
rect 517440 3602 517468 48758
rect 518820 4078 518848 48758
rect 520108 42090 520136 48758
rect 520096 42084 520148 42090
rect 520096 42026 520148 42032
rect 519084 5296 519136 5302
rect 519084 5238 519136 5244
rect 518808 4072 518860 4078
rect 518808 4014 518860 4020
rect 517428 3596 517480 3602
rect 517428 3538 517480 3544
rect 517888 3188 517940 3194
rect 517888 3130 517940 3136
rect 516784 604 516836 610
rect 516784 546 516836 552
rect 516796 480 516824 546
rect 517900 480 517928 3130
rect 519096 480 519124 5238
rect 520200 3369 520228 52020
rect 521410 52006 521608 52034
rect 520372 36576 520424 36582
rect 520372 36518 520424 36524
rect 520384 19666 520412 36518
rect 520384 19638 520504 19666
rect 520476 19394 520504 19638
rect 520384 19366 520504 19394
rect 520384 9654 520412 19366
rect 520372 9648 520424 9654
rect 520372 9590 520424 9596
rect 521580 4146 521608 52006
rect 523696 41410 523724 85303
rect 523788 77246 523816 111959
rect 523880 111790 523908 138615
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 523868 111784 523920 111790
rect 523868 111726 523920 111732
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 523866 98696 523922 98705
rect 523866 98631 523922 98640
rect 523776 77240 523828 77246
rect 523776 77182 523828 77188
rect 523774 72040 523830 72049
rect 523774 71975 523830 71984
rect 523684 41404 523736 41410
rect 523684 41346 523736 41352
rect 523788 30326 523816 71975
rect 523880 64870 523908 98631
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 523868 64864 523920 64870
rect 523868 64806 523920 64812
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 523866 58712 523922 58721
rect 523866 58647 523922 58656
rect 523776 30320 523828 30326
rect 523776 30262 523828 30268
rect 523880 17950 523908 58647
rect 542360 49224 542412 49230
rect 542360 49166 542412 49172
rect 535460 49156 535512 49162
rect 535460 49098 535512 49104
rect 528560 49020 528612 49026
rect 528560 48962 528612 48968
rect 527272 18624 527324 18630
rect 527272 18566 527324 18572
rect 523868 17944 523920 17950
rect 523868 17886 523920 17892
rect 523868 5364 523920 5370
rect 523868 5306 523920 5312
rect 522672 5228 522724 5234
rect 522672 5170 522724 5176
rect 521476 4140 521528 4146
rect 521476 4082 521528 4088
rect 521568 4140 521620 4146
rect 521568 4082 521620 4088
rect 520186 3360 520242 3369
rect 520186 3295 520242 3304
rect 520280 604 520332 610
rect 520280 546 520332 552
rect 520292 480 520320 546
rect 521488 480 521516 4082
rect 522684 480 522712 5170
rect 523880 480 523908 5306
rect 526260 5092 526312 5098
rect 526260 5034 526312 5040
rect 525064 3324 525116 3330
rect 525064 3266 525116 3272
rect 525076 480 525104 3266
rect 526272 480 526300 5034
rect 527284 610 527312 18566
rect 528572 7426 528600 48962
rect 535472 46918 535500 49098
rect 535460 46912 535512 46918
rect 535460 46854 535512 46860
rect 536840 39364 536892 39370
rect 536840 39306 536892 39312
rect 535460 37324 535512 37330
rect 535460 37266 535512 37272
rect 535472 27606 535500 37266
rect 535460 27600 535512 27606
rect 535460 27542 535512 27548
rect 534080 21412 534132 21418
rect 534080 21354 534132 21360
rect 529940 19984 529992 19990
rect 529940 19926 529992 19932
rect 528652 15904 528704 15910
rect 528652 15846 528704 15852
rect 528664 7614 528692 15846
rect 529952 12442 529980 19926
rect 534092 12442 534120 21354
rect 529940 12436 529992 12442
rect 529940 12378 529992 12384
rect 531044 12436 531096 12442
rect 531044 12378 531096 12384
rect 534080 12436 534132 12442
rect 534080 12378 534132 12384
rect 534540 12436 534592 12442
rect 534540 12378 534592 12384
rect 528652 7608 528704 7614
rect 528652 7550 528704 7556
rect 529848 7608 529900 7614
rect 529848 7550 529900 7556
rect 528572 7398 528692 7426
rect 527272 604 527324 610
rect 527272 546 527324 552
rect 527456 604 527508 610
rect 527456 546 527508 552
rect 527468 480 527496 546
rect 528664 480 528692 7398
rect 529860 480 529888 7550
rect 531056 480 531084 12378
rect 533436 5432 533488 5438
rect 533436 5374 533488 5380
rect 532240 3120 532292 3126
rect 532240 3062 532292 3068
rect 532252 480 532280 3062
rect 533448 480 533476 5374
rect 534552 480 534580 12378
rect 535736 9716 535788 9722
rect 535736 9658 535788 9664
rect 535748 480 535776 9658
rect 536852 7614 536880 39306
rect 542372 12442 542400 49166
rect 549260 49088 549312 49094
rect 549260 49030 549312 49036
rect 545120 37936 545172 37942
rect 545120 37878 545172 37884
rect 542360 12436 542412 12442
rect 542360 12378 542412 12384
rect 542912 12436 542964 12442
rect 542912 12378 542964 12384
rect 541716 7676 541768 7682
rect 541716 7618 541768 7624
rect 536840 7608 536892 7614
rect 536840 7550 536892 7556
rect 538128 7608 538180 7614
rect 538128 7550 538180 7556
rect 536932 4820 536984 4826
rect 536932 4762 536984 4768
rect 536944 480 536972 4762
rect 538140 480 538168 7550
rect 540520 4956 540572 4962
rect 540520 4898 540572 4904
rect 539324 3392 539376 3398
rect 539324 3334 539376 3340
rect 539336 480 539364 3334
rect 540532 480 540560 4898
rect 541728 480 541756 7618
rect 542924 480 542952 12378
rect 544108 5160 544160 5166
rect 544108 5102 544160 5108
rect 544120 480 544148 5102
rect 545132 3482 545160 37878
rect 547880 25560 547932 25566
rect 547880 25502 547932 25508
rect 547696 4888 547748 4894
rect 547696 4830 547748 4836
rect 546498 3632 546554 3641
rect 546498 3567 546554 3576
rect 545132 3454 545344 3482
rect 545316 480 545344 3454
rect 546512 480 546540 3567
rect 547708 480 547736 4830
rect 547892 3482 547920 25502
rect 549272 3482 549300 49030
rect 561680 47592 561732 47598
rect 561680 47534 561732 47540
rect 554780 44872 554832 44878
rect 554780 44814 554832 44820
rect 552020 26920 552072 26926
rect 552020 26862 552072 26868
rect 551192 8968 551244 8974
rect 551192 8910 551244 8916
rect 547892 3454 548932 3482
rect 549272 3454 550128 3482
rect 548904 480 548932 3454
rect 550100 480 550128 3454
rect 551204 480 551232 8910
rect 552032 3482 552060 26862
rect 553584 3528 553636 3534
rect 552032 3454 552428 3482
rect 553584 3470 553636 3476
rect 552400 480 552428 3454
rect 553596 480 553624 3470
rect 554792 480 554820 44814
rect 554872 28280 554924 28286
rect 554872 28222 554924 28228
rect 554884 3482 554912 28222
rect 558920 24132 558972 24138
rect 558920 24074 558972 24080
rect 557540 10328 557592 10334
rect 557540 10270 557592 10276
rect 557172 4004 557224 4010
rect 557172 3946 557224 3952
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3946
rect 557552 3482 557580 10270
rect 558932 3482 558960 24074
rect 560760 3664 560812 3670
rect 560760 3606 560812 3612
rect 557552 3454 558408 3482
rect 558932 3454 559604 3482
rect 558380 480 558408 3454
rect 559576 480 559604 3454
rect 560772 480 560800 3606
rect 561692 3482 561720 47534
rect 575480 46232 575532 46238
rect 575480 46174 575532 46180
rect 571432 43444 571484 43450
rect 571432 43386 571484 43392
rect 569960 32428 570012 32434
rect 569960 32370 570012 32376
rect 565820 31068 565872 31074
rect 565820 31010 565872 31016
rect 564440 13116 564492 13122
rect 564440 13058 564492 13064
rect 563152 11756 563204 11762
rect 563152 11698 563204 11704
rect 561692 3454 561996 3482
rect 561968 480 561996 3454
rect 563164 480 563192 11698
rect 564348 3732 564400 3738
rect 564348 3674 564400 3680
rect 564360 480 564388 3674
rect 564452 3482 564480 13058
rect 565832 3482 565860 31010
rect 568580 14476 568632 14482
rect 568580 14418 568632 14424
rect 567844 3800 567896 3806
rect 567844 3742 567896 3748
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3742
rect 568592 3482 568620 14418
rect 569972 3482 570000 32370
rect 571340 3868 571392 3874
rect 571340 3810 571392 3816
rect 568592 3454 569080 3482
rect 569972 3454 570276 3482
rect 569052 480 569080 3454
rect 570248 480 570276 3454
rect 571352 3346 571380 3810
rect 571444 3534 571472 43386
rect 575020 3936 575072 3942
rect 575020 3878 575072 3884
rect 571432 3528 571484 3534
rect 571432 3470 571484 3476
rect 572628 3528 572680 3534
rect 572628 3470 572680 3476
rect 571352 3318 571472 3346
rect 571444 480 571472 3318
rect 572640 480 572668 3470
rect 573824 3460 573876 3466
rect 573824 3402 573876 3408
rect 573836 480 573864 3402
rect 575032 480 575060 3878
rect 575492 3482 575520 46174
rect 579620 42084 579672 42090
rect 579620 42026 579672 42032
rect 578608 4072 578660 4078
rect 578608 4014 578660 4020
rect 577412 3596 577464 3602
rect 577412 3538 577464 3544
rect 575492 3454 576256 3482
rect 576228 480 576256 3454
rect 577424 480 577452 3538
rect 578620 480 578648 4014
rect 579632 610 579660 42026
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 580080 17944 580132 17950
rect 580080 17886 580132 17892
rect 580092 17649 580120 17886
rect 580078 17640 580134 17649
rect 580078 17575 580134 17584
rect 582196 4140 582248 4146
rect 582196 4082 582248 4088
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 579620 604 579672 610
rect 579620 546 579672 552
rect 579804 604 579856 610
rect 579804 546 579856 552
rect 579816 480 579844 546
rect 581012 480 581040 3295
rect 582208 480 582236 4082
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667936 3478 667992
rect 3606 653520 3662 653576
rect 3514 624824 3570 624880
rect 3422 610408 3478 610464
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 580170 697992 580226 698048
rect 59358 644680 59414 644736
rect 580170 686296 580226 686352
rect 580262 674600 580318 674656
rect 523774 645224 523830 645280
rect 580170 639376 580226 639432
rect 523682 631896 523738 631952
rect 59358 630400 59414 630456
rect 59358 616120 59414 616176
rect 523130 605240 523186 605296
rect 59358 601840 59414 601896
rect 3514 595992 3570 596048
rect 59358 587560 59414 587616
rect 59358 573280 59414 573336
rect 3422 567296 3478 567352
rect 523130 565256 523186 565312
rect 59358 559000 59414 559056
rect 3422 553016 3478 553072
rect 580446 651072 580502 651128
rect 580354 627680 580410 627736
rect 524326 618568 524382 618624
rect 579802 592456 579858 592512
rect 523774 591912 523830 591968
rect 580262 580760 580318 580816
rect 524326 578584 524382 578640
rect 580170 557232 580226 557288
rect 523682 551928 523738 551984
rect 59358 544720 59414 544776
rect 3422 538600 3478 538656
rect 523682 538600 523738 538656
rect 59358 530440 59414 530496
rect 59358 516180 59414 516216
rect 59358 516160 59360 516180
rect 59360 516160 59412 516180
rect 59412 516160 59414 516180
rect 580170 545536 580226 545592
rect 580446 604152 580502 604208
rect 580262 533840 580318 533896
rect 523774 525272 523830 525328
rect 523682 511944 523738 512000
rect 580170 510312 580226 510368
rect 3422 509904 3478 509960
rect 59358 501880 59414 501936
rect 523682 498616 523738 498672
rect 3330 495488 3386 495544
rect 59358 487600 59414 487656
rect 3422 481072 3478 481128
rect 59358 473356 59360 473376
rect 59360 473356 59412 473376
rect 59412 473356 59414 473376
rect 59358 473320 59414 473356
rect 580170 498616 580226 498672
rect 580262 486784 580318 486840
rect 523774 485288 523830 485344
rect 523682 471960 523738 472016
rect 580170 463392 580226 463448
rect 59358 459040 59414 459096
rect 3422 452376 3478 452432
rect 524326 458632 524382 458688
rect 580170 451696 580226 451752
rect 523682 445304 523738 445360
rect 59358 444760 59414 444816
rect 3514 437960 3570 438016
rect 59358 430480 59414 430536
rect 3422 423680 3478 423736
rect 3422 380568 3478 380624
rect 580170 439864 580226 439920
rect 523774 431976 523830 432032
rect 523682 418648 523738 418704
rect 580170 416472 580226 416528
rect 59358 416200 59414 416256
rect 523682 405320 523738 405376
rect 580170 404776 580226 404832
rect 59358 401920 59414 401976
rect 3606 394984 3662 395040
rect 580170 392944 580226 393000
rect 523774 391992 523830 392048
rect 60094 387640 60150 387696
rect 59358 373360 59414 373416
rect 3514 366152 3570 366208
rect 3330 337456 3386 337512
rect 3054 294344 3110 294400
rect 59358 359080 59414 359136
rect 60002 344664 60058 344720
rect 59358 330384 59414 330440
rect 3606 323040 3662 323096
rect 59358 316104 59414 316160
rect 3514 308760 3570 308816
rect 3422 280064 3478 280120
rect 3146 251232 3202 251288
rect 523682 378664 523738 378720
rect 580170 369552 580226 369608
rect 524234 365336 524290 365392
rect 580170 357856 580226 357912
rect 523682 351872 523738 351928
rect 580170 346024 580226 346080
rect 523774 338544 523830 338600
rect 524326 325216 524382 325272
rect 580170 322632 580226 322688
rect 524326 311888 524382 311944
rect 580170 310800 580226 310856
rect 60094 301824 60150 301880
rect 59358 287544 59414 287600
rect 59358 273284 59414 273320
rect 59358 273264 59360 273284
rect 59360 273264 59412 273284
rect 59412 273264 59414 273284
rect 3606 265648 3662 265704
rect 60002 258984 60058 259040
rect 59358 244704 59414 244760
rect 3514 236952 3570 237008
rect 3422 222536 3478 222592
rect 3146 208120 3202 208176
rect 3422 165008 3478 165064
rect 2962 122032 3018 122088
rect 59358 230424 59414 230480
rect 3606 193840 3662 193896
rect 3514 150728 3570 150784
rect 580170 299104 580226 299160
rect 524326 298560 524382 298616
rect 523682 285232 523738 285288
rect 580170 275712 580226 275768
rect 523682 271904 523738 271960
rect 580170 263880 580226 263936
rect 523682 258576 523738 258632
rect 579802 252184 579858 252240
rect 523682 245248 523738 245304
rect 523774 231920 523830 231976
rect 580170 228792 580226 228848
rect 523866 218592 523922 218648
rect 60094 216144 60150 216200
rect 59358 201864 59414 201920
rect 59358 187584 59414 187640
rect 3698 179424 3754 179480
rect 60002 173304 60058 173360
rect 59358 159024 59414 159080
rect 59358 144744 59414 144800
rect 3606 136312 3662 136368
rect 3422 107616 3478 107672
rect 3054 78920 3110 78976
rect 3330 35844 3332 35864
rect 3332 35844 3384 35864
rect 3384 35844 3386 35864
rect 3330 35808 3386 35844
rect 3514 64504 3570 64560
rect 3422 21392 3478 21448
rect 580170 216960 580226 217016
rect 523682 205264 523738 205320
rect 579802 205264 579858 205320
rect 523774 191936 523830 191992
rect 580170 181872 580226 181928
rect 523866 178608 523922 178664
rect 523682 165280 523738 165336
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 523774 151952 523830 152008
rect 60094 130464 60150 130520
rect 59358 116184 59414 116240
rect 59358 101904 59414 101960
rect 3698 93200 3754 93256
rect 60002 87624 60058 87680
rect 59358 73344 59414 73400
rect 59358 59064 59414 59120
rect 3606 50088 3662 50144
rect 523682 125296 523738 125352
rect 523866 138624 523922 138680
rect 523774 111968 523830 112024
rect 523682 85312 523738 85368
rect 3514 7112 3570 7168
rect 85486 3440 85542 3496
rect 92386 3304 92442 3360
rect 146850 3440 146906 3496
rect 153934 3304 153990 3360
rect 339406 3304 339462 3360
rect 364246 3440 364302 3496
rect 400218 3304 400274 3360
rect 407026 3304 407082 3360
rect 425150 3440 425206 3496
rect 449806 3440 449862 3496
rect 467930 3304 467986 3360
rect 485686 3576 485742 3632
rect 510802 3440 510858 3496
rect 515954 9696 516010 9752
rect 516138 9696 516194 9752
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 523866 98640 523922 98696
rect 523774 71984 523830 72040
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 523866 58656 523922 58712
rect 520186 3304 520242 3360
rect 546498 3576 546554 3632
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 580078 17584 580134 17640
rect 580998 3304 581054 3360
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3601 653578 3667 653581
rect -960 653576 3667 653578
rect -960 653520 3606 653576
rect 3662 653520 3667 653576
rect -960 653518 3667 653520
rect -960 653428 480 653518
rect 3601 653515 3667 653518
rect 580441 651130 580507 651133
rect 583520 651130 584960 651220
rect 580441 651128 584960 651130
rect 580441 651072 580446 651128
rect 580502 651072 584960 651128
rect 580441 651070 584960 651072
rect 580441 651067 580507 651070
rect 583520 650980 584960 651070
rect 523769 645282 523835 645285
rect 521916 645280 523835 645282
rect 521916 645224 523774 645280
rect 523830 645224 523835 645280
rect 521916 645222 523835 645224
rect 523769 645219 523835 645222
rect 59353 644738 59419 644741
rect 59353 644736 62100 644738
rect 59353 644680 59358 644736
rect 59414 644680 62100 644736
rect 59353 644678 62100 644680
rect 59353 644675 59419 644678
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 523677 631954 523743 631957
rect 521916 631952 523743 631954
rect 521916 631896 523682 631952
rect 523738 631896 523743 631952
rect 521916 631894 523743 631896
rect 523677 631891 523743 631894
rect 59353 630458 59419 630461
rect 59353 630456 62100 630458
rect 59353 630400 59358 630456
rect 59414 630400 62100 630456
rect 59353 630398 62100 630400
rect 59353 630395 59419 630398
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3509 624882 3575 624885
rect -960 624880 3575 624882
rect -960 624824 3514 624880
rect 3570 624824 3575 624880
rect -960 624822 3575 624824
rect -960 624732 480 624822
rect 3509 624819 3575 624822
rect 524321 618626 524387 618629
rect 521916 618624 524387 618626
rect 521916 618568 524326 618624
rect 524382 618568 524387 618624
rect 521916 618566 524387 618568
rect 524321 618563 524387 618566
rect 59353 616178 59419 616181
rect 59353 616176 62100 616178
rect 59353 616120 59358 616176
rect 59414 616120 62100 616176
rect 59353 616118 62100 616120
rect 59353 616115 59419 616118
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 523125 605298 523191 605301
rect 521916 605296 523191 605298
rect 521916 605240 523130 605296
rect 523186 605240 523191 605296
rect 521916 605238 523191 605240
rect 523125 605235 523191 605238
rect 580441 604210 580507 604213
rect 583520 604210 584960 604300
rect 580441 604208 584960 604210
rect 580441 604152 580446 604208
rect 580502 604152 584960 604208
rect 580441 604150 584960 604152
rect 580441 604147 580507 604150
rect 583520 604060 584960 604150
rect 59353 601898 59419 601901
rect 59353 601896 62100 601898
rect 59353 601840 59358 601896
rect 59414 601840 62100 601896
rect 59353 601838 62100 601840
rect 59353 601835 59419 601838
rect -960 596050 480 596140
rect 3509 596050 3575 596053
rect -960 596048 3575 596050
rect -960 595992 3514 596048
rect 3570 595992 3575 596048
rect -960 595990 3575 595992
rect -960 595900 480 595990
rect 3509 595987 3575 595990
rect 579797 592514 579863 592517
rect 583520 592514 584960 592604
rect 579797 592512 584960 592514
rect 579797 592456 579802 592512
rect 579858 592456 584960 592512
rect 579797 592454 584960 592456
rect 579797 592451 579863 592454
rect 583520 592364 584960 592454
rect 523769 591970 523835 591973
rect 521916 591968 523835 591970
rect 521916 591912 523774 591968
rect 523830 591912 523835 591968
rect 521916 591910 523835 591912
rect 523769 591907 523835 591910
rect 59353 587618 59419 587621
rect 59353 587616 62100 587618
rect 59353 587560 59358 587616
rect 59414 587560 62100 587616
rect 59353 587558 62100 587560
rect 59353 587555 59419 587558
rect -960 581620 480 581860
rect 580257 580818 580323 580821
rect 583520 580818 584960 580908
rect 580257 580816 584960 580818
rect 580257 580760 580262 580816
rect 580318 580760 584960 580816
rect 580257 580758 584960 580760
rect 580257 580755 580323 580758
rect 583520 580668 584960 580758
rect 524321 578642 524387 578645
rect 521916 578640 524387 578642
rect 521916 578584 524326 578640
rect 524382 578584 524387 578640
rect 521916 578582 524387 578584
rect 524321 578579 524387 578582
rect 59353 573338 59419 573341
rect 59353 573336 62100 573338
rect 59353 573280 59358 573336
rect 59414 573280 62100 573336
rect 59353 573278 62100 573280
rect 59353 573275 59419 573278
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 523125 565314 523191 565317
rect 521916 565312 523191 565314
rect 521916 565256 523130 565312
rect 523186 565256 523191 565312
rect 521916 565254 523191 565256
rect 523125 565251 523191 565254
rect 59353 559058 59419 559061
rect 59353 559056 62100 559058
rect 59353 559000 59358 559056
rect 59414 559000 62100 559056
rect 59353 558998 62100 559000
rect 59353 558995 59419 558998
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3417 553074 3483 553077
rect -960 553072 3483 553074
rect -960 553016 3422 553072
rect 3478 553016 3483 553072
rect -960 553014 3483 553016
rect -960 552924 480 553014
rect 3417 553011 3483 553014
rect 523677 551986 523743 551989
rect 521916 551984 523743 551986
rect 521916 551928 523682 551984
rect 523738 551928 523743 551984
rect 521916 551926 523743 551928
rect 523677 551923 523743 551926
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 59353 544778 59419 544781
rect 59353 544776 62100 544778
rect 59353 544720 59358 544776
rect 59414 544720 62100 544776
rect 59353 544718 62100 544720
rect 59353 544715 59419 544718
rect -960 538658 480 538748
rect 3417 538658 3483 538661
rect 523677 538658 523743 538661
rect -960 538656 3483 538658
rect -960 538600 3422 538656
rect 3478 538600 3483 538656
rect -960 538598 3483 538600
rect 521916 538656 523743 538658
rect 521916 538600 523682 538656
rect 523738 538600 523743 538656
rect 521916 538598 523743 538600
rect -960 538508 480 538598
rect 3417 538595 3483 538598
rect 523677 538595 523743 538598
rect 580257 533898 580323 533901
rect 583520 533898 584960 533988
rect 580257 533896 584960 533898
rect 580257 533840 580262 533896
rect 580318 533840 584960 533896
rect 580257 533838 584960 533840
rect 580257 533835 580323 533838
rect 583520 533748 584960 533838
rect 59353 530498 59419 530501
rect 59353 530496 62100 530498
rect 59353 530440 59358 530496
rect 59414 530440 62100 530496
rect 59353 530438 62100 530440
rect 59353 530435 59419 530438
rect 523769 525330 523835 525333
rect 521916 525328 523835 525330
rect 521916 525272 523774 525328
rect 523830 525272 523835 525328
rect 521916 525270 523835 525272
rect 523769 525267 523835 525270
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 59353 516218 59419 516221
rect 59353 516216 62100 516218
rect 59353 516160 59358 516216
rect 59414 516160 62100 516216
rect 59353 516158 62100 516160
rect 59353 516155 59419 516158
rect 523677 512002 523743 512005
rect 521916 512000 523743 512002
rect 521916 511944 523682 512000
rect 523738 511944 523743 512000
rect 521916 511942 523743 511944
rect 523677 511939 523743 511942
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3417 509962 3483 509965
rect -960 509960 3483 509962
rect -960 509904 3422 509960
rect 3478 509904 3483 509960
rect -960 509902 3483 509904
rect -960 509812 480 509902
rect 3417 509899 3483 509902
rect 59353 501938 59419 501941
rect 59353 501936 62100 501938
rect 59353 501880 59358 501936
rect 59414 501880 62100 501936
rect 59353 501878 62100 501880
rect 59353 501875 59419 501878
rect 523677 498674 523743 498677
rect 521916 498672 523743 498674
rect 521916 498616 523682 498672
rect 523738 498616 523743 498672
rect 521916 498614 523743 498616
rect 523677 498611 523743 498614
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 59353 487658 59419 487661
rect 59353 487656 62100 487658
rect 59353 487600 59358 487656
rect 59414 487600 62100 487656
rect 59353 487598 62100 487600
rect 59353 487595 59419 487598
rect 580257 486842 580323 486845
rect 583520 486842 584960 486932
rect 580257 486840 584960 486842
rect 580257 486784 580262 486840
rect 580318 486784 584960 486840
rect 580257 486782 584960 486784
rect 580257 486779 580323 486782
rect 583520 486692 584960 486782
rect 523769 485346 523835 485349
rect 521916 485344 523835 485346
rect 521916 485288 523774 485344
rect 523830 485288 523835 485344
rect 521916 485286 523835 485288
rect 523769 485283 523835 485286
rect -960 481130 480 481220
rect 3417 481130 3483 481133
rect -960 481128 3483 481130
rect -960 481072 3422 481128
rect 3478 481072 3483 481128
rect -960 481070 3483 481072
rect -960 480980 480 481070
rect 3417 481067 3483 481070
rect 583520 474996 584960 475236
rect 59353 473378 59419 473381
rect 59353 473376 62100 473378
rect 59353 473320 59358 473376
rect 59414 473320 62100 473376
rect 59353 473318 62100 473320
rect 59353 473315 59419 473318
rect 523677 472018 523743 472021
rect 521916 472016 523743 472018
rect 521916 471960 523682 472016
rect 523738 471960 523743 472016
rect 521916 471958 523743 471960
rect 523677 471955 523743 471958
rect -960 466700 480 466940
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 59353 459098 59419 459101
rect 59353 459096 62100 459098
rect 59353 459040 59358 459096
rect 59414 459040 62100 459096
rect 59353 459038 62100 459040
rect 59353 459035 59419 459038
rect 524321 458690 524387 458693
rect 521916 458688 524387 458690
rect 521916 458632 524326 458688
rect 524382 458632 524387 458688
rect 521916 458630 524387 458632
rect 524321 458627 524387 458630
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 523677 445362 523743 445365
rect 521916 445360 523743 445362
rect 521916 445304 523682 445360
rect 523738 445304 523743 445360
rect 521916 445302 523743 445304
rect 523677 445299 523743 445302
rect 59353 444818 59419 444821
rect 59353 444816 62100 444818
rect 59353 444760 59358 444816
rect 59414 444760 62100 444816
rect 59353 444758 62100 444760
rect 59353 444755 59419 444758
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3509 438018 3575 438021
rect -960 438016 3575 438018
rect -960 437960 3514 438016
rect 3570 437960 3575 438016
rect -960 437958 3575 437960
rect -960 437868 480 437958
rect 3509 437955 3575 437958
rect 523769 432034 523835 432037
rect 521916 432032 523835 432034
rect 521916 431976 523774 432032
rect 523830 431976 523835 432032
rect 521916 431974 523835 431976
rect 523769 431971 523835 431974
rect 59353 430538 59419 430541
rect 59353 430536 62100 430538
rect 59353 430480 59358 430536
rect 59414 430480 62100 430536
rect 59353 430478 62100 430480
rect 59353 430475 59419 430478
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3417 423738 3483 423741
rect -960 423736 3483 423738
rect -960 423680 3422 423736
rect 3478 423680 3483 423736
rect -960 423678 3483 423680
rect -960 423588 480 423678
rect 3417 423675 3483 423678
rect 523677 418706 523743 418709
rect 521916 418704 523743 418706
rect 521916 418648 523682 418704
rect 523738 418648 523743 418704
rect 521916 418646 523743 418648
rect 523677 418643 523743 418646
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 59353 416258 59419 416261
rect 59353 416256 62100 416258
rect 59353 416200 59358 416256
rect 59414 416200 62100 416256
rect 59353 416198 62100 416200
rect 59353 416195 59419 416198
rect -960 409172 480 409412
rect 523677 405378 523743 405381
rect 521916 405376 523743 405378
rect 521916 405320 523682 405376
rect 523738 405320 523743 405376
rect 521916 405318 523743 405320
rect 523677 405315 523743 405318
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 59353 401978 59419 401981
rect 59353 401976 62100 401978
rect 59353 401920 59358 401976
rect 59414 401920 62100 401976
rect 59353 401918 62100 401920
rect 59353 401915 59419 401918
rect -960 395042 480 395132
rect 3601 395042 3667 395045
rect -960 395040 3667 395042
rect -960 394984 3606 395040
rect 3662 394984 3667 395040
rect -960 394982 3667 394984
rect -960 394892 480 394982
rect 3601 394979 3667 394982
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 523769 392050 523835 392053
rect 521916 392048 523835 392050
rect 521916 391992 523774 392048
rect 523830 391992 523835 392048
rect 521916 391990 523835 391992
rect 523769 391987 523835 391990
rect 60089 387698 60155 387701
rect 60089 387696 62100 387698
rect 60089 387640 60094 387696
rect 60150 387640 62100 387696
rect 60089 387638 62100 387640
rect 60089 387635 60155 387638
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3417 380626 3483 380629
rect -960 380624 3483 380626
rect -960 380568 3422 380624
rect 3478 380568 3483 380624
rect -960 380566 3483 380568
rect -960 380476 480 380566
rect 3417 380563 3483 380566
rect 523677 378722 523743 378725
rect 521916 378720 523743 378722
rect 521916 378664 523682 378720
rect 523738 378664 523743 378720
rect 521916 378662 523743 378664
rect 523677 378659 523743 378662
rect 59353 373418 59419 373421
rect 59353 373416 62100 373418
rect 59353 373360 59358 373416
rect 59414 373360 62100 373416
rect 59353 373358 62100 373360
rect 59353 373355 59419 373358
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3509 366210 3575 366213
rect -960 366208 3575 366210
rect -960 366152 3514 366208
rect 3570 366152 3575 366208
rect -960 366150 3575 366152
rect -960 366060 480 366150
rect 3509 366147 3575 366150
rect 524229 365394 524295 365397
rect 521916 365392 524295 365394
rect 521916 365336 524234 365392
rect 524290 365336 524295 365392
rect 521916 365334 524295 365336
rect 524229 365331 524295 365334
rect 59353 359138 59419 359141
rect 59353 359136 62100 359138
rect 59353 359080 59358 359136
rect 59414 359080 62100 359136
rect 59353 359078 62100 359080
rect 59353 359075 59419 359078
rect 580165 357914 580231 357917
rect 583520 357914 584960 358004
rect 580165 357912 584960 357914
rect 580165 357856 580170 357912
rect 580226 357856 584960 357912
rect 580165 357854 584960 357856
rect 580165 357851 580231 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 523677 351930 523743 351933
rect 521916 351928 523743 351930
rect 521916 351872 523682 351928
rect 523738 351872 523743 351928
rect 521916 351870 523743 351872
rect 523677 351867 523743 351870
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 59997 344722 60063 344725
rect 59997 344720 62100 344722
rect 59997 344664 60002 344720
rect 60058 344664 62100 344720
rect 59997 344662 62100 344664
rect 59997 344659 60063 344662
rect 523769 338602 523835 338605
rect 521916 338600 523835 338602
rect 521916 338544 523774 338600
rect 523830 338544 523835 338600
rect 521916 338542 523835 338544
rect 523769 338539 523835 338542
rect -960 337514 480 337604
rect 3325 337514 3391 337517
rect -960 337512 3391 337514
rect -960 337456 3330 337512
rect 3386 337456 3391 337512
rect -960 337454 3391 337456
rect -960 337364 480 337454
rect 3325 337451 3391 337454
rect 583520 334236 584960 334476
rect 59353 330442 59419 330445
rect 59353 330440 62100 330442
rect 59353 330384 59358 330440
rect 59414 330384 62100 330440
rect 59353 330382 62100 330384
rect 59353 330379 59419 330382
rect 524321 325274 524387 325277
rect 521916 325272 524387 325274
rect 521916 325216 524326 325272
rect 524382 325216 524387 325272
rect 521916 325214 524387 325216
rect 524321 325211 524387 325214
rect -960 323098 480 323188
rect 3601 323098 3667 323101
rect -960 323096 3667 323098
rect -960 323040 3606 323096
rect 3662 323040 3667 323096
rect -960 323038 3667 323040
rect -960 322948 480 323038
rect 3601 323035 3667 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 59353 316162 59419 316165
rect 59353 316160 62100 316162
rect 59353 316104 59358 316160
rect 59414 316104 62100 316160
rect 59353 316102 62100 316104
rect 59353 316099 59419 316102
rect 524321 311946 524387 311949
rect 521916 311944 524387 311946
rect 521916 311888 524326 311944
rect 524382 311888 524387 311944
rect 521916 311886 524387 311888
rect 524321 311883 524387 311886
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3509 308818 3575 308821
rect -960 308816 3575 308818
rect -960 308760 3514 308816
rect 3570 308760 3575 308816
rect -960 308758 3575 308760
rect -960 308668 480 308758
rect 3509 308755 3575 308758
rect 60089 301882 60155 301885
rect 60089 301880 62100 301882
rect 60089 301824 60094 301880
rect 60150 301824 62100 301880
rect 60089 301822 62100 301824
rect 60089 301819 60155 301822
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect 524321 298618 524387 298621
rect 521916 298616 524387 298618
rect 521916 298560 524326 298616
rect 524382 298560 524387 298616
rect 521916 298558 524387 298560
rect 524321 298555 524387 298558
rect -960 294402 480 294492
rect 3049 294402 3115 294405
rect -960 294400 3115 294402
rect -960 294344 3054 294400
rect 3110 294344 3115 294400
rect -960 294342 3115 294344
rect -960 294252 480 294342
rect 3049 294339 3115 294342
rect 59353 287602 59419 287605
rect 59353 287600 62100 287602
rect 59353 287544 59358 287600
rect 59414 287544 62100 287600
rect 59353 287542 62100 287544
rect 59353 287539 59419 287542
rect 583520 287316 584960 287556
rect 523677 285290 523743 285293
rect 521916 285288 523743 285290
rect 521916 285232 523682 285288
rect 523738 285232 523743 285288
rect 521916 285230 523743 285232
rect 523677 285227 523743 285230
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 59353 273322 59419 273325
rect 59353 273320 62100 273322
rect 59353 273264 59358 273320
rect 59414 273264 62100 273320
rect 59353 273262 62100 273264
rect 59353 273259 59419 273262
rect 523677 271962 523743 271965
rect 521916 271960 523743 271962
rect 521916 271904 523682 271960
rect 523738 271904 523743 271960
rect 521916 271902 523743 271904
rect 523677 271899 523743 271902
rect -960 265706 480 265796
rect 3601 265706 3667 265709
rect -960 265704 3667 265706
rect -960 265648 3606 265704
rect 3662 265648 3667 265704
rect -960 265646 3667 265648
rect -960 265556 480 265646
rect 3601 265643 3667 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 59997 259042 60063 259045
rect 59997 259040 62100 259042
rect 59997 258984 60002 259040
rect 60058 258984 62100 259040
rect 59997 258982 62100 258984
rect 59997 258979 60063 258982
rect 523677 258634 523743 258637
rect 521916 258632 523743 258634
rect 521916 258576 523682 258632
rect 523738 258576 523743 258632
rect 521916 258574 523743 258576
rect 523677 258571 523743 258574
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 523677 245306 523743 245309
rect 521916 245304 523743 245306
rect 521916 245248 523682 245304
rect 523738 245248 523743 245304
rect 521916 245246 523743 245248
rect 523677 245243 523743 245246
rect 59353 244762 59419 244765
rect 59353 244760 62100 244762
rect 59353 244704 59358 244760
rect 59414 244704 62100 244760
rect 59353 244702 62100 244704
rect 59353 244699 59419 244702
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3509 237010 3575 237013
rect -960 237008 3575 237010
rect -960 236952 3514 237008
rect 3570 236952 3575 237008
rect -960 236950 3575 236952
rect -960 236860 480 236950
rect 3509 236947 3575 236950
rect 523769 231978 523835 231981
rect 521916 231976 523835 231978
rect 521916 231920 523774 231976
rect 523830 231920 523835 231976
rect 521916 231918 523835 231920
rect 523769 231915 523835 231918
rect 59353 230482 59419 230485
rect 59353 230480 62100 230482
rect 59353 230424 59358 230480
rect 59414 230424 62100 230480
rect 59353 230422 62100 230424
rect 59353 230419 59419 230422
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3417 222594 3483 222597
rect -960 222592 3483 222594
rect -960 222536 3422 222592
rect 3478 222536 3483 222592
rect -960 222534 3483 222536
rect -960 222444 480 222534
rect 3417 222531 3483 222534
rect 523861 218650 523927 218653
rect 521916 218648 523927 218650
rect 521916 218592 523866 218648
rect 523922 218592 523927 218648
rect 521916 218590 523927 218592
rect 523861 218587 523927 218590
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 60089 216202 60155 216205
rect 60089 216200 62100 216202
rect 60089 216144 60094 216200
rect 60150 216144 62100 216200
rect 60089 216142 62100 216144
rect 60089 216139 60155 216142
rect -960 208178 480 208268
rect 3141 208178 3207 208181
rect -960 208176 3207 208178
rect -960 208120 3146 208176
rect 3202 208120 3207 208176
rect -960 208118 3207 208120
rect -960 208028 480 208118
rect 3141 208115 3207 208118
rect 523677 205322 523743 205325
rect 521916 205320 523743 205322
rect 521916 205264 523682 205320
rect 523738 205264 523743 205320
rect 521916 205262 523743 205264
rect 523677 205259 523743 205262
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 59353 201922 59419 201925
rect 59353 201920 62100 201922
rect 59353 201864 59358 201920
rect 59414 201864 62100 201920
rect 59353 201862 62100 201864
rect 59353 201859 59419 201862
rect -960 193898 480 193988
rect 3601 193898 3667 193901
rect -960 193896 3667 193898
rect -960 193840 3606 193896
rect 3662 193840 3667 193896
rect -960 193838 3667 193840
rect -960 193748 480 193838
rect 3601 193835 3667 193838
rect 583520 193476 584960 193716
rect 523769 191994 523835 191997
rect 521916 191992 523835 191994
rect 521916 191936 523774 191992
rect 523830 191936 523835 191992
rect 521916 191934 523835 191936
rect 523769 191931 523835 191934
rect 59353 187642 59419 187645
rect 59353 187640 62100 187642
rect 59353 187584 59358 187640
rect 59414 187584 62100 187640
rect 59353 187582 62100 187584
rect 59353 187579 59419 187582
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3693 179482 3759 179485
rect -960 179480 3759 179482
rect -960 179424 3698 179480
rect 3754 179424 3759 179480
rect -960 179422 3759 179424
rect -960 179332 480 179422
rect 3693 179419 3759 179422
rect 523861 178666 523927 178669
rect 521916 178664 523927 178666
rect 521916 178608 523866 178664
rect 523922 178608 523927 178664
rect 521916 178606 523927 178608
rect 523861 178603 523927 178606
rect 59997 173362 60063 173365
rect 59997 173360 62100 173362
rect 59997 173304 60002 173360
rect 60058 173304 62100 173360
rect 59997 173302 62100 173304
rect 59997 173299 60063 173302
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 523677 165338 523743 165341
rect 521916 165336 523743 165338
rect 521916 165280 523682 165336
rect 523738 165280 523743 165336
rect 521916 165278 523743 165280
rect 523677 165275 523743 165278
rect -960 165066 480 165156
rect 3417 165066 3483 165069
rect -960 165064 3483 165066
rect -960 165008 3422 165064
rect 3478 165008 3483 165064
rect -960 165006 3483 165008
rect -960 164916 480 165006
rect 3417 165003 3483 165006
rect 59353 159082 59419 159085
rect 59353 159080 62100 159082
rect 59353 159024 59358 159080
rect 59414 159024 62100 159080
rect 59353 159022 62100 159024
rect 59353 159019 59419 159022
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 523769 152010 523835 152013
rect 521916 152008 523835 152010
rect 521916 151952 523774 152008
rect 523830 151952 523835 152008
rect 521916 151950 523835 151952
rect 523769 151947 523835 151950
rect -960 150786 480 150876
rect 3509 150786 3575 150789
rect -960 150784 3575 150786
rect -960 150728 3514 150784
rect 3570 150728 3575 150784
rect -960 150726 3575 150728
rect -960 150636 480 150726
rect 3509 150723 3575 150726
rect 583520 146556 584960 146796
rect 59353 144802 59419 144805
rect 59353 144800 62100 144802
rect 59353 144744 59358 144800
rect 59414 144744 62100 144800
rect 59353 144742 62100 144744
rect 59353 144739 59419 144742
rect 523861 138682 523927 138685
rect 521916 138680 523927 138682
rect 521916 138624 523866 138680
rect 523922 138624 523927 138680
rect 521916 138622 523927 138624
rect 523861 138619 523927 138622
rect -960 136370 480 136460
rect 3601 136370 3667 136373
rect -960 136368 3667 136370
rect -960 136312 3606 136368
rect 3662 136312 3667 136368
rect -960 136310 3667 136312
rect -960 136220 480 136310
rect 3601 136307 3667 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 60089 130522 60155 130525
rect 60089 130520 62100 130522
rect 60089 130464 60094 130520
rect 60150 130464 62100 130520
rect 60089 130462 62100 130464
rect 60089 130459 60155 130462
rect 523677 125354 523743 125357
rect 521916 125352 523743 125354
rect 521916 125296 523682 125352
rect 523738 125296 523743 125352
rect 521916 125294 523743 125296
rect 523677 125291 523743 125294
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2957 122090 3023 122093
rect -960 122088 3023 122090
rect -960 122032 2962 122088
rect 3018 122032 3023 122088
rect -960 122030 3023 122032
rect -960 121940 480 122030
rect 2957 122027 3023 122030
rect 59353 116242 59419 116245
rect 59353 116240 62100 116242
rect 59353 116184 59358 116240
rect 59414 116184 62100 116240
rect 59353 116182 62100 116184
rect 59353 116179 59419 116182
rect 523769 112026 523835 112029
rect 521916 112024 523835 112026
rect 521916 111968 523774 112024
rect 523830 111968 523835 112024
rect 521916 111966 523835 111968
rect 523769 111963 523835 111966
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3417 107674 3483 107677
rect -960 107672 3483 107674
rect -960 107616 3422 107672
rect 3478 107616 3483 107672
rect -960 107614 3483 107616
rect -960 107524 480 107614
rect 3417 107611 3483 107614
rect 59353 101962 59419 101965
rect 59353 101960 62100 101962
rect 59353 101904 59358 101960
rect 59414 101904 62100 101960
rect 59353 101902 62100 101904
rect 59353 101899 59419 101902
rect 583520 99636 584960 99876
rect 523861 98698 523927 98701
rect 521916 98696 523927 98698
rect 521916 98640 523866 98696
rect 523922 98640 523927 98696
rect 521916 98638 523927 98640
rect 523861 98635 523927 98638
rect -960 93258 480 93348
rect 3693 93258 3759 93261
rect -960 93256 3759 93258
rect -960 93200 3698 93256
rect 3754 93200 3759 93256
rect -960 93198 3759 93200
rect -960 93108 480 93198
rect 3693 93195 3759 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 59997 87682 60063 87685
rect 59997 87680 62100 87682
rect 59997 87624 60002 87680
rect 60058 87624 62100 87680
rect 59997 87622 62100 87624
rect 59997 87619 60063 87622
rect 523677 85370 523743 85373
rect 521916 85368 523743 85370
rect 521916 85312 523682 85368
rect 523738 85312 523743 85368
rect 521916 85310 523743 85312
rect 523677 85307 523743 85310
rect -960 78978 480 79068
rect 3049 78978 3115 78981
rect -960 78976 3115 78978
rect -960 78920 3054 78976
rect 3110 78920 3115 78976
rect -960 78918 3115 78920
rect -960 78828 480 78918
rect 3049 78915 3115 78918
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 59353 73402 59419 73405
rect 59353 73400 62100 73402
rect 59353 73344 59358 73400
rect 59414 73344 62100 73400
rect 59353 73342 62100 73344
rect 59353 73339 59419 73342
rect 523769 72042 523835 72045
rect 521916 72040 523835 72042
rect 521916 71984 523774 72040
rect 523830 71984 523835 72040
rect 521916 71982 523835 71984
rect 523769 71979 523835 71982
rect -960 64562 480 64652
rect 3509 64562 3575 64565
rect -960 64560 3575 64562
rect -960 64504 3514 64560
rect 3570 64504 3575 64560
rect -960 64502 3575 64504
rect -960 64412 480 64502
rect 3509 64499 3575 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 59353 59122 59419 59125
rect 59353 59120 62100 59122
rect 59353 59064 59358 59120
rect 59414 59064 62100 59120
rect 59353 59062 62100 59064
rect 59353 59059 59419 59062
rect 523861 58714 523927 58717
rect 521916 58712 523927 58714
rect 521916 58656 523866 58712
rect 523922 58656 523927 58712
rect 521916 58654 523927 58656
rect 523861 58651 523927 58654
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3601 50146 3667 50149
rect -960 50144 3667 50146
rect -960 50088 3606 50144
rect 3662 50088 3667 50144
rect -960 50086 3667 50088
rect -960 49996 480 50086
rect 3601 50083 3667 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3325 35866 3391 35869
rect -960 35864 3391 35866
rect -960 35808 3330 35864
rect 3386 35808 3391 35864
rect -960 35806 3391 35808
rect -960 35716 480 35806
rect 3325 35803 3391 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3417 21450 3483 21453
rect -960 21448 3483 21450
rect -960 21392 3422 21448
rect 3478 21392 3483 21448
rect -960 21390 3483 21392
rect -960 21300 480 21390
rect 3417 21387 3483 21390
rect 580073 17642 580139 17645
rect 583520 17642 584960 17732
rect 580073 17640 584960 17642
rect 580073 17584 580078 17640
rect 580134 17584 584960 17640
rect 580073 17582 584960 17584
rect 580073 17579 580139 17582
rect 583520 17492 584960 17582
rect 515949 9754 516015 9757
rect 516133 9754 516199 9757
rect 515949 9752 516199 9754
rect 515949 9696 515954 9752
rect 516010 9696 516138 9752
rect 516194 9696 516199 9752
rect 515949 9694 516199 9696
rect 515949 9691 516015 9694
rect 516133 9691 516199 9694
rect -960 7170 480 7260
rect 3509 7170 3575 7173
rect -960 7168 3575 7170
rect -960 7112 3514 7168
rect 3570 7112 3575 7168
rect -960 7110 3575 7112
rect -960 7020 480 7110
rect 3509 7107 3575 7110
rect 583520 5796 584960 6036
rect 485681 3634 485747 3637
rect 546493 3634 546559 3637
rect 485681 3632 546559 3634
rect 485681 3576 485686 3632
rect 485742 3576 546498 3632
rect 546554 3576 546559 3632
rect 485681 3574 546559 3576
rect 485681 3571 485747 3574
rect 546493 3571 546559 3574
rect 85481 3498 85547 3501
rect 146845 3498 146911 3501
rect 85481 3496 146911 3498
rect 85481 3440 85486 3496
rect 85542 3440 146850 3496
rect 146906 3440 146911 3496
rect 85481 3438 146911 3440
rect 85481 3435 85547 3438
rect 146845 3435 146911 3438
rect 364241 3498 364307 3501
rect 425145 3498 425211 3501
rect 364241 3496 425211 3498
rect 364241 3440 364246 3496
rect 364302 3440 425150 3496
rect 425206 3440 425211 3496
rect 364241 3438 425211 3440
rect 364241 3435 364307 3438
rect 425145 3435 425211 3438
rect 449801 3498 449867 3501
rect 510797 3498 510863 3501
rect 449801 3496 510863 3498
rect 449801 3440 449806 3496
rect 449862 3440 510802 3496
rect 510858 3440 510863 3496
rect 449801 3438 510863 3440
rect 449801 3435 449867 3438
rect 510797 3435 510863 3438
rect 92381 3362 92447 3365
rect 153929 3362 153995 3365
rect 92381 3360 153995 3362
rect 92381 3304 92386 3360
rect 92442 3304 153934 3360
rect 153990 3304 153995 3360
rect 92381 3302 153995 3304
rect 92381 3299 92447 3302
rect 153929 3299 153995 3302
rect 339401 3362 339467 3365
rect 400213 3362 400279 3365
rect 339401 3360 400279 3362
rect 339401 3304 339406 3360
rect 339462 3304 400218 3360
rect 400274 3304 400279 3360
rect 339401 3302 400279 3304
rect 339401 3299 339467 3302
rect 400213 3299 400279 3302
rect 407021 3362 407087 3365
rect 467925 3362 467991 3365
rect 407021 3360 467991 3362
rect 407021 3304 407026 3360
rect 407082 3304 467930 3360
rect 467986 3304 467991 3360
rect 407021 3302 467991 3304
rect 407021 3299 407087 3302
rect 467925 3299 467991 3302
rect 520181 3362 520247 3365
rect 580993 3362 581059 3365
rect 520181 3360 581059 3362
rect 520181 3304 520186 3360
rect 520242 3304 580998 3360
rect 581054 3304 581059 3360
rect 520181 3302 581059 3304
rect 520181 3299 520247 3302
rect 580993 3299 581059 3302
<< metal4 >>
rect -2956 705798 -2356 705820
rect -2956 705562 -2774 705798
rect -2538 705562 -2356 705798
rect -2956 705478 -2356 705562
rect -2956 705242 -2774 705478
rect -2538 705242 -2356 705478
rect -2956 668454 -2356 705242
rect -2956 668218 -2774 668454
rect -2538 668218 -2356 668454
rect -2956 668134 -2356 668218
rect -2956 667898 -2774 668134
rect -2538 667898 -2356 668134
rect -2956 632454 -2356 667898
rect -2956 632218 -2774 632454
rect -2538 632218 -2356 632454
rect -2956 632134 -2356 632218
rect -2956 631898 -2774 632134
rect -2538 631898 -2356 632134
rect -2956 596454 -2356 631898
rect -2956 596218 -2774 596454
rect -2538 596218 -2356 596454
rect -2956 596134 -2356 596218
rect -2956 595898 -2774 596134
rect -2538 595898 -2356 596134
rect -2956 560454 -2356 595898
rect -2956 560218 -2774 560454
rect -2538 560218 -2356 560454
rect -2956 560134 -2356 560218
rect -2956 559898 -2774 560134
rect -2538 559898 -2356 560134
rect -2956 524454 -2356 559898
rect -2956 524218 -2774 524454
rect -2538 524218 -2356 524454
rect -2956 524134 -2356 524218
rect -2956 523898 -2774 524134
rect -2538 523898 -2356 524134
rect -2956 488454 -2356 523898
rect -2956 488218 -2774 488454
rect -2538 488218 -2356 488454
rect -2956 488134 -2356 488218
rect -2956 487898 -2774 488134
rect -2538 487898 -2356 488134
rect -2956 452454 -2356 487898
rect -2956 452218 -2774 452454
rect -2538 452218 -2356 452454
rect -2956 452134 -2356 452218
rect -2956 451898 -2774 452134
rect -2538 451898 -2356 452134
rect -2956 416454 -2356 451898
rect -2956 416218 -2774 416454
rect -2538 416218 -2356 416454
rect -2956 416134 -2356 416218
rect -2956 415898 -2774 416134
rect -2538 415898 -2356 416134
rect -2956 380454 -2356 415898
rect -2956 380218 -2774 380454
rect -2538 380218 -2356 380454
rect -2956 380134 -2356 380218
rect -2956 379898 -2774 380134
rect -2538 379898 -2356 380134
rect -2956 344454 -2356 379898
rect -2956 344218 -2774 344454
rect -2538 344218 -2356 344454
rect -2956 344134 -2356 344218
rect -2956 343898 -2774 344134
rect -2538 343898 -2356 344134
rect -2956 308454 -2356 343898
rect -2956 308218 -2774 308454
rect -2538 308218 -2356 308454
rect -2956 308134 -2356 308218
rect -2956 307898 -2774 308134
rect -2538 307898 -2356 308134
rect -2956 272454 -2356 307898
rect -2956 272218 -2774 272454
rect -2538 272218 -2356 272454
rect -2956 272134 -2356 272218
rect -2956 271898 -2774 272134
rect -2538 271898 -2356 272134
rect -2956 236454 -2356 271898
rect -2956 236218 -2774 236454
rect -2538 236218 -2356 236454
rect -2956 236134 -2356 236218
rect -2956 235898 -2774 236134
rect -2538 235898 -2356 236134
rect -2956 200454 -2356 235898
rect -2956 200218 -2774 200454
rect -2538 200218 -2356 200454
rect -2956 200134 -2356 200218
rect -2956 199898 -2774 200134
rect -2538 199898 -2356 200134
rect -2956 164454 -2356 199898
rect -2956 164218 -2774 164454
rect -2538 164218 -2356 164454
rect -2956 164134 -2356 164218
rect -2956 163898 -2774 164134
rect -2538 163898 -2356 164134
rect -2956 128454 -2356 163898
rect -2956 128218 -2774 128454
rect -2538 128218 -2356 128454
rect -2956 128134 -2356 128218
rect -2956 127898 -2774 128134
rect -2538 127898 -2356 128134
rect -2956 92454 -2356 127898
rect -2956 92218 -2774 92454
rect -2538 92218 -2356 92454
rect -2956 92134 -2356 92218
rect -2956 91898 -2774 92134
rect -2538 91898 -2356 92134
rect -2956 56454 -2356 91898
rect -2956 56218 -2774 56454
rect -2538 56218 -2356 56454
rect -2956 56134 -2356 56218
rect -2956 55898 -2774 56134
rect -2538 55898 -2356 56134
rect -2956 20454 -2356 55898
rect -2956 20218 -2774 20454
rect -2538 20218 -2356 20454
rect -2956 20134 -2356 20218
rect -2956 19898 -2774 20134
rect -2538 19898 -2356 20134
rect -2956 -1306 -2356 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705820
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2956 -1542 -2774 -1306
rect -2538 -1542 -2356 -1306
rect -2956 -1626 -2356 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 -2356 -1626
rect -2956 -1884 -2356 -1862
rect 804 -1884 1404 -902
rect 18804 705798 19404 705820
rect 18804 705562 18986 705798
rect 19222 705562 19404 705798
rect 18804 705478 19404 705562
rect 18804 705242 18986 705478
rect 19222 705242 19404 705478
rect 18804 668454 19404 705242
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1306 19404 19898
rect 18804 -1542 18986 -1306
rect 19222 -1542 19404 -1306
rect 18804 -1626 19404 -1542
rect 18804 -1862 18986 -1626
rect 19222 -1862 19404 -1626
rect 18804 -1884 19404 -1862
rect 36804 704838 37404 705820
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1884 37404 -902
rect 54804 705798 55404 705820
rect 54804 705562 54986 705798
rect 55222 705562 55404 705798
rect 54804 705478 55404 705562
rect 54804 705242 54986 705478
rect 55222 705242 55404 705478
rect 54804 668454 55404 705242
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 72804 704838 73404 705820
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 652000 73404 685898
rect 90804 705798 91404 705820
rect 90804 705562 90986 705798
rect 91222 705562 91404 705798
rect 90804 705478 91404 705562
rect 90804 705242 90986 705478
rect 91222 705242 91404 705478
rect 90804 668454 91404 705242
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 652000 91404 667898
rect 108804 704838 109404 705820
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 652000 109404 685898
rect 126804 705798 127404 705820
rect 126804 705562 126986 705798
rect 127222 705562 127404 705798
rect 126804 705478 127404 705562
rect 126804 705242 126986 705478
rect 127222 705242 127404 705478
rect 126804 668454 127404 705242
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 652000 127404 667898
rect 144804 704838 145404 705820
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 652000 145404 685898
rect 162804 705798 163404 705820
rect 162804 705562 162986 705798
rect 163222 705562 163404 705798
rect 162804 705478 163404 705562
rect 162804 705242 162986 705478
rect 163222 705242 163404 705478
rect 162804 668454 163404 705242
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 652000 163404 667898
rect 180804 704838 181404 705820
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 652000 181404 685898
rect 198804 705798 199404 705820
rect 198804 705562 198986 705798
rect 199222 705562 199404 705798
rect 198804 705478 199404 705562
rect 198804 705242 198986 705478
rect 199222 705242 199404 705478
rect 198804 668454 199404 705242
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 652000 199404 667898
rect 216804 704838 217404 705820
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 652000 217404 685898
rect 234804 705798 235404 705820
rect 234804 705562 234986 705798
rect 235222 705562 235404 705798
rect 234804 705478 235404 705562
rect 234804 705242 234986 705478
rect 235222 705242 235404 705478
rect 234804 668454 235404 705242
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 652000 235404 667898
rect 252804 704838 253404 705820
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 652000 253404 685898
rect 270804 705798 271404 705820
rect 270804 705562 270986 705798
rect 271222 705562 271404 705798
rect 270804 705478 271404 705562
rect 270804 705242 270986 705478
rect 271222 705242 271404 705478
rect 270804 668454 271404 705242
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 652000 271404 667898
rect 288804 704838 289404 705820
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 652000 289404 685898
rect 306804 705798 307404 705820
rect 306804 705562 306986 705798
rect 307222 705562 307404 705798
rect 306804 705478 307404 705562
rect 306804 705242 306986 705478
rect 307222 705242 307404 705478
rect 306804 668454 307404 705242
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 652000 307404 667898
rect 324804 704838 325404 705820
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 652000 325404 685898
rect 342804 705798 343404 705820
rect 342804 705562 342986 705798
rect 343222 705562 343404 705798
rect 342804 705478 343404 705562
rect 342804 705242 342986 705478
rect 343222 705242 343404 705478
rect 342804 668454 343404 705242
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 652000 343404 667898
rect 360804 704838 361404 705820
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 652000 361404 685898
rect 378804 705798 379404 705820
rect 378804 705562 378986 705798
rect 379222 705562 379404 705798
rect 378804 705478 379404 705562
rect 378804 705242 378986 705478
rect 379222 705242 379404 705478
rect 378804 668454 379404 705242
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 652000 379404 667898
rect 396804 704838 397404 705820
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 652000 397404 685898
rect 414804 705798 415404 705820
rect 414804 705562 414986 705798
rect 415222 705562 415404 705798
rect 414804 705478 415404 705562
rect 414804 705242 414986 705478
rect 415222 705242 415404 705478
rect 414804 668454 415404 705242
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 652000 415404 667898
rect 432804 704838 433404 705820
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 652000 433404 685898
rect 450804 705798 451404 705820
rect 450804 705562 450986 705798
rect 451222 705562 451404 705798
rect 450804 705478 451404 705562
rect 450804 705242 450986 705478
rect 451222 705242 451404 705478
rect 450804 668454 451404 705242
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 652000 451404 667898
rect 468804 704838 469404 705820
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 652000 469404 685898
rect 486804 705798 487404 705820
rect 486804 705562 486986 705798
rect 487222 705562 487404 705798
rect 486804 705478 487404 705562
rect 486804 705242 486986 705478
rect 487222 705242 487404 705478
rect 486804 668454 487404 705242
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 652000 487404 667898
rect 504804 704838 505404 705820
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 652000 505404 685898
rect 522804 705798 523404 705820
rect 522804 705562 522986 705798
rect 523222 705562 523404 705798
rect 522804 705478 523404 705562
rect 522804 705242 522986 705478
rect 523222 705242 523404 705478
rect 522804 668454 523404 705242
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 81568 632454 81888 632476
rect 81568 632218 81610 632454
rect 81846 632218 81888 632454
rect 81568 632134 81888 632218
rect 81568 631898 81610 632134
rect 81846 631898 81888 632134
rect 81568 631876 81888 631898
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 66208 614454 66528 614476
rect 66208 614218 66250 614454
rect 66486 614218 66528 614454
rect 66208 614134 66528 614218
rect 66208 613898 66250 614134
rect 66486 613898 66528 614134
rect 66208 613876 66528 613898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 81568 596454 81888 596476
rect 81568 596218 81610 596454
rect 81846 596218 81888 596454
rect 81568 596134 81888 596218
rect 81568 595898 81610 596134
rect 81846 595898 81888 596134
rect 81568 595876 81888 595898
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 66208 578454 66528 578476
rect 66208 578218 66250 578454
rect 66486 578218 66528 578454
rect 66208 578134 66528 578218
rect 66208 577898 66250 578134
rect 66486 577898 66528 578134
rect 66208 577876 66528 577898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 81568 560454 81888 560476
rect 81568 560218 81610 560454
rect 81846 560218 81888 560454
rect 81568 560134 81888 560218
rect 81568 559898 81610 560134
rect 81846 559898 81888 560134
rect 81568 559876 81888 559898
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 66208 542454 66528 542476
rect 66208 542218 66250 542454
rect 66486 542218 66528 542454
rect 66208 542134 66528 542218
rect 66208 541898 66250 542134
rect 66486 541898 66528 542134
rect 66208 541876 66528 541898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 81568 524454 81888 524476
rect 81568 524218 81610 524454
rect 81846 524218 81888 524454
rect 81568 524134 81888 524218
rect 81568 523898 81610 524134
rect 81846 523898 81888 524134
rect 81568 523876 81888 523898
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 66208 506454 66528 506476
rect 66208 506218 66250 506454
rect 66486 506218 66528 506454
rect 66208 506134 66528 506218
rect 66208 505898 66250 506134
rect 66486 505898 66528 506134
rect 66208 505876 66528 505898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 81568 488454 81888 488476
rect 81568 488218 81610 488454
rect 81846 488218 81888 488454
rect 81568 488134 81888 488218
rect 81568 487898 81610 488134
rect 81846 487898 81888 488134
rect 81568 487876 81888 487898
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 66208 470454 66528 470476
rect 66208 470218 66250 470454
rect 66486 470218 66528 470454
rect 66208 470134 66528 470218
rect 66208 469898 66250 470134
rect 66486 469898 66528 470134
rect 66208 469876 66528 469898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 81568 452454 81888 452476
rect 81568 452218 81610 452454
rect 81846 452218 81888 452454
rect 81568 452134 81888 452218
rect 81568 451898 81610 452134
rect 81846 451898 81888 452134
rect 81568 451876 81888 451898
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 66208 434454 66528 434476
rect 66208 434218 66250 434454
rect 66486 434218 66528 434454
rect 66208 434134 66528 434218
rect 66208 433898 66250 434134
rect 66486 433898 66528 434134
rect 66208 433876 66528 433898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 81568 416454 81888 416476
rect 81568 416218 81610 416454
rect 81846 416218 81888 416454
rect 81568 416134 81888 416218
rect 81568 415898 81610 416134
rect 81846 415898 81888 416134
rect 81568 415876 81888 415898
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 66208 398454 66528 398476
rect 66208 398218 66250 398454
rect 66486 398218 66528 398454
rect 66208 398134 66528 398218
rect 66208 397898 66250 398134
rect 66486 397898 66528 398134
rect 66208 397876 66528 397898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 81568 380454 81888 380476
rect 81568 380218 81610 380454
rect 81846 380218 81888 380454
rect 81568 380134 81888 380218
rect 81568 379898 81610 380134
rect 81846 379898 81888 380134
rect 81568 379876 81888 379898
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 66208 362454 66528 362476
rect 66208 362218 66250 362454
rect 66486 362218 66528 362454
rect 66208 362134 66528 362218
rect 66208 361898 66250 362134
rect 66486 361898 66528 362134
rect 66208 361876 66528 361898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 81568 344454 81888 344476
rect 81568 344218 81610 344454
rect 81846 344218 81888 344454
rect 81568 344134 81888 344218
rect 81568 343898 81610 344134
rect 81846 343898 81888 344134
rect 81568 343876 81888 343898
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 66208 326454 66528 326476
rect 66208 326218 66250 326454
rect 66486 326218 66528 326454
rect 66208 326134 66528 326218
rect 66208 325898 66250 326134
rect 66486 325898 66528 326134
rect 66208 325876 66528 325898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 81568 308454 81888 308476
rect 81568 308218 81610 308454
rect 81846 308218 81888 308454
rect 81568 308134 81888 308218
rect 81568 307898 81610 308134
rect 81846 307898 81888 308134
rect 81568 307876 81888 307898
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 66208 290454 66528 290476
rect 66208 290218 66250 290454
rect 66486 290218 66528 290454
rect 66208 290134 66528 290218
rect 66208 289898 66250 290134
rect 66486 289898 66528 290134
rect 66208 289876 66528 289898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 81568 272454 81888 272476
rect 81568 272218 81610 272454
rect 81846 272218 81888 272454
rect 81568 272134 81888 272218
rect 81568 271898 81610 272134
rect 81846 271898 81888 272134
rect 81568 271876 81888 271898
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 66208 254454 66528 254476
rect 66208 254218 66250 254454
rect 66486 254218 66528 254454
rect 66208 254134 66528 254218
rect 66208 253898 66250 254134
rect 66486 253898 66528 254134
rect 66208 253876 66528 253898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 81568 236454 81888 236476
rect 81568 236218 81610 236454
rect 81846 236218 81888 236454
rect 81568 236134 81888 236218
rect 81568 235898 81610 236134
rect 81846 235898 81888 236134
rect 81568 235876 81888 235898
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 66208 218454 66528 218476
rect 66208 218218 66250 218454
rect 66486 218218 66528 218454
rect 66208 218134 66528 218218
rect 66208 217898 66250 218134
rect 66486 217898 66528 218134
rect 66208 217876 66528 217898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 81568 200454 81888 200476
rect 81568 200218 81610 200454
rect 81846 200218 81888 200454
rect 81568 200134 81888 200218
rect 81568 199898 81610 200134
rect 81846 199898 81888 200134
rect 81568 199876 81888 199898
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 66208 182454 66528 182476
rect 66208 182218 66250 182454
rect 66486 182218 66528 182454
rect 66208 182134 66528 182218
rect 66208 181898 66250 182134
rect 66486 181898 66528 182134
rect 66208 181876 66528 181898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 81568 164454 81888 164476
rect 81568 164218 81610 164454
rect 81846 164218 81888 164454
rect 81568 164134 81888 164218
rect 81568 163898 81610 164134
rect 81846 163898 81888 164134
rect 81568 163876 81888 163898
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 66208 146454 66528 146476
rect 66208 146218 66250 146454
rect 66486 146218 66528 146454
rect 66208 146134 66528 146218
rect 66208 145898 66250 146134
rect 66486 145898 66528 146134
rect 66208 145876 66528 145898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 81568 128454 81888 128476
rect 81568 128218 81610 128454
rect 81846 128218 81888 128454
rect 81568 128134 81888 128218
rect 81568 127898 81610 128134
rect 81846 127898 81888 128134
rect 81568 127876 81888 127898
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 66208 110454 66528 110476
rect 66208 110218 66250 110454
rect 66486 110218 66528 110454
rect 66208 110134 66528 110218
rect 66208 109898 66250 110134
rect 66486 109898 66528 110134
rect 66208 109876 66528 109898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 81568 92454 81888 92476
rect 81568 92218 81610 92454
rect 81846 92218 81888 92454
rect 81568 92134 81888 92218
rect 81568 91898 81610 92134
rect 81846 91898 81888 92134
rect 81568 91876 81888 91898
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 66208 74454 66528 74476
rect 66208 74218 66250 74454
rect 66486 74218 66528 74454
rect 66208 74134 66528 74218
rect 66208 73898 66250 74134
rect 66486 73898 66528 74134
rect 66208 73876 66528 73898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 81568 56454 81888 56476
rect 81568 56218 81610 56454
rect 81846 56218 81888 56454
rect 81568 56134 81888 56218
rect 81568 55898 81610 56134
rect 81846 55898 81888 56134
rect 81568 55876 81888 55898
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1306 55404 19898
rect 54804 -1542 54986 -1306
rect 55222 -1542 55404 -1306
rect 54804 -1626 55404 -1542
rect 54804 -1862 54986 -1626
rect 55222 -1862 55404 -1626
rect 54804 -1884 55404 -1862
rect 72804 38454 73404 52000
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1884 73404 -902
rect 90804 20454 91404 52000
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1306 91404 19898
rect 90804 -1542 90986 -1306
rect 91222 -1542 91404 -1306
rect 90804 -1626 91404 -1542
rect 90804 -1862 90986 -1626
rect 91222 -1862 91404 -1626
rect 90804 -1884 91404 -1862
rect 108804 38454 109404 52000
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1884 109404 -902
rect 126804 20454 127404 52000
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1306 127404 19898
rect 126804 -1542 126986 -1306
rect 127222 -1542 127404 -1306
rect 126804 -1626 127404 -1542
rect 126804 -1862 126986 -1626
rect 127222 -1862 127404 -1626
rect 126804 -1884 127404 -1862
rect 144804 38454 145404 52000
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1884 145404 -902
rect 162804 20454 163404 52000
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1306 163404 19898
rect 162804 -1542 162986 -1306
rect 163222 -1542 163404 -1306
rect 162804 -1626 163404 -1542
rect 162804 -1862 162986 -1626
rect 163222 -1862 163404 -1626
rect 162804 -1884 163404 -1862
rect 180804 38454 181404 52000
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1884 181404 -902
rect 198804 20454 199404 52000
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1306 199404 19898
rect 198804 -1542 198986 -1306
rect 199222 -1542 199404 -1306
rect 198804 -1626 199404 -1542
rect 198804 -1862 198986 -1626
rect 199222 -1862 199404 -1626
rect 198804 -1884 199404 -1862
rect 216804 38454 217404 52000
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1884 217404 -902
rect 234804 20454 235404 52000
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1306 235404 19898
rect 234804 -1542 234986 -1306
rect 235222 -1542 235404 -1306
rect 234804 -1626 235404 -1542
rect 234804 -1862 234986 -1626
rect 235222 -1862 235404 -1626
rect 234804 -1884 235404 -1862
rect 252804 38454 253404 52000
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1884 253404 -902
rect 270804 20454 271404 52000
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1306 271404 19898
rect 270804 -1542 270986 -1306
rect 271222 -1542 271404 -1306
rect 270804 -1626 271404 -1542
rect 270804 -1862 270986 -1626
rect 271222 -1862 271404 -1626
rect 270804 -1884 271404 -1862
rect 288804 38454 289404 52000
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1884 289404 -902
rect 306804 20454 307404 52000
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1306 307404 19898
rect 306804 -1542 306986 -1306
rect 307222 -1542 307404 -1306
rect 306804 -1626 307404 -1542
rect 306804 -1862 306986 -1626
rect 307222 -1862 307404 -1626
rect 306804 -1884 307404 -1862
rect 324804 38454 325404 52000
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1884 325404 -902
rect 342804 20454 343404 52000
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1306 343404 19898
rect 342804 -1542 342986 -1306
rect 343222 -1542 343404 -1306
rect 342804 -1626 343404 -1542
rect 342804 -1862 342986 -1626
rect 343222 -1862 343404 -1626
rect 342804 -1884 343404 -1862
rect 360804 38454 361404 52000
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1884 361404 -902
rect 378804 20454 379404 52000
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1306 379404 19898
rect 378804 -1542 378986 -1306
rect 379222 -1542 379404 -1306
rect 378804 -1626 379404 -1542
rect 378804 -1862 378986 -1626
rect 379222 -1862 379404 -1626
rect 378804 -1884 379404 -1862
rect 396804 38454 397404 52000
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1884 397404 -902
rect 414804 20454 415404 52000
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1306 415404 19898
rect 414804 -1542 414986 -1306
rect 415222 -1542 415404 -1306
rect 414804 -1626 415404 -1542
rect 414804 -1862 414986 -1626
rect 415222 -1862 415404 -1626
rect 414804 -1884 415404 -1862
rect 432804 38454 433404 52000
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1884 433404 -902
rect 450804 20454 451404 52000
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1306 451404 19898
rect 450804 -1542 450986 -1306
rect 451222 -1542 451404 -1306
rect 450804 -1626 451404 -1542
rect 450804 -1862 450986 -1626
rect 451222 -1862 451404 -1626
rect 450804 -1884 451404 -1862
rect 468804 38454 469404 52000
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1884 469404 -902
rect 486804 20454 487404 52000
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1306 487404 19898
rect 486804 -1542 486986 -1306
rect 487222 -1542 487404 -1306
rect 486804 -1626 487404 -1542
rect 486804 -1862 486986 -1626
rect 487222 -1862 487404 -1626
rect 486804 -1884 487404 -1862
rect 504804 38454 505404 52000
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1884 505404 -902
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1306 523404 19898
rect 522804 -1542 522986 -1306
rect 523222 -1542 523404 -1306
rect 522804 -1626 523404 -1542
rect 522804 -1862 522986 -1626
rect 523222 -1862 523404 -1626
rect 522804 -1884 523404 -1862
rect 540804 704838 541404 705820
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1884 541404 -902
rect 558804 705798 559404 705820
rect 558804 705562 558986 705798
rect 559222 705562 559404 705798
rect 558804 705478 559404 705562
rect 558804 705242 558986 705478
rect 559222 705242 559404 705478
rect 558804 668454 559404 705242
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1306 559404 19898
rect 558804 -1542 558986 -1306
rect 559222 -1542 559404 -1306
rect 558804 -1626 559404 -1542
rect 558804 -1862 558986 -1626
rect 559222 -1862 559404 -1626
rect 558804 -1884 559404 -1862
rect 576804 704838 577404 705820
rect 586280 705798 586880 705820
rect 586280 705562 586462 705798
rect 586698 705562 586880 705798
rect 586280 705478 586880 705562
rect 586280 705242 586462 705478
rect 586698 705242 586880 705478
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1884 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586280 668454 586880 705242
rect 586280 668218 586462 668454
rect 586698 668218 586880 668454
rect 586280 668134 586880 668218
rect 586280 667898 586462 668134
rect 586698 667898 586880 668134
rect 586280 632454 586880 667898
rect 586280 632218 586462 632454
rect 586698 632218 586880 632454
rect 586280 632134 586880 632218
rect 586280 631898 586462 632134
rect 586698 631898 586880 632134
rect 586280 596454 586880 631898
rect 586280 596218 586462 596454
rect 586698 596218 586880 596454
rect 586280 596134 586880 596218
rect 586280 595898 586462 596134
rect 586698 595898 586880 596134
rect 586280 560454 586880 595898
rect 586280 560218 586462 560454
rect 586698 560218 586880 560454
rect 586280 560134 586880 560218
rect 586280 559898 586462 560134
rect 586698 559898 586880 560134
rect 586280 524454 586880 559898
rect 586280 524218 586462 524454
rect 586698 524218 586880 524454
rect 586280 524134 586880 524218
rect 586280 523898 586462 524134
rect 586698 523898 586880 524134
rect 586280 488454 586880 523898
rect 586280 488218 586462 488454
rect 586698 488218 586880 488454
rect 586280 488134 586880 488218
rect 586280 487898 586462 488134
rect 586698 487898 586880 488134
rect 586280 452454 586880 487898
rect 586280 452218 586462 452454
rect 586698 452218 586880 452454
rect 586280 452134 586880 452218
rect 586280 451898 586462 452134
rect 586698 451898 586880 452134
rect 586280 416454 586880 451898
rect 586280 416218 586462 416454
rect 586698 416218 586880 416454
rect 586280 416134 586880 416218
rect 586280 415898 586462 416134
rect 586698 415898 586880 416134
rect 586280 380454 586880 415898
rect 586280 380218 586462 380454
rect 586698 380218 586880 380454
rect 586280 380134 586880 380218
rect 586280 379898 586462 380134
rect 586698 379898 586880 380134
rect 586280 344454 586880 379898
rect 586280 344218 586462 344454
rect 586698 344218 586880 344454
rect 586280 344134 586880 344218
rect 586280 343898 586462 344134
rect 586698 343898 586880 344134
rect 586280 308454 586880 343898
rect 586280 308218 586462 308454
rect 586698 308218 586880 308454
rect 586280 308134 586880 308218
rect 586280 307898 586462 308134
rect 586698 307898 586880 308134
rect 586280 272454 586880 307898
rect 586280 272218 586462 272454
rect 586698 272218 586880 272454
rect 586280 272134 586880 272218
rect 586280 271898 586462 272134
rect 586698 271898 586880 272134
rect 586280 236454 586880 271898
rect 586280 236218 586462 236454
rect 586698 236218 586880 236454
rect 586280 236134 586880 236218
rect 586280 235898 586462 236134
rect 586698 235898 586880 236134
rect 586280 200454 586880 235898
rect 586280 200218 586462 200454
rect 586698 200218 586880 200454
rect 586280 200134 586880 200218
rect 586280 199898 586462 200134
rect 586698 199898 586880 200134
rect 586280 164454 586880 199898
rect 586280 164218 586462 164454
rect 586698 164218 586880 164454
rect 586280 164134 586880 164218
rect 586280 163898 586462 164134
rect 586698 163898 586880 164134
rect 586280 128454 586880 163898
rect 586280 128218 586462 128454
rect 586698 128218 586880 128454
rect 586280 128134 586880 128218
rect 586280 127898 586462 128134
rect 586698 127898 586880 128134
rect 586280 92454 586880 127898
rect 586280 92218 586462 92454
rect 586698 92218 586880 92454
rect 586280 92134 586880 92218
rect 586280 91898 586462 92134
rect 586698 91898 586880 92134
rect 586280 56454 586880 91898
rect 586280 56218 586462 56454
rect 586698 56218 586880 56454
rect 586280 56134 586880 56218
rect 586280 55898 586462 56134
rect 586698 55898 586880 56134
rect 586280 20454 586880 55898
rect 586280 20218 586462 20454
rect 586698 20218 586880 20454
rect 586280 20134 586880 20218
rect 586280 19898 586462 20134
rect 586698 19898 586880 20134
rect 586280 -1306 586880 19898
rect 586280 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect 586280 -1626 586880 -1542
rect 586280 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect 586280 -1884 586880 -1862
<< via4 >>
rect -2774 705562 -2538 705798
rect -2774 705242 -2538 705478
rect -2774 668218 -2538 668454
rect -2774 667898 -2538 668134
rect -2774 632218 -2538 632454
rect -2774 631898 -2538 632134
rect -2774 596218 -2538 596454
rect -2774 595898 -2538 596134
rect -2774 560218 -2538 560454
rect -2774 559898 -2538 560134
rect -2774 524218 -2538 524454
rect -2774 523898 -2538 524134
rect -2774 488218 -2538 488454
rect -2774 487898 -2538 488134
rect -2774 452218 -2538 452454
rect -2774 451898 -2538 452134
rect -2774 416218 -2538 416454
rect -2774 415898 -2538 416134
rect -2774 380218 -2538 380454
rect -2774 379898 -2538 380134
rect -2774 344218 -2538 344454
rect -2774 343898 -2538 344134
rect -2774 308218 -2538 308454
rect -2774 307898 -2538 308134
rect -2774 272218 -2538 272454
rect -2774 271898 -2538 272134
rect -2774 236218 -2538 236454
rect -2774 235898 -2538 236134
rect -2774 200218 -2538 200454
rect -2774 199898 -2538 200134
rect -2774 164218 -2538 164454
rect -2774 163898 -2538 164134
rect -2774 128218 -2538 128454
rect -2774 127898 -2538 128134
rect -2774 92218 -2538 92454
rect -2774 91898 -2538 92134
rect -2774 56218 -2538 56454
rect -2774 55898 -2538 56134
rect -2774 20218 -2538 20454
rect -2774 19898 -2538 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2774 -1542 -2538 -1306
rect -2774 -1862 -2538 -1626
rect 18986 705562 19222 705798
rect 18986 705242 19222 705478
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1542 19222 -1306
rect 18986 -1862 19222 -1626
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 705562 55222 705798
rect 54986 705242 55222 705478
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 90986 705562 91222 705798
rect 90986 705242 91222 705478
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 126986 705562 127222 705798
rect 126986 705242 127222 705478
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 162986 705562 163222 705798
rect 162986 705242 163222 705478
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 198986 705562 199222 705798
rect 198986 705242 199222 705478
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 234986 705562 235222 705798
rect 234986 705242 235222 705478
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 270986 705562 271222 705798
rect 270986 705242 271222 705478
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 306986 705562 307222 705798
rect 306986 705242 307222 705478
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 342986 705562 343222 705798
rect 342986 705242 343222 705478
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 378986 705562 379222 705798
rect 378986 705242 379222 705478
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 414986 705562 415222 705798
rect 414986 705242 415222 705478
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 450986 705562 451222 705798
rect 450986 705242 451222 705478
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 486986 705562 487222 705798
rect 486986 705242 487222 705478
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 522986 705562 523222 705798
rect 522986 705242 523222 705478
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 81610 632218 81846 632454
rect 81610 631898 81846 632134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 66250 614218 66486 614454
rect 66250 613898 66486 614134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 81610 596218 81846 596454
rect 81610 595898 81846 596134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 66250 578218 66486 578454
rect 66250 577898 66486 578134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 81610 560218 81846 560454
rect 81610 559898 81846 560134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 66250 542218 66486 542454
rect 66250 541898 66486 542134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 81610 524218 81846 524454
rect 81610 523898 81846 524134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 66250 506218 66486 506454
rect 66250 505898 66486 506134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 81610 488218 81846 488454
rect 81610 487898 81846 488134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 66250 470218 66486 470454
rect 66250 469898 66486 470134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 81610 452218 81846 452454
rect 81610 451898 81846 452134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 66250 434218 66486 434454
rect 66250 433898 66486 434134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 81610 416218 81846 416454
rect 81610 415898 81846 416134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 66250 398218 66486 398454
rect 66250 397898 66486 398134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 81610 380218 81846 380454
rect 81610 379898 81846 380134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 66250 362218 66486 362454
rect 66250 361898 66486 362134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 81610 344218 81846 344454
rect 81610 343898 81846 344134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 66250 326218 66486 326454
rect 66250 325898 66486 326134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 81610 308218 81846 308454
rect 81610 307898 81846 308134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 66250 290218 66486 290454
rect 66250 289898 66486 290134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 81610 272218 81846 272454
rect 81610 271898 81846 272134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 66250 254218 66486 254454
rect 66250 253898 66486 254134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 81610 236218 81846 236454
rect 81610 235898 81846 236134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 66250 218218 66486 218454
rect 66250 217898 66486 218134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 81610 200218 81846 200454
rect 81610 199898 81846 200134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 66250 182218 66486 182454
rect 66250 181898 66486 182134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 81610 164218 81846 164454
rect 81610 163898 81846 164134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 66250 146218 66486 146454
rect 66250 145898 66486 146134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 81610 128218 81846 128454
rect 81610 127898 81846 128134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 66250 110218 66486 110454
rect 66250 109898 66486 110134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 81610 92218 81846 92454
rect 81610 91898 81846 92134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 66250 74218 66486 74454
rect 66250 73898 66486 74134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 81610 56218 81846 56454
rect 81610 55898 81846 56134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1542 55222 -1306
rect 54986 -1862 55222 -1626
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1542 91222 -1306
rect 90986 -1862 91222 -1626
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1542 127222 -1306
rect 126986 -1862 127222 -1626
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1542 163222 -1306
rect 162986 -1862 163222 -1626
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1542 199222 -1306
rect 198986 -1862 199222 -1626
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1542 235222 -1306
rect 234986 -1862 235222 -1626
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1542 271222 -1306
rect 270986 -1862 271222 -1626
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1542 307222 -1306
rect 306986 -1862 307222 -1626
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1542 343222 -1306
rect 342986 -1862 343222 -1626
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1542 379222 -1306
rect 378986 -1862 379222 -1626
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1542 415222 -1306
rect 414986 -1862 415222 -1626
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1542 451222 -1306
rect 450986 -1862 451222 -1626
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1542 487222 -1306
rect 486986 -1862 487222 -1626
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1542 523222 -1306
rect 522986 -1862 523222 -1626
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 705562 559222 705798
rect 558986 705242 559222 705478
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1542 559222 -1306
rect 558986 -1862 559222 -1626
rect 586462 705562 586698 705798
rect 586462 705242 586698 705478
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586462 668218 586698 668454
rect 586462 667898 586698 668134
rect 586462 632218 586698 632454
rect 586462 631898 586698 632134
rect 586462 596218 586698 596454
rect 586462 595898 586698 596134
rect 586462 560218 586698 560454
rect 586462 559898 586698 560134
rect 586462 524218 586698 524454
rect 586462 523898 586698 524134
rect 586462 488218 586698 488454
rect 586462 487898 586698 488134
rect 586462 452218 586698 452454
rect 586462 451898 586698 452134
rect 586462 416218 586698 416454
rect 586462 415898 586698 416134
rect 586462 380218 586698 380454
rect 586462 379898 586698 380134
rect 586462 344218 586698 344454
rect 586462 343898 586698 344134
rect 586462 308218 586698 308454
rect 586462 307898 586698 308134
rect 586462 272218 586698 272454
rect 586462 271898 586698 272134
rect 586462 236218 586698 236454
rect 586462 235898 586698 236134
rect 586462 200218 586698 200454
rect 586462 199898 586698 200134
rect 586462 164218 586698 164454
rect 586462 163898 586698 164134
rect 586462 128218 586698 128454
rect 586462 127898 586698 128134
rect 586462 92218 586698 92454
rect 586462 91898 586698 92134
rect 586462 56218 586698 56454
rect 586462 55898 586698 56134
rect 586462 20218 586698 20454
rect 586462 19898 586698 20134
rect 586462 -1542 586698 -1306
rect 586462 -1862 586698 -1626
<< metal5 >>
rect -2956 705820 -2356 705822
rect 18804 705820 19404 705822
rect 54804 705820 55404 705822
rect 90804 705820 91404 705822
rect 126804 705820 127404 705822
rect 162804 705820 163404 705822
rect 198804 705820 199404 705822
rect 234804 705820 235404 705822
rect 270804 705820 271404 705822
rect 306804 705820 307404 705822
rect 342804 705820 343404 705822
rect 378804 705820 379404 705822
rect 414804 705820 415404 705822
rect 450804 705820 451404 705822
rect 486804 705820 487404 705822
rect 522804 705820 523404 705822
rect 558804 705820 559404 705822
rect 586280 705820 586880 705822
rect -2956 705798 586880 705820
rect -2956 705562 -2774 705798
rect -2538 705562 18986 705798
rect 19222 705562 54986 705798
rect 55222 705562 90986 705798
rect 91222 705562 126986 705798
rect 127222 705562 162986 705798
rect 163222 705562 198986 705798
rect 199222 705562 234986 705798
rect 235222 705562 270986 705798
rect 271222 705562 306986 705798
rect 307222 705562 342986 705798
rect 343222 705562 378986 705798
rect 379222 705562 414986 705798
rect 415222 705562 450986 705798
rect 451222 705562 486986 705798
rect 487222 705562 522986 705798
rect 523222 705562 558986 705798
rect 559222 705562 586462 705798
rect 586698 705562 586880 705798
rect -2956 705478 586880 705562
rect -2956 705242 -2774 705478
rect -2538 705242 18986 705478
rect 19222 705242 54986 705478
rect 55222 705242 90986 705478
rect 91222 705242 126986 705478
rect 127222 705242 162986 705478
rect 163222 705242 198986 705478
rect 199222 705242 234986 705478
rect 235222 705242 270986 705478
rect 271222 705242 306986 705478
rect 307222 705242 342986 705478
rect 343222 705242 378986 705478
rect 379222 705242 414986 705478
rect 415222 705242 450986 705478
rect 451222 705242 486986 705478
rect 487222 705242 522986 705478
rect 523222 705242 558986 705478
rect 559222 705242 586462 705478
rect 586698 705242 586880 705478
rect -2956 705220 586880 705242
rect -2956 705218 -2356 705220
rect 18804 705218 19404 705220
rect 54804 705218 55404 705220
rect 90804 705218 91404 705220
rect 126804 705218 127404 705220
rect 162804 705218 163404 705220
rect 198804 705218 199404 705220
rect 234804 705218 235404 705220
rect 270804 705218 271404 705220
rect 306804 705218 307404 705220
rect 342804 705218 343404 705220
rect 378804 705218 379404 705220
rect 414804 705218 415404 705220
rect 450804 705218 451404 705220
rect 486804 705218 487404 705220
rect 522804 705218 523404 705220
rect 558804 705218 559404 705220
rect 586280 705218 586880 705220
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2956 686454 586880 686476
rect -2956 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586880 686454
rect -2956 686134 586880 686218
rect -2956 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586880 686134
rect -2956 685876 586880 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2956 668476 -2356 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586280 668476 586880 668478
rect -2956 668454 586880 668476
rect -2956 668218 -2774 668454
rect -2538 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586462 668454
rect 586698 668218 586880 668454
rect -2956 668134 586880 668218
rect -2956 667898 -2774 668134
rect -2538 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586462 668134
rect 586698 667898 586880 668134
rect -2956 667876 586880 667898
rect -2956 667874 -2356 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586280 667874 586880 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2956 650454 586880 650476
rect -2956 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586880 650454
rect -2956 650134 586880 650218
rect -2956 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586880 650134
rect -2956 649876 586880 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2956 632476 -2356 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 81568 632476 81888 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586280 632476 586880 632478
rect -2956 632454 586880 632476
rect -2956 632218 -2774 632454
rect -2538 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 81610 632454
rect 81846 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586462 632454
rect 586698 632218 586880 632454
rect -2956 632134 586880 632218
rect -2956 631898 -2774 632134
rect -2538 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 81610 632134
rect 81846 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586462 632134
rect 586698 631898 586880 632134
rect -2956 631876 586880 631898
rect -2956 631874 -2356 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 81568 631874 81888 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586280 631874 586880 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 66208 614476 66528 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2956 614454 586880 614476
rect -2956 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 66250 614454
rect 66486 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586880 614454
rect -2956 614134 586880 614218
rect -2956 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 66250 614134
rect 66486 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586880 614134
rect -2956 613876 586880 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 66208 613874 66528 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2956 596476 -2356 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 81568 596476 81888 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586280 596476 586880 596478
rect -2956 596454 586880 596476
rect -2956 596218 -2774 596454
rect -2538 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 81610 596454
rect 81846 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586462 596454
rect 586698 596218 586880 596454
rect -2956 596134 586880 596218
rect -2956 595898 -2774 596134
rect -2538 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 81610 596134
rect 81846 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586462 596134
rect 586698 595898 586880 596134
rect -2956 595876 586880 595898
rect -2956 595874 -2356 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 81568 595874 81888 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586280 595874 586880 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 66208 578476 66528 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2956 578454 586880 578476
rect -2956 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 66250 578454
rect 66486 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586880 578454
rect -2956 578134 586880 578218
rect -2956 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 66250 578134
rect 66486 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586880 578134
rect -2956 577876 586880 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 66208 577874 66528 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2956 560476 -2356 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 81568 560476 81888 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586280 560476 586880 560478
rect -2956 560454 586880 560476
rect -2956 560218 -2774 560454
rect -2538 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 81610 560454
rect 81846 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586462 560454
rect 586698 560218 586880 560454
rect -2956 560134 586880 560218
rect -2956 559898 -2774 560134
rect -2538 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 81610 560134
rect 81846 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586462 560134
rect 586698 559898 586880 560134
rect -2956 559876 586880 559898
rect -2956 559874 -2356 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 81568 559874 81888 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586280 559874 586880 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 66208 542476 66528 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2956 542454 586880 542476
rect -2956 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 66250 542454
rect 66486 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586880 542454
rect -2956 542134 586880 542218
rect -2956 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 66250 542134
rect 66486 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586880 542134
rect -2956 541876 586880 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 66208 541874 66528 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2956 524476 -2356 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 81568 524476 81888 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586280 524476 586880 524478
rect -2956 524454 586880 524476
rect -2956 524218 -2774 524454
rect -2538 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 81610 524454
rect 81846 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586462 524454
rect 586698 524218 586880 524454
rect -2956 524134 586880 524218
rect -2956 523898 -2774 524134
rect -2538 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 81610 524134
rect 81846 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586462 524134
rect 586698 523898 586880 524134
rect -2956 523876 586880 523898
rect -2956 523874 -2356 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 81568 523874 81888 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586280 523874 586880 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 66208 506476 66528 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2956 506454 586880 506476
rect -2956 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 66250 506454
rect 66486 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586880 506454
rect -2956 506134 586880 506218
rect -2956 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 66250 506134
rect 66486 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586880 506134
rect -2956 505876 586880 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 66208 505874 66528 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -2956 488476 -2356 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 81568 488476 81888 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586280 488476 586880 488478
rect -2956 488454 586880 488476
rect -2956 488218 -2774 488454
rect -2538 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 81610 488454
rect 81846 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586462 488454
rect 586698 488218 586880 488454
rect -2956 488134 586880 488218
rect -2956 487898 -2774 488134
rect -2538 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 81610 488134
rect 81846 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586462 488134
rect 586698 487898 586880 488134
rect -2956 487876 586880 487898
rect -2956 487874 -2356 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 81568 487874 81888 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586280 487874 586880 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 66208 470476 66528 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2956 470454 586880 470476
rect -2956 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 66250 470454
rect 66486 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586880 470454
rect -2956 470134 586880 470218
rect -2956 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 66250 470134
rect 66486 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586880 470134
rect -2956 469876 586880 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 66208 469874 66528 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2956 452476 -2356 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 81568 452476 81888 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586280 452476 586880 452478
rect -2956 452454 586880 452476
rect -2956 452218 -2774 452454
rect -2538 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 81610 452454
rect 81846 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586462 452454
rect 586698 452218 586880 452454
rect -2956 452134 586880 452218
rect -2956 451898 -2774 452134
rect -2538 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 81610 452134
rect 81846 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586462 452134
rect 586698 451898 586880 452134
rect -2956 451876 586880 451898
rect -2956 451874 -2356 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 81568 451874 81888 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586280 451874 586880 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 66208 434476 66528 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2956 434454 586880 434476
rect -2956 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 66250 434454
rect 66486 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586880 434454
rect -2956 434134 586880 434218
rect -2956 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 66250 434134
rect 66486 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586880 434134
rect -2956 433876 586880 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 66208 433874 66528 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -2956 416476 -2356 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 81568 416476 81888 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586280 416476 586880 416478
rect -2956 416454 586880 416476
rect -2956 416218 -2774 416454
rect -2538 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 81610 416454
rect 81846 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586462 416454
rect 586698 416218 586880 416454
rect -2956 416134 586880 416218
rect -2956 415898 -2774 416134
rect -2538 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 81610 416134
rect 81846 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586462 416134
rect 586698 415898 586880 416134
rect -2956 415876 586880 415898
rect -2956 415874 -2356 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 81568 415874 81888 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586280 415874 586880 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 66208 398476 66528 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2956 398454 586880 398476
rect -2956 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 66250 398454
rect 66486 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586880 398454
rect -2956 398134 586880 398218
rect -2956 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 66250 398134
rect 66486 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586880 398134
rect -2956 397876 586880 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 66208 397874 66528 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2956 380476 -2356 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 81568 380476 81888 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586280 380476 586880 380478
rect -2956 380454 586880 380476
rect -2956 380218 -2774 380454
rect -2538 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 81610 380454
rect 81846 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586462 380454
rect 586698 380218 586880 380454
rect -2956 380134 586880 380218
rect -2956 379898 -2774 380134
rect -2538 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 81610 380134
rect 81846 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586462 380134
rect 586698 379898 586880 380134
rect -2956 379876 586880 379898
rect -2956 379874 -2356 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 81568 379874 81888 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586280 379874 586880 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 66208 362476 66528 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2956 362454 586880 362476
rect -2956 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 66250 362454
rect 66486 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586880 362454
rect -2956 362134 586880 362218
rect -2956 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 66250 362134
rect 66486 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586880 362134
rect -2956 361876 586880 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 66208 361874 66528 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2956 344476 -2356 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 81568 344476 81888 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586280 344476 586880 344478
rect -2956 344454 586880 344476
rect -2956 344218 -2774 344454
rect -2538 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 81610 344454
rect 81846 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586462 344454
rect 586698 344218 586880 344454
rect -2956 344134 586880 344218
rect -2956 343898 -2774 344134
rect -2538 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 81610 344134
rect 81846 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586462 344134
rect 586698 343898 586880 344134
rect -2956 343876 586880 343898
rect -2956 343874 -2356 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 81568 343874 81888 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586280 343874 586880 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 66208 326476 66528 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2956 326454 586880 326476
rect -2956 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 66250 326454
rect 66486 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586880 326454
rect -2956 326134 586880 326218
rect -2956 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 66250 326134
rect 66486 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586880 326134
rect -2956 325876 586880 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 66208 325874 66528 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2956 308476 -2356 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 81568 308476 81888 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586280 308476 586880 308478
rect -2956 308454 586880 308476
rect -2956 308218 -2774 308454
rect -2538 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 81610 308454
rect 81846 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586462 308454
rect 586698 308218 586880 308454
rect -2956 308134 586880 308218
rect -2956 307898 -2774 308134
rect -2538 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 81610 308134
rect 81846 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586462 308134
rect 586698 307898 586880 308134
rect -2956 307876 586880 307898
rect -2956 307874 -2356 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 81568 307874 81888 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586280 307874 586880 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 66208 290476 66528 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2956 290454 586880 290476
rect -2956 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 66250 290454
rect 66486 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586880 290454
rect -2956 290134 586880 290218
rect -2956 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 66250 290134
rect 66486 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586880 290134
rect -2956 289876 586880 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 66208 289874 66528 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2956 272476 -2356 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 81568 272476 81888 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586280 272476 586880 272478
rect -2956 272454 586880 272476
rect -2956 272218 -2774 272454
rect -2538 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 81610 272454
rect 81846 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586462 272454
rect 586698 272218 586880 272454
rect -2956 272134 586880 272218
rect -2956 271898 -2774 272134
rect -2538 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 81610 272134
rect 81846 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586462 272134
rect 586698 271898 586880 272134
rect -2956 271876 586880 271898
rect -2956 271874 -2356 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 81568 271874 81888 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586280 271874 586880 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 66208 254476 66528 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2956 254454 586880 254476
rect -2956 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 66250 254454
rect 66486 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586880 254454
rect -2956 254134 586880 254218
rect -2956 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 66250 254134
rect 66486 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586880 254134
rect -2956 253876 586880 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 66208 253874 66528 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -2956 236476 -2356 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 81568 236476 81888 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586280 236476 586880 236478
rect -2956 236454 586880 236476
rect -2956 236218 -2774 236454
rect -2538 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 81610 236454
rect 81846 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586462 236454
rect 586698 236218 586880 236454
rect -2956 236134 586880 236218
rect -2956 235898 -2774 236134
rect -2538 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 81610 236134
rect 81846 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586462 236134
rect 586698 235898 586880 236134
rect -2956 235876 586880 235898
rect -2956 235874 -2356 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 81568 235874 81888 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586280 235874 586880 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 66208 218476 66528 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2956 218454 586880 218476
rect -2956 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 66250 218454
rect 66486 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586880 218454
rect -2956 218134 586880 218218
rect -2956 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 66250 218134
rect 66486 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586880 218134
rect -2956 217876 586880 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 66208 217874 66528 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2956 200476 -2356 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 81568 200476 81888 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586280 200476 586880 200478
rect -2956 200454 586880 200476
rect -2956 200218 -2774 200454
rect -2538 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 81610 200454
rect 81846 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586462 200454
rect 586698 200218 586880 200454
rect -2956 200134 586880 200218
rect -2956 199898 -2774 200134
rect -2538 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 81610 200134
rect 81846 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586462 200134
rect 586698 199898 586880 200134
rect -2956 199876 586880 199898
rect -2956 199874 -2356 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 81568 199874 81888 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586280 199874 586880 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 66208 182476 66528 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2956 182454 586880 182476
rect -2956 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 66250 182454
rect 66486 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586880 182454
rect -2956 182134 586880 182218
rect -2956 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 66250 182134
rect 66486 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586880 182134
rect -2956 181876 586880 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 66208 181874 66528 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2956 164476 -2356 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 81568 164476 81888 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586280 164476 586880 164478
rect -2956 164454 586880 164476
rect -2956 164218 -2774 164454
rect -2538 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 81610 164454
rect 81846 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586462 164454
rect 586698 164218 586880 164454
rect -2956 164134 586880 164218
rect -2956 163898 -2774 164134
rect -2538 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 81610 164134
rect 81846 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586462 164134
rect 586698 163898 586880 164134
rect -2956 163876 586880 163898
rect -2956 163874 -2356 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 81568 163874 81888 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586280 163874 586880 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 66208 146476 66528 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2956 146454 586880 146476
rect -2956 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 66250 146454
rect 66486 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586880 146454
rect -2956 146134 586880 146218
rect -2956 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 66250 146134
rect 66486 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586880 146134
rect -2956 145876 586880 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 66208 145874 66528 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2956 128476 -2356 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 81568 128476 81888 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586280 128476 586880 128478
rect -2956 128454 586880 128476
rect -2956 128218 -2774 128454
rect -2538 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 81610 128454
rect 81846 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586462 128454
rect 586698 128218 586880 128454
rect -2956 128134 586880 128218
rect -2956 127898 -2774 128134
rect -2538 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 81610 128134
rect 81846 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586462 128134
rect 586698 127898 586880 128134
rect -2956 127876 586880 127898
rect -2956 127874 -2356 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 81568 127874 81888 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586280 127874 586880 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 66208 110476 66528 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2956 110454 586880 110476
rect -2956 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 66250 110454
rect 66486 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586880 110454
rect -2956 110134 586880 110218
rect -2956 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 66250 110134
rect 66486 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586880 110134
rect -2956 109876 586880 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 66208 109874 66528 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2956 92476 -2356 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 81568 92476 81888 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586280 92476 586880 92478
rect -2956 92454 586880 92476
rect -2956 92218 -2774 92454
rect -2538 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 81610 92454
rect 81846 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586462 92454
rect 586698 92218 586880 92454
rect -2956 92134 586880 92218
rect -2956 91898 -2774 92134
rect -2538 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 81610 92134
rect 81846 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586462 92134
rect 586698 91898 586880 92134
rect -2956 91876 586880 91898
rect -2956 91874 -2356 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 81568 91874 81888 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586280 91874 586880 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 66208 74476 66528 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2956 74454 586880 74476
rect -2956 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 66250 74454
rect 66486 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586880 74454
rect -2956 74134 586880 74218
rect -2956 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 66250 74134
rect 66486 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586880 74134
rect -2956 73876 586880 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 66208 73874 66528 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2956 56476 -2356 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 81568 56476 81888 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586280 56476 586880 56478
rect -2956 56454 586880 56476
rect -2956 56218 -2774 56454
rect -2538 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 81610 56454
rect 81846 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586462 56454
rect 586698 56218 586880 56454
rect -2956 56134 586880 56218
rect -2956 55898 -2774 56134
rect -2538 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 81610 56134
rect 81846 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586462 56134
rect 586698 55898 586880 56134
rect -2956 55876 586880 55898
rect -2956 55874 -2356 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 81568 55874 81888 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586280 55874 586880 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2956 38454 586880 38476
rect -2956 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586880 38454
rect -2956 38134 586880 38218
rect -2956 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586880 38134
rect -2956 37876 586880 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2956 20476 -2356 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586280 20476 586880 20478
rect -2956 20454 586880 20476
rect -2956 20218 -2774 20454
rect -2538 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586462 20454
rect 586698 20218 586880 20454
rect -2956 20134 586880 20218
rect -2956 19898 -2774 20134
rect -2538 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586462 20134
rect 586698 19898 586880 20134
rect -2956 19876 586880 19898
rect -2956 19874 -2356 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586280 19874 586880 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2956 2454 586880 2476
rect -2956 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586880 2454
rect -2956 2134 586880 2218
rect -2956 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586880 2134
rect -2956 1876 586880 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2956 -1284 -2356 -1282
rect 18804 -1284 19404 -1282
rect 54804 -1284 55404 -1282
rect 90804 -1284 91404 -1282
rect 126804 -1284 127404 -1282
rect 162804 -1284 163404 -1282
rect 198804 -1284 199404 -1282
rect 234804 -1284 235404 -1282
rect 270804 -1284 271404 -1282
rect 306804 -1284 307404 -1282
rect 342804 -1284 343404 -1282
rect 378804 -1284 379404 -1282
rect 414804 -1284 415404 -1282
rect 450804 -1284 451404 -1282
rect 486804 -1284 487404 -1282
rect 522804 -1284 523404 -1282
rect 558804 -1284 559404 -1282
rect 586280 -1284 586880 -1282
rect -2956 -1306 586880 -1284
rect -2956 -1542 -2774 -1306
rect -2538 -1542 18986 -1306
rect 19222 -1542 54986 -1306
rect 55222 -1542 90986 -1306
rect 91222 -1542 126986 -1306
rect 127222 -1542 162986 -1306
rect 163222 -1542 198986 -1306
rect 199222 -1542 234986 -1306
rect 235222 -1542 270986 -1306
rect 271222 -1542 306986 -1306
rect 307222 -1542 342986 -1306
rect 343222 -1542 378986 -1306
rect 379222 -1542 414986 -1306
rect 415222 -1542 450986 -1306
rect 451222 -1542 486986 -1306
rect 487222 -1542 522986 -1306
rect 523222 -1542 558986 -1306
rect 559222 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect -2956 -1626 586880 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 18986 -1626
rect 19222 -1862 54986 -1626
rect 55222 -1862 90986 -1626
rect 91222 -1862 126986 -1626
rect 127222 -1862 162986 -1626
rect 163222 -1862 198986 -1626
rect 199222 -1862 234986 -1626
rect 235222 -1862 270986 -1626
rect 271222 -1862 306986 -1626
rect 307222 -1862 342986 -1626
rect 343222 -1862 378986 -1626
rect 379222 -1862 414986 -1626
rect 415222 -1862 450986 -1626
rect 451222 -1862 486986 -1626
rect 487222 -1862 522986 -1626
rect 523222 -1862 558986 -1626
rect 559222 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect -2956 -1884 586880 -1862
rect -2956 -1886 -2356 -1884
rect 18804 -1886 19404 -1884
rect 54804 -1886 55404 -1884
rect 90804 -1886 91404 -1884
rect 126804 -1886 127404 -1884
rect 162804 -1886 163404 -1884
rect 198804 -1886 199404 -1884
rect 234804 -1886 235404 -1884
rect 270804 -1886 271404 -1884
rect 306804 -1886 307404 -1884
rect 342804 -1886 343404 -1884
rect 378804 -1886 379404 -1884
rect 414804 -1886 415404 -1884
rect 450804 -1886 451404 -1884
rect 486804 -1886 487404 -1884
rect 522804 -1886 523404 -1884
rect 558804 -1886 559404 -1884
rect 586280 -1886 586880 -1884
use ghazi_top_dffram_csv  mprj
timestamp 1608285900
transform 1 0 62000 0 1 52000
box 0 0 460000 600000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2956 -1884 586880 -1284 8 vssd1
port 637 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
