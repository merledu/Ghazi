VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ghazi_top_dffram_csv
  CLASS BLOCK ;
  FOREIGN ghazi_top_dffram_csv ;
  ORIGIN 0.000 0.000 ;
  SIZE 2300.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 33.360 2300.000 33.960 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2033.240 2300.000 2033.840 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2233.160 2300.000 2233.760 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2433.080 2300.000 2433.680 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2633.000 2300.000 2633.600 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2832.920 2300.000 2833.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.850 2996.000 2257.130 3000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2001.550 2996.000 2001.830 3000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1745.790 2996.000 1746.070 3000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1490.490 2996.000 1490.770 3000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.730 2996.000 1235.010 3000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 233.280 2300.000 233.880 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.430 2996.000 979.710 3000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.670 2996.000 723.950 3000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.910 2996.000 468.190 3000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.610 2996.000 212.890 3000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2963.480 4.000 2964.080 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2749.280 4.000 2749.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2535.080 4.000 2535.680 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2320.880 4.000 2321.480 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2106.680 4.000 2107.280 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1892.480 4.000 1893.080 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 433.200 2300.000 433.800 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1678.280 4.000 1678.880 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1463.400 4.000 1464.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1249.200 4.000 1249.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.000 4.000 1035.600 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 633.120 2300.000 633.720 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 833.040 2300.000 833.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1032.960 2300.000 1033.560 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1232.880 2300.000 1233.480 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1432.800 2300.000 1433.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1633.400 2300.000 1634.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1833.320 2300.000 1833.920 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 166.640 2300.000 167.240 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2166.520 2300.000 2167.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2366.440 2300.000 2367.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2566.360 2300.000 2566.960 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2766.280 2300.000 2766.880 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2966.200 2300.000 2966.800 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2086.650 2996.000 2086.930 3000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1830.890 2996.000 1831.170 3000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1575.590 2996.000 1575.870 3000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1319.830 2996.000 1320.110 3000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1064.530 2996.000 1064.810 3000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 366.560 2300.000 367.160 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 808.770 2996.000 809.050 3000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 553.470 2996.000 553.750 3000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 297.710 2996.000 297.990 3000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 2996.000 42.690 3000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2820.680 4.000 2821.280 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2606.480 4.000 2607.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2392.280 4.000 2392.880 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2178.080 4.000 2178.680 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1963.880 4.000 1964.480 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1749.680 4.000 1750.280 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 566.480 2300.000 567.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1535.480 4.000 1536.080 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1320.600 4.000 1321.200 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1106.400 4.000 1107.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 766.400 2300.000 767.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 966.320 2300.000 966.920 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1166.240 2300.000 1166.840 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1366.160 2300.000 1366.760 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1566.760 2300.000 1567.360 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1766.680 2300.000 1767.280 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1966.600 2300.000 1967.200 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 100.000 2300.000 100.600 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2099.880 2300.000 2100.480 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2299.800 2300.000 2300.400 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2499.720 2300.000 2500.320 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2699.640 2300.000 2700.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 2899.560 2300.000 2900.160 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2171.750 2996.000 2172.030 3000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1916.450 2996.000 1916.730 3000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1660.690 2996.000 1660.970 3000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1404.930 2996.000 1405.210 3000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1149.630 2996.000 1149.910 3000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 299.920 2300.000 300.520 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.870 2996.000 894.150 3000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.570 2996.000 638.850 3000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.810 2996.000 383.090 3000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 2996.000 127.790 3000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2892.080 4.000 2892.680 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2677.880 4.000 2678.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2463.680 4.000 2464.280 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2249.480 4.000 2250.080 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2035.280 4.000 2035.880 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1821.080 4.000 1821.680 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 499.840 2300.000 500.440 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1606.880 4.000 1607.480 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.000 4.000 1392.600 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.800 4.000 1178.400 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 699.760 2300.000 700.360 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 899.680 2300.000 900.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1099.600 2300.000 1100.200 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1299.520 2300.000 1300.120 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1499.440 2300.000 1500.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1700.040 2300.000 1700.640 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2296.000 1899.960 2300.000 1900.560 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1801.910 0.000 1802.190 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1819.850 0.000 1820.130 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1837.790 0.000 1838.070 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1855.730 0.000 1856.010 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1873.670 0.000 1873.950 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1891.610 0.000 1891.890 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1927.030 0.000 1927.310 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1944.970 0.000 1945.250 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1962.910 0.000 1963.190 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1980.850 0.000 1981.130 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1998.790 0.000 1999.070 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2016.730 0.000 2017.010 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2034.670 0.000 2034.950 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2052.150 0.000 2052.430 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2070.090 0.000 2070.370 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2088.030 0.000 2088.310 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2123.910 0.000 2124.190 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2141.850 0.000 2142.130 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2159.790 0.000 2160.070 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2177.270 0.000 2177.550 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2195.210 0.000 2195.490 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2213.150 0.000 2213.430 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2231.090 0.000 2231.370 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2249.030 0.000 2249.310 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2266.970 0.000 2267.250 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2284.910 0.000 2285.190 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.530 0.000 765.810 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 818.890 0.000 819.170 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 836.830 0.000 837.110 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 890.650 0.000 890.930 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.890 0.000 980.170 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 997.830 0.000 998.110 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.770 0.000 1016.050 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1105.010 0.000 1105.290 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.950 0.000 1123.230 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1140.890 0.000 1141.170 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1158.370 0.000 1158.650 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1176.310 0.000 1176.590 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1212.190 0.000 1212.470 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1230.130 0.000 1230.410 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1248.070 0.000 1248.350 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1283.490 0.000 1283.770 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1319.370 0.000 1319.650 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1337.310 0.000 1337.590 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1355.250 0.000 1355.530 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1373.190 0.000 1373.470 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1408.610 0.000 1408.890 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1426.550 0.000 1426.830 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.490 0.000 1444.770 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1462.430 0.000 1462.710 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1480.370 0.000 1480.650 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.310 0.000 1498.590 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1516.250 0.000 1516.530 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1551.670 0.000 1551.950 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1569.610 0.000 1569.890 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1587.550 0.000 1587.830 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1605.490 0.000 1605.770 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1623.430 0.000 1623.710 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1641.370 0.000 1641.650 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1659.310 0.000 1659.590 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1676.790 0.000 1677.070 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1694.730 0.000 1695.010 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1712.670 0.000 1712.950 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1730.610 0.000 1730.890 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1748.550 0.000 1748.830 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1766.490 0.000 1766.770 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1784.430 0.000 1784.710 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1825.830 0.000 1826.110 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1843.770 0.000 1844.050 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1861.710 0.000 1861.990 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1879.650 0.000 1879.930 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1897.590 0.000 1897.870 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1915.530 0.000 1915.810 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1933.010 0.000 1933.290 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1950.950 0.000 1951.230 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1968.890 0.000 1969.170 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1986.830 0.000 1987.110 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2004.770 0.000 2005.050 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2022.710 0.000 2022.990 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2040.650 0.000 2040.930 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2058.130 0.000 2058.410 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2076.070 0.000 2076.350 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2094.010 0.000 2094.290 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2111.950 0.000 2112.230 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2129.890 0.000 2130.170 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2147.830 0.000 2148.110 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2165.770 0.000 2166.050 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2183.250 0.000 2183.530 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2201.190 0.000 2201.470 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2219.130 0.000 2219.410 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2237.070 0.000 2237.350 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2255.010 0.000 2255.290 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2272.950 0.000 2273.230 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2290.890 0.000 2291.170 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.930 0.000 807.210 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 914.110 0.000 914.390 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1003.810 0.000 1004.090 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1021.750 0.000 1022.030 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1039.230 0.000 1039.510 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1057.170 0.000 1057.450 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1146.870 0.000 1147.150 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1182.290 0.000 1182.570 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1200.230 0.000 1200.510 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1236.110 0.000 1236.390 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1254.050 0.000 1254.330 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1289.470 0.000 1289.750 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1343.290 0.000 1343.570 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1361.230 0.000 1361.510 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1397.110 0.000 1397.390 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1414.590 0.000 1414.870 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1432.530 0.000 1432.810 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1450.470 0.000 1450.750 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1486.350 0.000 1486.630 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1504.290 0.000 1504.570 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1522.230 0.000 1522.510 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1539.710 0.000 1539.990 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1557.650 0.000 1557.930 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1575.590 0.000 1575.870 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1593.530 0.000 1593.810 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1629.410 0.000 1629.690 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1647.350 0.000 1647.630 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1664.830 0.000 1665.110 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1682.770 0.000 1683.050 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1700.710 0.000 1700.990 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1718.650 0.000 1718.930 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1736.590 0.000 1736.870 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1754.530 0.000 1754.810 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1772.470 0.000 1772.750 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1790.410 0.000 1790.690 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1813.870 0.000 1814.150 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1831.810 0.000 1832.090 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1849.750 0.000 1850.030 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1885.630 0.000 1885.910 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1921.050 0.000 1921.330 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1938.990 0.000 1939.270 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1956.930 0.000 1957.210 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1974.870 0.000 1975.150 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1992.810 0.000 1993.090 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2010.750 0.000 2011.030 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2028.690 0.000 2028.970 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2046.630 0.000 2046.910 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2082.050 0.000 2082.330 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2099.990 0.000 2100.270 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2117.930 0.000 2118.210 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2135.870 0.000 2136.150 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2153.810 0.000 2154.090 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2171.750 0.000 2172.030 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2189.230 0.000 2189.510 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2207.170 0.000 2207.450 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2225.110 0.000 2225.390 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2243.050 0.000 2243.330 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2260.990 0.000 2261.270 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2278.930 0.000 2279.210 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2296.870 0.000 2297.150 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.970 0.000 795.250 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.910 0.000 813.190 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.670 0.000 884.950 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.150 0.000 902.430 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.090 0.000 920.370 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 955.970 0.000 956.250 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.910 0.000 974.190 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.150 0.000 1063.430 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1081.090 0.000 1081.370 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1099.030 0.000 1099.310 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.970 0.000 1117.250 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1170.330 0.000 1170.610 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1206.210 0.000 1206.490 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1242.090 0.000 1242.370 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1260.030 0.000 1260.310 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.970 0.000 1278.250 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1295.450 0.000 1295.730 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1313.390 0.000 1313.670 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1331.330 0.000 1331.610 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1367.210 0.000 1367.490 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1420.570 0.000 1420.850 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1438.510 0.000 1438.790 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1456.450 0.000 1456.730 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1474.390 0.000 1474.670 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1528.210 0.000 1528.490 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1545.690 0.000 1545.970 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1581.570 0.000 1581.850 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1599.510 0.000 1599.790 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1617.450 0.000 1617.730 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1635.390 0.000 1635.670 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1653.330 0.000 1653.610 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1670.810 0.000 1671.090 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1688.750 0.000 1689.030 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1706.690 0.000 1706.970 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1724.630 0.000 1724.910 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1742.570 0.000 1742.850 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1760.510 0.000 1760.790 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1778.450 0.000 1778.730 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1795.930 0.000 1796.210 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wb_rst_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2294.480 2986.645 ;
      LAYER met1 ;
        RECT 5.520 9.220 2294.480 2995.700 ;
      LAYER met2 ;
        RECT 2.850 2995.720 42.130 2996.000 ;
        RECT 42.970 2995.720 127.230 2996.000 ;
        RECT 128.070 2995.720 212.330 2996.000 ;
        RECT 213.170 2995.720 297.430 2996.000 ;
        RECT 298.270 2995.720 382.530 2996.000 ;
        RECT 383.370 2995.720 467.630 2996.000 ;
        RECT 468.470 2995.720 553.190 2996.000 ;
        RECT 554.030 2995.720 638.290 2996.000 ;
        RECT 639.130 2995.720 723.390 2996.000 ;
        RECT 724.230 2995.720 808.490 2996.000 ;
        RECT 809.330 2995.720 893.590 2996.000 ;
        RECT 894.430 2995.720 979.150 2996.000 ;
        RECT 979.990 2995.720 1064.250 2996.000 ;
        RECT 1065.090 2995.720 1149.350 2996.000 ;
        RECT 1150.190 2995.720 1234.450 2996.000 ;
        RECT 1235.290 2995.720 1319.550 2996.000 ;
        RECT 1320.390 2995.720 1404.650 2996.000 ;
        RECT 1405.490 2995.720 1490.210 2996.000 ;
        RECT 1491.050 2995.720 1575.310 2996.000 ;
        RECT 1576.150 2995.720 1660.410 2996.000 ;
        RECT 1661.250 2995.720 1745.510 2996.000 ;
        RECT 1746.350 2995.720 1830.610 2996.000 ;
        RECT 1831.450 2995.720 1916.170 2996.000 ;
        RECT 1917.010 2995.720 2001.270 2996.000 ;
        RECT 2002.110 2995.720 2086.370 2996.000 ;
        RECT 2087.210 2995.720 2171.470 2996.000 ;
        RECT 2172.310 2995.720 2256.570 2996.000 ;
        RECT 2257.410 2995.720 2291.160 2996.000 ;
        RECT 2.850 4.280 2291.160 2995.720 ;
        RECT 3.410 4.000 8.090 4.280 ;
        RECT 8.930 4.000 14.070 4.280 ;
        RECT 14.910 4.000 20.050 4.280 ;
        RECT 20.890 4.000 26.030 4.280 ;
        RECT 26.870 4.000 32.010 4.280 ;
        RECT 32.850 4.000 37.990 4.280 ;
        RECT 38.830 4.000 43.970 4.280 ;
        RECT 44.810 4.000 49.950 4.280 ;
        RECT 50.790 4.000 55.930 4.280 ;
        RECT 56.770 4.000 61.910 4.280 ;
        RECT 62.750 4.000 67.890 4.280 ;
        RECT 68.730 4.000 73.870 4.280 ;
        RECT 74.710 4.000 79.850 4.280 ;
        RECT 80.690 4.000 85.830 4.280 ;
        RECT 86.670 4.000 91.810 4.280 ;
        RECT 92.650 4.000 97.790 4.280 ;
        RECT 98.630 4.000 103.770 4.280 ;
        RECT 104.610 4.000 109.750 4.280 ;
        RECT 110.590 4.000 115.730 4.280 ;
        RECT 116.570 4.000 121.710 4.280 ;
        RECT 122.550 4.000 127.690 4.280 ;
        RECT 128.530 4.000 133.210 4.280 ;
        RECT 134.050 4.000 139.190 4.280 ;
        RECT 140.030 4.000 145.170 4.280 ;
        RECT 146.010 4.000 151.150 4.280 ;
        RECT 151.990 4.000 157.130 4.280 ;
        RECT 157.970 4.000 163.110 4.280 ;
        RECT 163.950 4.000 169.090 4.280 ;
        RECT 169.930 4.000 175.070 4.280 ;
        RECT 175.910 4.000 181.050 4.280 ;
        RECT 181.890 4.000 187.030 4.280 ;
        RECT 187.870 4.000 193.010 4.280 ;
        RECT 193.850 4.000 198.990 4.280 ;
        RECT 199.830 4.000 204.970 4.280 ;
        RECT 205.810 4.000 210.950 4.280 ;
        RECT 211.790 4.000 216.930 4.280 ;
        RECT 217.770 4.000 222.910 4.280 ;
        RECT 223.750 4.000 228.890 4.280 ;
        RECT 229.730 4.000 234.870 4.280 ;
        RECT 235.710 4.000 240.850 4.280 ;
        RECT 241.690 4.000 246.830 4.280 ;
        RECT 247.670 4.000 252.810 4.280 ;
        RECT 253.650 4.000 258.330 4.280 ;
        RECT 259.170 4.000 264.310 4.280 ;
        RECT 265.150 4.000 270.290 4.280 ;
        RECT 271.130 4.000 276.270 4.280 ;
        RECT 277.110 4.000 282.250 4.280 ;
        RECT 283.090 4.000 288.230 4.280 ;
        RECT 289.070 4.000 294.210 4.280 ;
        RECT 295.050 4.000 300.190 4.280 ;
        RECT 301.030 4.000 306.170 4.280 ;
        RECT 307.010 4.000 312.150 4.280 ;
        RECT 312.990 4.000 318.130 4.280 ;
        RECT 318.970 4.000 324.110 4.280 ;
        RECT 324.950 4.000 330.090 4.280 ;
        RECT 330.930 4.000 336.070 4.280 ;
        RECT 336.910 4.000 342.050 4.280 ;
        RECT 342.890 4.000 348.030 4.280 ;
        RECT 348.870 4.000 354.010 4.280 ;
        RECT 354.850 4.000 359.990 4.280 ;
        RECT 360.830 4.000 365.970 4.280 ;
        RECT 366.810 4.000 371.950 4.280 ;
        RECT 372.790 4.000 377.930 4.280 ;
        RECT 378.770 4.000 383.910 4.280 ;
        RECT 384.750 4.000 389.430 4.280 ;
        RECT 390.270 4.000 395.410 4.280 ;
        RECT 396.250 4.000 401.390 4.280 ;
        RECT 402.230 4.000 407.370 4.280 ;
        RECT 408.210 4.000 413.350 4.280 ;
        RECT 414.190 4.000 419.330 4.280 ;
        RECT 420.170 4.000 425.310 4.280 ;
        RECT 426.150 4.000 431.290 4.280 ;
        RECT 432.130 4.000 437.270 4.280 ;
        RECT 438.110 4.000 443.250 4.280 ;
        RECT 444.090 4.000 449.230 4.280 ;
        RECT 450.070 4.000 455.210 4.280 ;
        RECT 456.050 4.000 461.190 4.280 ;
        RECT 462.030 4.000 467.170 4.280 ;
        RECT 468.010 4.000 473.150 4.280 ;
        RECT 473.990 4.000 479.130 4.280 ;
        RECT 479.970 4.000 485.110 4.280 ;
        RECT 485.950 4.000 491.090 4.280 ;
        RECT 491.930 4.000 497.070 4.280 ;
        RECT 497.910 4.000 503.050 4.280 ;
        RECT 503.890 4.000 509.030 4.280 ;
        RECT 509.870 4.000 514.550 4.280 ;
        RECT 515.390 4.000 520.530 4.280 ;
        RECT 521.370 4.000 526.510 4.280 ;
        RECT 527.350 4.000 532.490 4.280 ;
        RECT 533.330 4.000 538.470 4.280 ;
        RECT 539.310 4.000 544.450 4.280 ;
        RECT 545.290 4.000 550.430 4.280 ;
        RECT 551.270 4.000 556.410 4.280 ;
        RECT 557.250 4.000 562.390 4.280 ;
        RECT 563.230 4.000 568.370 4.280 ;
        RECT 569.210 4.000 574.350 4.280 ;
        RECT 575.190 4.000 580.330 4.280 ;
        RECT 581.170 4.000 586.310 4.280 ;
        RECT 587.150 4.000 592.290 4.280 ;
        RECT 593.130 4.000 598.270 4.280 ;
        RECT 599.110 4.000 604.250 4.280 ;
        RECT 605.090 4.000 610.230 4.280 ;
        RECT 611.070 4.000 616.210 4.280 ;
        RECT 617.050 4.000 622.190 4.280 ;
        RECT 623.030 4.000 628.170 4.280 ;
        RECT 629.010 4.000 634.150 4.280 ;
        RECT 634.990 4.000 640.130 4.280 ;
        RECT 640.970 4.000 645.650 4.280 ;
        RECT 646.490 4.000 651.630 4.280 ;
        RECT 652.470 4.000 657.610 4.280 ;
        RECT 658.450 4.000 663.590 4.280 ;
        RECT 664.430 4.000 669.570 4.280 ;
        RECT 670.410 4.000 675.550 4.280 ;
        RECT 676.390 4.000 681.530 4.280 ;
        RECT 682.370 4.000 687.510 4.280 ;
        RECT 688.350 4.000 693.490 4.280 ;
        RECT 694.330 4.000 699.470 4.280 ;
        RECT 700.310 4.000 705.450 4.280 ;
        RECT 706.290 4.000 711.430 4.280 ;
        RECT 712.270 4.000 717.410 4.280 ;
        RECT 718.250 4.000 723.390 4.280 ;
        RECT 724.230 4.000 729.370 4.280 ;
        RECT 730.210 4.000 735.350 4.280 ;
        RECT 736.190 4.000 741.330 4.280 ;
        RECT 742.170 4.000 747.310 4.280 ;
        RECT 748.150 4.000 753.290 4.280 ;
        RECT 754.130 4.000 759.270 4.280 ;
        RECT 760.110 4.000 765.250 4.280 ;
        RECT 766.090 4.000 770.770 4.280 ;
        RECT 771.610 4.000 776.750 4.280 ;
        RECT 777.590 4.000 782.730 4.280 ;
        RECT 783.570 4.000 788.710 4.280 ;
        RECT 789.550 4.000 794.690 4.280 ;
        RECT 795.530 4.000 800.670 4.280 ;
        RECT 801.510 4.000 806.650 4.280 ;
        RECT 807.490 4.000 812.630 4.280 ;
        RECT 813.470 4.000 818.610 4.280 ;
        RECT 819.450 4.000 824.590 4.280 ;
        RECT 825.430 4.000 830.570 4.280 ;
        RECT 831.410 4.000 836.550 4.280 ;
        RECT 837.390 4.000 842.530 4.280 ;
        RECT 843.370 4.000 848.510 4.280 ;
        RECT 849.350 4.000 854.490 4.280 ;
        RECT 855.330 4.000 860.470 4.280 ;
        RECT 861.310 4.000 866.450 4.280 ;
        RECT 867.290 4.000 872.430 4.280 ;
        RECT 873.270 4.000 878.410 4.280 ;
        RECT 879.250 4.000 884.390 4.280 ;
        RECT 885.230 4.000 890.370 4.280 ;
        RECT 891.210 4.000 896.350 4.280 ;
        RECT 897.190 4.000 901.870 4.280 ;
        RECT 902.710 4.000 907.850 4.280 ;
        RECT 908.690 4.000 913.830 4.280 ;
        RECT 914.670 4.000 919.810 4.280 ;
        RECT 920.650 4.000 925.790 4.280 ;
        RECT 926.630 4.000 931.770 4.280 ;
        RECT 932.610 4.000 937.750 4.280 ;
        RECT 938.590 4.000 943.730 4.280 ;
        RECT 944.570 4.000 949.710 4.280 ;
        RECT 950.550 4.000 955.690 4.280 ;
        RECT 956.530 4.000 961.670 4.280 ;
        RECT 962.510 4.000 967.650 4.280 ;
        RECT 968.490 4.000 973.630 4.280 ;
        RECT 974.470 4.000 979.610 4.280 ;
        RECT 980.450 4.000 985.590 4.280 ;
        RECT 986.430 4.000 991.570 4.280 ;
        RECT 992.410 4.000 997.550 4.280 ;
        RECT 998.390 4.000 1003.530 4.280 ;
        RECT 1004.370 4.000 1009.510 4.280 ;
        RECT 1010.350 4.000 1015.490 4.280 ;
        RECT 1016.330 4.000 1021.470 4.280 ;
        RECT 1022.310 4.000 1026.990 4.280 ;
        RECT 1027.830 4.000 1032.970 4.280 ;
        RECT 1033.810 4.000 1038.950 4.280 ;
        RECT 1039.790 4.000 1044.930 4.280 ;
        RECT 1045.770 4.000 1050.910 4.280 ;
        RECT 1051.750 4.000 1056.890 4.280 ;
        RECT 1057.730 4.000 1062.870 4.280 ;
        RECT 1063.710 4.000 1068.850 4.280 ;
        RECT 1069.690 4.000 1074.830 4.280 ;
        RECT 1075.670 4.000 1080.810 4.280 ;
        RECT 1081.650 4.000 1086.790 4.280 ;
        RECT 1087.630 4.000 1092.770 4.280 ;
        RECT 1093.610 4.000 1098.750 4.280 ;
        RECT 1099.590 4.000 1104.730 4.280 ;
        RECT 1105.570 4.000 1110.710 4.280 ;
        RECT 1111.550 4.000 1116.690 4.280 ;
        RECT 1117.530 4.000 1122.670 4.280 ;
        RECT 1123.510 4.000 1128.650 4.280 ;
        RECT 1129.490 4.000 1134.630 4.280 ;
        RECT 1135.470 4.000 1140.610 4.280 ;
        RECT 1141.450 4.000 1146.590 4.280 ;
        RECT 1147.430 4.000 1152.570 4.280 ;
        RECT 1153.410 4.000 1158.090 4.280 ;
        RECT 1158.930 4.000 1164.070 4.280 ;
        RECT 1164.910 4.000 1170.050 4.280 ;
        RECT 1170.890 4.000 1176.030 4.280 ;
        RECT 1176.870 4.000 1182.010 4.280 ;
        RECT 1182.850 4.000 1187.990 4.280 ;
        RECT 1188.830 4.000 1193.970 4.280 ;
        RECT 1194.810 4.000 1199.950 4.280 ;
        RECT 1200.790 4.000 1205.930 4.280 ;
        RECT 1206.770 4.000 1211.910 4.280 ;
        RECT 1212.750 4.000 1217.890 4.280 ;
        RECT 1218.730 4.000 1223.870 4.280 ;
        RECT 1224.710 4.000 1229.850 4.280 ;
        RECT 1230.690 4.000 1235.830 4.280 ;
        RECT 1236.670 4.000 1241.810 4.280 ;
        RECT 1242.650 4.000 1247.790 4.280 ;
        RECT 1248.630 4.000 1253.770 4.280 ;
        RECT 1254.610 4.000 1259.750 4.280 ;
        RECT 1260.590 4.000 1265.730 4.280 ;
        RECT 1266.570 4.000 1271.710 4.280 ;
        RECT 1272.550 4.000 1277.690 4.280 ;
        RECT 1278.530 4.000 1283.210 4.280 ;
        RECT 1284.050 4.000 1289.190 4.280 ;
        RECT 1290.030 4.000 1295.170 4.280 ;
        RECT 1296.010 4.000 1301.150 4.280 ;
        RECT 1301.990 4.000 1307.130 4.280 ;
        RECT 1307.970 4.000 1313.110 4.280 ;
        RECT 1313.950 4.000 1319.090 4.280 ;
        RECT 1319.930 4.000 1325.070 4.280 ;
        RECT 1325.910 4.000 1331.050 4.280 ;
        RECT 1331.890 4.000 1337.030 4.280 ;
        RECT 1337.870 4.000 1343.010 4.280 ;
        RECT 1343.850 4.000 1348.990 4.280 ;
        RECT 1349.830 4.000 1354.970 4.280 ;
        RECT 1355.810 4.000 1360.950 4.280 ;
        RECT 1361.790 4.000 1366.930 4.280 ;
        RECT 1367.770 4.000 1372.910 4.280 ;
        RECT 1373.750 4.000 1378.890 4.280 ;
        RECT 1379.730 4.000 1384.870 4.280 ;
        RECT 1385.710 4.000 1390.850 4.280 ;
        RECT 1391.690 4.000 1396.830 4.280 ;
        RECT 1397.670 4.000 1402.810 4.280 ;
        RECT 1403.650 4.000 1408.330 4.280 ;
        RECT 1409.170 4.000 1414.310 4.280 ;
        RECT 1415.150 4.000 1420.290 4.280 ;
        RECT 1421.130 4.000 1426.270 4.280 ;
        RECT 1427.110 4.000 1432.250 4.280 ;
        RECT 1433.090 4.000 1438.230 4.280 ;
        RECT 1439.070 4.000 1444.210 4.280 ;
        RECT 1445.050 4.000 1450.190 4.280 ;
        RECT 1451.030 4.000 1456.170 4.280 ;
        RECT 1457.010 4.000 1462.150 4.280 ;
        RECT 1462.990 4.000 1468.130 4.280 ;
        RECT 1468.970 4.000 1474.110 4.280 ;
        RECT 1474.950 4.000 1480.090 4.280 ;
        RECT 1480.930 4.000 1486.070 4.280 ;
        RECT 1486.910 4.000 1492.050 4.280 ;
        RECT 1492.890 4.000 1498.030 4.280 ;
        RECT 1498.870 4.000 1504.010 4.280 ;
        RECT 1504.850 4.000 1509.990 4.280 ;
        RECT 1510.830 4.000 1515.970 4.280 ;
        RECT 1516.810 4.000 1521.950 4.280 ;
        RECT 1522.790 4.000 1527.930 4.280 ;
        RECT 1528.770 4.000 1533.910 4.280 ;
        RECT 1534.750 4.000 1539.430 4.280 ;
        RECT 1540.270 4.000 1545.410 4.280 ;
        RECT 1546.250 4.000 1551.390 4.280 ;
        RECT 1552.230 4.000 1557.370 4.280 ;
        RECT 1558.210 4.000 1563.350 4.280 ;
        RECT 1564.190 4.000 1569.330 4.280 ;
        RECT 1570.170 4.000 1575.310 4.280 ;
        RECT 1576.150 4.000 1581.290 4.280 ;
        RECT 1582.130 4.000 1587.270 4.280 ;
        RECT 1588.110 4.000 1593.250 4.280 ;
        RECT 1594.090 4.000 1599.230 4.280 ;
        RECT 1600.070 4.000 1605.210 4.280 ;
        RECT 1606.050 4.000 1611.190 4.280 ;
        RECT 1612.030 4.000 1617.170 4.280 ;
        RECT 1618.010 4.000 1623.150 4.280 ;
        RECT 1623.990 4.000 1629.130 4.280 ;
        RECT 1629.970 4.000 1635.110 4.280 ;
        RECT 1635.950 4.000 1641.090 4.280 ;
        RECT 1641.930 4.000 1647.070 4.280 ;
        RECT 1647.910 4.000 1653.050 4.280 ;
        RECT 1653.890 4.000 1659.030 4.280 ;
        RECT 1659.870 4.000 1664.550 4.280 ;
        RECT 1665.390 4.000 1670.530 4.280 ;
        RECT 1671.370 4.000 1676.510 4.280 ;
        RECT 1677.350 4.000 1682.490 4.280 ;
        RECT 1683.330 4.000 1688.470 4.280 ;
        RECT 1689.310 4.000 1694.450 4.280 ;
        RECT 1695.290 4.000 1700.430 4.280 ;
        RECT 1701.270 4.000 1706.410 4.280 ;
        RECT 1707.250 4.000 1712.390 4.280 ;
        RECT 1713.230 4.000 1718.370 4.280 ;
        RECT 1719.210 4.000 1724.350 4.280 ;
        RECT 1725.190 4.000 1730.330 4.280 ;
        RECT 1731.170 4.000 1736.310 4.280 ;
        RECT 1737.150 4.000 1742.290 4.280 ;
        RECT 1743.130 4.000 1748.270 4.280 ;
        RECT 1749.110 4.000 1754.250 4.280 ;
        RECT 1755.090 4.000 1760.230 4.280 ;
        RECT 1761.070 4.000 1766.210 4.280 ;
        RECT 1767.050 4.000 1772.190 4.280 ;
        RECT 1773.030 4.000 1778.170 4.280 ;
        RECT 1779.010 4.000 1784.150 4.280 ;
        RECT 1784.990 4.000 1790.130 4.280 ;
        RECT 1790.970 4.000 1795.650 4.280 ;
        RECT 1796.490 4.000 1801.630 4.280 ;
        RECT 1802.470 4.000 1807.610 4.280 ;
        RECT 1808.450 4.000 1813.590 4.280 ;
        RECT 1814.430 4.000 1819.570 4.280 ;
        RECT 1820.410 4.000 1825.550 4.280 ;
        RECT 1826.390 4.000 1831.530 4.280 ;
        RECT 1832.370 4.000 1837.510 4.280 ;
        RECT 1838.350 4.000 1843.490 4.280 ;
        RECT 1844.330 4.000 1849.470 4.280 ;
        RECT 1850.310 4.000 1855.450 4.280 ;
        RECT 1856.290 4.000 1861.430 4.280 ;
        RECT 1862.270 4.000 1867.410 4.280 ;
        RECT 1868.250 4.000 1873.390 4.280 ;
        RECT 1874.230 4.000 1879.370 4.280 ;
        RECT 1880.210 4.000 1885.350 4.280 ;
        RECT 1886.190 4.000 1891.330 4.280 ;
        RECT 1892.170 4.000 1897.310 4.280 ;
        RECT 1898.150 4.000 1903.290 4.280 ;
        RECT 1904.130 4.000 1909.270 4.280 ;
        RECT 1910.110 4.000 1915.250 4.280 ;
        RECT 1916.090 4.000 1920.770 4.280 ;
        RECT 1921.610 4.000 1926.750 4.280 ;
        RECT 1927.590 4.000 1932.730 4.280 ;
        RECT 1933.570 4.000 1938.710 4.280 ;
        RECT 1939.550 4.000 1944.690 4.280 ;
        RECT 1945.530 4.000 1950.670 4.280 ;
        RECT 1951.510 4.000 1956.650 4.280 ;
        RECT 1957.490 4.000 1962.630 4.280 ;
        RECT 1963.470 4.000 1968.610 4.280 ;
        RECT 1969.450 4.000 1974.590 4.280 ;
        RECT 1975.430 4.000 1980.570 4.280 ;
        RECT 1981.410 4.000 1986.550 4.280 ;
        RECT 1987.390 4.000 1992.530 4.280 ;
        RECT 1993.370 4.000 1998.510 4.280 ;
        RECT 1999.350 4.000 2004.490 4.280 ;
        RECT 2005.330 4.000 2010.470 4.280 ;
        RECT 2011.310 4.000 2016.450 4.280 ;
        RECT 2017.290 4.000 2022.430 4.280 ;
        RECT 2023.270 4.000 2028.410 4.280 ;
        RECT 2029.250 4.000 2034.390 4.280 ;
        RECT 2035.230 4.000 2040.370 4.280 ;
        RECT 2041.210 4.000 2046.350 4.280 ;
        RECT 2047.190 4.000 2051.870 4.280 ;
        RECT 2052.710 4.000 2057.850 4.280 ;
        RECT 2058.690 4.000 2063.830 4.280 ;
        RECT 2064.670 4.000 2069.810 4.280 ;
        RECT 2070.650 4.000 2075.790 4.280 ;
        RECT 2076.630 4.000 2081.770 4.280 ;
        RECT 2082.610 4.000 2087.750 4.280 ;
        RECT 2088.590 4.000 2093.730 4.280 ;
        RECT 2094.570 4.000 2099.710 4.280 ;
        RECT 2100.550 4.000 2105.690 4.280 ;
        RECT 2106.530 4.000 2111.670 4.280 ;
        RECT 2112.510 4.000 2117.650 4.280 ;
        RECT 2118.490 4.000 2123.630 4.280 ;
        RECT 2124.470 4.000 2129.610 4.280 ;
        RECT 2130.450 4.000 2135.590 4.280 ;
        RECT 2136.430 4.000 2141.570 4.280 ;
        RECT 2142.410 4.000 2147.550 4.280 ;
        RECT 2148.390 4.000 2153.530 4.280 ;
        RECT 2154.370 4.000 2159.510 4.280 ;
        RECT 2160.350 4.000 2165.490 4.280 ;
        RECT 2166.330 4.000 2171.470 4.280 ;
        RECT 2172.310 4.000 2176.990 4.280 ;
        RECT 2177.830 4.000 2182.970 4.280 ;
        RECT 2183.810 4.000 2188.950 4.280 ;
        RECT 2189.790 4.000 2194.930 4.280 ;
        RECT 2195.770 4.000 2200.910 4.280 ;
        RECT 2201.750 4.000 2206.890 4.280 ;
        RECT 2207.730 4.000 2212.870 4.280 ;
        RECT 2213.710 4.000 2218.850 4.280 ;
        RECT 2219.690 4.000 2224.830 4.280 ;
        RECT 2225.670 4.000 2230.810 4.280 ;
        RECT 2231.650 4.000 2236.790 4.280 ;
        RECT 2237.630 4.000 2242.770 4.280 ;
        RECT 2243.610 4.000 2248.750 4.280 ;
        RECT 2249.590 4.000 2254.730 4.280 ;
        RECT 2255.570 4.000 2260.710 4.280 ;
        RECT 2261.550 4.000 2266.690 4.280 ;
        RECT 2267.530 4.000 2272.670 4.280 ;
        RECT 2273.510 4.000 2278.650 4.280 ;
        RECT 2279.490 4.000 2284.630 4.280 ;
        RECT 2285.470 4.000 2290.610 4.280 ;
      LAYER met3 ;
        RECT 2.825 2967.200 2296.010 2986.725 ;
        RECT 2.825 2965.800 2295.600 2967.200 ;
        RECT 2.825 2964.480 2296.010 2965.800 ;
        RECT 4.400 2963.080 2296.010 2964.480 ;
        RECT 2.825 2900.560 2296.010 2963.080 ;
        RECT 2.825 2899.160 2295.600 2900.560 ;
        RECT 2.825 2893.080 2296.010 2899.160 ;
        RECT 4.400 2891.680 2296.010 2893.080 ;
        RECT 2.825 2833.920 2296.010 2891.680 ;
        RECT 2.825 2832.520 2295.600 2833.920 ;
        RECT 2.825 2821.680 2296.010 2832.520 ;
        RECT 4.400 2820.280 2296.010 2821.680 ;
        RECT 2.825 2767.280 2296.010 2820.280 ;
        RECT 2.825 2765.880 2295.600 2767.280 ;
        RECT 2.825 2750.280 2296.010 2765.880 ;
        RECT 4.400 2748.880 2296.010 2750.280 ;
        RECT 2.825 2700.640 2296.010 2748.880 ;
        RECT 2.825 2699.240 2295.600 2700.640 ;
        RECT 2.825 2678.880 2296.010 2699.240 ;
        RECT 4.400 2677.480 2296.010 2678.880 ;
        RECT 2.825 2634.000 2296.010 2677.480 ;
        RECT 2.825 2632.600 2295.600 2634.000 ;
        RECT 2.825 2607.480 2296.010 2632.600 ;
        RECT 4.400 2606.080 2296.010 2607.480 ;
        RECT 2.825 2567.360 2296.010 2606.080 ;
        RECT 2.825 2565.960 2295.600 2567.360 ;
        RECT 2.825 2536.080 2296.010 2565.960 ;
        RECT 4.400 2534.680 2296.010 2536.080 ;
        RECT 2.825 2500.720 2296.010 2534.680 ;
        RECT 2.825 2499.320 2295.600 2500.720 ;
        RECT 2.825 2464.680 2296.010 2499.320 ;
        RECT 4.400 2463.280 2296.010 2464.680 ;
        RECT 2.825 2434.080 2296.010 2463.280 ;
        RECT 2.825 2432.680 2295.600 2434.080 ;
        RECT 2.825 2393.280 2296.010 2432.680 ;
        RECT 4.400 2391.880 2296.010 2393.280 ;
        RECT 2.825 2367.440 2296.010 2391.880 ;
        RECT 2.825 2366.040 2295.600 2367.440 ;
        RECT 2.825 2321.880 2296.010 2366.040 ;
        RECT 4.400 2320.480 2296.010 2321.880 ;
        RECT 2.825 2300.800 2296.010 2320.480 ;
        RECT 2.825 2299.400 2295.600 2300.800 ;
        RECT 2.825 2250.480 2296.010 2299.400 ;
        RECT 4.400 2249.080 2296.010 2250.480 ;
        RECT 2.825 2234.160 2296.010 2249.080 ;
        RECT 2.825 2232.760 2295.600 2234.160 ;
        RECT 2.825 2179.080 2296.010 2232.760 ;
        RECT 4.400 2177.680 2296.010 2179.080 ;
        RECT 2.825 2167.520 2296.010 2177.680 ;
        RECT 2.825 2166.120 2295.600 2167.520 ;
        RECT 2.825 2107.680 2296.010 2166.120 ;
        RECT 4.400 2106.280 2296.010 2107.680 ;
        RECT 2.825 2100.880 2296.010 2106.280 ;
        RECT 2.825 2099.480 2295.600 2100.880 ;
        RECT 2.825 2036.280 2296.010 2099.480 ;
        RECT 4.400 2034.880 2296.010 2036.280 ;
        RECT 2.825 2034.240 2296.010 2034.880 ;
        RECT 2.825 2032.840 2295.600 2034.240 ;
        RECT 2.825 1967.600 2296.010 2032.840 ;
        RECT 2.825 1966.200 2295.600 1967.600 ;
        RECT 2.825 1964.880 2296.010 1966.200 ;
        RECT 4.400 1963.480 2296.010 1964.880 ;
        RECT 2.825 1900.960 2296.010 1963.480 ;
        RECT 2.825 1899.560 2295.600 1900.960 ;
        RECT 2.825 1893.480 2296.010 1899.560 ;
        RECT 4.400 1892.080 2296.010 1893.480 ;
        RECT 2.825 1834.320 2296.010 1892.080 ;
        RECT 2.825 1832.920 2295.600 1834.320 ;
        RECT 2.825 1822.080 2296.010 1832.920 ;
        RECT 4.400 1820.680 2296.010 1822.080 ;
        RECT 2.825 1767.680 2296.010 1820.680 ;
        RECT 2.825 1766.280 2295.600 1767.680 ;
        RECT 2.825 1750.680 2296.010 1766.280 ;
        RECT 4.400 1749.280 2296.010 1750.680 ;
        RECT 2.825 1701.040 2296.010 1749.280 ;
        RECT 2.825 1699.640 2295.600 1701.040 ;
        RECT 2.825 1679.280 2296.010 1699.640 ;
        RECT 4.400 1677.880 2296.010 1679.280 ;
        RECT 2.825 1634.400 2296.010 1677.880 ;
        RECT 2.825 1633.000 2295.600 1634.400 ;
        RECT 2.825 1607.880 2296.010 1633.000 ;
        RECT 4.400 1606.480 2296.010 1607.880 ;
        RECT 2.825 1567.760 2296.010 1606.480 ;
        RECT 2.825 1566.360 2295.600 1567.760 ;
        RECT 2.825 1536.480 2296.010 1566.360 ;
        RECT 4.400 1535.080 2296.010 1536.480 ;
        RECT 2.825 1500.440 2296.010 1535.080 ;
        RECT 2.825 1499.040 2295.600 1500.440 ;
        RECT 2.825 1464.400 2296.010 1499.040 ;
        RECT 4.400 1463.000 2296.010 1464.400 ;
        RECT 2.825 1433.800 2296.010 1463.000 ;
        RECT 2.825 1432.400 2295.600 1433.800 ;
        RECT 2.825 1393.000 2296.010 1432.400 ;
        RECT 4.400 1391.600 2296.010 1393.000 ;
        RECT 2.825 1367.160 2296.010 1391.600 ;
        RECT 2.825 1365.760 2295.600 1367.160 ;
        RECT 2.825 1321.600 2296.010 1365.760 ;
        RECT 4.400 1320.200 2296.010 1321.600 ;
        RECT 2.825 1300.520 2296.010 1320.200 ;
        RECT 2.825 1299.120 2295.600 1300.520 ;
        RECT 2.825 1250.200 2296.010 1299.120 ;
        RECT 4.400 1248.800 2296.010 1250.200 ;
        RECT 2.825 1233.880 2296.010 1248.800 ;
        RECT 2.825 1232.480 2295.600 1233.880 ;
        RECT 2.825 1178.800 2296.010 1232.480 ;
        RECT 4.400 1177.400 2296.010 1178.800 ;
        RECT 2.825 1167.240 2296.010 1177.400 ;
        RECT 2.825 1165.840 2295.600 1167.240 ;
        RECT 2.825 1107.400 2296.010 1165.840 ;
        RECT 4.400 1106.000 2296.010 1107.400 ;
        RECT 2.825 1100.600 2296.010 1106.000 ;
        RECT 2.825 1099.200 2295.600 1100.600 ;
        RECT 2.825 1036.000 2296.010 1099.200 ;
        RECT 4.400 1034.600 2296.010 1036.000 ;
        RECT 2.825 1033.960 2296.010 1034.600 ;
        RECT 2.825 1032.560 2295.600 1033.960 ;
        RECT 2.825 967.320 2296.010 1032.560 ;
        RECT 2.825 965.920 2295.600 967.320 ;
        RECT 2.825 964.600 2296.010 965.920 ;
        RECT 4.400 963.200 2296.010 964.600 ;
        RECT 2.825 900.680 2296.010 963.200 ;
        RECT 2.825 899.280 2295.600 900.680 ;
        RECT 2.825 893.200 2296.010 899.280 ;
        RECT 4.400 891.800 2296.010 893.200 ;
        RECT 2.825 834.040 2296.010 891.800 ;
        RECT 2.825 832.640 2295.600 834.040 ;
        RECT 2.825 821.800 2296.010 832.640 ;
        RECT 4.400 820.400 2296.010 821.800 ;
        RECT 2.825 767.400 2296.010 820.400 ;
        RECT 2.825 766.000 2295.600 767.400 ;
        RECT 2.825 750.400 2296.010 766.000 ;
        RECT 4.400 749.000 2296.010 750.400 ;
        RECT 2.825 700.760 2296.010 749.000 ;
        RECT 2.825 699.360 2295.600 700.760 ;
        RECT 2.825 679.000 2296.010 699.360 ;
        RECT 4.400 677.600 2296.010 679.000 ;
        RECT 2.825 634.120 2296.010 677.600 ;
        RECT 2.825 632.720 2295.600 634.120 ;
        RECT 2.825 607.600 2296.010 632.720 ;
        RECT 4.400 606.200 2296.010 607.600 ;
        RECT 2.825 567.480 2296.010 606.200 ;
        RECT 2.825 566.080 2295.600 567.480 ;
        RECT 2.825 536.200 2296.010 566.080 ;
        RECT 4.400 534.800 2296.010 536.200 ;
        RECT 2.825 500.840 2296.010 534.800 ;
        RECT 2.825 499.440 2295.600 500.840 ;
        RECT 2.825 464.800 2296.010 499.440 ;
        RECT 4.400 463.400 2296.010 464.800 ;
        RECT 2.825 434.200 2296.010 463.400 ;
        RECT 2.825 432.800 2295.600 434.200 ;
        RECT 2.825 393.400 2296.010 432.800 ;
        RECT 4.400 392.000 2296.010 393.400 ;
        RECT 2.825 367.560 2296.010 392.000 ;
        RECT 2.825 366.160 2295.600 367.560 ;
        RECT 2.825 322.000 2296.010 366.160 ;
        RECT 4.400 320.600 2296.010 322.000 ;
        RECT 2.825 300.920 2296.010 320.600 ;
        RECT 2.825 299.520 2295.600 300.920 ;
        RECT 2.825 250.600 2296.010 299.520 ;
        RECT 4.400 249.200 2296.010 250.600 ;
        RECT 2.825 234.280 2296.010 249.200 ;
        RECT 2.825 232.880 2295.600 234.280 ;
        RECT 2.825 179.200 2296.010 232.880 ;
        RECT 4.400 177.800 2296.010 179.200 ;
        RECT 2.825 167.640 2296.010 177.800 ;
        RECT 2.825 166.240 2295.600 167.640 ;
        RECT 2.825 107.800 2296.010 166.240 ;
        RECT 4.400 106.400 2296.010 107.800 ;
        RECT 2.825 101.000 2296.010 106.400 ;
        RECT 2.825 99.600 2295.600 101.000 ;
        RECT 2.825 36.400 2296.010 99.600 ;
        RECT 4.400 35.000 2296.010 36.400 ;
        RECT 2.825 34.360 2296.010 35.000 ;
        RECT 2.825 32.960 2295.600 34.360 ;
        RECT 2.825 4.255 2296.010 32.960 ;
      LAYER met4 ;
        RECT 76.655 10.640 97.440 2986.800 ;
        RECT 99.840 10.640 2254.625 2986.800 ;
  END
END ghazi_top_dffram_csv
END LIBRARY

