magic
tech sky130A
magscale 1 2
timestamp 1607663363
<< locali >>
rect 8125 685899 8159 695453
rect 72525 683247 72559 692733
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72709 678895 72743 683077
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 72801 656931 72835 666485
rect 219081 656931 219115 666485
rect 278973 48331 279007 49045
rect 427921 48331 427955 49113
rect 434821 48331 434855 49045
rect 285781 37315 285815 46869
rect 427921 29019 427955 38573
rect 434821 29019 434855 38573
rect 248429 9707 248463 19261
rect 259469 9707 259503 19261
rect 269129 9707 269163 19261
rect 278973 9707 279007 19261
rect 284309 9707 284343 19261
rect 285781 9707 285815 27557
rect 301421 9707 301455 13141
rect 427921 9707 427955 19261
rect 434821 9707 434855 19261
rect 249809 5083 249843 5185
rect 259377 5015 259411 5185
rect 260849 5015 260883 5117
rect 270509 5015 270543 5117
rect 278789 4879 278823 5117
rect 287069 4743 287103 4845
rect 296637 4743 296671 4981
rect 393329 4743 393363 4845
rect 402989 4743 403023 4845
rect 419273 4743 419307 4913
rect 425069 4675 425103 4913
rect 350491 3417 350641 3451
rect 431141 595 431175 9605
rect 434637 4675 434671 4845
rect 434729 4743 434763 4913
rect 437029 595 437063 9605
rect 444297 4743 444331 4845
rect 445125 2975 445159 4845
rect 528569 3315 528603 3553
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 692733 72559 692767
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 72525 683213 72559 683247
rect 154313 685797 154347 685831
rect 72709 683077 72743 683111
rect 72709 678861 72743 678895
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 284033 676209 284067 676243
rect 72801 666485 72835 666519
rect 72801 656897 72835 656931
rect 219081 666485 219115 666519
rect 219081 656897 219115 656931
rect 427921 49113 427955 49147
rect 278973 49045 279007 49079
rect 278973 48297 279007 48331
rect 427921 48297 427955 48331
rect 434821 49045 434855 49079
rect 434821 48297 434855 48331
rect 285781 46869 285815 46903
rect 285781 37281 285815 37315
rect 427921 38573 427955 38607
rect 427921 28985 427955 29019
rect 434821 38573 434855 38607
rect 434821 28985 434855 29019
rect 285781 27557 285815 27591
rect 248429 19261 248463 19295
rect 248429 9673 248463 9707
rect 259469 19261 259503 19295
rect 259469 9673 259503 9707
rect 269129 19261 269163 19295
rect 269129 9673 269163 9707
rect 278973 19261 279007 19295
rect 278973 9673 279007 9707
rect 284309 19261 284343 19295
rect 284309 9673 284343 9707
rect 427921 19261 427955 19295
rect 285781 9673 285815 9707
rect 301421 13141 301455 13175
rect 301421 9673 301455 9707
rect 427921 9673 427955 9707
rect 434821 19261 434855 19295
rect 434821 9673 434855 9707
rect 431141 9605 431175 9639
rect 249809 5185 249843 5219
rect 249809 5049 249843 5083
rect 259377 5185 259411 5219
rect 259377 4981 259411 5015
rect 260849 5117 260883 5151
rect 260849 4981 260883 5015
rect 270509 5117 270543 5151
rect 270509 4981 270543 5015
rect 278789 5117 278823 5151
rect 296637 4981 296671 5015
rect 278789 4845 278823 4879
rect 287069 4845 287103 4879
rect 287069 4709 287103 4743
rect 419273 4913 419307 4947
rect 296637 4709 296671 4743
rect 393329 4845 393363 4879
rect 393329 4709 393363 4743
rect 402989 4845 403023 4879
rect 402989 4709 403023 4743
rect 419273 4709 419307 4743
rect 425069 4913 425103 4947
rect 425069 4641 425103 4675
rect 350457 3417 350491 3451
rect 350641 3417 350675 3451
rect 437029 9605 437063 9639
rect 434729 4913 434763 4947
rect 434637 4845 434671 4879
rect 434729 4709 434763 4743
rect 434637 4641 434671 4675
rect 431141 561 431175 595
rect 444297 4845 444331 4879
rect 444297 4709 444331 4743
rect 445125 4845 445159 4879
rect 528569 3553 528603 3587
rect 528569 3281 528603 3315
rect 445125 2941 445159 2975
rect 437029 561 437063 595
<< metal1 >>
rect 411162 700408 411168 700460
rect 411220 700448 411226 700460
rect 429838 700448 429844 700460
rect 411220 700420 429844 700448
rect 411220 700408 411226 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 463602 700408 463608 700460
rect 463660 700448 463666 700460
rect 494790 700448 494796 700460
rect 463660 700420 494796 700448
rect 463660 700408 463666 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 514662 700408 514668 700460
rect 514720 700448 514726 700460
rect 559650 700448 559656 700460
rect 514720 700420 559656 700448
rect 514720 700408 514726 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 394602 700340 394608 700392
rect 394660 700380 394666 700392
rect 413646 700380 413652 700392
rect 394660 700352 413652 700380
rect 394660 700340 394666 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 445662 700340 445668 700392
rect 445720 700380 445726 700392
rect 478506 700380 478512 700392
rect 445720 700352 478512 700380
rect 445720 700340 445726 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 496722 700340 496728 700392
rect 496780 700380 496786 700392
rect 543458 700380 543464 700392
rect 496780 700352 543464 700380
rect 496780 700340 496786 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 343542 700272 343548 700324
rect 343600 700312 343606 700324
rect 348786 700312 348792 700324
rect 343600 700284 348792 700312
rect 343600 700272 343606 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 378042 700272 378048 700324
rect 378100 700312 378106 700324
rect 397454 700312 397460 700324
rect 378100 700284 397460 700312
rect 378100 700272 378106 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 429102 700272 429108 700324
rect 429160 700312 429166 700324
rect 462314 700312 462320 700324
rect 429160 700284 462320 700312
rect 429160 700272 429166 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 480162 700272 480168 700324
rect 480220 700312 480226 700324
rect 527174 700312 527180 700324
rect 480220 700284 527180 700312
rect 480220 700272 480226 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 326982 699660 326988 699712
rect 327040 699700 327046 699712
rect 332502 699700 332508 699712
rect 327040 699672 332508 699700
rect 327040 699660 327046 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 360102 699660 360108 699712
rect 360160 699700 360166 699712
rect 364978 699700 364984 699712
rect 360160 699672 364984 699700
rect 360160 699660 360166 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 523770 696940 523776 696992
rect 523828 696980 523834 696992
rect 580166 696980 580172 696992
rect 523828 696952 580172 696980
rect 523828 696940 523834 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 692767 72571 692773
rect 72513 692733 72525 692767
rect 72559 692764 72571 692767
rect 72694 692764 72700 692776
rect 72559 692736 72700 692764
rect 72559 692733 72571 692736
rect 72513 692727 72571 692733
rect 72694 692724 72700 692736
rect 72752 692724 72758 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 523678 685856 523684 685908
rect 523736 685896 523742 685908
rect 580166 685896 580172 685908
rect 523736 685868 580172 685896
rect 523736 685856 523742 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 683244 72516 683256
rect 72471 683216 72516 683244
rect 72510 683204 72516 683216
rect 72568 683204 72574 683256
rect 72510 683068 72516 683120
rect 72568 683108 72574 683120
rect 72697 683111 72755 683117
rect 72697 683108 72709 683111
rect 72568 683080 72709 683108
rect 72568 683068 72574 683080
rect 72697 683077 72709 683080
rect 72743 683077 72755 683111
rect 72697 683071 72755 683077
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 219066 679028 219072 679040
rect 218992 679000 219072 679028
rect 218992 678972 219020 679000
rect 219066 678988 219072 679000
rect 219124 678988 219130 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 218974 678920 218980 678972
rect 219032 678920 219038 678972
rect 72694 678892 72700 678904
rect 72655 678864 72700 678892
rect 72694 678852 72700 678864
rect 72752 678852 72758 678904
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 72694 669264 72700 669316
rect 72752 669304 72758 669316
rect 72878 669304 72884 669316
rect 72752 669276 72884 669304
rect 72752 669264 72758 669276
rect 72878 669264 72884 669276
rect 72936 669264 72942 669316
rect 218974 669264 218980 669316
rect 219032 669304 219038 669316
rect 219158 669304 219164 669316
rect 219032 669276 219164 669304
rect 219032 669264 219038 669276
rect 219158 669264 219164 669276
rect 219216 669264 219222 669316
rect 72789 666519 72847 666525
rect 72789 666485 72801 666519
rect 72835 666516 72847 666519
rect 72878 666516 72884 666528
rect 72835 666488 72884 666516
rect 72835 666485 72847 666488
rect 72789 666479 72847 666485
rect 72878 666476 72884 666488
rect 72936 666476 72942 666528
rect 219069 666519 219127 666525
rect 219069 666485 219081 666519
rect 219115 666516 219127 666519
rect 219158 666516 219164 666528
rect 219115 666488 219164 666516
rect 219115 666485 219127 666488
rect 219069 666479 219127 666485
rect 219158 666476 219164 666488
rect 219216 666476 219222 666528
rect 72786 656928 72792 656940
rect 72747 656900 72792 656928
rect 72786 656888 72792 656900
rect 72844 656888 72850 656940
rect 219066 656928 219072 656940
rect 219027 656900 219072 656928
rect 219066 656888 219072 656900
rect 219124 656888 219130 656940
rect 377122 655460 377128 655512
rect 377180 655500 377186 655512
rect 378042 655500 378048 655512
rect 377180 655472 378048 655500
rect 377180 655460 377186 655472
rect 378042 655460 378048 655472
rect 378100 655460 378106 655512
rect 428182 655460 428188 655512
rect 428240 655500 428246 655512
rect 429102 655500 429108 655512
rect 428240 655472 429108 655500
rect 428240 655460 428246 655472
rect 429102 655460 429108 655472
rect 429160 655460 429166 655512
rect 462314 655460 462320 655512
rect 462372 655500 462378 655512
rect 463602 655500 463608 655512
rect 462372 655472 463608 655500
rect 462372 655460 462378 655472
rect 463602 655460 463608 655472
rect 463660 655460 463666 655512
rect 479334 655460 479340 655512
rect 479392 655500 479398 655512
rect 480162 655500 480168 655512
rect 479392 655472 480168 655500
rect 479392 655460 479398 655472
rect 480162 655460 480168 655472
rect 480220 655460 480226 655512
rect 513374 655256 513380 655308
rect 513432 655296 513438 655308
rect 514662 655296 514668 655308
rect 513432 655268 514668 655296
rect 513432 655256 513438 655268
rect 514662 655256 514668 655268
rect 514720 655256 514726 655308
rect 325970 655120 325976 655172
rect 326028 655160 326034 655172
rect 326982 655160 326988 655172
rect 326028 655132 326988 655160
rect 326028 655120 326034 655132
rect 326982 655120 326988 655132
rect 327040 655120 327046 655172
rect 154298 654984 154304 655036
rect 154356 655024 154362 655036
rect 189718 655024 189724 655036
rect 154356 654996 189724 655024
rect 154356 654984 154362 654996
rect 189718 654984 189724 654996
rect 189776 654984 189782 655036
rect 41322 654916 41328 654968
rect 41380 654956 41386 654968
rect 104526 654956 104532 654968
rect 41380 654928 104532 654956
rect 41380 654916 41386 654928
rect 104526 654916 104532 654928
rect 104584 654916 104590 654968
rect 106182 654916 106188 654968
rect 106240 654956 106246 654968
rect 155586 654956 155592 654968
rect 106240 654928 155592 654956
rect 106240 654916 106246 654928
rect 155586 654916 155592 654928
rect 155644 654916 155650 654968
rect 24762 654848 24768 654900
rect 24820 654888 24826 654900
rect 87506 654888 87512 654900
rect 24820 654860 87512 654888
rect 24820 654848 24826 654860
rect 87506 654848 87512 654860
rect 87564 654848 87570 654900
rect 89622 654848 89628 654900
rect 89680 654888 89686 654900
rect 138566 654888 138572 654900
rect 89680 654860 138572 654888
rect 89680 654848 89686 654860
rect 138566 654848 138572 654860
rect 138624 654848 138630 654900
rect 171042 654848 171048 654900
rect 171100 654888 171106 654900
rect 206738 654888 206744 654900
rect 171100 654860 206744 654888
rect 171100 654848 171106 654860
rect 206738 654848 206744 654860
rect 206796 654848 206802 654900
rect 219066 654848 219072 654900
rect 219124 654888 219130 654900
rect 240778 654888 240784 654900
rect 219124 654860 240784 654888
rect 219124 654848 219130 654860
rect 240778 654848 240784 654860
rect 240836 654848 240842 654900
rect 8018 654780 8024 654832
rect 8076 654820 8082 654832
rect 70486 654820 70492 654832
rect 8076 654792 70492 654820
rect 8076 654780 8082 654792
rect 70486 654780 70492 654792
rect 70544 654780 70550 654832
rect 72786 654780 72792 654832
rect 72844 654820 72850 654832
rect 121546 654820 121552 654832
rect 72844 654792 121552 654820
rect 72844 654780 72850 654792
rect 121546 654780 121552 654792
rect 121604 654780 121610 654832
rect 137738 654780 137744 654832
rect 137796 654820 137802 654832
rect 172698 654820 172704 654832
rect 137796 654792 172704 654820
rect 137796 654780 137802 654792
rect 172698 654780 172704 654792
rect 172756 654780 172762 654832
rect 202782 654780 202788 654832
rect 202840 654820 202846 654832
rect 223758 654820 223764 654832
rect 202840 654792 223764 654820
rect 202840 654780 202846 654792
rect 223758 654780 223764 654792
rect 223816 654780 223822 654832
rect 235902 654780 235908 654832
rect 235960 654820 235966 654832
rect 257890 654820 257896 654832
rect 235960 654792 257896 654820
rect 235960 654780 235966 654792
rect 257890 654780 257896 654792
rect 257948 654780 257954 654832
rect 267642 654780 267648 654832
rect 267700 654820 267706 654832
rect 274910 654820 274916 654832
rect 267700 654792 274916 654820
rect 267700 654780 267706 654792
rect 274910 654780 274916 654792
rect 274968 654780 274974 654832
rect 284018 654780 284024 654832
rect 284076 654820 284082 654832
rect 291930 654820 291936 654832
rect 284076 654792 291936 654820
rect 284076 654780 284082 654792
rect 291930 654780 291936 654792
rect 291988 654780 291994 654832
rect 300762 654100 300768 654152
rect 300820 654140 300826 654152
rect 308950 654140 308956 654152
rect 300820 654112 308956 654140
rect 300820 654100 300826 654112
rect 308950 654100 308956 654112
rect 309008 654100 309014 654152
rect 3510 645804 3516 645856
rect 3568 645844 3574 645856
rect 59354 645844 59360 645856
rect 3568 645816 59360 645844
rect 3568 645804 3574 645816
rect 59354 645804 59360 645816
rect 59412 645804 59418 645856
rect 523770 638936 523776 638988
rect 523828 638976 523834 638988
rect 580166 638976 580172 638988
rect 523828 638948 580172 638976
rect 523828 638936 523834 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 3418 630572 3424 630624
rect 3476 630612 3482 630624
rect 59354 630612 59360 630624
rect 3476 630584 59360 630612
rect 3476 630572 3482 630584
rect 59354 630572 59360 630584
rect 59412 630572 59418 630624
rect 524322 619556 524328 619608
rect 524380 619596 524386 619608
rect 580258 619596 580264 619608
rect 524380 619568 580264 619596
rect 524380 619556 524386 619568
rect 580258 619556 580264 619568
rect 580316 619556 580322 619608
rect 3602 616768 3608 616820
rect 3660 616808 3666 616820
rect 59354 616808 59360 616820
rect 3660 616780 59360 616808
rect 3660 616768 3666 616780
rect 59354 616768 59360 616780
rect 59412 616768 59418 616820
rect 523126 605752 523132 605804
rect 523184 605792 523190 605804
rect 580442 605792 580448 605804
rect 523184 605764 580448 605792
rect 523184 605752 523190 605764
rect 580442 605752 580448 605764
rect 580500 605752 580506 605804
rect 3510 603032 3516 603084
rect 3568 603072 3574 603084
rect 59354 603072 59360 603084
rect 3568 603044 59360 603072
rect 3568 603032 3574 603044
rect 59354 603032 59360 603044
rect 59412 603032 59418 603084
rect 523678 592016 523684 592068
rect 523736 592056 523742 592068
rect 579798 592056 579804 592068
rect 523736 592028 579804 592056
rect 523736 592016 523742 592028
rect 579798 592016 579804 592028
rect 579856 592016 579862 592068
rect 3418 587800 3424 587852
rect 3476 587840 3482 587852
rect 59354 587840 59360 587852
rect 3476 587812 59360 587840
rect 3476 587800 3482 587812
rect 59354 587800 59360 587812
rect 59412 587800 59418 587852
rect 524322 579572 524328 579624
rect 524380 579612 524386 579624
rect 580350 579612 580356 579624
rect 524380 579584 580356 579612
rect 524380 579572 524386 579584
rect 580350 579572 580356 579584
rect 580408 579572 580414 579624
rect 3510 573996 3516 574048
rect 3568 574036 3574 574048
rect 59354 574036 59360 574048
rect 3568 574008 59360 574036
rect 3568 573996 3574 574008
rect 59354 573996 59360 574008
rect 59412 573996 59418 574048
rect 523126 565768 523132 565820
rect 523184 565808 523190 565820
rect 580442 565808 580448 565820
rect 523184 565780 580448 565808
rect 523184 565768 523190 565780
rect 580442 565768 580448 565780
rect 580500 565768 580506 565820
rect 3418 560192 3424 560244
rect 3476 560232 3482 560244
rect 59354 560232 59360 560244
rect 3476 560204 59360 560232
rect 3476 560192 3482 560204
rect 59354 560192 59360 560204
rect 59412 560192 59418 560244
rect 523770 556180 523776 556232
rect 523828 556220 523834 556232
rect 580166 556220 580172 556232
rect 523828 556192 580172 556220
rect 523828 556180 523834 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 523494 545096 523500 545148
rect 523552 545136 523558 545148
rect 580166 545136 580172 545148
rect 523552 545108 580172 545136
rect 523552 545096 523558 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 3418 545028 3424 545080
rect 3476 545068 3482 545080
rect 59354 545068 59360 545080
rect 3476 545040 59360 545068
rect 3476 545028 3482 545040
rect 59354 545028 59360 545040
rect 59412 545028 59418 545080
rect 523678 539520 523684 539572
rect 523736 539560 523742 539572
rect 580258 539560 580264 539572
rect 523736 539532 580264 539560
rect 523736 539520 523742 539532
rect 580258 539520 580264 539532
rect 580316 539520 580322 539572
rect 3418 531224 3424 531276
rect 3476 531264 3482 531276
rect 59354 531264 59360 531276
rect 3476 531236 59360 531264
rect 3476 531224 3482 531236
rect 59354 531224 59360 531236
rect 59412 531224 59418 531276
rect 3142 510552 3148 510604
rect 3200 510592 3206 510604
rect 59354 510592 59360 510604
rect 3200 510564 59360 510592
rect 3200 510552 3206 510564
rect 59354 510552 59360 510564
rect 59412 510552 59418 510604
rect 523770 509260 523776 509312
rect 523828 509300 523834 509312
rect 580166 509300 580172 509312
rect 523828 509272 580172 509300
rect 523828 509260 523834 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 523678 499468 523684 499520
rect 523736 499508 523742 499520
rect 580258 499508 580264 499520
rect 523736 499480 580264 499508
rect 523736 499468 523742 499480
rect 580258 499468 580264 499480
rect 580316 499468 580322 499520
rect 523678 498176 523684 498228
rect 523736 498216 523742 498228
rect 580166 498216 580172 498228
rect 523736 498188 580172 498216
rect 523736 498176 523742 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3418 496748 3424 496800
rect 3476 496788 3482 496800
rect 59998 496788 60004 496800
rect 3476 496760 60004 496788
rect 3476 496748 3482 496760
rect 59998 496748 60004 496760
rect 60056 496748 60062 496800
rect 3510 481584 3516 481636
rect 3568 481624 3574 481636
rect 59354 481624 59360 481636
rect 3568 481596 59360 481624
rect 3568 481584 3574 481596
rect 59354 481584 59360 481596
rect 59412 481584 59418 481636
rect 523678 462340 523684 462392
rect 523736 462380 523742 462392
rect 580166 462380 580172 462392
rect 523736 462352 580172 462380
rect 523736 462340 523742 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 524322 459484 524328 459536
rect 524380 459524 524386 459536
rect 580258 459524 580264 459536
rect 524380 459496 580264 459524
rect 524380 459484 524386 459496
rect 580258 459484 580264 459496
rect 580316 459484 580322 459536
rect 3418 452548 3424 452600
rect 3476 452588 3482 452600
rect 59998 452588 60004 452600
rect 3476 452560 60004 452588
rect 3476 452548 3482 452560
rect 59998 452548 60004 452560
rect 60056 452548 60062 452600
rect 523770 451256 523776 451308
rect 523828 451296 523834 451308
rect 580166 451296 580172 451308
rect 523828 451268 580172 451296
rect 523828 451256 523834 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 523678 438880 523684 438932
rect 523736 438920 523742 438932
rect 580166 438920 580172 438932
rect 523736 438892 580172 438920
rect 523736 438880 523742 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3142 438812 3148 438864
rect 3200 438852 3206 438864
rect 60090 438852 60096 438864
rect 3200 438824 60096 438852
rect 3200 438812 3206 438824
rect 60090 438812 60096 438824
rect 60148 438812 60154 438864
rect 3234 425008 3240 425060
rect 3292 425048 3298 425060
rect 59998 425048 60004 425060
rect 3292 425020 60004 425048
rect 3292 425008 3298 425020
rect 59998 425008 60004 425020
rect 60056 425008 60062 425060
rect 523678 415420 523684 415472
rect 523736 415460 523742 415472
rect 580166 415460 580172 415472
rect 523736 415432 580172 415460
rect 523736 415420 523742 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 523770 404336 523776 404388
rect 523828 404376 523834 404388
rect 580166 404376 580172 404388
rect 523828 404348 580172 404376
rect 523828 404336 523834 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 60090 396012 60096 396024
rect 3200 395984 60096 396012
rect 3200 395972 3206 395984
rect 60090 395972 60096 395984
rect 60148 395972 60154 396024
rect 523678 391960 523684 392012
rect 523736 392000 523742 392012
rect 580166 392000 580172 392012
rect 523736 391972 580172 392000
rect 523736 391960 523742 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 60182 380848 60188 380860
rect 3292 380820 60188 380848
rect 3292 380808 3298 380820
rect 60182 380808 60188 380820
rect 60240 380808 60246 380860
rect 524230 368500 524236 368552
rect 524288 368540 524294 368552
rect 580166 368540 580172 368552
rect 524288 368512 580172 368540
rect 524288 368500 524294 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 59998 367044 60004 367056
rect 3200 367016 60004 367044
rect 3200 367004 3206 367016
rect 59998 367004 60004 367016
rect 60056 367004 60062 367056
rect 523678 357416 523684 357468
rect 523736 357456 523742 357468
rect 580166 357456 580172 357468
rect 523736 357428 580172 357456
rect 523736 357416 523742 357428
rect 580166 357416 580172 357428
rect 580224 357416 580230 357468
rect 523770 345040 523776 345092
rect 523828 345080 523834 345092
rect 580166 345080 580172 345092
rect 523828 345052 580172 345080
rect 523828 345040 523834 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 60090 338076 60096 338088
rect 3476 338048 60096 338076
rect 3476 338036 3482 338048
rect 60090 338036 60096 338048
rect 60148 338036 60154 338088
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 60182 324272 60188 324284
rect 3292 324244 60188 324272
rect 3292 324232 3298 324244
rect 60182 324232 60188 324244
rect 60240 324232 60246 324284
rect 524322 322872 524328 322924
rect 524380 322912 524386 322924
rect 580166 322912 580172 322924
rect 524380 322884 580172 322912
rect 524380 322872 524386 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 524322 311788 524328 311840
rect 524380 311828 524386 311840
rect 580166 311828 580172 311840
rect 524380 311800 580172 311828
rect 524380 311788 524386 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 59998 309108 60004 309120
rect 3384 309080 60004 309108
rect 3384 309068 3390 309080
rect 59998 309068 60004 309080
rect 60056 309068 60062 309120
rect 524322 298732 524328 298784
rect 524380 298772 524386 298784
rect 580166 298772 580172 298784
rect 524380 298744 580172 298772
rect 524380 298732 524386 298744
rect 580166 298732 580172 298744
rect 580224 298732 580230 298784
rect 3418 295264 3424 295316
rect 3476 295304 3482 295316
rect 60366 295304 60372 295316
rect 3476 295276 60372 295304
rect 3476 295264 3482 295276
rect 60366 295264 60372 295276
rect 60424 295264 60430 295316
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 60090 280140 60096 280152
rect 3476 280112 60096 280140
rect 3476 280100 3482 280112
rect 60090 280100 60096 280112
rect 60148 280100 60154 280152
rect 523678 275952 523684 276004
rect 523736 275992 523742 276004
rect 580166 275992 580172 276004
rect 523736 275964 580172 275992
rect 523736 275952 523742 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 3142 266296 3148 266348
rect 3200 266336 3206 266348
rect 60274 266336 60280 266348
rect 3200 266308 60280 266336
rect 3200 266296 3206 266308
rect 60274 266296 60280 266308
rect 60332 266296 60338 266348
rect 523678 264868 523684 264920
rect 523736 264908 523742 264920
rect 580166 264908 580172 264920
rect 523736 264880 580172 264908
rect 523736 264868 523742 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 3418 252492 3424 252544
rect 3476 252532 3482 252544
rect 60458 252532 60464 252544
rect 3476 252504 60464 252532
rect 3476 252492 3482 252504
rect 60458 252492 60464 252504
rect 60516 252492 60522 252544
rect 523678 252492 523684 252544
rect 523736 252532 523742 252544
rect 579798 252532 579804 252544
rect 523736 252504 579804 252532
rect 523736 252492 523742 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 59998 237368 60004 237380
rect 3476 237340 60004 237368
rect 3476 237328 3482 237340
rect 59998 237328 60004 237340
rect 60056 237328 60062 237380
rect 523678 229032 523684 229084
rect 523736 229072 523742 229084
rect 580166 229072 580172 229084
rect 523736 229044 580172 229072
rect 523736 229032 523742 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 60182 223564 60188 223576
rect 3200 223536 60188 223564
rect 3200 223524 3206 223536
rect 60182 223524 60188 223536
rect 60240 223524 60246 223576
rect 523770 217948 523776 218000
rect 523828 217988 523834 218000
rect 580166 217988 580172 218000
rect 523828 217960 580172 217988
rect 523828 217948 523834 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 60090 208332 60096 208344
rect 3476 208304 60096 208332
rect 3476 208292 3482 208304
rect 60090 208292 60096 208304
rect 60148 208292 60154 208344
rect 523862 205572 523868 205624
rect 523920 205612 523926 205624
rect 579798 205612 579804 205624
rect 523920 205584 579804 205612
rect 523920 205572 523926 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 60274 194528 60280 194540
rect 3200 194500 60280 194528
rect 3200 194488 3206 194500
rect 60274 194488 60280 194500
rect 60332 194488 60338 194540
rect 523678 182112 523684 182164
rect 523736 182152 523742 182164
rect 580166 182152 580172 182164
rect 523736 182124 580172 182152
rect 523736 182112 523742 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 60366 180792 60372 180804
rect 3292 180764 60372 180792
rect 3292 180752 3298 180764
rect 60366 180752 60372 180764
rect 60424 180752 60430 180804
rect 523770 171028 523776 171080
rect 523828 171068 523834 171080
rect 580166 171068 580172 171080
rect 523828 171040 580172 171068
rect 523828 171028 523834 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 60182 165560 60188 165572
rect 3568 165532 60188 165560
rect 3568 165520 3574 165532
rect 60182 165520 60188 165532
rect 60240 165520 60246 165572
rect 523862 158652 523868 158704
rect 523920 158692 523926 158704
rect 579798 158692 579804 158704
rect 523920 158664 579804 158692
rect 523920 158652 523926 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 60090 151756 60096 151768
rect 3200 151728 60096 151756
rect 3200 151716 3206 151728
rect 60090 151716 60096 151728
rect 60148 151716 60154 151768
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 59998 136592 60004 136604
rect 3292 136564 60004 136592
rect 3292 136552 3298 136564
rect 59998 136552 60004 136564
rect 60056 136552 60062 136604
rect 523678 135192 523684 135244
rect 523736 135232 523742 135244
rect 580166 135232 580172 135244
rect 523736 135204 580172 135232
rect 523736 135192 523742 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 523770 124108 523776 124160
rect 523828 124148 523834 124160
rect 580166 124148 580172 124160
rect 523828 124120 580172 124148
rect 523828 124108 523834 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 3418 122748 3424 122800
rect 3476 122788 3482 122800
rect 60366 122788 60372 122800
rect 3476 122760 60372 122788
rect 3476 122748 3482 122760
rect 60366 122748 60372 122760
rect 60424 122748 60430 122800
rect 523862 111732 523868 111784
rect 523920 111772 523926 111784
rect 579798 111772 579804 111784
rect 523920 111744 579804 111772
rect 523920 111732 523926 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 60274 108984 60280 108996
rect 3292 108956 60280 108984
rect 3292 108944 3298 108956
rect 60274 108944 60280 108956
rect 60332 108944 60338 108996
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 60182 93820 60188 93832
rect 3476 93792 60188 93820
rect 3476 93780 3482 93792
rect 60182 93780 60188 93792
rect 60240 93780 60246 93832
rect 523678 88272 523684 88324
rect 523736 88312 523742 88324
rect 580166 88312 580172 88324
rect 523736 88284 580172 88312
rect 523736 88272 523742 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 3418 79976 3424 80028
rect 3476 80016 3482 80028
rect 59998 80016 60004 80028
rect 3476 79988 60004 80016
rect 3476 79976 3482 79988
rect 59998 79976 60004 79988
rect 60056 79976 60062 80028
rect 523770 77188 523776 77240
rect 523828 77228 523834 77240
rect 580166 77228 580172 77240
rect 523828 77200 580172 77228
rect 523828 77188 523834 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 60090 64852 60096 64864
rect 3384 64824 60096 64852
rect 3384 64812 3390 64824
rect 60090 64812 60096 64824
rect 60148 64812 60154 64864
rect 523862 64812 523868 64864
rect 523920 64852 523926 64864
rect 579798 64852 579804 64864
rect 523920 64824 579804 64852
rect 523920 64812 523926 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 60274 51048 60280 51060
rect 3476 51020 60280 51048
rect 3476 51008 3482 51020
rect 60274 51008 60280 51020
rect 60332 51008 60338 51060
rect 82814 49648 82820 49700
rect 82872 49688 82878 49700
rect 84838 49688 84844 49700
rect 82872 49660 84844 49688
rect 82872 49648 82878 49660
rect 84838 49648 84844 49660
rect 84896 49648 84902 49700
rect 169754 49648 169760 49700
rect 169812 49688 169818 49700
rect 172330 49688 172336 49700
rect 169812 49660 172336 49688
rect 169812 49648 169818 49660
rect 172330 49648 172336 49660
rect 172388 49648 172394 49700
rect 354490 49648 354496 49700
rect 354548 49688 354554 49700
rect 355318 49688 355324 49700
rect 354548 49660 355324 49688
rect 354548 49648 354554 49660
rect 355318 49648 355324 49660
rect 355376 49648 355382 49700
rect 383102 49648 383108 49700
rect 383160 49688 383166 49700
rect 384298 49688 384304 49700
rect 383160 49660 384304 49688
rect 383160 49648 383166 49660
rect 384298 49648 384304 49660
rect 384356 49648 384362 49700
rect 400950 49648 400956 49700
rect 401008 49688 401014 49700
rect 403618 49688 403624 49700
rect 401008 49660 403624 49688
rect 401008 49648 401014 49660
rect 403618 49648 403624 49660
rect 403676 49648 403682 49700
rect 440326 49648 440332 49700
rect 440384 49688 440390 49700
rect 442258 49688 442264 49700
rect 440384 49660 442264 49688
rect 440384 49648 440390 49660
rect 442258 49648 442264 49660
rect 442316 49648 442322 49700
rect 477218 49648 477224 49700
rect 477276 49688 477282 49700
rect 482278 49688 482284 49700
rect 477276 49660 482284 49688
rect 477276 49648 477282 49660
rect 482278 49648 482284 49660
rect 482336 49648 482342 49700
rect 81618 49308 81624 49360
rect 81676 49348 81682 49360
rect 142246 49348 142252 49360
rect 81676 49320 142252 49348
rect 81676 49308 81682 49320
rect 142246 49308 142252 49320
rect 142304 49308 142310 49360
rect 74442 49240 74448 49292
rect 74500 49280 74506 49292
rect 135438 49280 135444 49292
rect 74500 49252 135444 49280
rect 74500 49240 74506 49252
rect 135438 49240 135444 49252
rect 135496 49240 135502 49292
rect 396166 49240 396172 49292
rect 396224 49280 396230 49292
rect 456886 49280 456892 49292
rect 396224 49252 456892 49280
rect 396224 49240 396230 49252
rect 456886 49240 456892 49252
rect 456944 49240 456950 49292
rect 88702 49172 88708 49224
rect 88760 49212 88766 49224
rect 150618 49212 150624 49224
rect 88760 49184 150624 49212
rect 88760 49172 88766 49184
rect 150618 49172 150624 49184
rect 150676 49172 150682 49224
rect 210326 49172 210332 49224
rect 210384 49212 210390 49224
rect 270494 49212 270500 49224
rect 210384 49184 270500 49212
rect 210384 49172 210390 49184
rect 270494 49172 270500 49184
rect 270552 49172 270558 49224
rect 281810 49172 281816 49224
rect 281868 49212 281874 49224
rect 308398 49212 308404 49224
rect 281868 49184 308404 49212
rect 281868 49172 281874 49184
rect 308398 49172 308404 49184
rect 308456 49172 308462 49224
rect 309226 49172 309232 49224
rect 309284 49212 309290 49224
rect 319438 49212 319444 49224
rect 309284 49184 319444 49212
rect 309284 49172 309290 49184
rect 319438 49172 319444 49184
rect 319496 49172 319502 49224
rect 403342 49172 403348 49224
rect 403400 49212 403406 49224
rect 463786 49212 463792 49224
rect 403400 49184 463792 49212
rect 403400 49172 403406 49184
rect 463786 49172 463792 49184
rect 463844 49172 463850 49224
rect 489178 49172 489184 49224
rect 489236 49212 489242 49224
rect 549254 49212 549260 49224
rect 489236 49184 549260 49212
rect 489236 49172 489242 49184
rect 549254 49172 549260 49184
rect 549312 49172 549318 49224
rect 95878 49104 95884 49156
rect 95936 49144 95942 49156
rect 157426 49144 157432 49156
rect 95936 49116 157432 49144
rect 95936 49104 95942 49116
rect 157426 49104 157432 49116
rect 157484 49104 157490 49156
rect 167362 49104 167368 49156
rect 167420 49144 167426 49156
rect 227898 49144 227904 49156
rect 167420 49116 227904 49144
rect 167420 49104 167426 49116
rect 227898 49104 227904 49116
rect 227956 49104 227962 49156
rect 253198 49104 253204 49156
rect 253256 49144 253262 49156
rect 313458 49144 313464 49156
rect 253256 49116 313464 49144
rect 253256 49104 253262 49116
rect 313458 49104 313464 49116
rect 313516 49104 313522 49156
rect 367646 49104 367652 49156
rect 367704 49144 367710 49156
rect 427909 49147 427967 49153
rect 427909 49144 427921 49147
rect 367704 49116 427921 49144
rect 367704 49104 367710 49116
rect 427909 49113 427921 49116
rect 427955 49113 427967 49147
rect 427909 49107 427967 49113
rect 474826 49104 474832 49156
rect 474884 49144 474890 49156
rect 535454 49144 535460 49156
rect 474884 49116 535460 49144
rect 474884 49104 474890 49116
rect 535454 49104 535460 49116
rect 535512 49104 535518 49156
rect 103054 49036 103060 49088
rect 103112 49076 103118 49088
rect 164326 49076 164332 49088
rect 103112 49048 164332 49076
rect 103112 49036 103118 49048
rect 164326 49036 164332 49048
rect 164384 49036 164390 49088
rect 217410 49036 217416 49088
rect 217468 49076 217474 49088
rect 278961 49079 279019 49085
rect 278961 49076 278973 49079
rect 217468 49048 278973 49076
rect 217468 49036 217474 49048
rect 278961 49045 278973 49048
rect 279007 49045 279019 49079
rect 278961 49039 279019 49045
rect 296070 49036 296076 49088
rect 296128 49076 296134 49088
rect 333238 49076 333244 49088
rect 296128 49048 333244 49076
rect 296128 49036 296134 49048
rect 333238 49036 333244 49048
rect 333296 49036 333302 49088
rect 374730 49036 374736 49088
rect 374788 49076 374794 49088
rect 434809 49079 434867 49085
rect 434809 49076 434821 49079
rect 374788 49048 434821 49076
rect 374788 49036 374794 49048
rect 434809 49045 434821 49048
rect 434855 49045 434867 49079
rect 434809 49039 434867 49045
rect 450998 49036 451004 49088
rect 451056 49076 451062 49088
rect 451918 49076 451924 49088
rect 451056 49048 451924 49076
rect 451056 49036 451062 49048
rect 451918 49036 451924 49048
rect 451976 49036 451982 49088
rect 482002 49036 482008 49088
rect 482060 49076 482066 49088
rect 542354 49076 542360 49088
rect 482060 49048 542360 49076
rect 482060 49036 482066 49048
rect 542354 49036 542360 49048
rect 542412 49036 542418 49088
rect 67266 48968 67272 49020
rect 67324 49008 67330 49020
rect 128446 49008 128452 49020
rect 67324 48980 128452 49008
rect 67324 48968 67330 48980
rect 128446 48968 128452 48980
rect 128504 48968 128510 49020
rect 145926 48968 145932 49020
rect 145984 49008 145990 49020
rect 207106 49008 207112 49020
rect 145984 48980 207112 49008
rect 145984 48968 145990 48980
rect 207106 48968 207112 48980
rect 207164 48968 207170 49020
rect 224586 48968 224592 49020
rect 224644 49008 224650 49020
rect 285766 49008 285772 49020
rect 224644 48980 285772 49008
rect 224644 48968 224650 48980
rect 285766 48968 285772 48980
rect 285824 48968 285830 49020
rect 318702 48968 318708 49020
rect 318760 49008 318766 49020
rect 374638 49008 374644 49020
rect 318760 48980 374644 49008
rect 318760 48968 318766 48980
rect 374638 48968 374644 48980
rect 374696 48968 374702 49020
rect 389082 48968 389088 49020
rect 389140 49008 389146 49020
rect 449894 49008 449900 49020
rect 389140 48980 449900 49008
rect 389140 48968 389146 48980
rect 449894 48968 449900 48980
rect 449952 48968 449958 49020
rect 467742 48968 467748 49020
rect 467800 49008 467806 49020
rect 528554 49008 528560 49020
rect 467800 48980 528560 49008
rect 467800 48968 467806 48980
rect 528554 48968 528560 48980
rect 528612 48968 528618 49020
rect 66070 48764 66076 48816
rect 66128 48804 66134 48816
rect 66898 48804 66904 48816
rect 66128 48776 66904 48804
rect 66128 48764 66134 48776
rect 66898 48764 66904 48776
rect 66956 48764 66962 48816
rect 70854 48764 70860 48816
rect 70912 48804 70918 48816
rect 71682 48804 71688 48816
rect 70912 48776 71688 48804
rect 70912 48764 70918 48776
rect 71682 48764 71688 48776
rect 71740 48764 71746 48816
rect 72050 48764 72056 48816
rect 72108 48804 72114 48816
rect 73062 48804 73068 48816
rect 72108 48776 73068 48804
rect 72108 48764 72114 48776
rect 73062 48764 73068 48776
rect 73120 48764 73126 48816
rect 73246 48764 73252 48816
rect 73304 48804 73310 48816
rect 74442 48804 74448 48816
rect 73304 48776 74448 48804
rect 73304 48764 73310 48776
rect 74442 48764 74448 48776
rect 74500 48764 74506 48816
rect 76834 48764 76840 48816
rect 76892 48804 76898 48816
rect 77938 48804 77944 48816
rect 76892 48776 77944 48804
rect 76892 48764 76898 48776
rect 77938 48764 77944 48776
rect 77996 48764 78002 48816
rect 80422 48764 80428 48816
rect 80480 48804 80486 48816
rect 82078 48804 82084 48816
rect 80480 48776 82084 48804
rect 80480 48764 80486 48776
rect 82078 48764 82084 48776
rect 82136 48764 82142 48816
rect 89898 48764 89904 48816
rect 89956 48804 89962 48816
rect 91002 48804 91008 48816
rect 89956 48776 91008 48804
rect 89956 48764 89962 48776
rect 91002 48764 91008 48776
rect 91060 48764 91066 48816
rect 91094 48764 91100 48816
rect 91152 48804 91158 48816
rect 92290 48804 92296 48816
rect 91152 48776 92296 48804
rect 91152 48764 91158 48776
rect 92290 48764 92296 48776
rect 92348 48764 92354 48816
rect 97074 48764 97080 48816
rect 97132 48804 97138 48816
rect 97902 48804 97908 48816
rect 97132 48776 97908 48804
rect 97132 48764 97138 48776
rect 97902 48764 97908 48776
rect 97960 48764 97966 48816
rect 98270 48764 98276 48816
rect 98328 48804 98334 48816
rect 99282 48804 99288 48816
rect 98328 48776 99288 48804
rect 98328 48764 98334 48776
rect 99282 48764 99288 48776
rect 99340 48764 99346 48816
rect 99466 48764 99472 48816
rect 99524 48804 99530 48816
rect 100662 48804 100668 48816
rect 99524 48776 100668 48804
rect 99524 48764 99530 48776
rect 100662 48764 100668 48776
rect 100720 48764 100726 48816
rect 105446 48764 105452 48816
rect 105504 48804 105510 48816
rect 106182 48804 106188 48816
rect 105504 48776 106188 48804
rect 105504 48764 105510 48776
rect 106182 48764 106188 48776
rect 106240 48764 106246 48816
rect 106642 48764 106648 48816
rect 106700 48804 106706 48816
rect 107562 48804 107568 48816
rect 106700 48776 107568 48804
rect 106700 48764 106706 48776
rect 107562 48764 107568 48776
rect 107620 48764 107626 48816
rect 107838 48764 107844 48816
rect 107896 48804 107902 48816
rect 108942 48804 108948 48816
rect 107896 48776 108948 48804
rect 107896 48764 107902 48776
rect 108942 48764 108948 48776
rect 109000 48764 109006 48816
rect 109034 48764 109040 48816
rect 109092 48804 109098 48816
rect 110230 48804 110236 48816
rect 109092 48776 110236 48804
rect 109092 48764 109098 48776
rect 110230 48764 110236 48776
rect 110288 48764 110294 48816
rect 113726 48764 113732 48816
rect 113784 48804 113790 48816
rect 114462 48804 114468 48816
rect 113784 48776 114468 48804
rect 113784 48764 113790 48776
rect 114462 48764 114468 48776
rect 114520 48764 114526 48816
rect 114922 48764 114928 48816
rect 114980 48804 114986 48816
rect 115842 48804 115848 48816
rect 114980 48776 115848 48804
rect 114980 48764 114986 48776
rect 115842 48764 115848 48776
rect 115900 48764 115906 48816
rect 116118 48764 116124 48816
rect 116176 48804 116182 48816
rect 117222 48804 117228 48816
rect 116176 48776 117228 48804
rect 116176 48764 116182 48776
rect 117222 48764 117228 48776
rect 117280 48764 117286 48816
rect 117314 48764 117320 48816
rect 117372 48804 117378 48816
rect 118602 48804 118608 48816
rect 117372 48776 118608 48804
rect 117372 48764 117378 48776
rect 118602 48764 118608 48776
rect 118660 48764 118666 48816
rect 124490 48764 124496 48816
rect 124548 48804 124554 48816
rect 125502 48804 125508 48816
rect 124548 48776 125508 48804
rect 124548 48764 124554 48776
rect 125502 48764 125508 48776
rect 125560 48764 125566 48816
rect 132862 48764 132868 48816
rect 132920 48804 132926 48816
rect 133782 48804 133788 48816
rect 132920 48776 133788 48804
rect 132920 48764 132926 48776
rect 133782 48764 133788 48776
rect 133840 48764 133846 48816
rect 134058 48764 134064 48816
rect 134116 48804 134122 48816
rect 135162 48804 135168 48816
rect 134116 48776 135168 48804
rect 134116 48764 134122 48776
rect 135162 48764 135168 48776
rect 135220 48764 135226 48816
rect 135254 48764 135260 48816
rect 135312 48804 135318 48816
rect 136450 48804 136456 48816
rect 135312 48776 136456 48804
rect 135312 48764 135318 48776
rect 136450 48764 136456 48776
rect 136508 48764 136514 48816
rect 141142 48764 141148 48816
rect 141200 48804 141206 48816
rect 142062 48804 142068 48816
rect 141200 48776 142068 48804
rect 141200 48764 141206 48776
rect 142062 48764 142068 48776
rect 142120 48764 142126 48816
rect 142338 48764 142344 48816
rect 142396 48804 142402 48816
rect 143442 48804 143448 48816
rect 142396 48776 143448 48804
rect 142396 48764 142402 48776
rect 143442 48764 143448 48776
rect 143500 48764 143506 48816
rect 143534 48764 143540 48816
rect 143592 48804 143598 48816
rect 144822 48804 144828 48816
rect 143592 48776 144828 48804
rect 143592 48764 143598 48776
rect 144822 48764 144828 48776
rect 144880 48764 144886 48816
rect 149514 48764 149520 48816
rect 149572 48804 149578 48816
rect 150342 48804 150348 48816
rect 149572 48776 150348 48804
rect 149572 48764 149578 48776
rect 150342 48764 150348 48776
rect 150400 48764 150406 48816
rect 150710 48764 150716 48816
rect 150768 48804 150774 48816
rect 151722 48804 151728 48816
rect 150768 48776 151728 48804
rect 150768 48764 150774 48776
rect 151722 48764 151728 48776
rect 151780 48764 151786 48816
rect 151906 48764 151912 48816
rect 151964 48804 151970 48816
rect 153838 48804 153844 48816
rect 151964 48776 153844 48804
rect 151964 48764 151970 48776
rect 153838 48764 153844 48776
rect 153896 48764 153902 48816
rect 157886 48764 157892 48816
rect 157944 48804 157950 48816
rect 158622 48804 158628 48816
rect 157944 48776 158628 48804
rect 157944 48764 157950 48776
rect 158622 48764 158628 48776
rect 158680 48764 158686 48816
rect 159082 48764 159088 48816
rect 159140 48804 159146 48816
rect 160002 48804 160008 48816
rect 159140 48776 160008 48804
rect 159140 48764 159146 48776
rect 160002 48764 160008 48776
rect 160060 48764 160066 48816
rect 160278 48764 160284 48816
rect 160336 48804 160342 48816
rect 161382 48804 161388 48816
rect 160336 48776 161388 48804
rect 160336 48764 160342 48776
rect 161382 48764 161388 48776
rect 161440 48764 161446 48816
rect 166166 48764 166172 48816
rect 166224 48804 166230 48816
rect 167730 48804 167736 48816
rect 166224 48776 167736 48804
rect 166224 48764 166230 48776
rect 167730 48764 167736 48776
rect 167788 48764 167794 48816
rect 168558 48764 168564 48816
rect 168616 48804 168622 48816
rect 169662 48804 169668 48816
rect 168616 48776 169668 48804
rect 168616 48764 168622 48776
rect 169662 48764 169668 48776
rect 169720 48764 169726 48816
rect 176930 48764 176936 48816
rect 176988 48804 176994 48816
rect 177942 48804 177948 48816
rect 176988 48776 177948 48804
rect 176988 48764 176994 48776
rect 177942 48764 177948 48776
rect 178000 48764 178006 48816
rect 178126 48764 178132 48816
rect 178184 48804 178190 48816
rect 179322 48804 179328 48816
rect 178184 48776 179328 48804
rect 178184 48764 178190 48776
rect 179322 48764 179328 48776
rect 179380 48764 179386 48816
rect 185302 48764 185308 48816
rect 185360 48804 185366 48816
rect 186222 48804 186228 48816
rect 185360 48776 186228 48804
rect 185360 48764 185366 48776
rect 186222 48764 186228 48776
rect 186280 48764 186286 48816
rect 186498 48764 186504 48816
rect 186556 48804 186562 48816
rect 187602 48804 187608 48816
rect 186556 48776 187608 48804
rect 186556 48764 186562 48776
rect 187602 48764 187608 48776
rect 187660 48764 187666 48816
rect 187694 48764 187700 48816
rect 187752 48804 187758 48816
rect 189718 48804 189724 48816
rect 187752 48776 189724 48804
rect 187752 48764 187758 48776
rect 189718 48764 189724 48776
rect 189776 48764 189782 48816
rect 193582 48764 193588 48816
rect 193640 48804 193646 48816
rect 194502 48804 194508 48816
rect 193640 48776 194508 48804
rect 193640 48764 193646 48776
rect 194502 48764 194508 48776
rect 194560 48764 194566 48816
rect 201954 48764 201960 48816
rect 202012 48804 202018 48816
rect 202782 48804 202788 48816
rect 202012 48776 202788 48804
rect 202012 48764 202018 48776
rect 202782 48764 202788 48776
rect 202840 48764 202846 48816
rect 203150 48764 203156 48816
rect 203208 48804 203214 48816
rect 204162 48804 204168 48816
rect 203208 48776 204168 48804
rect 203208 48764 203214 48776
rect 204162 48764 204168 48776
rect 204220 48764 204226 48816
rect 204346 48764 204352 48816
rect 204404 48804 204410 48816
rect 205542 48804 205548 48816
rect 204404 48776 205548 48804
rect 204404 48764 204410 48776
rect 205542 48764 205548 48776
rect 205600 48764 205606 48816
rect 212718 48764 212724 48816
rect 212776 48804 212782 48816
rect 213822 48804 213828 48816
rect 212776 48776 213828 48804
rect 212776 48764 212782 48776
rect 213822 48764 213828 48776
rect 213880 48764 213886 48816
rect 213914 48764 213920 48816
rect 213972 48804 213978 48816
rect 215202 48804 215208 48816
rect 213972 48776 215208 48804
rect 213972 48764 213978 48776
rect 215202 48764 215208 48776
rect 215260 48764 215266 48816
rect 218606 48764 218612 48816
rect 218664 48804 218670 48816
rect 219342 48804 219348 48816
rect 218664 48776 219348 48804
rect 218664 48764 218670 48776
rect 219342 48764 219348 48776
rect 219400 48764 219406 48816
rect 219802 48764 219808 48816
rect 219860 48804 219866 48816
rect 220722 48804 220728 48816
rect 219860 48776 220728 48804
rect 219860 48764 219866 48776
rect 220722 48764 220728 48776
rect 220780 48764 220786 48816
rect 220998 48764 221004 48816
rect 221056 48804 221062 48816
rect 222102 48804 222108 48816
rect 221056 48776 222108 48804
rect 221056 48764 221062 48776
rect 222102 48764 222108 48776
rect 222160 48764 222166 48816
rect 222194 48764 222200 48816
rect 222252 48804 222258 48816
rect 223482 48804 223488 48816
rect 222252 48776 223488 48804
rect 222252 48764 222258 48776
rect 223482 48764 223488 48776
rect 223540 48764 223546 48816
rect 228174 48764 228180 48816
rect 228232 48804 228238 48816
rect 229002 48804 229008 48816
rect 228232 48776 229008 48804
rect 228232 48764 228238 48776
rect 229002 48764 229008 48776
rect 229060 48764 229066 48816
rect 229370 48764 229376 48816
rect 229428 48804 229434 48816
rect 230382 48804 230388 48816
rect 229428 48776 230388 48804
rect 229428 48764 229434 48776
rect 230382 48764 230388 48776
rect 230440 48764 230446 48816
rect 235350 48764 235356 48816
rect 235408 48804 235414 48816
rect 236638 48804 236644 48816
rect 235408 48776 236644 48804
rect 235408 48764 235414 48776
rect 236638 48764 236644 48776
rect 236696 48764 236702 48816
rect 237742 48764 237748 48816
rect 237800 48804 237806 48816
rect 238662 48804 238668 48816
rect 237800 48776 238668 48804
rect 237800 48764 237806 48776
rect 238662 48764 238668 48776
rect 238720 48764 238726 48816
rect 238938 48764 238944 48816
rect 238996 48804 239002 48816
rect 240042 48804 240048 48816
rect 238996 48776 240048 48804
rect 238996 48764 239002 48776
rect 240042 48764 240048 48776
rect 240100 48764 240106 48816
rect 240134 48764 240140 48816
rect 240192 48804 240198 48816
rect 241422 48804 241428 48816
rect 240192 48776 241428 48804
rect 240192 48764 240198 48776
rect 241422 48764 241428 48776
rect 241480 48764 241486 48816
rect 246022 48764 246028 48816
rect 246080 48804 246086 48816
rect 246942 48804 246948 48816
rect 246080 48776 246948 48804
rect 246080 48764 246086 48776
rect 246942 48764 246948 48776
rect 247000 48764 247006 48816
rect 247218 48764 247224 48816
rect 247276 48804 247282 48816
rect 248322 48804 248328 48816
rect 247276 48776 248328 48804
rect 247276 48764 247282 48776
rect 248322 48764 248328 48776
rect 248380 48764 248386 48816
rect 254394 48764 254400 48816
rect 254452 48804 254458 48816
rect 255222 48804 255228 48816
rect 254452 48776 255228 48804
rect 254452 48764 254458 48776
rect 255222 48764 255228 48776
rect 255280 48764 255286 48816
rect 255590 48764 255596 48816
rect 255648 48804 255654 48816
rect 256602 48804 256608 48816
rect 255648 48776 256608 48804
rect 255648 48764 255654 48776
rect 256602 48764 256608 48776
rect 256660 48764 256666 48816
rect 256786 48764 256792 48816
rect 256844 48804 256850 48816
rect 257982 48804 257988 48816
rect 256844 48776 257988 48804
rect 256844 48764 256850 48776
rect 257982 48764 257988 48776
rect 258040 48764 258046 48816
rect 260374 48764 260380 48816
rect 260432 48804 260438 48816
rect 261478 48804 261484 48816
rect 260432 48776 261484 48804
rect 260432 48764 260438 48776
rect 261478 48764 261484 48776
rect 261536 48764 261542 48816
rect 265158 48764 265164 48816
rect 265216 48804 265222 48816
rect 266262 48804 266268 48816
rect 265216 48776 266268 48804
rect 265216 48764 265222 48776
rect 266262 48764 266268 48776
rect 266320 48764 266326 48816
rect 266354 48764 266360 48816
rect 266412 48804 266418 48816
rect 267550 48804 267556 48816
rect 266412 48776 267556 48804
rect 266412 48764 266418 48776
rect 267550 48764 267556 48776
rect 267608 48764 267614 48816
rect 272242 48764 272248 48816
rect 272300 48804 272306 48816
rect 273162 48804 273168 48816
rect 272300 48776 273168 48804
rect 272300 48764 272306 48776
rect 273162 48764 273168 48776
rect 273220 48764 273226 48816
rect 273438 48764 273444 48816
rect 273496 48804 273502 48816
rect 274542 48804 274548 48816
rect 273496 48776 274548 48804
rect 273496 48764 273502 48776
rect 274542 48764 274548 48776
rect 274600 48764 274606 48816
rect 274634 48764 274640 48816
rect 274692 48804 274698 48816
rect 276658 48804 276664 48816
rect 274692 48776 276664 48804
rect 274692 48764 274698 48776
rect 276658 48764 276664 48776
rect 276716 48764 276722 48816
rect 280614 48764 280620 48816
rect 280672 48804 280678 48816
rect 281442 48804 281448 48816
rect 280672 48776 281448 48804
rect 280672 48764 280678 48776
rect 281442 48764 281448 48776
rect 281500 48764 281506 48816
rect 283006 48764 283012 48816
rect 283064 48804 283070 48816
rect 284202 48804 284208 48816
rect 283064 48776 284208 48804
rect 283064 48764 283070 48776
rect 284202 48764 284208 48776
rect 284260 48764 284266 48816
rect 290182 48764 290188 48816
rect 290240 48804 290246 48816
rect 291102 48804 291108 48816
rect 290240 48776 291108 48804
rect 290240 48764 290246 48776
rect 291102 48764 291108 48776
rect 291160 48764 291166 48816
rect 298462 48764 298468 48816
rect 298520 48804 298526 48816
rect 299382 48804 299388 48816
rect 298520 48776 299388 48804
rect 298520 48764 298526 48776
rect 299382 48764 299388 48776
rect 299440 48764 299446 48816
rect 299658 48764 299664 48816
rect 299716 48804 299722 48816
rect 301498 48804 301504 48816
rect 299716 48776 301504 48804
rect 299716 48764 299722 48776
rect 301498 48764 301504 48776
rect 301556 48764 301562 48816
rect 308030 48764 308036 48816
rect 308088 48804 308094 48816
rect 309042 48804 309048 48816
rect 308088 48776 309048 48804
rect 308088 48764 308094 48776
rect 309042 48764 309048 48776
rect 309100 48764 309106 48816
rect 316402 48764 316408 48816
rect 316460 48804 316466 48816
rect 317322 48804 317328 48816
rect 316460 48776 317328 48804
rect 316460 48764 316466 48776
rect 317322 48764 317328 48776
rect 317380 48764 317386 48816
rect 323486 48764 323492 48816
rect 323544 48804 323550 48816
rect 324222 48804 324228 48816
rect 323544 48776 324228 48804
rect 323544 48764 323550 48776
rect 324222 48764 324228 48776
rect 324280 48764 324286 48816
rect 324682 48764 324688 48816
rect 324740 48804 324746 48816
rect 325602 48804 325608 48816
rect 324740 48776 325608 48804
rect 324740 48764 324746 48776
rect 325602 48764 325608 48776
rect 325660 48764 325666 48816
rect 325878 48764 325884 48816
rect 325936 48804 325942 48816
rect 326982 48804 326988 48816
rect 325936 48776 326988 48804
rect 325936 48764 325942 48776
rect 326982 48764 326988 48776
rect 327040 48764 327046 48816
rect 327074 48764 327080 48816
rect 327132 48804 327138 48816
rect 328270 48804 328276 48816
rect 327132 48776 328276 48804
rect 327132 48764 327138 48776
rect 328270 48764 328276 48776
rect 328328 48764 328334 48816
rect 329466 48764 329472 48816
rect 329524 48804 329530 48816
rect 330478 48804 330484 48816
rect 329524 48776 330484 48804
rect 329524 48764 329530 48776
rect 330478 48764 330484 48776
rect 330536 48764 330542 48816
rect 333054 48764 333060 48816
rect 333112 48804 333118 48816
rect 333882 48804 333888 48816
rect 333112 48776 333888 48804
rect 333112 48764 333118 48776
rect 333882 48764 333888 48776
rect 333940 48764 333946 48816
rect 335446 48764 335452 48816
rect 335504 48804 335510 48816
rect 336642 48804 336648 48816
rect 335504 48776 336648 48804
rect 335504 48764 335510 48776
rect 336642 48764 336648 48776
rect 336700 48764 336706 48816
rect 343726 48764 343732 48816
rect 343784 48804 343790 48816
rect 344922 48804 344928 48816
rect 343784 48776 344928 48804
rect 343784 48764 343790 48776
rect 344922 48764 344928 48776
rect 344980 48764 344986 48816
rect 347314 48764 347320 48816
rect 347372 48804 347378 48816
rect 348418 48804 348424 48816
rect 347372 48776 348424 48804
rect 347372 48764 347378 48776
rect 348418 48764 348424 48776
rect 348476 48764 348482 48816
rect 350902 48764 350908 48816
rect 350960 48804 350966 48816
rect 351822 48804 351828 48816
rect 350960 48776 351828 48804
rect 350960 48764 350966 48776
rect 351822 48764 351828 48776
rect 351880 48764 351886 48816
rect 353294 48764 353300 48816
rect 353352 48804 353358 48816
rect 354582 48804 354588 48816
rect 353352 48776 354588 48804
rect 353352 48764 353358 48776
rect 354582 48764 354588 48776
rect 354640 48764 354646 48816
rect 359274 48764 359280 48816
rect 359332 48804 359338 48816
rect 360102 48804 360108 48816
rect 359332 48776 360108 48804
rect 359332 48764 359338 48776
rect 360102 48764 360108 48776
rect 360160 48764 360166 48816
rect 361666 48764 361672 48816
rect 361724 48804 361730 48816
rect 362862 48804 362868 48816
rect 361724 48776 362868 48804
rect 361724 48764 361730 48776
rect 362862 48764 362868 48776
rect 362920 48764 362926 48816
rect 369946 48764 369952 48816
rect 370004 48804 370010 48816
rect 371050 48804 371056 48816
rect 370004 48776 371056 48804
rect 370004 48764 370010 48776
rect 371050 48764 371056 48776
rect 371108 48764 371114 48816
rect 375926 48764 375932 48816
rect 375984 48804 375990 48816
rect 376662 48804 376668 48816
rect 375984 48776 376668 48804
rect 375984 48764 375990 48776
rect 376662 48764 376668 48776
rect 376720 48764 376726 48816
rect 378318 48764 378324 48816
rect 378376 48804 378382 48816
rect 379422 48804 379428 48816
rect 378376 48776 379428 48804
rect 378376 48764 378382 48776
rect 379422 48764 379428 48776
rect 379480 48764 379486 48816
rect 379514 48764 379520 48816
rect 379572 48804 379578 48816
rect 380802 48804 380808 48816
rect 379572 48776 380808 48804
rect 379572 48764 379578 48776
rect 380802 48764 380808 48776
rect 380860 48764 380866 48816
rect 385494 48764 385500 48816
rect 385552 48804 385558 48816
rect 386322 48804 386328 48816
rect 385552 48776 386328 48804
rect 385552 48764 385558 48776
rect 386322 48764 386328 48776
rect 386380 48764 386386 48816
rect 386690 48764 386696 48816
rect 386748 48804 386754 48816
rect 387702 48804 387708 48816
rect 386748 48776 387708 48804
rect 386748 48764 386754 48776
rect 387702 48764 387708 48776
rect 387760 48764 387766 48816
rect 387886 48764 387892 48816
rect 387944 48804 387950 48816
rect 389082 48804 389088 48816
rect 387944 48776 389088 48804
rect 387944 48764 387950 48776
rect 389082 48764 389088 48776
rect 389140 48764 389146 48816
rect 394970 48764 394976 48816
rect 395028 48804 395034 48816
rect 395982 48804 395988 48816
rect 395028 48776 395988 48804
rect 395028 48764 395034 48776
rect 395982 48764 395988 48776
rect 396040 48764 396046 48816
rect 404538 48764 404544 48816
rect 404596 48804 404602 48816
rect 405642 48804 405648 48816
rect 404596 48776 405648 48804
rect 404596 48764 404602 48776
rect 405642 48764 405648 48776
rect 405700 48764 405706 48816
rect 412910 48764 412916 48816
rect 412968 48804 412974 48816
rect 413922 48804 413928 48816
rect 412968 48776 413928 48804
rect 412968 48764 412974 48776
rect 413922 48764 413928 48776
rect 413980 48764 413986 48816
rect 414106 48764 414112 48816
rect 414164 48804 414170 48816
rect 415302 48804 415308 48816
rect 414164 48776 415308 48804
rect 414164 48764 414170 48776
rect 415302 48764 415308 48776
rect 415360 48764 415366 48816
rect 420086 48764 420092 48816
rect 420144 48804 420150 48816
rect 420822 48804 420828 48816
rect 420144 48776 420828 48804
rect 420144 48764 420150 48776
rect 420822 48764 420828 48776
rect 420880 48764 420886 48816
rect 421190 48764 421196 48816
rect 421248 48804 421254 48816
rect 422202 48804 422208 48816
rect 421248 48776 422208 48804
rect 421248 48764 421254 48776
rect 422202 48764 422208 48776
rect 422260 48764 422266 48816
rect 422386 48764 422392 48816
rect 422444 48804 422450 48816
rect 423582 48804 423588 48816
rect 422444 48776 423588 48804
rect 422444 48764 422450 48776
rect 423582 48764 423588 48776
rect 423640 48764 423646 48816
rect 428366 48764 428372 48816
rect 428424 48804 428430 48816
rect 429102 48804 429108 48816
rect 428424 48776 429108 48804
rect 428424 48764 428430 48776
rect 429102 48764 429108 48776
rect 429160 48764 429166 48816
rect 429562 48764 429568 48816
rect 429620 48804 429626 48816
rect 430482 48804 430488 48816
rect 429620 48776 430488 48804
rect 429620 48764 429626 48776
rect 430482 48764 430488 48776
rect 430540 48764 430546 48816
rect 430758 48764 430764 48816
rect 430816 48804 430822 48816
rect 431862 48804 431868 48816
rect 430816 48776 431868 48804
rect 430816 48764 430822 48776
rect 431862 48764 431868 48776
rect 431920 48764 431926 48816
rect 433150 48764 433156 48816
rect 433208 48804 433214 48816
rect 433978 48804 433984 48816
rect 433208 48776 433984 48804
rect 433208 48764 433214 48776
rect 433978 48764 433984 48776
rect 434036 48764 434042 48816
rect 437934 48764 437940 48816
rect 437992 48804 437998 48816
rect 438762 48804 438768 48816
rect 437992 48776 438768 48804
rect 437992 48764 437998 48776
rect 438762 48764 438768 48776
rect 438820 48764 438826 48816
rect 439130 48764 439136 48816
rect 439188 48804 439194 48816
rect 440142 48804 440148 48816
rect 439188 48776 440148 48804
rect 439188 48764 439194 48776
rect 440142 48764 440148 48776
rect 440200 48764 440206 48816
rect 446214 48764 446220 48816
rect 446272 48804 446278 48816
rect 447042 48804 447048 48816
rect 446272 48776 447048 48804
rect 446272 48764 446278 48776
rect 447042 48764 447048 48776
rect 447100 48764 447106 48816
rect 447410 48764 447416 48816
rect 447468 48804 447474 48816
rect 448422 48804 448428 48816
rect 447468 48776 448428 48804
rect 447468 48764 447474 48776
rect 448422 48764 448428 48776
rect 448480 48764 448486 48816
rect 448606 48764 448612 48816
rect 448664 48804 448670 48816
rect 449710 48804 449716 48816
rect 448664 48776 449716 48804
rect 448664 48764 448670 48776
rect 449710 48764 449716 48776
rect 449768 48764 449774 48816
rect 455782 48764 455788 48816
rect 455840 48804 455846 48816
rect 456702 48804 456708 48816
rect 455840 48776 456708 48804
rect 455840 48764 455846 48776
rect 456702 48764 456708 48776
rect 456760 48764 456766 48816
rect 456978 48764 456984 48816
rect 457036 48804 457042 48816
rect 458082 48804 458088 48816
rect 457036 48776 458088 48804
rect 457036 48764 457042 48776
rect 458082 48764 458088 48776
rect 458140 48764 458146 48816
rect 459370 48764 459376 48816
rect 459428 48804 459434 48816
rect 460198 48804 460204 48816
rect 459428 48776 460204 48804
rect 459428 48764 459434 48776
rect 460198 48764 460204 48776
rect 460256 48764 460262 48816
rect 464154 48764 464160 48816
rect 464212 48804 464218 48816
rect 464982 48804 464988 48816
rect 464212 48776 464988 48804
rect 464212 48764 464218 48776
rect 464982 48764 464988 48776
rect 465040 48764 465046 48816
rect 465350 48764 465356 48816
rect 465408 48804 465414 48816
rect 466362 48804 466368 48816
rect 465408 48776 466368 48804
rect 465408 48764 465414 48776
rect 466362 48764 466368 48776
rect 466420 48764 466426 48816
rect 466546 48764 466552 48816
rect 466604 48804 466610 48816
rect 467742 48804 467748 48816
rect 466604 48776 467748 48804
rect 466604 48764 466610 48776
rect 467742 48764 467748 48776
rect 467800 48764 467806 48816
rect 473630 48764 473636 48816
rect 473688 48804 473694 48816
rect 474642 48804 474648 48816
rect 473688 48776 474648 48804
rect 473688 48764 473694 48776
rect 474642 48764 474648 48776
rect 474700 48764 474706 48816
rect 480806 48764 480812 48816
rect 480864 48804 480870 48816
rect 481542 48804 481548 48816
rect 480864 48776 481548 48804
rect 480864 48764 480870 48776
rect 481542 48764 481548 48776
rect 481600 48764 481606 48816
rect 483198 48764 483204 48816
rect 483256 48804 483262 48816
rect 484302 48804 484308 48816
rect 483256 48776 484308 48804
rect 483256 48764 483262 48776
rect 484302 48764 484308 48776
rect 484360 48764 484366 48816
rect 484394 48764 484400 48816
rect 484452 48804 484458 48816
rect 485590 48804 485596 48816
rect 484452 48776 485596 48804
rect 484452 48764 484458 48776
rect 485590 48764 485596 48776
rect 485648 48764 485654 48816
rect 491570 48764 491576 48816
rect 491628 48804 491634 48816
rect 492582 48804 492588 48816
rect 491628 48776 492588 48804
rect 491628 48764 491634 48776
rect 492582 48764 492588 48776
rect 492640 48764 492646 48816
rect 492766 48764 492772 48816
rect 492824 48804 492830 48816
rect 493962 48804 493968 48816
rect 492824 48776 493968 48804
rect 492824 48764 492830 48776
rect 493962 48764 493968 48776
rect 494020 48764 494026 48816
rect 495158 48764 495164 48816
rect 495216 48804 495222 48816
rect 496078 48804 496084 48816
rect 495216 48776 496084 48804
rect 495216 48764 495222 48776
rect 496078 48764 496084 48776
rect 496136 48764 496142 48816
rect 498654 48764 498660 48816
rect 498712 48804 498718 48816
rect 499482 48804 499488 48816
rect 498712 48776 499488 48804
rect 498712 48764 498718 48776
rect 499482 48764 499488 48776
rect 499540 48764 499546 48816
rect 499850 48764 499856 48816
rect 499908 48804 499914 48816
rect 500862 48804 500868 48816
rect 499908 48776 500868 48804
rect 499908 48764 499914 48776
rect 500862 48764 500868 48776
rect 500920 48764 500926 48816
rect 501046 48764 501052 48816
rect 501104 48804 501110 48816
rect 502242 48804 502248 48816
rect 501104 48776 502248 48804
rect 501104 48764 501110 48776
rect 502242 48764 502248 48776
rect 502300 48764 502306 48816
rect 508222 48764 508228 48816
rect 508280 48804 508286 48816
rect 509142 48804 509148 48816
rect 508280 48776 509148 48804
rect 508280 48764 508286 48776
rect 509142 48764 509148 48776
rect 509200 48764 509206 48816
rect 509418 48764 509424 48816
rect 509476 48804 509482 48816
rect 510522 48804 510528 48816
rect 509476 48776 510528 48804
rect 509476 48764 509482 48776
rect 510522 48764 510528 48776
rect 510580 48764 510586 48816
rect 516594 48764 516600 48816
rect 516652 48804 516658 48816
rect 517422 48804 517428 48816
rect 516652 48776 517428 48804
rect 516652 48764 516658 48776
rect 517422 48764 517428 48776
rect 517480 48764 517486 48816
rect 517790 48764 517796 48816
rect 517848 48804 517854 48816
rect 518802 48804 518808 48816
rect 517848 48776 518808 48804
rect 517848 48764 517854 48776
rect 518802 48764 518808 48776
rect 518860 48764 518866 48816
rect 518986 48764 518992 48816
rect 519044 48804 519050 48816
rect 520090 48804 520096 48816
rect 519044 48776 520096 48804
rect 519044 48764 519050 48776
rect 520090 48764 520096 48776
rect 520148 48764 520154 48816
rect 64874 48696 64880 48748
rect 64932 48736 64938 48748
rect 66162 48736 66168 48748
rect 64932 48708 66168 48736
rect 64932 48696 64938 48708
rect 66162 48696 66168 48708
rect 66220 48696 66226 48748
rect 123294 48696 123300 48748
rect 123352 48736 123358 48748
rect 124122 48736 124128 48748
rect 123352 48708 124128 48736
rect 123352 48696 123358 48708
rect 124122 48696 124128 48708
rect 124180 48696 124186 48748
rect 161474 48696 161480 48748
rect 161532 48736 161538 48748
rect 167638 48736 167644 48748
rect 161532 48708 167644 48736
rect 161532 48696 161538 48708
rect 167638 48696 167644 48708
rect 167696 48696 167702 48748
rect 262766 48696 262772 48748
rect 262824 48736 262830 48748
rect 263502 48736 263508 48748
rect 262824 48708 263508 48736
rect 262824 48696 262830 48708
rect 263502 48696 263508 48708
rect 263560 48696 263566 48748
rect 263962 48696 263968 48748
rect 264020 48736 264026 48748
rect 265618 48736 265624 48748
rect 264020 48708 265624 48736
rect 264020 48696 264026 48708
rect 265618 48696 265624 48708
rect 265676 48696 265682 48748
rect 271046 48696 271052 48748
rect 271104 48736 271110 48748
rect 272518 48736 272524 48748
rect 271104 48708 272524 48736
rect 271104 48696 271110 48708
rect 272518 48696 272524 48708
rect 272576 48696 272582 48748
rect 288986 48696 288992 48748
rect 289044 48736 289050 48748
rect 290458 48736 290464 48748
rect 289044 48708 290464 48736
rect 289044 48696 289050 48708
rect 290458 48696 290464 48708
rect 290516 48696 290522 48748
rect 306834 48696 306840 48748
rect 306892 48736 306898 48748
rect 312538 48736 312544 48748
rect 306892 48708 312544 48736
rect 306892 48696 306898 48708
rect 312538 48696 312544 48708
rect 312596 48696 312602 48748
rect 334250 48696 334256 48748
rect 334308 48736 334314 48748
rect 335262 48736 335268 48748
rect 334308 48708 335268 48736
rect 334308 48696 334314 48708
rect 335262 48696 335268 48708
rect 335320 48696 335326 48748
rect 360470 48696 360476 48748
rect 360528 48736 360534 48748
rect 361482 48736 361488 48748
rect 360528 48708 361488 48736
rect 360528 48696 360534 48708
rect 361482 48696 361488 48708
rect 361540 48696 361546 48748
rect 431954 48696 431960 48748
rect 432012 48736 432018 48748
rect 433242 48736 433248 48748
rect 432012 48708 433248 48736
rect 432012 48696 432018 48708
rect 433242 48696 433248 48708
rect 433300 48696 433306 48748
rect 436738 48696 436744 48748
rect 436796 48736 436802 48748
rect 438118 48736 438124 48748
rect 436796 48708 438124 48736
rect 436796 48696 436802 48708
rect 438118 48696 438124 48708
rect 438176 48696 438182 48748
rect 458174 48696 458180 48748
rect 458232 48736 458238 48748
rect 459462 48736 459468 48748
rect 458232 48708 459468 48736
rect 458232 48696 458238 48708
rect 459462 48696 459468 48708
rect 459520 48696 459526 48748
rect 472434 48696 472440 48748
rect 472492 48736 472498 48748
rect 473998 48736 474004 48748
rect 472492 48708 474004 48736
rect 472492 48696 472498 48708
rect 473998 48696 474004 48708
rect 474056 48696 474062 48748
rect 487982 48696 487988 48748
rect 488040 48736 488046 48748
rect 489178 48736 489184 48748
rect 488040 48708 489184 48736
rect 488040 48696 488046 48708
rect 489178 48696 489184 48708
rect 489236 48696 489242 48748
rect 125686 48628 125692 48680
rect 125744 48668 125750 48680
rect 126790 48668 126796 48680
rect 125744 48640 126796 48668
rect 125744 48628 125750 48640
rect 126790 48628 126796 48640
rect 126848 48628 126854 48680
rect 195974 48628 195980 48680
rect 196032 48668 196038 48680
rect 197262 48668 197268 48680
rect 196032 48640 197268 48668
rect 196032 48628 196038 48640
rect 197262 48628 197268 48640
rect 197320 48628 197326 48680
rect 278222 48628 278228 48680
rect 278280 48668 278286 48680
rect 280798 48668 280804 48680
rect 278280 48640 280804 48668
rect 278280 48628 278286 48640
rect 280798 48628 280804 48640
rect 280856 48628 280862 48680
rect 292574 48628 292580 48680
rect 292632 48668 292638 48680
rect 293862 48668 293868 48680
rect 292632 48640 293868 48668
rect 292632 48628 292638 48640
rect 293862 48628 293868 48640
rect 293920 48628 293926 48680
rect 365254 48628 365260 48680
rect 365312 48668 365318 48680
rect 367738 48668 367744 48680
rect 365312 48640 367744 48668
rect 365312 48628 365318 48640
rect 367738 48628 367744 48640
rect 367796 48628 367802 48680
rect 175734 48560 175740 48612
rect 175792 48600 175798 48612
rect 176562 48600 176568 48612
rect 175792 48572 176568 48600
rect 175792 48560 175798 48572
rect 176562 48560 176568 48572
rect 176620 48560 176626 48612
rect 315206 48560 315212 48612
rect 315264 48600 315270 48612
rect 315942 48600 315948 48612
rect 315264 48572 315948 48600
rect 315264 48560 315270 48572
rect 315942 48560 315948 48572
rect 316000 48560 316006 48612
rect 248414 48492 248420 48544
rect 248472 48532 248478 48544
rect 249610 48532 249616 48544
rect 248472 48504 249616 48532
rect 248472 48492 248478 48504
rect 249610 48492 249616 48504
rect 249668 48492 249674 48544
rect 300854 48492 300860 48544
rect 300912 48532 300918 48544
rect 302142 48532 302148 48544
rect 300912 48504 302148 48532
rect 300912 48492 300918 48504
rect 302142 48492 302148 48504
rect 302200 48492 302206 48544
rect 342622 48492 342628 48544
rect 342680 48532 342686 48544
rect 343542 48532 343548 48544
rect 342680 48504 343548 48532
rect 342680 48492 342686 48504
rect 343542 48492 343548 48504
rect 343600 48492 343606 48544
rect 510614 48492 510620 48544
rect 510672 48532 510678 48544
rect 511902 48532 511908 48544
rect 510672 48504 511908 48532
rect 510672 48492 510678 48504
rect 511902 48492 511908 48504
rect 511960 48492 511966 48544
rect 352098 48424 352104 48476
rect 352156 48464 352162 48476
rect 353202 48464 353208 48476
rect 352156 48436 353208 48464
rect 352156 48424 352162 48436
rect 353202 48424 353208 48436
rect 353260 48424 353266 48476
rect 411714 48424 411720 48476
rect 411772 48464 411778 48476
rect 412542 48464 412548 48476
rect 411772 48436 412548 48464
rect 411772 48424 411778 48436
rect 412542 48424 412548 48436
rect 412600 48424 412606 48476
rect 293678 48356 293684 48408
rect 293736 48396 293742 48408
rect 294598 48396 294604 48408
rect 293736 48368 294604 48396
rect 293736 48356 293742 48368
rect 294598 48356 294604 48368
rect 294656 48356 294662 48408
rect 211522 48288 211528 48340
rect 211580 48328 211586 48340
rect 212442 48328 212448 48340
rect 211580 48300 212448 48328
rect 211580 48288 211586 48300
rect 212442 48288 212448 48300
rect 212500 48288 212506 48340
rect 278958 48328 278964 48340
rect 278919 48300 278964 48328
rect 278958 48288 278964 48300
rect 279016 48288 279022 48340
rect 317598 48288 317604 48340
rect 317656 48328 317662 48340
rect 318702 48328 318708 48340
rect 317656 48300 318708 48328
rect 317656 48288 317662 48300
rect 318702 48288 318708 48300
rect 318760 48288 318766 48340
rect 368842 48288 368848 48340
rect 368900 48328 368906 48340
rect 369762 48328 369768 48340
rect 368900 48300 369768 48328
rect 368900 48288 368906 48300
rect 369762 48288 369768 48300
rect 369820 48288 369826 48340
rect 377122 48288 377128 48340
rect 377180 48328 377186 48340
rect 378042 48328 378048 48340
rect 377180 48300 378048 48328
rect 377180 48288 377186 48300
rect 378042 48288 378048 48300
rect 378100 48288 378106 48340
rect 427906 48328 427912 48340
rect 427867 48300 427912 48328
rect 427906 48288 427912 48300
rect 427964 48288 427970 48340
rect 434806 48328 434812 48340
rect 434767 48300 434812 48328
rect 434806 48288 434812 48300
rect 434864 48288 434870 48340
rect 194778 47676 194784 47728
rect 194836 47716 194842 47728
rect 255314 47716 255320 47728
rect 194836 47688 255320 47716
rect 194836 47676 194842 47688
rect 255314 47676 255320 47688
rect 255372 47676 255378 47728
rect 136542 47608 136548 47660
rect 136600 47648 136606 47660
rect 197354 47648 197360 47660
rect 136600 47620 197360 47648
rect 136600 47608 136606 47620
rect 197354 47608 197360 47620
rect 197412 47608 197418 47660
rect 275830 47608 275836 47660
rect 275888 47648 275894 47660
rect 336734 47648 336740 47660
rect 275888 47620 336740 47648
rect 275888 47608 275894 47620
rect 336734 47608 336740 47620
rect 336792 47608 336798 47660
rect 94682 47540 94688 47592
rect 94740 47580 94746 47592
rect 155954 47580 155960 47592
rect 94740 47552 155960 47580
rect 94740 47540 94746 47552
rect 155954 47540 155960 47552
rect 156012 47540 156018 47592
rect 242434 47540 242440 47592
rect 242492 47580 242498 47592
rect 303614 47580 303620 47592
rect 242492 47552 303620 47580
rect 242492 47540 242498 47552
rect 303614 47540 303620 47552
rect 303672 47540 303678 47592
rect 336826 47540 336832 47592
rect 336884 47580 336890 47592
rect 397454 47580 397460 47592
rect 336884 47552 397460 47580
rect 336884 47540 336890 47552
rect 397454 47540 397460 47552
rect 397512 47540 397518 47592
rect 425974 47540 425980 47592
rect 426032 47580 426038 47592
rect 485774 47580 485780 47592
rect 426032 47552 485780 47580
rect 426032 47540 426038 47552
rect 485774 47540 485780 47552
rect 485832 47540 485838 47592
rect 490374 47540 490380 47592
rect 490432 47580 490438 47592
rect 550634 47580 550640 47592
rect 490432 47552 550640 47580
rect 490432 47540 490438 47552
rect 550634 47540 550640 47552
rect 550692 47540 550698 47592
rect 285766 46900 285772 46912
rect 285727 46872 285772 46900
rect 285766 46860 285772 46872
rect 285824 46860 285830 46912
rect 172330 46248 172336 46300
rect 172388 46288 172394 46300
rect 230474 46288 230480 46300
rect 172388 46260 230480 46288
rect 172388 46248 172394 46260
rect 230474 46248 230480 46260
rect 230532 46248 230538 46300
rect 291378 46248 291384 46300
rect 291436 46288 291442 46300
rect 351914 46288 351920 46300
rect 291436 46260 351920 46288
rect 291436 46248 291442 46260
rect 351914 46248 351920 46260
rect 351972 46248 351978 46300
rect 443914 46248 443920 46300
rect 443972 46288 443978 46300
rect 503714 46288 503720 46300
rect 443972 46260 503720 46288
rect 443972 46248 443978 46260
rect 503714 46248 503720 46260
rect 503772 46248 503778 46300
rect 112622 46180 112628 46232
rect 112680 46220 112686 46232
rect 173894 46220 173900 46232
rect 112680 46192 173900 46220
rect 112680 46180 112686 46192
rect 173894 46180 173900 46192
rect 173952 46180 173958 46232
rect 230566 46180 230572 46232
rect 230624 46220 230630 46232
rect 291194 46220 291200 46232
rect 230624 46192 291200 46220
rect 230624 46180 230630 46192
rect 291194 46180 291200 46192
rect 291252 46180 291258 46232
rect 344830 46180 344836 46232
rect 344888 46220 344894 46232
rect 405734 46220 405740 46232
rect 344888 46192 405740 46220
rect 344888 46180 344894 46192
rect 405734 46180 405740 46192
rect 405792 46180 405798 46232
rect 406010 46180 406016 46232
rect 406068 46220 406074 46232
rect 466454 46220 466460 46232
rect 406068 46192 466460 46220
rect 406068 46180 406074 46192
rect 466454 46180 466460 46192
rect 466512 46180 466518 46232
rect 504634 46180 504640 46232
rect 504692 46220 504698 46232
rect 564434 46220 564440 46232
rect 504692 46192 564440 46220
rect 504692 46180 504698 46192
rect 564434 46180 564440 46192
rect 564492 46180 564498 46232
rect 238662 44888 238668 44940
rect 238720 44928 238726 44940
rect 298094 44928 298100 44940
rect 238720 44900 298100 44928
rect 238720 44888 238726 44900
rect 298094 44888 298100 44900
rect 298152 44888 298158 44940
rect 349062 44888 349068 44940
rect 349120 44928 349126 44940
rect 408494 44928 408500 44940
rect 349120 44900 408500 44928
rect 349120 44888 349126 44900
rect 408494 44888 408500 44900
rect 408552 44888 408558 44940
rect 117222 44820 117228 44872
rect 117280 44860 117286 44872
rect 176654 44860 176660 44872
rect 117280 44832 176660 44860
rect 117280 44820 117286 44832
rect 176654 44820 176660 44832
rect 176712 44820 176718 44872
rect 177942 44820 177948 44872
rect 178000 44860 178006 44872
rect 237374 44860 237380 44872
rect 178000 44832 237380 44860
rect 178000 44820 178006 44832
rect 237374 44820 237380 44832
rect 237432 44820 237438 44872
rect 295242 44820 295248 44872
rect 295300 44860 295306 44872
rect 356054 44860 356060 44872
rect 295300 44832 356060 44860
rect 295300 44820 295306 44832
rect 356054 44820 356060 44832
rect 356112 44820 356118 44872
rect 415210 44820 415216 44872
rect 415268 44860 415274 44872
rect 476114 44860 476120 44872
rect 415268 44832 476120 44860
rect 415268 44820 415274 44832
rect 476114 44820 476120 44832
rect 476172 44820 476178 44872
rect 480162 44820 480168 44872
rect 480220 44860 480226 44872
rect 539594 44860 539600 44872
rect 480220 44832 539600 44860
rect 480220 44820 480226 44832
rect 539594 44820 539600 44832
rect 539652 44820 539658 44872
rect 135162 43460 135168 43512
rect 135220 43500 135226 43512
rect 194594 43500 194600 43512
rect 135220 43472 194600 43500
rect 135220 43460 135226 43472
rect 194594 43460 194600 43472
rect 194652 43460 194658 43512
rect 249610 43460 249616 43512
rect 249668 43500 249674 43512
rect 309134 43500 309140 43512
rect 249668 43472 309140 43500
rect 249668 43460 249674 43472
rect 309134 43460 309140 43472
rect 309192 43460 309198 43512
rect 355962 43460 355968 43512
rect 356020 43500 356026 43512
rect 416866 43500 416872 43512
rect 356020 43472 416872 43500
rect 356020 43460 356026 43472
rect 416866 43460 416872 43472
rect 416924 43460 416930 43512
rect 191742 43392 191748 43444
rect 191800 43432 191806 43444
rect 252646 43432 252652 43444
rect 191800 43404 252652 43432
rect 191800 43392 191806 43404
rect 252646 43392 252652 43404
rect 252704 43392 252710 43444
rect 302050 43392 302056 43444
rect 302108 43432 302114 43444
rect 362954 43432 362960 43444
rect 302108 43404 362960 43432
rect 302108 43392 302114 43404
rect 362954 43392 362960 43404
rect 363012 43392 363018 43444
rect 402882 43392 402888 43444
rect 402940 43432 402946 43444
rect 462314 43432 462320 43444
rect 402940 43404 462320 43432
rect 402940 43392 402946 43404
rect 462314 43392 462320 43404
rect 462372 43392 462378 43444
rect 493870 43392 493876 43444
rect 493928 43432 493934 43444
rect 554774 43432 554780 43444
rect 493928 43404 554780 43432
rect 493928 43392 493934 43404
rect 554774 43392 554780 43404
rect 554832 43392 554838 43444
rect 202782 42100 202788 42152
rect 202840 42140 202846 42152
rect 262214 42140 262220 42152
rect 202840 42112 262220 42140
rect 202840 42100 202846 42112
rect 262214 42100 262220 42112
rect 262272 42100 262278 42152
rect 263502 42100 263508 42152
rect 263560 42140 263566 42152
rect 322934 42140 322940 42152
rect 263560 42112 322940 42140
rect 263560 42100 263566 42112
rect 322934 42100 322940 42112
rect 322992 42100 322998 42152
rect 84102 42032 84108 42084
rect 84160 42072 84166 42084
rect 144914 42072 144920 42084
rect 84160 42044 144920 42072
rect 84160 42032 84166 42044
rect 144914 42032 144920 42044
rect 144972 42032 144978 42084
rect 148962 42032 148968 42084
rect 149020 42072 149026 42084
rect 209866 42072 209872 42084
rect 149020 42044 209872 42072
rect 149020 42032 149026 42044
rect 209866 42032 209872 42044
rect 209924 42032 209930 42084
rect 320082 42032 320088 42084
rect 320140 42072 320146 42084
rect 380894 42072 380900 42084
rect 320140 42044 380900 42072
rect 320140 42032 320146 42044
rect 380894 42032 380900 42044
rect 380952 42032 380958 42084
rect 419442 42032 419448 42084
rect 419500 42072 419506 42084
rect 478874 42072 478880 42084
rect 419500 42044 478880 42072
rect 419500 42032 419506 42044
rect 478874 42032 478880 42044
rect 478932 42032 478938 42084
rect 498102 42032 498108 42084
rect 498160 42072 498166 42084
rect 557534 42072 557540 42084
rect 498160 42044 557540 42072
rect 498160 42032 498166 42044
rect 557534 42032 557540 42044
rect 557592 42032 557598 42084
rect 523678 41352 523684 41404
rect 523736 41392 523742 41404
rect 580166 41392 580172 41404
rect 523736 41364 580172 41392
rect 523736 41352 523742 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 220722 40740 220728 40792
rect 220780 40780 220786 40792
rect 280154 40780 280160 40792
rect 220780 40752 280160 40780
rect 220780 40740 220786 40752
rect 280154 40740 280160 40752
rect 280212 40740 280218 40792
rect 331122 40740 331128 40792
rect 331180 40780 331186 40792
rect 390554 40780 390560 40792
rect 331180 40752 390560 40780
rect 331180 40740 331186 40752
rect 390554 40740 390560 40752
rect 390612 40740 390618 40792
rect 88242 40672 88248 40724
rect 88300 40712 88306 40724
rect 149054 40712 149060 40724
rect 88300 40684 149060 40712
rect 88300 40672 88306 40684
rect 149054 40672 149060 40684
rect 149112 40672 149118 40724
rect 162762 40672 162768 40724
rect 162820 40712 162826 40724
rect 223574 40712 223580 40724
rect 162820 40684 223580 40712
rect 162820 40672 162826 40684
rect 223574 40672 223580 40684
rect 223632 40672 223638 40724
rect 277302 40672 277308 40724
rect 277360 40712 277366 40724
rect 338114 40712 338120 40724
rect 277360 40684 338120 40712
rect 277360 40672 277366 40684
rect 338114 40672 338120 40684
rect 338172 40672 338178 40724
rect 391842 40672 391848 40724
rect 391900 40712 391906 40724
rect 451274 40712 451280 40724
rect 391900 40684 451280 40712
rect 391900 40672 391906 40684
rect 451274 40672 451280 40684
rect 451332 40672 451338 40724
rect 274542 39380 274548 39432
rect 274600 39420 274606 39432
rect 333974 39420 333980 39432
rect 274600 39392 333980 39420
rect 274600 39380 274606 39392
rect 333974 39380 333980 39392
rect 334032 39380 334038 39432
rect 384942 39380 384948 39432
rect 385000 39420 385006 39432
rect 444374 39420 444380 39432
rect 385000 39392 444380 39420
rect 385000 39380 385006 39392
rect 444374 39380 444380 39392
rect 444432 39380 444438 39432
rect 82078 39312 82084 39364
rect 82136 39352 82142 39364
rect 140774 39352 140780 39364
rect 82136 39324 140780 39352
rect 82136 39312 82142 39324
rect 140774 39312 140780 39324
rect 140832 39312 140838 39364
rect 153838 39312 153844 39364
rect 153896 39352 153902 39364
rect 212534 39352 212540 39364
rect 153896 39324 212540 39352
rect 153896 39312 153902 39324
rect 212534 39312 212540 39324
rect 212592 39312 212598 39364
rect 213822 39312 213828 39364
rect 213880 39352 213886 39364
rect 273254 39352 273260 39364
rect 213880 39324 273260 39352
rect 213880 39312 213886 39324
rect 273254 39312 273260 39324
rect 273312 39312 273318 39364
rect 328270 39312 328276 39364
rect 328328 39352 328334 39364
rect 387794 39352 387800 39364
rect 328328 39324 387800 39352
rect 328328 39312 328334 39324
rect 387794 39312 387800 39324
rect 387852 39312 387858 39364
rect 420822 39312 420828 39364
rect 420880 39352 420886 39364
rect 480254 39352 480260 39364
rect 420880 39324 480260 39352
rect 420880 39312 420886 39324
rect 480254 39312 480260 39324
rect 480312 39312 480318 39364
rect 509142 39312 509148 39364
rect 509200 39352 509206 39364
rect 568574 39352 568580 39364
rect 509200 39324 568580 39352
rect 509200 39312 509206 39324
rect 568574 39312 568580 39324
rect 568632 39312 568638 39364
rect 427906 38604 427912 38616
rect 427867 38576 427912 38604
rect 427906 38564 427912 38576
rect 427964 38564 427970 38616
rect 434806 38604 434812 38616
rect 434767 38576 434812 38604
rect 434806 38564 434812 38576
rect 434864 38564 434870 38616
rect 142062 37952 142068 38004
rect 142120 37992 142126 38004
rect 201494 37992 201500 38004
rect 142120 37964 201500 37992
rect 142120 37952 142126 37964
rect 201494 37952 201500 37964
rect 201552 37952 201558 38004
rect 256602 37952 256608 38004
rect 256660 37992 256666 38004
rect 316034 37992 316040 38004
rect 256660 37964 316040 37992
rect 256660 37952 256666 37964
rect 316034 37952 316040 37964
rect 316092 37952 316098 38004
rect 413922 37952 413928 38004
rect 413980 37992 413986 38004
rect 473354 37992 473360 38004
rect 413980 37964 473360 37992
rect 413980 37952 413986 37964
rect 473354 37952 473360 37964
rect 473412 37952 473418 38004
rect 77938 37884 77944 37936
rect 77996 37924 78002 37936
rect 138014 37924 138020 37936
rect 77996 37896 138020 37924
rect 77996 37884 78002 37896
rect 138014 37884 138020 37896
rect 138072 37884 138078 37936
rect 198642 37884 198648 37936
rect 198700 37924 198706 37936
rect 259454 37924 259460 37936
rect 198700 37896 259460 37924
rect 198700 37884 198706 37896
rect 259454 37884 259460 37896
rect 259512 37884 259518 37936
rect 313182 37884 313188 37936
rect 313240 37924 313246 37936
rect 374086 37924 374092 37936
rect 313240 37896 374092 37924
rect 313240 37884 313246 37896
rect 374086 37884 374092 37896
rect 374144 37884 374150 37936
rect 380710 37884 380716 37936
rect 380768 37924 380774 37936
rect 441614 37924 441620 37936
rect 380768 37896 441620 37924
rect 380768 37884 380774 37896
rect 441614 37884 441620 37896
rect 441672 37884 441678 37936
rect 511810 37884 511816 37936
rect 511868 37924 511874 37936
rect 571426 37924 571432 37936
rect 511868 37896 571432 37924
rect 511868 37884 511874 37896
rect 571426 37884 571432 37896
rect 571484 37884 571490 37936
rect 285766 37312 285772 37324
rect 285727 37284 285772 37312
rect 285766 37272 285772 37284
rect 285824 37272 285830 37324
rect 353202 36660 353208 36712
rect 353260 36700 353266 36712
rect 412634 36700 412640 36712
rect 353260 36672 412640 36700
rect 353260 36660 353266 36672
rect 412634 36660 412640 36672
rect 412692 36660 412698 36712
rect 189718 36592 189724 36644
rect 189776 36632 189782 36644
rect 248414 36632 248420 36644
rect 189776 36604 248420 36632
rect 189776 36592 189782 36604
rect 248414 36592 248420 36604
rect 248472 36592 248478 36644
rect 299382 36592 299388 36644
rect 299440 36632 299446 36644
rect 358814 36632 358820 36644
rect 299440 36604 358820 36632
rect 299440 36592 299446 36604
rect 358814 36592 358820 36604
rect 358872 36592 358878 36644
rect 137922 36524 137928 36576
rect 137980 36564 137986 36576
rect 198734 36564 198740 36576
rect 137980 36536 198740 36564
rect 137980 36524 137986 36536
rect 198734 36524 198740 36536
rect 198792 36524 198798 36576
rect 245562 36524 245568 36576
rect 245620 36564 245626 36576
rect 304994 36564 305000 36576
rect 245620 36536 305000 36564
rect 245620 36524 245626 36536
rect 304994 36524 305000 36536
rect 305052 36524 305058 36576
rect 398742 36524 398748 36576
rect 398800 36564 398806 36576
rect 459646 36564 459652 36576
rect 398800 36536 459652 36564
rect 398800 36524 398806 36536
rect 459646 36524 459652 36536
rect 459704 36524 459710 36576
rect 516042 36524 516048 36576
rect 516100 36564 516106 36576
rect 574738 36564 574744 36576
rect 516100 36536 574744 36564
rect 516100 36524 516106 36536
rect 574738 36524 574744 36536
rect 574796 36524 574802 36576
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 60182 35884 60188 35896
rect 3476 35856 60188 35884
rect 3476 35844 3482 35856
rect 60182 35844 60188 35856
rect 60240 35844 60246 35896
rect 184842 35232 184848 35284
rect 184900 35272 184906 35284
rect 244274 35272 244280 35284
rect 184900 35244 244280 35272
rect 184900 35232 184906 35244
rect 244274 35232 244280 35244
rect 244332 35232 244338 35284
rect 288342 35232 288348 35284
rect 288400 35272 288406 35284
rect 347774 35272 347780 35284
rect 288400 35244 347780 35272
rect 288400 35232 288406 35244
rect 347774 35232 347780 35244
rect 347832 35232 347838 35284
rect 395982 35232 395988 35284
rect 396040 35272 396046 35284
rect 455414 35272 455420 35284
rect 396040 35244 455420 35272
rect 396040 35232 396046 35244
rect 455414 35232 455420 35244
rect 455472 35232 455478 35284
rect 131022 35164 131028 35216
rect 131080 35204 131086 35216
rect 191834 35204 191840 35216
rect 131080 35176 191840 35204
rect 131080 35164 131086 35176
rect 191834 35164 191840 35176
rect 191892 35164 191898 35216
rect 241330 35164 241336 35216
rect 241388 35204 241394 35216
rect 302234 35204 302240 35216
rect 241388 35176 302240 35204
rect 241388 35164 241394 35176
rect 302234 35164 302240 35176
rect 302292 35164 302298 35216
rect 342162 35164 342168 35216
rect 342220 35204 342226 35216
rect 401594 35204 401600 35216
rect 342220 35176 401600 35204
rect 342220 35164 342226 35176
rect 401594 35164 401600 35176
rect 401652 35164 401658 35216
rect 460198 35164 460204 35216
rect 460256 35204 460262 35216
rect 520366 35204 520372 35216
rect 460256 35176 520372 35204
rect 460256 35164 460262 35176
rect 520366 35164 520372 35176
rect 520424 35164 520430 35216
rect 124122 33804 124128 33856
rect 124180 33844 124186 33856
rect 183554 33844 183560 33856
rect 124180 33816 183560 33844
rect 124180 33804 124186 33816
rect 183554 33804 183560 33816
rect 183612 33804 183618 33856
rect 227622 33804 227628 33856
rect 227680 33844 227686 33856
rect 287054 33844 287060 33856
rect 227680 33816 287060 33844
rect 227680 33804 227686 33816
rect 287054 33804 287060 33816
rect 287112 33804 287118 33856
rect 338022 33804 338028 33856
rect 338080 33844 338086 33856
rect 398834 33844 398840 33856
rect 338080 33816 398840 33844
rect 338080 33804 338086 33816
rect 398834 33804 398840 33816
rect 398892 33804 398898 33856
rect 441522 33804 441528 33856
rect 441580 33844 441586 33856
rect 502426 33844 502432 33856
rect 441580 33816 502432 33844
rect 441580 33804 441586 33816
rect 502426 33804 502432 33816
rect 502484 33804 502490 33856
rect 173802 33736 173808 33788
rect 173860 33776 173866 33788
rect 234614 33776 234620 33788
rect 173860 33748 234620 33776
rect 173860 33736 173866 33748
rect 234614 33736 234620 33748
rect 234672 33736 234678 33788
rect 284110 33736 284116 33788
rect 284168 33776 284174 33788
rect 345014 33776 345020 33788
rect 284168 33748 345020 33776
rect 284168 33736 284174 33748
rect 345014 33736 345020 33748
rect 345072 33736 345078 33788
rect 409782 33736 409788 33788
rect 409840 33776 409846 33788
rect 469214 33776 469220 33788
rect 409840 33748 469220 33776
rect 409840 33736 409846 33748
rect 469214 33736 469220 33748
rect 469272 33736 469278 33788
rect 502150 33736 502156 33788
rect 502208 33776 502214 33788
rect 563146 33776 563152 33788
rect 502208 33748 563152 33776
rect 502208 33736 502214 33748
rect 563146 33736 563152 33748
rect 563204 33736 563210 33788
rect 167730 32444 167736 32496
rect 167788 32484 167794 32496
rect 227806 32484 227812 32496
rect 167788 32456 227812 32484
rect 167788 32444 167794 32456
rect 227806 32444 227812 32456
rect 227864 32444 227870 32496
rect 281442 32444 281448 32496
rect 281500 32484 281506 32496
rect 340874 32484 340880 32496
rect 281500 32456 340880 32484
rect 281500 32444 281506 32456
rect 340874 32444 340880 32456
rect 340932 32444 340938 32496
rect 389082 32444 389088 32496
rect 389140 32484 389146 32496
rect 448514 32484 448520 32496
rect 389140 32456 448520 32484
rect 389140 32444 389146 32456
rect 448514 32444 448520 32456
rect 448572 32444 448578 32496
rect 119982 32376 119988 32428
rect 120040 32416 120046 32428
rect 180794 32416 180800 32428
rect 120040 32388 180800 32416
rect 120040 32376 120046 32388
rect 180794 32376 180800 32388
rect 180852 32376 180858 32428
rect 223390 32376 223396 32428
rect 223448 32416 223454 32428
rect 284294 32416 284300 32428
rect 223448 32388 284300 32416
rect 223448 32376 223454 32388
rect 284294 32376 284300 32388
rect 284352 32376 284358 32428
rect 335262 32376 335268 32428
rect 335320 32416 335326 32428
rect 394694 32416 394700 32428
rect 335320 32388 394700 32416
rect 335320 32376 335326 32388
rect 394694 32376 394700 32388
rect 394752 32376 394758 32428
rect 467742 32376 467748 32428
rect 467800 32416 467806 32428
rect 527174 32416 527180 32428
rect 467800 32388 527180 32416
rect 467800 32376 467806 32388
rect 527174 32376 527180 32388
rect 527232 32376 527238 32428
rect 160002 31084 160008 31136
rect 160060 31124 160066 31136
rect 219434 31124 219440 31136
rect 160060 31096 219440 31124
rect 160060 31084 160066 31096
rect 219434 31084 219440 31096
rect 219492 31084 219498 31136
rect 267550 31084 267556 31136
rect 267608 31124 267614 31136
rect 327074 31124 327080 31136
rect 267608 31096 327080 31124
rect 267608 31084 267614 31096
rect 327074 31084 327080 31096
rect 327132 31084 327138 31136
rect 378042 31084 378048 31136
rect 378100 31124 378106 31136
rect 437474 31124 437480 31136
rect 378100 31096 437480 31124
rect 378100 31084 378106 31096
rect 437474 31084 437480 31096
rect 437532 31084 437538 31136
rect 106182 31016 106188 31068
rect 106240 31056 106246 31068
rect 167086 31056 167092 31068
rect 106240 31028 167092 31056
rect 106240 31016 106246 31028
rect 167086 31016 167092 31028
rect 167144 31016 167150 31068
rect 216582 31016 216588 31068
rect 216640 31056 216646 31068
rect 277394 31056 277400 31068
rect 216640 31028 277400 31056
rect 216640 31016 216646 31028
rect 277394 31016 277400 31028
rect 277452 31016 277458 31068
rect 324222 31016 324228 31068
rect 324280 31056 324286 31068
rect 383654 31056 383660 31068
rect 324280 31028 383660 31056
rect 324280 31016 324286 31028
rect 383654 31016 383660 31028
rect 383712 31016 383718 31068
rect 449710 31016 449716 31068
rect 449768 31056 449774 31068
rect 509234 31056 509240 31068
rect 449768 31028 509240 31056
rect 449768 31016 449774 31028
rect 509234 31016 509240 31028
rect 509292 31016 509298 31068
rect 510522 31016 510528 31068
rect 510580 31056 510586 31068
rect 569954 31056 569960 31068
rect 510580 31028 569960 31056
rect 510580 31016 510586 31028
rect 569954 31016 569960 31028
rect 570012 31016 570018 31068
rect 523770 30268 523776 30320
rect 523828 30308 523834 30320
rect 580166 30308 580172 30320
rect 523828 30280 580172 30308
rect 523828 30268 523834 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 155862 29656 155868 29708
rect 155920 29696 155926 29708
rect 216674 29696 216680 29708
rect 155920 29668 216680 29696
rect 155920 29656 155926 29668
rect 216674 29656 216680 29668
rect 216732 29656 216738 29708
rect 259362 29656 259368 29708
rect 259420 29696 259426 29708
rect 320174 29696 320180 29708
rect 259420 29668 320180 29696
rect 259420 29656 259426 29668
rect 320174 29656 320180 29668
rect 320232 29656 320238 29708
rect 373902 29656 373908 29708
rect 373960 29696 373966 29708
rect 433334 29696 433340 29708
rect 373960 29668 433340 29696
rect 373960 29656 373966 29668
rect 433334 29656 433340 29668
rect 433392 29656 433398 29708
rect 102042 29588 102048 29640
rect 102100 29628 102106 29640
rect 162854 29628 162860 29640
rect 102100 29600 162860 29628
rect 102100 29588 102106 29600
rect 162854 29588 162860 29600
rect 162912 29588 162918 29640
rect 205450 29588 205456 29640
rect 205508 29628 205514 29640
rect 266354 29628 266360 29640
rect 205508 29600 266360 29628
rect 205508 29588 205514 29600
rect 266354 29588 266360 29600
rect 266412 29588 266418 29640
rect 317322 29588 317328 29640
rect 317380 29628 317386 29640
rect 376754 29628 376760 29640
rect 317380 29600 376760 29628
rect 317380 29588 317386 29600
rect 376754 29588 376760 29600
rect 376812 29588 376818 29640
rect 438762 29588 438768 29640
rect 438820 29628 438826 29640
rect 498194 29628 498200 29640
rect 438820 29600 498200 29628
rect 438820 29588 438826 29600
rect 498194 29588 498200 29600
rect 498252 29588 498258 29640
rect 427906 29016 427912 29028
rect 427867 28988 427912 29016
rect 427906 28976 427912 28988
rect 427964 28976 427970 29028
rect 434806 29016 434812 29028
rect 434767 28988 434812 29016
rect 434806 28976 434812 28988
rect 434864 28976 434870 29028
rect 248414 28908 248420 28960
rect 248472 28948 248478 28960
rect 248506 28948 248512 28960
rect 248472 28920 248512 28948
rect 248472 28908 248478 28920
rect 248506 28908 248512 28920
rect 248564 28908 248570 28960
rect 280798 28364 280804 28416
rect 280856 28404 280862 28416
rect 339494 28404 339500 28416
rect 280856 28376 339500 28404
rect 280856 28364 280862 28376
rect 339494 28364 339500 28376
rect 339552 28364 339558 28416
rect 97902 28296 97908 28348
rect 97960 28336 97966 28348
rect 158806 28336 158812 28348
rect 97960 28308 158812 28336
rect 97960 28296 97966 28308
rect 158806 28296 158812 28308
rect 158864 28296 158870 28348
rect 236638 28296 236644 28348
rect 236696 28336 236702 28348
rect 296714 28336 296720 28348
rect 236696 28308 296720 28336
rect 236696 28296 236702 28308
rect 296714 28296 296720 28308
rect 296772 28296 296778 28348
rect 371050 28296 371056 28348
rect 371108 28336 371114 28348
rect 430574 28336 430580 28348
rect 371108 28308 430580 28336
rect 371108 28296 371114 28308
rect 430574 28296 430580 28308
rect 430632 28296 430638 28348
rect 144730 28228 144736 28280
rect 144788 28268 144794 28280
rect 205634 28268 205640 28280
rect 144788 28240 205640 28268
rect 144788 28228 144794 28240
rect 205634 28228 205640 28240
rect 205692 28228 205698 28280
rect 208302 28228 208308 28280
rect 208360 28268 208366 28280
rect 269114 28268 269120 28280
rect 208360 28240 269120 28268
rect 208360 28228 208366 28240
rect 269114 28228 269120 28240
rect 269172 28228 269178 28280
rect 311802 28228 311808 28280
rect 311860 28268 311866 28280
rect 372614 28268 372620 28280
rect 311860 28240 372620 28268
rect 311860 28228 311866 28240
rect 372614 28228 372620 28240
rect 372672 28228 372678 28280
rect 445662 28228 445668 28280
rect 445720 28268 445726 28280
rect 505094 28268 505100 28280
rect 445720 28240 505100 28268
rect 445720 28228 445726 28240
rect 505094 28228 505100 28240
rect 505152 28228 505158 28280
rect 285766 27588 285772 27600
rect 285727 27560 285772 27588
rect 285766 27548 285772 27560
rect 285824 27548 285830 27600
rect 319438 26936 319444 26988
rect 319496 26976 319502 26988
rect 369854 26976 369860 26988
rect 319496 26948 369860 26976
rect 319496 26936 319502 26948
rect 369854 26936 369860 26948
rect 369912 26936 369918 26988
rect 492582 26936 492588 26988
rect 492640 26976 492646 26988
rect 552014 26976 552020 26988
rect 492640 26948 552020 26976
rect 492640 26936 492646 26948
rect 552014 26936 552020 26948
rect 552072 26936 552078 26988
rect 93762 26868 93768 26920
rect 93820 26908 93826 26920
rect 154574 26908 154580 26920
rect 93820 26880 154580 26908
rect 93820 26868 93826 26880
rect 154574 26868 154580 26880
rect 154632 26868 154638 26920
rect 165522 26868 165528 26920
rect 165580 26908 165586 26920
rect 226334 26908 226340 26920
rect 165580 26880 226340 26908
rect 165580 26868 165586 26880
rect 226334 26868 226340 26880
rect 226392 26868 226398 26920
rect 257890 26868 257896 26920
rect 257948 26908 257954 26920
rect 318794 26908 318800 26920
rect 257948 26880 318800 26908
rect 257948 26868 257954 26880
rect 318794 26868 318800 26880
rect 318852 26868 318858 26920
rect 367002 26868 367008 26920
rect 367060 26908 367066 26920
rect 426434 26908 426440 26920
rect 367060 26880 426440 26908
rect 367060 26868 367066 26880
rect 426434 26868 426440 26880
rect 426492 26868 426498 26920
rect 434622 26868 434628 26920
rect 434680 26908 434686 26920
rect 494054 26908 494060 26920
rect 434680 26880 494060 26908
rect 434680 26868 434686 26880
rect 494054 26868 494060 26880
rect 494112 26868 494118 26920
rect 306282 25576 306288 25628
rect 306340 25616 306346 25628
rect 365714 25616 365720 25628
rect 306340 25588 365720 25616
rect 306340 25576 306346 25588
rect 365714 25576 365720 25588
rect 365772 25576 365778 25628
rect 431862 25576 431868 25628
rect 431920 25616 431926 25628
rect 491294 25616 491300 25628
rect 431920 25588 491300 25616
rect 431920 25576 431926 25588
rect 491294 25576 491300 25588
rect 491352 25576 491358 25628
rect 91002 25508 91008 25560
rect 91060 25548 91066 25560
rect 150526 25548 150532 25560
rect 91060 25520 150532 25548
rect 91060 25508 91066 25520
rect 150526 25508 150532 25520
rect 150584 25508 150590 25560
rect 158622 25508 158628 25560
rect 158680 25548 158686 25560
rect 218054 25548 218060 25560
rect 158680 25520 218060 25548
rect 158680 25508 158686 25520
rect 218054 25508 218060 25520
rect 218112 25508 218118 25560
rect 251082 25508 251088 25560
rect 251140 25548 251146 25560
rect 311894 25548 311900 25560
rect 251140 25520 311900 25548
rect 251140 25508 251146 25520
rect 311894 25508 311900 25520
rect 311952 25508 311958 25560
rect 360102 25508 360108 25560
rect 360160 25548 360166 25560
rect 419534 25548 419540 25560
rect 360160 25520 419540 25548
rect 360160 25508 360166 25520
rect 419534 25508 419540 25520
rect 419592 25508 419598 25560
rect 485590 25508 485596 25560
rect 485648 25548 485654 25560
rect 545114 25548 545120 25560
rect 485648 25520 545120 25548
rect 485648 25508 485654 25520
rect 545114 25508 545120 25520
rect 545172 25508 545178 25560
rect 309042 24216 309048 24268
rect 309100 24256 309106 24268
rect 368474 24256 368480 24268
rect 309100 24228 368480 24256
rect 309100 24216 309106 24228
rect 368474 24216 368480 24228
rect 368532 24216 368538 24268
rect 249702 24148 249708 24200
rect 249760 24188 249766 24200
rect 310514 24188 310520 24200
rect 249760 24160 310520 24188
rect 249760 24148 249766 24160
rect 310514 24148 310520 24160
rect 310572 24148 310578 24200
rect 481542 24148 481548 24200
rect 481600 24188 481606 24200
rect 540974 24188 540980 24200
rect 481600 24160 540980 24188
rect 481600 24148 481606 24160
rect 540974 24148 540980 24160
rect 541032 24148 541038 24200
rect 86862 24080 86868 24132
rect 86920 24120 86926 24132
rect 147674 24120 147680 24132
rect 86920 24092 147680 24120
rect 86920 24080 86926 24092
rect 147674 24080 147680 24092
rect 147732 24080 147738 24132
rect 154482 24080 154488 24132
rect 154540 24120 154546 24132
rect 215294 24120 215300 24132
rect 154540 24092 215300 24120
rect 154540 24080 154546 24092
rect 215294 24080 215300 24092
rect 215352 24080 215358 24132
rect 226242 24080 226248 24132
rect 226300 24120 226306 24132
rect 287146 24120 287152 24132
rect 226300 24092 287152 24120
rect 226300 24080 226306 24092
rect 287146 24080 287152 24092
rect 287204 24080 287210 24132
rect 362770 24080 362776 24132
rect 362828 24120 362834 24132
rect 423674 24120 423680 24132
rect 362828 24092 423680 24120
rect 362828 24080 362834 24092
rect 423674 24080 423680 24092
rect 423732 24080 423738 24132
rect 427722 24080 427728 24132
rect 427780 24120 427786 24132
rect 487154 24120 487160 24132
rect 427780 24092 487160 24120
rect 427780 24080 427786 24092
rect 487154 24080 487160 24092
rect 487212 24080 487218 24132
rect 261478 22788 261484 22840
rect 261536 22828 261542 22840
rect 321554 22828 321560 22840
rect 261536 22800 321560 22828
rect 261536 22788 261542 22800
rect 321554 22788 321560 22800
rect 321612 22788 321618 22840
rect 482278 22788 482284 22840
rect 482336 22828 482342 22840
rect 536834 22828 536840 22840
rect 482336 22800 536840 22828
rect 482336 22788 482342 22800
rect 536834 22788 536840 22800
rect 536892 22788 536898 22840
rect 84838 22720 84844 22772
rect 84896 22760 84902 22772
rect 143534 22760 143540 22772
rect 84896 22732 143540 22760
rect 84896 22720 84902 22732
rect 143534 22720 143540 22732
rect 143592 22720 143598 22772
rect 151722 22720 151728 22772
rect 151780 22760 151786 22772
rect 211154 22760 211160 22772
rect 151780 22732 211160 22760
rect 151780 22720 151786 22732
rect 211154 22720 211160 22732
rect 211212 22720 211218 22772
rect 215110 22720 215116 22772
rect 215168 22760 215174 22772
rect 276014 22760 276020 22772
rect 215168 22732 276020 22760
rect 215168 22720 215174 22732
rect 276014 22720 276020 22732
rect 276072 22720 276078 22772
rect 286962 22720 286968 22772
rect 287020 22760 287026 22772
rect 347866 22760 347872 22772
rect 287020 22732 347872 22760
rect 287020 22720 287026 22732
rect 347866 22720 347872 22732
rect 347924 22720 347930 22772
rect 348418 22720 348424 22772
rect 348476 22760 348482 22772
rect 408586 22760 408592 22772
rect 348476 22732 408592 22760
rect 348476 22720 348482 22732
rect 408586 22720 408592 22732
rect 408644 22720 408650 22772
rect 423490 22720 423496 22772
rect 423548 22760 423554 22772
rect 484394 22760 484400 22772
rect 423548 22732 484400 22760
rect 423548 22720 423554 22732
rect 484394 22720 484400 22732
rect 484452 22720 484458 22772
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 59998 22080 60004 22092
rect 3200 22052 60004 22080
rect 3200 22040 3206 22052
rect 59998 22040 60004 22052
rect 60056 22040 60062 22092
rect 79962 21360 79968 21412
rect 80020 21400 80026 21412
rect 140866 21400 140872 21412
rect 80020 21372 140872 21400
rect 80020 21360 80026 21372
rect 140866 21360 140872 21372
rect 140924 21360 140930 21412
rect 147582 21360 147588 21412
rect 147640 21400 147646 21412
rect 208394 21400 208400 21412
rect 147640 21372 208400 21400
rect 147640 21360 147646 21372
rect 208394 21360 208400 21372
rect 208452 21360 208458 21412
rect 212442 21360 212448 21412
rect 212500 21400 212506 21412
rect 271874 21400 271880 21412
rect 212500 21372 271880 21400
rect 212500 21360 212506 21372
rect 271874 21360 271880 21372
rect 271932 21360 271938 21412
rect 273162 21360 273168 21412
rect 273220 21400 273226 21412
rect 332594 21400 332600 21412
rect 273220 21372 332600 21400
rect 273220 21360 273226 21372
rect 332594 21360 332600 21372
rect 332652 21360 332658 21412
rect 333882 21360 333888 21412
rect 333940 21400 333946 21412
rect 393314 21400 393320 21412
rect 333940 21372 393320 21400
rect 333940 21360 333946 21372
rect 393314 21360 393320 21372
rect 393372 21360 393378 21412
rect 412542 21360 412548 21412
rect 412600 21400 412606 21412
rect 471974 21400 471980 21412
rect 412600 21372 471980 21400
rect 412600 21360 412606 21372
rect 471974 21360 471980 21372
rect 472032 21360 472038 21412
rect 474642 21360 474648 21412
rect 474700 21400 474706 21412
rect 534074 21400 534080 21412
rect 474700 21372 534080 21400
rect 474700 21360 474706 21372
rect 534074 21360 534080 21372
rect 534132 21360 534138 21412
rect 312538 20000 312544 20052
rect 312596 20040 312602 20052
rect 367094 20040 367100 20052
rect 312596 20012 367100 20040
rect 312596 20000 312602 20012
rect 367094 20000 367100 20012
rect 367152 20000 367158 20052
rect 75822 19932 75828 19984
rect 75880 19972 75886 19984
rect 136634 19972 136640 19984
rect 75880 19944 136640 19972
rect 75880 19932 75886 19944
rect 136634 19932 136640 19944
rect 136692 19932 136698 19984
rect 144822 19932 144828 19984
rect 144880 19972 144886 19984
rect 204254 19972 204260 19984
rect 144880 19944 204260 19972
rect 144880 19932 144886 19944
rect 204254 19932 204260 19944
rect 204312 19932 204318 19984
rect 205542 19932 205548 19984
rect 205600 19972 205606 19984
rect 264974 19972 264980 19984
rect 205600 19944 264980 19972
rect 205600 19932 205606 19944
rect 264974 19932 264980 19944
rect 265032 19932 265038 19984
rect 269022 19932 269028 19984
rect 269080 19972 269086 19984
rect 329834 19972 329840 19984
rect 269080 19944 329840 19972
rect 269080 19932 269086 19944
rect 329834 19932 329840 19944
rect 329892 19932 329898 19984
rect 330478 19932 330484 19984
rect 330536 19972 330542 19984
rect 390646 19972 390652 19984
rect 330536 19944 390652 19972
rect 330536 19932 330542 19944
rect 390646 19932 390652 19944
rect 390704 19932 390710 19984
rect 408402 19932 408408 19984
rect 408460 19972 408466 19984
rect 467834 19972 467840 19984
rect 408460 19944 467840 19972
rect 408460 19932 408466 19944
rect 467834 19932 467840 19944
rect 467892 19932 467898 19984
rect 470502 19932 470508 19984
rect 470560 19972 470566 19984
rect 529934 19972 529940 19984
rect 470560 19944 529940 19972
rect 470560 19932 470566 19944
rect 529934 19932 529940 19944
rect 529992 19932 529998 19984
rect 248414 19292 248420 19304
rect 248375 19264 248420 19292
rect 248414 19252 248420 19264
rect 248472 19252 248478 19304
rect 259454 19292 259460 19304
rect 259415 19264 259460 19292
rect 259454 19252 259460 19264
rect 259512 19252 259518 19304
rect 269114 19292 269120 19304
rect 269075 19264 269120 19292
rect 269114 19252 269120 19264
rect 269172 19252 269178 19304
rect 277394 19252 277400 19304
rect 277452 19292 277458 19304
rect 277762 19292 277768 19304
rect 277452 19264 277768 19292
rect 277452 19252 277458 19264
rect 277762 19252 277768 19264
rect 277820 19252 277826 19304
rect 278958 19292 278964 19304
rect 278919 19264 278964 19292
rect 278958 19252 278964 19264
rect 279016 19252 279022 19304
rect 284294 19292 284300 19304
rect 284255 19264 284300 19292
rect 284294 19252 284300 19264
rect 284352 19252 284358 19304
rect 427906 19292 427912 19304
rect 427867 19264 427912 19292
rect 427906 19252 427912 19264
rect 427964 19252 427970 19304
rect 434806 19292 434812 19304
rect 434767 19264 434812 19292
rect 434806 19252 434812 19264
rect 434864 19252 434870 19304
rect 201402 18640 201408 18692
rect 201460 18680 201466 18692
rect 262306 18680 262312 18692
rect 201460 18652 262312 18680
rect 201460 18640 201466 18652
rect 262306 18640 262312 18652
rect 262364 18640 262370 18692
rect 266262 18640 266268 18692
rect 266320 18680 266326 18692
rect 325694 18680 325700 18692
rect 266320 18652 325700 18680
rect 266320 18640 266326 18652
rect 325694 18640 325700 18652
rect 325752 18640 325758 18692
rect 326982 18640 326988 18692
rect 327040 18680 327046 18692
rect 386414 18680 386420 18692
rect 327040 18652 386420 18680
rect 327040 18640 327046 18652
rect 386414 18640 386420 18652
rect 386472 18640 386478 18692
rect 73062 18572 73068 18624
rect 73120 18612 73126 18624
rect 132586 18612 132592 18624
rect 73120 18584 132592 18612
rect 73120 18572 73126 18584
rect 132586 18572 132592 18584
rect 132644 18572 132650 18624
rect 140682 18572 140688 18624
rect 140740 18612 140746 18624
rect 201586 18612 201592 18624
rect 140740 18584 201592 18612
rect 140740 18572 140746 18584
rect 201586 18572 201592 18584
rect 201644 18572 201650 18624
rect 303522 18572 303528 18624
rect 303580 18612 303586 18624
rect 364334 18612 364340 18624
rect 303580 18584 364340 18612
rect 303580 18572 303586 18584
rect 364334 18572 364340 18584
rect 364392 18572 364398 18624
rect 405642 18572 405648 18624
rect 405700 18612 405706 18624
rect 465074 18612 465080 18624
rect 405700 18584 465080 18612
rect 405700 18572 405706 18584
rect 465074 18572 465080 18584
rect 465132 18572 465138 18624
rect 473998 18572 474004 18624
rect 474056 18612 474062 18624
rect 532694 18612 532700 18624
rect 474056 18584 532700 18612
rect 474056 18572 474062 18584
rect 532694 18572 532700 18584
rect 532752 18572 532758 18624
rect 523862 17892 523868 17944
rect 523920 17932 523926 17944
rect 579798 17932 579804 17944
rect 523920 17904 579804 17932
rect 523920 17892 523926 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 129642 17280 129648 17332
rect 129700 17320 129706 17332
rect 190454 17320 190460 17332
rect 129700 17292 190460 17320
rect 129700 17280 129706 17292
rect 190454 17280 190460 17292
rect 190512 17280 190518 17332
rect 290458 17280 290464 17332
rect 290516 17320 290522 17332
rect 349154 17320 349160 17332
rect 290516 17292 349160 17320
rect 290516 17280 290522 17292
rect 349154 17280 349160 17292
rect 349212 17280 349218 17332
rect 403618 17280 403624 17332
rect 403676 17320 403682 17332
rect 460934 17320 460940 17332
rect 403676 17292 460940 17320
rect 403676 17280 403682 17292
rect 460934 17280 460940 17292
rect 460992 17280 460998 17332
rect 70302 17212 70308 17264
rect 70360 17252 70366 17264
rect 131114 17252 131120 17264
rect 70360 17224 131120 17252
rect 70360 17212 70366 17224
rect 131114 17212 131120 17224
rect 131172 17212 131178 17264
rect 197170 17212 197176 17264
rect 197228 17252 197234 17264
rect 258074 17252 258080 17264
rect 197228 17224 258080 17252
rect 197228 17212 197234 17224
rect 258074 17212 258080 17224
rect 258132 17212 258138 17264
rect 262122 17212 262128 17264
rect 262180 17252 262186 17264
rect 321646 17252 321652 17264
rect 262180 17224 321652 17252
rect 262180 17212 262186 17224
rect 321646 17212 321652 17224
rect 321704 17212 321710 17264
rect 322842 17212 322848 17264
rect 322900 17252 322906 17264
rect 382366 17252 382372 17264
rect 322900 17224 382372 17252
rect 322900 17212 322906 17224
rect 382366 17212 382372 17224
rect 382424 17212 382430 17264
rect 456702 17212 456708 17264
rect 456760 17252 456766 17264
rect 516134 17252 516140 17264
rect 456760 17224 516140 17252
rect 456760 17212 456766 17224
rect 516134 17212 516140 17224
rect 516192 17212 516198 17264
rect 126790 15920 126796 15972
rect 126848 15960 126854 15972
rect 186314 15960 186320 15972
rect 126848 15932 186320 15960
rect 126848 15920 126854 15932
rect 186314 15920 186320 15932
rect 186372 15920 186378 15972
rect 255222 15920 255228 15972
rect 255280 15960 255286 15972
rect 314654 15960 314660 15972
rect 255280 15932 314660 15960
rect 255280 15920 255286 15932
rect 314654 15920 314660 15932
rect 314712 15920 314718 15972
rect 315942 15920 315948 15972
rect 316000 15960 316006 15972
rect 375374 15960 375380 15972
rect 316000 15932 375380 15960
rect 316000 15920 316006 15932
rect 375374 15920 375380 15932
rect 375432 15920 375438 15972
rect 66898 15852 66904 15904
rect 66956 15892 66962 15904
rect 126974 15892 126980 15904
rect 66956 15864 126980 15892
rect 66956 15852 66962 15864
rect 126974 15852 126980 15864
rect 127032 15852 127038 15904
rect 194502 15852 194508 15904
rect 194560 15892 194566 15904
rect 253934 15892 253940 15904
rect 194560 15864 253940 15892
rect 194560 15852 194566 15864
rect 253934 15852 253940 15864
rect 253992 15852 253998 15904
rect 285582 15852 285588 15904
rect 285640 15892 285646 15904
rect 346394 15892 346400 15904
rect 285640 15864 346400 15892
rect 285640 15852 285646 15864
rect 346394 15852 346400 15864
rect 346452 15852 346458 15904
rect 397362 15852 397368 15904
rect 397420 15892 397426 15904
rect 458174 15892 458180 15904
rect 397420 15864 458180 15892
rect 397420 15852 397426 15864
rect 458174 15852 458180 15864
rect 458232 15852 458238 15904
rect 469122 15852 469128 15904
rect 469180 15892 469186 15904
rect 528646 15892 528652 15904
rect 469180 15864 528652 15892
rect 469180 15852 469186 15864
rect 528646 15852 528652 15864
rect 528704 15852 528710 15904
rect 276658 14560 276664 14612
rect 276716 14600 276722 14612
rect 335354 14600 335360 14612
rect 276716 14572 335360 14600
rect 276716 14560 276722 14572
rect 335354 14560 335360 14572
rect 335412 14560 335418 14612
rect 74442 14492 74448 14544
rect 74500 14532 74506 14544
rect 133874 14532 133880 14544
rect 74500 14504 133880 14532
rect 74500 14492 74506 14504
rect 133874 14492 133880 14504
rect 133932 14492 133938 14544
rect 187602 14492 187608 14544
rect 187660 14532 187666 14544
rect 247034 14532 247040 14544
rect 187660 14504 247040 14532
rect 187660 14492 187666 14504
rect 247034 14492 247040 14504
rect 247092 14492 247098 14544
rect 304902 14492 304908 14544
rect 304960 14532 304966 14544
rect 365806 14532 365812 14544
rect 304960 14504 365812 14532
rect 304960 14492 304966 14504
rect 365806 14492 365812 14504
rect 365864 14492 365870 14544
rect 122742 14424 122748 14476
rect 122800 14464 122806 14476
rect 183646 14464 183652 14476
rect 122800 14436 183652 14464
rect 122800 14424 122806 14436
rect 183646 14424 183652 14436
rect 183704 14424 183710 14476
rect 244182 14424 244188 14476
rect 244240 14464 244246 14476
rect 305086 14464 305092 14476
rect 244240 14436 305092 14464
rect 244240 14424 244246 14436
rect 305086 14424 305092 14436
rect 305144 14424 305150 14476
rect 384298 14424 384304 14476
rect 384356 14464 384362 14476
rect 443086 14464 443092 14476
rect 384356 14436 443092 14464
rect 384356 14424 384362 14436
rect 443086 14424 443092 14436
rect 443144 14424 443150 14476
rect 451918 14424 451924 14476
rect 451976 14464 451982 14476
rect 511994 14464 512000 14476
rect 451976 14436 512000 14464
rect 451976 14424 451982 14436
rect 511994 14424 512000 14436
rect 512052 14424 512058 14476
rect 272518 13200 272524 13252
rect 272576 13240 272582 13252
rect 331214 13240 331220 13252
rect 272576 13212 331220 13240
rect 272576 13200 272582 13212
rect 331214 13200 331220 13212
rect 331272 13200 331278 13252
rect 92290 13132 92296 13184
rect 92348 13172 92354 13184
rect 151814 13172 151820 13184
rect 92348 13144 151820 13172
rect 92348 13132 92354 13144
rect 151814 13132 151820 13144
rect 151872 13132 151878 13184
rect 241422 13132 241428 13184
rect 241480 13172 241486 13184
rect 301409 13175 301467 13181
rect 301409 13172 301421 13175
rect 241480 13144 301421 13172
rect 241480 13132 241486 13144
rect 301409 13141 301421 13144
rect 301455 13141 301467 13175
rect 301409 13135 301467 13141
rect 506382 13132 506388 13184
rect 506440 13172 506446 13184
rect 565814 13172 565820 13184
rect 506440 13144 565820 13172
rect 506440 13132 506446 13144
rect 565814 13132 565820 13144
rect 565872 13132 565878 13184
rect 118510 13064 118516 13116
rect 118568 13104 118574 13116
rect 179414 13104 179420 13116
rect 118568 13076 179420 13104
rect 118568 13064 118574 13076
rect 179414 13064 179420 13076
rect 179472 13064 179478 13116
rect 183462 13064 183468 13116
rect 183520 13104 183526 13116
rect 244366 13104 244372 13116
rect 183520 13076 244372 13104
rect 183520 13064 183526 13076
rect 244366 13064 244372 13076
rect 244424 13064 244430 13116
rect 302142 13064 302148 13116
rect 302200 13104 302206 13116
rect 361574 13104 361580 13116
rect 302200 13076 361580 13104
rect 302200 13064 302206 13076
rect 361574 13064 361580 13076
rect 361632 13064 361638 13116
rect 376662 13064 376668 13116
rect 376720 13104 376726 13116
rect 436094 13104 436100 13116
rect 376720 13076 436100 13104
rect 376720 13064 376726 13076
rect 436094 13064 436100 13076
rect 436152 13064 436158 13116
rect 448422 13064 448428 13116
rect 448480 13104 448486 13116
rect 507854 13104 507860 13116
rect 448480 13076 507860 13104
rect 448480 13064 448486 13076
rect 507854 13064 507860 13076
rect 507912 13064 507918 13116
rect 276014 12452 276020 12504
rect 276072 12452 276078 12504
rect 247034 12384 247040 12436
rect 247092 12424 247098 12436
rect 247954 12424 247960 12436
rect 247092 12396 247960 12424
rect 247092 12384 247098 12396
rect 247954 12384 247960 12396
rect 248012 12384 248018 12436
rect 253934 12384 253940 12436
rect 253992 12424 253998 12436
rect 255038 12424 255044 12436
rect 253992 12396 255044 12424
rect 253992 12384 253998 12396
rect 255038 12384 255044 12396
rect 255096 12384 255102 12436
rect 255314 12384 255320 12436
rect 255372 12424 255378 12436
rect 256234 12424 256240 12436
rect 255372 12396 256240 12424
rect 255372 12384 255378 12396
rect 256234 12384 256240 12396
rect 256292 12384 256298 12436
rect 258074 12384 258080 12436
rect 258132 12424 258138 12436
rect 258626 12424 258632 12436
rect 258132 12396 258632 12424
rect 258132 12384 258138 12396
rect 258626 12384 258632 12396
rect 258684 12384 258690 12436
rect 264974 12384 264980 12436
rect 265032 12424 265038 12436
rect 265802 12424 265808 12436
rect 265032 12396 265808 12424
rect 265032 12384 265038 12396
rect 265802 12384 265808 12396
rect 265860 12384 265866 12436
rect 266354 12384 266360 12436
rect 266412 12424 266418 12436
rect 266998 12424 267004 12436
rect 266412 12396 267004 12424
rect 266412 12384 266418 12396
rect 266998 12384 267004 12396
rect 267056 12384 267062 12436
rect 271874 12384 271880 12436
rect 271932 12424 271938 12436
rect 272886 12424 272892 12436
rect 271932 12396 272892 12424
rect 271932 12384 271938 12396
rect 272886 12384 272892 12396
rect 272944 12384 272950 12436
rect 273254 12384 273260 12436
rect 273312 12424 273318 12436
rect 274082 12424 274088 12436
rect 273312 12396 274088 12424
rect 273312 12384 273318 12396
rect 274082 12384 274088 12396
rect 274140 12384 274146 12436
rect 276032 12356 276060 12452
rect 280154 12384 280160 12436
rect 280212 12424 280218 12436
rect 281258 12424 281264 12436
rect 280212 12396 281264 12424
rect 280212 12384 280218 12396
rect 281258 12384 281264 12396
rect 281316 12384 281322 12436
rect 291194 12384 291200 12436
rect 291252 12424 291258 12436
rect 291930 12424 291936 12436
rect 291252 12396 291936 12424
rect 291252 12384 291258 12396
rect 291930 12384 291936 12396
rect 291988 12384 291994 12436
rect 298094 12384 298100 12436
rect 298152 12424 298158 12436
rect 299106 12424 299112 12436
rect 298152 12396 299112 12424
rect 298152 12384 298158 12396
rect 299106 12384 299112 12396
rect 299164 12384 299170 12436
rect 276474 12356 276480 12368
rect 276032 12328 276480 12356
rect 276474 12316 276480 12328
rect 276532 12316 276538 12368
rect 237282 11772 237288 11824
rect 237340 11812 237346 11824
rect 297910 11812 297916 11824
rect 237340 11784 297916 11812
rect 237340 11772 237346 11784
rect 297910 11772 297916 11784
rect 297968 11772 297974 11824
rect 298002 11772 298008 11824
rect 298060 11812 298066 11824
rect 357434 11812 357440 11824
rect 298060 11784 357440 11812
rect 298060 11772 298066 11784
rect 357434 11772 357440 11784
rect 357492 11772 357498 11824
rect 367738 11772 367744 11824
rect 367796 11812 367802 11824
rect 425054 11812 425060 11824
rect 367796 11784 425060 11812
rect 367796 11772 367802 11784
rect 425054 11772 425060 11784
rect 425112 11772 425118 11824
rect 442258 11772 442264 11824
rect 442316 11812 442322 11824
rect 500954 11812 500960 11824
rect 442316 11784 500960 11812
rect 442316 11772 442322 11784
rect 500954 11772 500960 11784
rect 501012 11772 501018 11824
rect 115842 11704 115848 11756
rect 115900 11744 115906 11756
rect 175366 11744 175372 11756
rect 115900 11716 175372 11744
rect 115900 11704 115906 11716
rect 175366 11704 175372 11716
rect 175424 11704 175430 11756
rect 179230 11704 179236 11756
rect 179288 11744 179294 11756
rect 240134 11744 240140 11756
rect 179288 11716 240140 11744
rect 179288 11704 179294 11716
rect 240134 11704 240140 11716
rect 240192 11704 240198 11756
rect 267642 11704 267648 11756
rect 267700 11744 267706 11756
rect 328454 11744 328460 11756
rect 267700 11716 328460 11744
rect 267700 11704 267706 11716
rect 328454 11704 328460 11716
rect 328512 11704 328518 11756
rect 424962 11704 424968 11756
rect 425020 11744 425026 11756
rect 485866 11744 485872 11756
rect 425020 11716 485872 11744
rect 425020 11704 425026 11716
rect 485866 11704 485872 11716
rect 485924 11704 485930 11756
rect 499482 11704 499488 11756
rect 499540 11744 499546 11756
rect 558914 11744 558920 11756
rect 499540 11716 558920 11744
rect 499540 11704 499546 11716
rect 558914 11704 558920 11716
rect 558972 11704 558978 11756
rect 176562 10344 176568 10396
rect 176620 10384 176626 10396
rect 236086 10384 236092 10396
rect 176620 10356 236092 10384
rect 176620 10344 176626 10356
rect 236086 10344 236092 10356
rect 236144 10344 236150 10396
rect 265618 10344 265624 10396
rect 265676 10384 265682 10396
rect 324314 10384 324320 10396
rect 265676 10356 324320 10384
rect 265676 10344 265682 10356
rect 324314 10344 324320 10356
rect 324372 10344 324378 10396
rect 438118 10344 438124 10396
rect 438176 10384 438182 10396
rect 496814 10384 496820 10396
rect 438176 10356 496820 10384
rect 438176 10344 438182 10356
rect 496814 10344 496820 10356
rect 496872 10344 496878 10396
rect 111702 10276 111708 10328
rect 111760 10316 111766 10328
rect 172514 10316 172520 10328
rect 111760 10288 172520 10316
rect 111760 10276 111766 10288
rect 172514 10276 172520 10288
rect 172572 10276 172578 10328
rect 233142 10276 233148 10328
rect 233200 10316 233206 10328
rect 294322 10316 294328 10328
rect 233200 10288 294328 10316
rect 233200 10276 233206 10288
rect 294322 10276 294328 10288
rect 294380 10276 294386 10328
rect 294598 10276 294604 10328
rect 294656 10316 294662 10328
rect 354674 10316 354680 10328
rect 294656 10288 354680 10316
rect 294656 10276 294662 10288
rect 354674 10276 354680 10288
rect 354732 10276 354738 10328
rect 355318 10276 355324 10328
rect 355376 10316 355382 10328
rect 415394 10316 415400 10328
rect 355376 10288 415400 10316
rect 355376 10276 355382 10288
rect 415394 10276 415400 10288
rect 415452 10276 415458 10328
rect 416682 10276 416688 10328
rect 416740 10316 416746 10328
rect 477586 10316 477592 10328
rect 416740 10288 477592 10316
rect 416740 10276 416746 10288
rect 477586 10276 477592 10288
rect 477644 10276 477650 10328
rect 496078 10276 496084 10328
rect 496136 10316 496142 10328
rect 554866 10316 554872 10328
rect 496136 10288 554872 10316
rect 496136 10276 496142 10288
rect 554866 10276 554872 10288
rect 554924 10276 554930 10328
rect 248417 9707 248475 9713
rect 248417 9673 248429 9707
rect 248463 9704 248475 9707
rect 249150 9704 249156 9716
rect 248463 9676 249156 9704
rect 248463 9673 248475 9676
rect 248417 9667 248475 9673
rect 249150 9664 249156 9676
rect 249208 9664 249214 9716
rect 259457 9707 259515 9713
rect 259457 9673 259469 9707
rect 259503 9704 259515 9707
rect 259822 9704 259828 9716
rect 259503 9676 259828 9704
rect 259503 9673 259515 9676
rect 259457 9667 259515 9673
rect 259822 9664 259828 9676
rect 259880 9664 259886 9716
rect 269117 9707 269175 9713
rect 269117 9673 269129 9707
rect 269163 9704 269175 9707
rect 269298 9704 269304 9716
rect 269163 9676 269304 9704
rect 269163 9673 269175 9676
rect 269117 9667 269175 9673
rect 269298 9664 269304 9676
rect 269356 9664 269362 9716
rect 278958 9704 278964 9716
rect 278919 9676 278964 9704
rect 278958 9664 278964 9676
rect 279016 9664 279022 9716
rect 284297 9707 284355 9713
rect 284297 9673 284309 9707
rect 284343 9704 284355 9707
rect 284754 9704 284760 9716
rect 284343 9676 284760 9704
rect 284343 9673 284355 9676
rect 284297 9667 284355 9673
rect 284754 9664 284760 9676
rect 284812 9664 284818 9716
rect 285769 9707 285827 9713
rect 285769 9673 285781 9707
rect 285815 9704 285827 9707
rect 285950 9704 285956 9716
rect 285815 9676 285956 9704
rect 285815 9673 285827 9676
rect 285769 9667 285827 9673
rect 285950 9664 285956 9676
rect 286008 9664 286014 9716
rect 301406 9704 301412 9716
rect 301367 9676 301412 9704
rect 301406 9664 301412 9676
rect 301464 9664 301470 9716
rect 427906 9704 427912 9716
rect 427867 9676 427912 9704
rect 427906 9664 427912 9676
rect 427964 9664 427970 9716
rect 434806 9704 434812 9716
rect 434767 9676 434812 9704
rect 434806 9664 434812 9676
rect 434864 9664 434870 9716
rect 276474 9596 276480 9648
rect 276532 9596 276538 9648
rect 430574 9596 430580 9648
rect 430632 9636 430638 9648
rect 431129 9639 431187 9645
rect 431129 9636 431141 9639
rect 430632 9608 431141 9636
rect 430632 9596 430638 9608
rect 431129 9605 431141 9608
rect 431175 9605 431187 9639
rect 431129 9599 431187 9605
rect 436094 9596 436100 9648
rect 436152 9636 436158 9648
rect 437017 9639 437075 9645
rect 437017 9636 437029 9639
rect 436152 9608 437029 9636
rect 436152 9596 436158 9608
rect 437017 9605 437029 9608
rect 437063 9605 437075 9639
rect 437017 9599 437075 9605
rect 276492 9512 276520 9596
rect 276474 9460 276480 9512
rect 276532 9460 276538 9512
rect 230382 9052 230388 9104
rect 230440 9092 230446 9104
rect 290734 9092 290740 9104
rect 230440 9064 290740 9092
rect 230440 9052 230446 9064
rect 290734 9052 290740 9064
rect 290792 9052 290798 9104
rect 291102 9052 291108 9104
rect 291160 9092 291166 9104
rect 351362 9092 351368 9104
rect 291160 9064 351368 9092
rect 291160 9052 291166 9064
rect 351362 9052 351368 9064
rect 351420 9052 351426 9104
rect 257982 8984 257988 9036
rect 258040 9024 258046 9036
rect 318058 9024 318064 9036
rect 258040 8996 318064 9024
rect 258040 8984 258046 8996
rect 318058 8984 318064 8996
rect 318116 8984 318122 9036
rect 351822 8984 351828 9036
rect 351880 9024 351886 9036
rect 412082 9024 412088 9036
rect 351880 8996 412088 9024
rect 351880 8984 351886 8996
rect 412082 8984 412088 8996
rect 412140 8984 412146 9036
rect 489178 8984 489184 9036
rect 489236 9024 489242 9036
rect 548886 9024 548892 9036
rect 489236 8996 548892 9024
rect 489236 8984 489242 8996
rect 548886 8984 548892 8996
rect 548944 8984 548950 9036
rect 108942 8916 108948 8968
rect 109000 8956 109006 8968
rect 169386 8956 169392 8968
rect 109000 8928 169392 8956
rect 109000 8916 109006 8928
rect 169386 8916 169392 8928
rect 169444 8916 169450 8968
rect 172422 8916 172428 8968
rect 172480 8956 172486 8968
rect 233694 8956 233700 8968
rect 172480 8928 233700 8956
rect 172480 8916 172486 8928
rect 233694 8916 233700 8928
rect 233752 8916 233758 8968
rect 310422 8916 310428 8968
rect 310480 8956 310486 8968
rect 371602 8956 371608 8968
rect 310480 8928 371608 8956
rect 310480 8916 310486 8928
rect 371602 8916 371608 8928
rect 371660 8916 371666 8968
rect 433978 8916 433984 8968
rect 434036 8956 434042 8968
rect 494146 8956 494152 8968
rect 434036 8928 494152 8956
rect 434036 8916 434042 8928
rect 494146 8916 494152 8928
rect 494204 8916 494210 8968
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 60090 8276 60096 8288
rect 3476 8248 60096 8276
rect 3476 8236 3482 8248
rect 60090 8236 60096 8248
rect 60148 8236 60154 8288
rect 284202 7760 284208 7812
rect 284260 7800 284266 7812
rect 284260 7772 288480 7800
rect 284260 7760 284266 7772
rect 223482 7624 223488 7676
rect 223540 7664 223546 7676
rect 283650 7664 283656 7676
rect 223540 7636 283656 7664
rect 223540 7624 223546 7636
rect 283650 7624 283656 7636
rect 283708 7624 283714 7676
rect 287054 7624 287060 7676
rect 287112 7664 287118 7676
rect 288342 7664 288348 7676
rect 287112 7636 288348 7664
rect 287112 7624 287118 7636
rect 288342 7624 288348 7636
rect 288400 7624 288406 7676
rect 288452 7664 288480 7772
rect 293862 7692 293868 7744
rect 293920 7732 293926 7744
rect 353754 7732 353760 7744
rect 293920 7704 353760 7732
rect 293920 7692 293926 7704
rect 353754 7692 353760 7704
rect 353812 7692 353818 7744
rect 344278 7664 344284 7676
rect 288452 7636 344284 7664
rect 344278 7624 344284 7636
rect 344336 7624 344342 7676
rect 423582 7624 423588 7676
rect 423640 7664 423646 7676
rect 483474 7664 483480 7676
rect 423640 7636 483480 7664
rect 423640 7624 423646 7636
rect 483474 7624 483480 7636
rect 483532 7624 483538 7676
rect 104802 7556 104808 7608
rect 104860 7596 104866 7608
rect 165890 7596 165896 7608
rect 104860 7568 165896 7596
rect 104860 7556 104866 7568
rect 165890 7556 165896 7568
rect 165948 7556 165954 7608
rect 169662 7556 169668 7608
rect 169720 7596 169726 7608
rect 230106 7596 230112 7608
rect 169720 7568 230112 7596
rect 169720 7556 169726 7568
rect 230106 7556 230112 7568
rect 230164 7556 230170 7608
rect 234522 7556 234528 7608
rect 234580 7596 234586 7608
rect 295518 7596 295524 7608
rect 234580 7568 295524 7596
rect 234580 7556 234586 7568
rect 295518 7556 295524 7568
rect 295576 7556 295582 7608
rect 344922 7556 344928 7608
rect 344980 7596 344986 7608
rect 404906 7596 404912 7608
rect 344980 7568 404912 7596
rect 344980 7556 344986 7568
rect 404906 7556 404912 7568
rect 404964 7556 404970 7608
rect 433334 7556 433340 7608
rect 433392 7596 433398 7608
rect 434622 7596 434628 7608
rect 433392 7568 434628 7596
rect 433392 7556 433398 7568
rect 434622 7556 434628 7568
rect 434680 7556 434686 7608
rect 452562 7556 452568 7608
rect 452620 7596 452626 7608
rect 513190 7596 513196 7608
rect 452620 7568 513196 7596
rect 452620 7556 452626 7568
rect 513190 7556 513196 7568
rect 513248 7556 513254 7608
rect 520090 7556 520096 7608
rect 520148 7596 520154 7608
rect 579798 7596 579804 7608
rect 520148 7568 579804 7596
rect 520148 7556 520154 7568
rect 579798 7556 579804 7568
rect 579856 7556 579862 7608
rect 244274 7488 244280 7540
rect 244332 7528 244338 7540
rect 245562 7528 245568 7540
rect 244332 7500 245568 7528
rect 244332 7488 244338 7500
rect 245562 7488 245568 7500
rect 245620 7488 245626 7540
rect 262214 7488 262220 7540
rect 262272 7528 262278 7540
rect 263410 7528 263416 7540
rect 262272 7500 263416 7528
rect 262272 7488 262278 7500
rect 263410 7488 263416 7500
rect 263468 7488 263474 7540
rect 270494 7488 270500 7540
rect 270552 7528 270558 7540
rect 271690 7528 271696 7540
rect 270552 7500 271696 7528
rect 270552 7488 270558 7500
rect 271690 7488 271696 7500
rect 271748 7488 271754 7540
rect 167638 6264 167644 6316
rect 167696 6304 167702 6316
rect 222930 6304 222936 6316
rect 167696 6276 222936 6304
rect 167696 6264 167702 6276
rect 222930 6264 222936 6276
rect 222988 6264 222994 6316
rect 301498 6264 301504 6316
rect 301556 6304 301562 6316
rect 360930 6304 360936 6316
rect 301556 6276 360936 6304
rect 301556 6264 301562 6276
rect 360930 6264 360936 6276
rect 360988 6264 360994 6316
rect 110230 6196 110236 6248
rect 110288 6236 110294 6248
rect 170582 6236 170588 6248
rect 110288 6208 170588 6236
rect 110288 6196 110294 6208
rect 170582 6196 170588 6208
rect 170640 6196 170646 6248
rect 219342 6196 219348 6248
rect 219400 6236 219406 6248
rect 279970 6236 279976 6248
rect 219400 6208 279976 6236
rect 219400 6196 219406 6208
rect 279970 6196 279976 6208
rect 280028 6196 280034 6248
rect 280062 6196 280068 6248
rect 280120 6236 280126 6248
rect 340690 6236 340696 6248
rect 280120 6208 340696 6236
rect 280120 6196 280126 6208
rect 340690 6196 340696 6208
rect 340748 6196 340754 6248
rect 100570 6128 100576 6180
rect 100628 6168 100634 6180
rect 162302 6168 162308 6180
rect 100628 6140 162308 6168
rect 100628 6128 100634 6140
rect 162302 6128 162308 6140
rect 162360 6128 162366 6180
rect 180702 6128 180708 6180
rect 180760 6168 180766 6180
rect 241974 6168 241980 6180
rect 180760 6140 241980 6168
rect 180760 6128 180766 6140
rect 241974 6128 241980 6140
rect 242032 6128 242038 6180
rect 252462 6128 252468 6180
rect 252520 6168 252526 6180
rect 313366 6168 313372 6180
rect 252520 6140 313372 6168
rect 252520 6128 252526 6140
rect 313366 6128 313372 6140
rect 313424 6128 313430 6180
rect 340782 6128 340788 6180
rect 340840 6168 340846 6180
rect 401318 6168 401324 6180
rect 340840 6140 401324 6168
rect 340840 6128 340846 6140
rect 401318 6128 401324 6140
rect 401376 6128 401382 6180
rect 430482 6128 430488 6180
rect 430540 6168 430546 6180
rect 490558 6168 490564 6180
rect 430540 6140 490564 6168
rect 430540 6128 430546 6140
rect 490558 6128 490564 6140
rect 490616 6128 490622 6180
rect 502242 6128 502248 6180
rect 502300 6168 502306 6180
rect 561950 6168 561956 6180
rect 502300 6140 561956 6168
rect 502300 6128 502306 6140
rect 561950 6128 561956 6140
rect 562008 6128 562014 6180
rect 374638 5516 374644 5568
rect 374696 5556 374702 5568
rect 379974 5556 379980 5568
rect 374696 5528 379980 5556
rect 374696 5516 374702 5528
rect 379974 5516 379980 5528
rect 380032 5516 380038 5568
rect 362862 5244 362868 5296
rect 362920 5284 362926 5296
rect 422754 5284 422760 5296
rect 362920 5256 422760 5284
rect 362920 5244 362926 5256
rect 422754 5244 422760 5256
rect 422812 5244 422818 5296
rect 463602 5244 463608 5296
rect 463660 5284 463666 5296
rect 523862 5284 523868 5296
rect 463660 5256 523868 5284
rect 463660 5244 463666 5256
rect 523862 5244 523868 5256
rect 523920 5244 523926 5296
rect 249797 5219 249855 5225
rect 249797 5185 249809 5219
rect 249843 5216 249855 5219
rect 259365 5219 259423 5225
rect 259365 5216 259377 5219
rect 249843 5188 259377 5216
rect 249843 5185 249855 5188
rect 249797 5179 249855 5185
rect 259365 5185 259377 5188
rect 259411 5185 259423 5219
rect 259365 5179 259423 5185
rect 380802 5176 380808 5228
rect 380860 5216 380866 5228
rect 440602 5216 440608 5228
rect 380860 5188 440608 5216
rect 380860 5176 380866 5188
rect 440602 5176 440608 5188
rect 440660 5176 440666 5228
rect 462222 5176 462228 5228
rect 462280 5216 462286 5228
rect 522666 5216 522672 5228
rect 462280 5188 522672 5216
rect 462280 5176 462286 5188
rect 522666 5176 522672 5188
rect 522724 5176 522730 5228
rect 260837 5151 260895 5157
rect 260837 5117 260849 5151
rect 260883 5148 260895 5151
rect 270497 5151 270555 5157
rect 260883 5120 262444 5148
rect 260883 5117 260895 5120
rect 260837 5111 260895 5117
rect 248322 5040 248328 5092
rect 248380 5080 248386 5092
rect 249797 5083 249855 5089
rect 249797 5080 249809 5083
rect 248380 5052 249809 5080
rect 248380 5040 248386 5052
rect 249797 5049 249809 5052
rect 249843 5049 249855 5083
rect 249797 5043 249855 5049
rect 259365 5015 259423 5021
rect 259365 4981 259377 5015
rect 259411 5012 259423 5015
rect 260837 5015 260895 5021
rect 260837 5012 260849 5015
rect 259411 4984 260849 5012
rect 259411 4981 259423 4984
rect 259365 4975 259423 4981
rect 260837 4981 260849 4984
rect 260883 4981 260895 5015
rect 262416 5012 262444 5120
rect 270497 5117 270509 5151
rect 270543 5148 270555 5151
rect 278777 5151 278835 5157
rect 278777 5148 278789 5151
rect 270543 5120 278789 5148
rect 270543 5117 270555 5120
rect 270497 5111 270555 5117
rect 278777 5117 278789 5120
rect 278823 5117 278835 5151
rect 278777 5111 278835 5117
rect 394602 5108 394608 5160
rect 394660 5148 394666 5160
rect 454862 5148 454868 5160
rect 394660 5120 454868 5148
rect 394660 5108 394666 5120
rect 454862 5108 454868 5120
rect 454920 5108 454926 5160
rect 487062 5108 487068 5160
rect 487120 5148 487126 5160
rect 547690 5148 547696 5160
rect 487120 5120 547696 5148
rect 487120 5108 487126 5120
rect 547690 5108 547696 5120
rect 547748 5108 547754 5160
rect 387702 5040 387708 5092
rect 387760 5080 387766 5092
rect 447778 5080 447784 5092
rect 387760 5052 447784 5080
rect 387760 5040 387766 5052
rect 447778 5040 447784 5052
rect 447836 5040 447842 5092
rect 484302 5040 484308 5092
rect 484360 5080 484366 5092
rect 544102 5080 544108 5092
rect 484360 5052 544108 5080
rect 484360 5040 484366 5052
rect 544102 5040 544108 5052
rect 544160 5040 544166 5092
rect 270497 5015 270555 5021
rect 270497 5012 270509 5015
rect 262416 4984 270509 5012
rect 260837 4975 260895 4981
rect 270497 4981 270509 4984
rect 270543 4981 270555 5015
rect 270497 4975 270555 4981
rect 296625 5015 296683 5021
rect 296625 4981 296637 5015
rect 296671 5012 296683 5015
rect 296671 4984 298048 5012
rect 296671 4981 296683 4984
rect 296625 4975 296683 4981
rect 298020 4944 298048 4984
rect 358722 4972 358728 5024
rect 358780 5012 358786 5024
rect 358780 4984 369164 5012
rect 358780 4972 358786 4984
rect 308582 4944 308588 4956
rect 298020 4916 308588 4944
rect 308582 4904 308588 4916
rect 308640 4904 308646 4956
rect 369136 4944 369164 4984
rect 369762 4972 369768 5024
rect 369820 5012 369826 5024
rect 429930 5012 429936 5024
rect 369820 4984 429936 5012
rect 369820 4972 369826 4984
rect 429930 4972 429936 4984
rect 429988 4972 429994 5024
rect 466362 4972 466368 5024
rect 466420 5012 466426 5024
rect 526254 5012 526260 5024
rect 466420 4984 526260 5012
rect 466420 4972 466426 4984
rect 526254 4972 526260 4984
rect 526312 4972 526318 5024
rect 419166 4944 419172 4956
rect 369136 4916 419172 4944
rect 419166 4904 419172 4916
rect 419224 4904 419230 4956
rect 419261 4947 419319 4953
rect 419261 4913 419273 4947
rect 419307 4944 419319 4947
rect 425057 4947 425115 4953
rect 425057 4944 425069 4947
rect 419307 4916 425069 4944
rect 419307 4913 419319 4916
rect 419261 4907 419319 4913
rect 425057 4913 425069 4916
rect 425103 4913 425115 4947
rect 434717 4947 434775 4953
rect 434717 4944 434729 4947
rect 425057 4907 425115 4913
rect 434640 4916 434729 4944
rect 68922 4836 68928 4888
rect 68980 4876 68986 4888
rect 130194 4876 130200 4888
rect 68980 4848 130200 4876
rect 68980 4836 68986 4848
rect 130194 4836 130200 4848
rect 130252 4836 130258 4888
rect 133782 4836 133788 4888
rect 133840 4876 133846 4888
rect 194410 4876 194416 4888
rect 133840 4848 194416 4876
rect 133840 4836 133846 4848
rect 194410 4836 194416 4848
rect 194468 4836 194474 4888
rect 209682 4836 209688 4888
rect 209740 4876 209746 4888
rect 270586 4876 270592 4888
rect 209740 4848 270592 4876
rect 209740 4836 209746 4848
rect 270586 4836 270592 4848
rect 270644 4836 270650 4888
rect 278777 4879 278835 4885
rect 278777 4845 278789 4879
rect 278823 4876 278835 4879
rect 287057 4879 287115 4885
rect 287057 4876 287069 4879
rect 278823 4848 287069 4876
rect 278823 4845 278835 4848
rect 278777 4839 278835 4845
rect 287057 4845 287069 4848
rect 287103 4845 287115 4879
rect 287057 4839 287115 4845
rect 308398 4836 308404 4888
rect 308456 4876 308462 4888
rect 343082 4876 343088 4888
rect 308456 4848 343088 4876
rect 308456 4836 308462 4848
rect 343082 4836 343088 4848
rect 343140 4836 343146 4888
rect 434640 4885 434668 4916
rect 434717 4913 434729 4916
rect 434763 4913 434775 4947
rect 434717 4907 434775 4913
rect 455322 4904 455328 4956
rect 455380 4944 455386 4956
rect 515582 4944 515588 4956
rect 455380 4916 515588 4944
rect 455380 4904 455386 4916
rect 515582 4904 515588 4916
rect 515640 4904 515646 4956
rect 393317 4879 393375 4885
rect 393317 4845 393329 4879
rect 393363 4876 393375 4879
rect 402977 4879 403035 4885
rect 402977 4876 402989 4879
rect 393363 4848 402989 4876
rect 393363 4845 393375 4848
rect 393317 4839 393375 4845
rect 402977 4845 402989 4848
rect 403023 4845 403035 4879
rect 402977 4839 403035 4845
rect 434625 4879 434683 4885
rect 434625 4845 434637 4879
rect 434671 4845 434683 4879
rect 434625 4839 434683 4845
rect 444285 4879 444343 4885
rect 444285 4845 444297 4879
rect 444331 4876 444343 4879
rect 445113 4879 445171 4885
rect 445113 4876 445125 4879
rect 444331 4848 445125 4876
rect 444331 4845 444343 4848
rect 444285 4839 444343 4845
rect 445113 4845 445125 4848
rect 445159 4845 445171 4879
rect 445113 4839 445171 4845
rect 459462 4836 459468 4888
rect 459520 4876 459526 4888
rect 519078 4876 519084 4888
rect 459520 4848 519084 4876
rect 459520 4836 459526 4848
rect 519078 4836 519084 4848
rect 519136 4836 519142 4888
rect 66162 4768 66168 4820
rect 66220 4808 66226 4820
rect 126606 4808 126612 4820
rect 66220 4780 126612 4808
rect 66220 4768 66226 4780
rect 126606 4768 126612 4780
rect 126664 4768 126670 4820
rect 126882 4768 126888 4820
rect 126940 4808 126946 4820
rect 188430 4808 188436 4820
rect 126940 4780 188436 4808
rect 126940 4768 126946 4780
rect 188430 4768 188436 4780
rect 188488 4768 188494 4820
rect 190362 4768 190368 4820
rect 190420 4808 190426 4820
rect 251450 4808 251456 4820
rect 190420 4780 251456 4808
rect 190420 4768 190426 4780
rect 251450 4768 251456 4780
rect 251508 4768 251514 4820
rect 270402 4768 270408 4820
rect 270460 4808 270466 4820
rect 331306 4808 331312 4820
rect 270460 4780 331312 4808
rect 270460 4768 270466 4780
rect 331306 4768 331312 4780
rect 331364 4768 331370 4820
rect 333238 4768 333244 4820
rect 333296 4808 333302 4820
rect 357250 4808 357256 4820
rect 333296 4780 357256 4808
rect 333296 4768 333302 4780
rect 357250 4768 357256 4780
rect 357308 4768 357314 4820
rect 372522 4768 372528 4820
rect 372580 4808 372586 4820
rect 433518 4808 433524 4820
rect 372580 4780 433524 4808
rect 372580 4768 372586 4780
rect 433518 4768 433524 4780
rect 433576 4768 433582 4820
rect 476022 4768 476028 4820
rect 476080 4808 476086 4820
rect 536926 4808 536932 4820
rect 476080 4780 536932 4808
rect 476080 4768 476086 4780
rect 536926 4768 536932 4780
rect 536984 4768 536990 4820
rect 287057 4743 287115 4749
rect 287057 4709 287069 4743
rect 287103 4740 287115 4743
rect 296625 4743 296683 4749
rect 296625 4740 296637 4743
rect 287103 4712 296637 4740
rect 287103 4709 287115 4712
rect 287057 4703 287115 4709
rect 296625 4709 296637 4712
rect 296671 4709 296683 4743
rect 296625 4703 296683 4709
rect 390462 4700 390468 4752
rect 390520 4740 390526 4752
rect 393317 4743 393375 4749
rect 393317 4740 393329 4743
rect 390520 4712 393329 4740
rect 390520 4700 390526 4712
rect 393317 4709 393329 4712
rect 393363 4709 393375 4743
rect 393317 4703 393375 4709
rect 402977 4743 403035 4749
rect 402977 4709 402989 4743
rect 403023 4740 403035 4743
rect 419261 4743 419319 4749
rect 419261 4740 419273 4743
rect 403023 4712 419273 4740
rect 403023 4709 403035 4712
rect 402977 4703 403035 4709
rect 419261 4709 419273 4712
rect 419307 4709 419319 4743
rect 419261 4703 419319 4709
rect 434717 4743 434775 4749
rect 434717 4709 434729 4743
rect 434763 4740 434775 4743
rect 444285 4743 444343 4749
rect 444285 4740 444297 4743
rect 434763 4712 444297 4740
rect 434763 4709 434775 4712
rect 434717 4703 434775 4709
rect 444285 4709 444297 4712
rect 444331 4709 444343 4743
rect 444285 4703 444343 4709
rect 425057 4675 425115 4681
rect 425057 4641 425069 4675
rect 425103 4672 425115 4675
rect 434625 4675 434683 4681
rect 434625 4672 434637 4675
rect 425103 4644 434637 4672
rect 425103 4641 425115 4644
rect 425057 4635 425115 4641
rect 434625 4641 434637 4644
rect 434671 4641 434683 4675
rect 434625 4635 434683 4641
rect 143442 4088 143448 4140
rect 143500 4128 143506 4140
rect 203886 4128 203892 4140
rect 143500 4100 203892 4128
rect 143500 4088 143506 4100
rect 203886 4088 203892 4100
rect 203944 4088 203950 4140
rect 222102 4088 222108 4140
rect 222160 4128 222166 4140
rect 282454 4128 282460 4140
rect 222160 4100 282460 4128
rect 222160 4088 222166 4100
rect 282454 4088 282460 4100
rect 282512 4088 282518 4140
rect 336642 4088 336648 4140
rect 336700 4128 336706 4140
rect 396626 4128 396632 4140
rect 336700 4100 396632 4128
rect 336700 4088 336706 4100
rect 396626 4088 396632 4100
rect 396684 4088 396690 4140
rect 433242 4088 433248 4140
rect 433300 4128 433306 4140
rect 492950 4128 492956 4140
rect 433300 4100 492956 4128
rect 433300 4088 433306 4100
rect 492950 4088 492956 4100
rect 493008 4088 493014 4140
rect 496722 4088 496728 4140
rect 496780 4128 496786 4140
rect 557166 4128 557172 4140
rect 496780 4100 557172 4128
rect 496780 4088 496786 4100
rect 557166 4088 557172 4100
rect 557224 4088 557230 4140
rect 125502 4020 125508 4072
rect 125560 4060 125566 4072
rect 186038 4060 186044 4072
rect 125560 4032 186044 4060
rect 125560 4020 125566 4032
rect 186038 4020 186044 4032
rect 186096 4020 186102 4072
rect 193122 4020 193128 4072
rect 193180 4060 193186 4072
rect 253842 4060 253848 4072
rect 193180 4032 253848 4060
rect 193180 4020 193186 4032
rect 253842 4020 253848 4032
rect 253900 4020 253906 4072
rect 357342 4020 357348 4072
rect 357400 4060 357406 4072
rect 417970 4060 417976 4072
rect 357400 4032 417976 4060
rect 357400 4020 357406 4032
rect 417970 4020 417976 4032
rect 418028 4020 418034 4072
rect 464982 4020 464988 4072
rect 465040 4060 465046 4072
rect 525058 4060 525064 4072
rect 465040 4032 525064 4060
rect 465040 4020 465046 4032
rect 525058 4020 525064 4032
rect 525116 4020 525122 4072
rect 78582 3952 78588 4004
rect 78640 3992 78646 4004
rect 139670 3992 139676 4004
rect 78640 3964 139676 3992
rect 78640 3952 78646 3964
rect 139670 3952 139676 3964
rect 139728 3952 139734 4004
rect 161382 3952 161388 4004
rect 161440 3992 161446 4004
rect 221734 3992 221740 4004
rect 161440 3964 221740 3992
rect 161440 3952 161446 3964
rect 221734 3952 221740 3964
rect 221792 3952 221798 4004
rect 229002 3952 229008 4004
rect 229060 3992 229066 4004
rect 289538 3992 289544 4004
rect 229060 3964 289544 3992
rect 229060 3952 229066 3964
rect 289538 3952 289544 3964
rect 289596 3952 289602 4004
rect 343542 3952 343548 4004
rect 343600 3992 343606 4004
rect 403710 3992 403716 4004
rect 343600 3964 403716 3992
rect 343600 3952 343606 3964
rect 403710 3952 403716 3964
rect 403768 3952 403774 4004
rect 442902 3952 442908 4004
rect 442960 3992 442966 4004
rect 503622 3992 503628 4004
rect 442960 3964 503628 3992
rect 442960 3952 442966 3964
rect 503622 3952 503628 3964
rect 503680 3952 503686 4004
rect 514662 3952 514668 4004
rect 514720 3992 514726 4004
rect 575014 3992 575020 4004
rect 514720 3964 575020 3992
rect 514720 3952 514726 3964
rect 575014 3952 575020 3964
rect 575072 3952 575078 4004
rect 85482 3884 85488 3936
rect 85540 3924 85546 3936
rect 146846 3924 146852 3936
rect 85540 3896 146852 3924
rect 85540 3884 85546 3896
rect 146846 3884 146852 3896
rect 146904 3884 146910 3936
rect 150526 3884 150532 3936
rect 150584 3924 150590 3936
rect 151538 3924 151544 3936
rect 150584 3896 151544 3924
rect 150584 3884 150590 3896
rect 151538 3884 151544 3896
rect 151596 3884 151602 3936
rect 171042 3884 171048 3936
rect 171100 3924 171106 3936
rect 232498 3924 232504 3936
rect 171100 3896 232504 3924
rect 171100 3884 171106 3896
rect 232498 3884 232504 3896
rect 232556 3884 232562 3936
rect 361482 3884 361488 3936
rect 361540 3924 361546 3936
rect 421558 3924 421564 3936
rect 361540 3896 421564 3924
rect 361540 3884 361546 3896
rect 421558 3884 421564 3896
rect 421616 3884 421622 3936
rect 429102 3884 429108 3936
rect 429160 3924 429166 3936
rect 489362 3924 489368 3936
rect 429160 3896 489368 3924
rect 429160 3884 429166 3896
rect 489362 3884 489368 3896
rect 489420 3884 489426 3936
rect 500862 3884 500868 3936
rect 500920 3924 500926 3936
rect 560754 3924 560760 3936
rect 500920 3896 560760 3924
rect 500920 3884 500926 3896
rect 560754 3884 560760 3896
rect 560812 3884 560818 3936
rect 128262 3816 128268 3868
rect 128320 3856 128326 3868
rect 189626 3856 189632 3868
rect 128320 3828 189632 3856
rect 128320 3816 128326 3828
rect 189626 3816 189632 3828
rect 189684 3816 189690 3868
rect 201494 3816 201500 3868
rect 201552 3856 201558 3868
rect 202690 3856 202696 3868
rect 201552 3828 202696 3856
rect 201552 3816 201558 3828
rect 202690 3816 202696 3828
rect 202748 3816 202754 3868
rect 215202 3816 215208 3868
rect 215260 3856 215266 3868
rect 275278 3856 275284 3868
rect 215260 3828 275284 3856
rect 215260 3816 215266 3828
rect 275278 3816 275284 3828
rect 275336 3816 275342 3868
rect 332502 3816 332508 3868
rect 332560 3856 332566 3868
rect 393038 3856 393044 3868
rect 332560 3828 393044 3856
rect 332560 3816 332566 3828
rect 393038 3816 393044 3828
rect 393096 3816 393102 3868
rect 393222 3816 393228 3868
rect 393280 3856 393286 3868
rect 453666 3856 453672 3868
rect 393280 3828 453672 3856
rect 393280 3816 393286 3828
rect 453666 3816 453672 3828
rect 453724 3816 453730 3868
rect 493962 3816 493968 3868
rect 494020 3856 494026 3868
rect 553578 3856 553584 3868
rect 494020 3828 553584 3856
rect 494020 3816 494026 3828
rect 553578 3816 553584 3828
rect 553636 3816 553642 3868
rect 110322 3748 110328 3800
rect 110380 3788 110386 3800
rect 171778 3788 171784 3800
rect 110380 3760 171784 3788
rect 110380 3748 110386 3760
rect 171778 3748 171784 3760
rect 171836 3748 171842 3800
rect 175182 3748 175188 3800
rect 175240 3788 175246 3800
rect 235994 3788 236000 3800
rect 175240 3760 236000 3788
rect 175240 3748 175246 3760
rect 235994 3748 236000 3760
rect 236052 3748 236058 3800
rect 240042 3748 240048 3800
rect 240100 3788 240106 3800
rect 300302 3788 300308 3800
rect 240100 3760 300308 3788
rect 240100 3748 240106 3760
rect 300302 3748 300308 3760
rect 300360 3748 300366 3800
rect 350442 3748 350448 3800
rect 350500 3788 350506 3800
rect 410886 3788 410892 3800
rect 350500 3760 410892 3788
rect 350500 3748 350506 3760
rect 410886 3748 410892 3760
rect 410944 3748 410950 3800
rect 411162 3748 411168 3800
rect 411220 3788 411226 3800
rect 471514 3788 471520 3800
rect 411220 3760 471520 3788
rect 411220 3748 411226 3760
rect 471514 3748 471520 3760
rect 471572 3748 471578 3800
rect 478782 3748 478788 3800
rect 478840 3788 478846 3800
rect 539318 3788 539324 3800
rect 478840 3760 539324 3788
rect 478840 3748 478846 3760
rect 539318 3748 539324 3760
rect 539376 3748 539382 3800
rect 114462 3680 114468 3732
rect 114520 3720 114526 3732
rect 175274 3720 175280 3732
rect 114520 3692 175280 3720
rect 114520 3680 114526 3692
rect 175274 3680 175280 3692
rect 175332 3680 175338 3732
rect 175366 3680 175372 3732
rect 175424 3720 175430 3732
rect 176562 3720 176568 3732
rect 175424 3692 176568 3720
rect 175424 3680 175430 3692
rect 176562 3680 176568 3692
rect 176620 3680 176626 3732
rect 182082 3680 182088 3732
rect 182140 3720 182146 3732
rect 243170 3720 243176 3732
rect 182140 3692 243176 3720
rect 182140 3680 182146 3692
rect 243170 3680 243176 3692
rect 243228 3680 243234 3732
rect 328362 3680 328368 3732
rect 328420 3720 328426 3732
rect 389450 3720 389456 3732
rect 328420 3692 389456 3720
rect 328420 3680 328426 3692
rect 389450 3680 389456 3692
rect 389508 3680 389514 3732
rect 400122 3680 400128 3732
rect 400180 3720 400186 3732
rect 460842 3720 460848 3732
rect 400180 3692 460848 3720
rect 400180 3680 400186 3692
rect 460842 3680 460848 3692
rect 460900 3680 460906 3732
rect 460934 3680 460940 3732
rect 460992 3720 460998 3732
rect 521470 3720 521476 3732
rect 460992 3692 521476 3720
rect 460992 3680 460998 3692
rect 521470 3680 521476 3692
rect 521528 3680 521534 3732
rect 521562 3680 521568 3732
rect 521620 3720 521626 3732
rect 582190 3720 582196 3732
rect 521620 3692 582196 3720
rect 521620 3680 521626 3692
rect 582190 3680 582196 3692
rect 582248 3680 582254 3732
rect 121362 3612 121368 3664
rect 121420 3652 121426 3664
rect 182542 3652 182548 3664
rect 121420 3624 182548 3652
rect 121420 3612 121426 3624
rect 182542 3612 182548 3624
rect 182600 3612 182606 3664
rect 183554 3612 183560 3664
rect 183612 3652 183618 3664
rect 184842 3652 184848 3664
rect 183612 3624 184848 3652
rect 183612 3612 183618 3624
rect 184842 3612 184848 3624
rect 184900 3612 184906 3664
rect 188982 3612 188988 3664
rect 189040 3652 189046 3664
rect 250346 3652 250352 3664
rect 189040 3624 250352 3652
rect 189040 3612 189046 3624
rect 250346 3612 250352 3624
rect 250404 3612 250410 3664
rect 321462 3612 321468 3664
rect 321520 3652 321526 3664
rect 382274 3652 382280 3664
rect 321520 3624 382280 3652
rect 321520 3612 321526 3624
rect 382274 3612 382280 3624
rect 382332 3612 382338 3664
rect 382366 3612 382372 3664
rect 382424 3652 382430 3664
rect 383562 3652 383568 3664
rect 382424 3624 383568 3652
rect 382424 3612 382430 3624
rect 383562 3612 383568 3624
rect 383620 3612 383626 3664
rect 390554 3612 390560 3664
rect 390612 3652 390618 3664
rect 391842 3652 391848 3664
rect 390612 3624 391848 3652
rect 390612 3612 390618 3624
rect 391842 3612 391848 3624
rect 391900 3612 391906 3664
rect 408494 3612 408500 3664
rect 408552 3652 408558 3664
rect 409690 3652 409696 3664
rect 408552 3624 409696 3652
rect 408552 3612 408558 3624
rect 409690 3612 409696 3624
rect 409748 3612 409754 3664
rect 418062 3612 418068 3664
rect 418120 3652 418126 3664
rect 478690 3652 478696 3664
rect 418120 3624 478696 3652
rect 418120 3612 418126 3624
rect 478690 3612 478696 3624
rect 478748 3612 478754 3664
rect 485774 3612 485780 3664
rect 485832 3652 485838 3664
rect 486970 3652 486976 3664
rect 485832 3624 486976 3652
rect 485832 3612 485838 3624
rect 486970 3612 486976 3624
rect 487028 3612 487034 3664
rect 503438 3612 503444 3664
rect 503496 3652 503502 3664
rect 564342 3652 564348 3664
rect 503496 3624 564348 3652
rect 503496 3612 503502 3624
rect 564342 3612 564348 3624
rect 564400 3612 564406 3664
rect 132402 3544 132408 3596
rect 132460 3584 132466 3596
rect 193214 3584 193220 3596
rect 132460 3556 193220 3584
rect 132460 3544 132466 3556
rect 193214 3544 193220 3556
rect 193272 3544 193278 3596
rect 200022 3544 200028 3596
rect 200080 3584 200086 3596
rect 261018 3584 261024 3596
rect 200080 3556 261024 3584
rect 200080 3544 200086 3556
rect 261018 3544 261024 3556
rect 261076 3544 261082 3596
rect 321646 3544 321652 3596
rect 321704 3584 321710 3596
rect 322842 3584 322848 3596
rect 321704 3556 322848 3584
rect 321704 3544 321710 3556
rect 322842 3544 322848 3556
rect 322900 3544 322906 3596
rect 378778 3584 378784 3596
rect 322952 3556 378784 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 63494 3516 63500 3528
rect 1728 3488 63500 3516
rect 1728 3476 1734 3488
rect 63494 3476 63500 3488
rect 63552 3476 63558 3528
rect 132586 3476 132592 3528
rect 132644 3516 132650 3528
rect 133782 3516 133788 3528
rect 132644 3488 133788 3516
rect 132644 3476 132650 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 139302 3476 139308 3528
rect 139360 3516 139366 3528
rect 200390 3516 200396 3528
rect 139360 3488 200396 3516
rect 139360 3476 139366 3488
rect 200390 3476 200396 3488
rect 200448 3476 200454 3528
rect 206922 3476 206928 3528
rect 206980 3516 206986 3528
rect 268102 3516 268108 3528
rect 206980 3488 268108 3516
rect 206980 3476 206986 3488
rect 268102 3476 268108 3488
rect 268160 3476 268166 3528
rect 304994 3476 305000 3528
rect 305052 3516 305058 3528
rect 306190 3516 306196 3528
rect 305052 3488 306196 3516
rect 305052 3476 305058 3488
rect 306190 3476 306196 3488
rect 306248 3476 306254 3528
rect 318702 3476 318708 3528
rect 318760 3516 318766 3528
rect 322952 3516 322980 3556
rect 378778 3544 378784 3556
rect 378836 3544 378842 3596
rect 382182 3544 382188 3596
rect 382240 3584 382246 3596
rect 442994 3584 443000 3596
rect 382240 3556 443000 3584
rect 382240 3544 382246 3556
rect 442994 3544 443000 3556
rect 443052 3544 443058 3596
rect 451274 3544 451280 3596
rect 451332 3584 451338 3596
rect 452470 3584 452476 3596
rect 451332 3556 452476 3584
rect 451332 3544 451338 3556
rect 452470 3544 452476 3556
rect 452528 3544 452534 3596
rect 467834 3544 467840 3596
rect 467892 3584 467898 3596
rect 469122 3584 469128 3596
rect 467892 3556 469128 3584
rect 467892 3544 467898 3556
rect 469122 3544 469128 3556
rect 469180 3544 469186 3596
rect 471882 3544 471888 3596
rect 471940 3584 471946 3596
rect 528557 3587 528615 3593
rect 528557 3584 528569 3587
rect 471940 3556 528569 3584
rect 471940 3544 471946 3556
rect 528557 3553 528569 3556
rect 528603 3553 528615 3587
rect 528557 3547 528615 3553
rect 528646 3544 528652 3596
rect 528704 3584 528710 3596
rect 529842 3584 529848 3596
rect 528704 3556 529848 3584
rect 528704 3544 528710 3556
rect 529842 3544 529848 3556
rect 529900 3544 529906 3596
rect 536834 3544 536840 3596
rect 536892 3584 536898 3596
rect 538122 3584 538128 3596
rect 536892 3556 538128 3584
rect 536892 3544 536898 3556
rect 538122 3544 538128 3556
rect 538180 3544 538186 3596
rect 318760 3488 322980 3516
rect 318760 3476 318766 3488
rect 331214 3476 331220 3528
rect 331272 3516 331278 3528
rect 332410 3516 332416 3528
rect 331272 3488 332416 3516
rect 331272 3476 331278 3488
rect 332410 3476 332416 3488
rect 332468 3476 332474 3528
rect 347774 3476 347780 3528
rect 347832 3516 347838 3528
rect 349062 3516 349068 3528
rect 347832 3488 349068 3516
rect 347832 3476 347838 3488
rect 349062 3476 349068 3488
rect 349120 3476 349126 3528
rect 407298 3516 407304 3528
rect 350552 3488 407304 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 62114 3448 62120 3460
rect 624 3420 62120 3448
rect 624 3408 630 3420
rect 62114 3408 62120 3420
rect 62172 3408 62178 3460
rect 71682 3408 71688 3460
rect 71740 3448 71746 3460
rect 71740 3420 132632 3448
rect 71740 3408 71746 3420
rect 132604 3392 132632 3420
rect 140774 3408 140780 3460
rect 140832 3448 140838 3460
rect 142062 3448 142068 3460
rect 140832 3420 142068 3448
rect 140832 3408 140838 3420
rect 142062 3408 142068 3420
rect 142120 3408 142126 3460
rect 164142 3408 164148 3460
rect 164200 3448 164206 3460
rect 225322 3448 225328 3460
rect 164200 3420 225328 3448
rect 164200 3408 164206 3420
rect 225322 3408 225328 3420
rect 225380 3408 225386 3460
rect 246942 3408 246948 3460
rect 247000 3448 247006 3460
rect 307386 3448 307392 3460
rect 247000 3420 307392 3448
rect 247000 3408 247006 3420
rect 307386 3408 307392 3420
rect 307444 3408 307450 3460
rect 314562 3408 314568 3460
rect 314620 3448 314626 3460
rect 314620 3420 314700 3448
rect 314620 3408 314626 3420
rect 132586 3340 132592 3392
rect 132644 3340 132650 3392
rect 136450 3340 136456 3392
rect 136508 3380 136514 3392
rect 196802 3380 196808 3392
rect 136508 3352 196808 3380
rect 136508 3340 136514 3352
rect 196802 3340 196808 3352
rect 196860 3340 196866 3392
rect 197262 3340 197268 3392
rect 197320 3380 197326 3392
rect 257430 3380 257436 3392
rect 197320 3352 257436 3380
rect 197320 3340 197326 3352
rect 257430 3340 257436 3352
rect 257488 3340 257494 3392
rect 150342 3272 150348 3324
rect 150400 3312 150406 3324
rect 211062 3312 211068 3324
rect 150400 3284 211068 3312
rect 150400 3272 150406 3284
rect 211062 3272 211068 3284
rect 211120 3272 211126 3324
rect 218054 3272 218060 3324
rect 218112 3312 218118 3324
rect 219342 3312 219348 3324
rect 218112 3284 219348 3312
rect 218112 3272 218118 3284
rect 219342 3272 219348 3284
rect 219400 3272 219406 3324
rect 314672 3312 314700 3420
rect 339402 3408 339408 3460
rect 339460 3448 339466 3460
rect 350445 3451 350503 3457
rect 350445 3448 350457 3451
rect 339460 3420 350457 3448
rect 339460 3408 339466 3420
rect 350445 3417 350457 3420
rect 350491 3417 350503 3451
rect 350445 3411 350503 3417
rect 346302 3340 346308 3392
rect 346360 3380 346366 3392
rect 350552 3380 350580 3488
rect 407298 3476 407304 3488
rect 407356 3476 407362 3528
rect 415302 3476 415308 3528
rect 415360 3516 415366 3528
rect 475102 3516 475108 3528
rect 415360 3488 475108 3516
rect 415360 3476 415366 3488
rect 475102 3476 475108 3488
rect 475160 3476 475166 3528
rect 494054 3476 494060 3528
rect 494112 3516 494118 3528
rect 495342 3516 495348 3528
rect 494112 3488 495348 3516
rect 494112 3476 494118 3488
rect 495342 3476 495348 3488
rect 495400 3476 495406 3528
rect 507762 3476 507768 3528
rect 507820 3516 507826 3528
rect 567838 3516 567844 3528
rect 507820 3488 567844 3516
rect 507820 3476 507826 3488
rect 567838 3476 567844 3488
rect 567896 3476 567902 3528
rect 571426 3476 571432 3528
rect 571484 3516 571490 3528
rect 572622 3516 572628 3528
rect 571484 3488 572628 3516
rect 571484 3476 571490 3488
rect 572622 3476 572628 3488
rect 572680 3476 572686 3528
rect 574738 3476 574744 3528
rect 574796 3516 574802 3528
rect 576210 3516 576216 3528
rect 574796 3488 576216 3516
rect 574796 3476 574802 3488
rect 576210 3476 576216 3488
rect 576268 3476 576274 3528
rect 350629 3451 350687 3457
rect 350629 3417 350641 3451
rect 350675 3448 350687 3451
rect 400214 3448 400220 3460
rect 350675 3420 400220 3448
rect 350675 3417 350687 3420
rect 350629 3411 350687 3417
rect 400214 3408 400220 3420
rect 400272 3408 400278 3460
rect 422202 3408 422208 3460
rect 422260 3448 422266 3460
rect 482278 3448 482284 3460
rect 422260 3420 482284 3448
rect 422260 3408 422266 3420
rect 482278 3408 482284 3420
rect 482336 3408 482342 3460
rect 518802 3408 518808 3460
rect 518860 3448 518866 3460
rect 578602 3448 578608 3460
rect 518860 3420 578608 3448
rect 518860 3408 518866 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 346360 3352 350580 3380
rect 346360 3340 346366 3352
rect 354582 3340 354588 3392
rect 354640 3380 354646 3392
rect 414474 3380 414480 3392
rect 354640 3352 414480 3380
rect 354640 3340 354646 3352
rect 414474 3340 414480 3352
rect 414532 3340 414538 3392
rect 425054 3340 425060 3392
rect 425112 3380 425118 3392
rect 426342 3380 426348 3392
rect 425112 3352 426348 3380
rect 425112 3340 425118 3352
rect 426342 3340 426348 3352
rect 426400 3340 426406 3392
rect 453942 3340 453948 3392
rect 454000 3380 454006 3392
rect 514386 3380 514392 3392
rect 454000 3352 514392 3380
rect 454000 3340 454006 3352
rect 514386 3340 514392 3352
rect 514444 3340 514450 3392
rect 517422 3340 517428 3392
rect 517480 3380 517486 3392
rect 577406 3380 577412 3392
rect 517480 3352 577412 3380
rect 517480 3340 517486 3352
rect 577406 3340 577412 3352
rect 577464 3340 577470 3392
rect 375190 3312 375196 3324
rect 314672 3284 375196 3312
rect 375190 3272 375196 3284
rect 375248 3272 375254 3324
rect 386322 3272 386328 3324
rect 386380 3312 386386 3324
rect 446582 3312 446588 3324
rect 386380 3284 446588 3312
rect 386380 3272 386386 3284
rect 446582 3272 446588 3284
rect 446640 3272 446646 3324
rect 458082 3272 458088 3324
rect 458140 3312 458146 3324
rect 517882 3312 517888 3324
rect 458140 3284 517888 3312
rect 458140 3272 458146 3284
rect 517882 3272 517888 3284
rect 517940 3272 517946 3324
rect 528557 3315 528615 3321
rect 528557 3281 528569 3315
rect 528603 3312 528615 3315
rect 532234 3312 532240 3324
rect 528603 3284 532240 3312
rect 528603 3281 528615 3284
rect 528557 3275 528615 3281
rect 532234 3272 532240 3284
rect 532292 3272 532298 3324
rect 118602 3204 118608 3256
rect 118660 3244 118666 3256
rect 178954 3244 178960 3256
rect 118660 3216 178960 3244
rect 118660 3204 118666 3216
rect 178954 3204 178960 3216
rect 179012 3204 179018 3256
rect 179322 3204 179328 3256
rect 179380 3244 179386 3256
rect 239582 3244 239588 3256
rect 179380 3216 239588 3244
rect 179380 3204 179386 3216
rect 239582 3204 239588 3216
rect 239640 3204 239646 3256
rect 365714 3204 365720 3256
rect 365772 3244 365778 3256
rect 366910 3244 366916 3256
rect 365772 3216 366916 3244
rect 365772 3204 365778 3216
rect 366910 3204 366916 3216
rect 366968 3204 366974 3256
rect 379422 3204 379428 3256
rect 379480 3244 379486 3256
rect 439406 3244 439412 3256
rect 379480 3216 439412 3244
rect 379480 3204 379486 3216
rect 439406 3204 439412 3216
rect 439464 3204 439470 3256
rect 440142 3204 440148 3256
rect 440200 3244 440206 3256
rect 500126 3244 500132 3256
rect 440200 3216 500132 3244
rect 440200 3204 440206 3216
rect 500126 3204 500132 3216
rect 500184 3204 500190 3256
rect 511902 3204 511908 3256
rect 511960 3244 511966 3256
rect 571426 3244 571432 3256
rect 511960 3216 571432 3244
rect 511960 3204 511966 3216
rect 571426 3204 571432 3216
rect 571484 3204 571490 3256
rect 100662 3136 100668 3188
rect 100720 3176 100726 3188
rect 161106 3176 161112 3188
rect 100720 3148 161112 3176
rect 100720 3136 100726 3148
rect 161106 3136 161112 3148
rect 161164 3136 161170 3188
rect 204162 3136 204168 3188
rect 204220 3176 204226 3188
rect 264606 3176 264612 3188
rect 204220 3148 264612 3176
rect 204220 3136 204226 3148
rect 264606 3136 264612 3148
rect 264664 3136 264670 3188
rect 325602 3136 325608 3188
rect 325660 3176 325666 3188
rect 385862 3176 385868 3188
rect 325660 3148 385868 3176
rect 325660 3136 325666 3148
rect 385862 3136 385868 3148
rect 385920 3136 385926 3188
rect 436002 3136 436008 3188
rect 436060 3176 436066 3188
rect 496538 3176 496544 3188
rect 436060 3148 496544 3176
rect 436060 3136 436066 3148
rect 496538 3136 496544 3148
rect 496596 3136 496602 3188
rect 513282 3136 513288 3188
rect 513340 3176 513346 3188
rect 573818 3176 573824 3188
rect 513340 3148 573824 3176
rect 513340 3136 513346 3148
rect 573818 3136 573824 3148
rect 573876 3136 573882 3188
rect 107562 3068 107568 3120
rect 107620 3108 107626 3120
rect 168190 3108 168196 3120
rect 107620 3080 168196 3108
rect 107620 3068 107626 3080
rect 168190 3068 168196 3080
rect 168248 3068 168254 3120
rect 186222 3068 186228 3120
rect 186280 3108 186286 3120
rect 246758 3108 246764 3120
rect 186280 3080 246764 3108
rect 186280 3068 186286 3080
rect 246758 3068 246764 3080
rect 246816 3068 246822 3120
rect 447042 3068 447048 3120
rect 447100 3108 447106 3120
rect 507210 3108 507216 3120
rect 447100 3080 507216 3108
rect 447100 3068 447106 3080
rect 507210 3068 507216 3080
rect 507268 3068 507274 3120
rect 99282 3000 99288 3052
rect 99340 3040 99346 3052
rect 159910 3040 159916 3052
rect 99340 3012 159916 3040
rect 99340 3000 99346 3012
rect 159910 3000 159916 3012
rect 159968 3000 159974 3052
rect 445113 2975 445171 2981
rect 445113 2941 445125 2975
rect 445159 2972 445171 2975
rect 451274 2972 451280 2984
rect 445159 2944 451280 2972
rect 445159 2941 445171 2944
rect 445113 2935 445171 2941
rect 451274 2932 451280 2944
rect 451332 2932 451338 2984
rect 427906 2796 427912 2848
rect 427964 2836 427970 2848
rect 427964 2808 428780 2836
rect 427964 2796 427970 2808
rect 428752 2780 428780 2808
rect 434806 2796 434812 2848
rect 434864 2836 434870 2848
rect 434864 2808 435864 2836
rect 434864 2796 434870 2808
rect 435836 2780 435864 2808
rect 428734 2728 428740 2780
rect 428792 2728 428798 2780
rect 435818 2728 435824 2780
rect 435876 2728 435882 2780
rect 301314 552 301320 604
rect 301372 592 301378 604
rect 301406 592 301412 604
rect 301372 564 301412 592
rect 301372 552 301378 564
rect 301406 552 301412 564
rect 301464 552 301470 604
rect 354674 552 354680 604
rect 354732 592 354738 604
rect 354950 592 354956 604
rect 354732 564 354956 592
rect 354732 552 354738 564
rect 354950 552 354956 564
rect 355008 552 355014 604
rect 357434 552 357440 604
rect 357492 592 357498 604
rect 358538 592 358544 604
rect 357492 564 358544 592
rect 357492 552 357498 564
rect 358538 552 358544 564
rect 358596 552 358602 604
rect 358814 552 358820 604
rect 358872 592 358878 604
rect 359734 592 359740 604
rect 358872 564 359740 592
rect 358872 552 358878 564
rect 359734 552 359740 564
rect 359792 552 359798 604
rect 361574 552 361580 604
rect 361632 592 361638 604
rect 362126 592 362132 604
rect 361632 564 362132 592
rect 361632 552 361638 564
rect 362126 552 362132 564
rect 362184 552 362190 604
rect 431126 592 431132 604
rect 431087 564 431132 592
rect 431126 552 431132 564
rect 431184 552 431190 604
rect 437014 592 437020 604
rect 436975 564 437020 592
rect 437014 552 437020 564
rect 437072 552 437078 604
rect 461026 552 461032 604
rect 461084 592 461090 604
rect 462038 592 462044 604
rect 461084 564 462044 592
rect 461084 552 461090 564
rect 462038 552 462044 564
rect 462096 552 462102 604
rect 462314 552 462320 604
rect 462372 592 462378 604
rect 463234 592 463240 604
rect 462372 564 463240 592
rect 462372 552 462378 564
rect 463234 552 463240 564
rect 463292 552 463298 604
rect 463786 552 463792 604
rect 463844 592 463850 604
rect 464430 592 464436 604
rect 463844 564 464436 592
rect 463844 552 463850 564
rect 464430 552 464436 564
rect 464488 552 464494 604
rect 465074 552 465080 604
rect 465132 592 465138 604
rect 465626 592 465632 604
rect 465132 564 465632 592
rect 465132 552 465138 564
rect 465626 552 465632 564
rect 465684 552 465690 604
rect 466454 552 466460 604
rect 466512 592 466518 604
rect 466822 592 466828 604
rect 466512 564 466828 592
rect 466512 552 466518 564
rect 466822 552 466828 564
rect 466880 552 466886 604
rect 469214 552 469220 604
rect 469272 592 469278 604
rect 470318 592 470324 604
rect 469272 564 470324 592
rect 469272 552 469278 564
rect 470318 552 470324 564
rect 470376 552 470382 604
<< via1 >>
rect 411168 700408 411220 700460
rect 429844 700408 429896 700460
rect 463608 700408 463660 700460
rect 494796 700408 494848 700460
rect 514668 700408 514720 700460
rect 559656 700408 559708 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 394608 700340 394660 700392
rect 413652 700340 413704 700392
rect 445668 700340 445720 700392
rect 478512 700340 478564 700392
rect 496728 700340 496780 700392
rect 543464 700340 543516 700392
rect 343548 700272 343600 700324
rect 348792 700272 348844 700324
rect 378048 700272 378100 700324
rect 397460 700272 397512 700324
rect 429108 700272 429160 700324
rect 462320 700272 462372 700324
rect 480168 700272 480220 700324
rect 527180 700272 527232 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 326988 699660 327040 699712
rect 332508 699660 332560 699712
rect 360108 699660 360160 699712
rect 364984 699660 365036 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 523776 696940 523828 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 692724 72752 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 523684 685856 523736 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 683247 72568 683256
rect 72516 683213 72525 683247
rect 72525 683213 72559 683247
rect 72559 683213 72568 683247
rect 72516 683204 72568 683213
rect 72516 683068 72568 683120
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 219072 678988 219124 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 218980 678920 219032 678972
rect 72700 678895 72752 678904
rect 72700 678861 72709 678895
rect 72709 678861 72743 678895
rect 72743 678861 72752 678895
rect 72700 678852 72752 678861
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 72700 669264 72752 669316
rect 72884 669264 72936 669316
rect 218980 669264 219032 669316
rect 219164 669264 219216 669316
rect 72884 666476 72936 666528
rect 219164 666476 219216 666528
rect 72792 656931 72844 656940
rect 72792 656897 72801 656931
rect 72801 656897 72835 656931
rect 72835 656897 72844 656931
rect 72792 656888 72844 656897
rect 219072 656931 219124 656940
rect 219072 656897 219081 656931
rect 219081 656897 219115 656931
rect 219115 656897 219124 656931
rect 219072 656888 219124 656897
rect 377128 655460 377180 655512
rect 378048 655460 378100 655512
rect 428188 655460 428240 655512
rect 429108 655460 429160 655512
rect 462320 655460 462372 655512
rect 463608 655460 463660 655512
rect 479340 655460 479392 655512
rect 480168 655460 480220 655512
rect 513380 655256 513432 655308
rect 514668 655256 514720 655308
rect 325976 655120 326028 655172
rect 326988 655120 327040 655172
rect 154304 654984 154356 655036
rect 189724 654984 189776 655036
rect 41328 654916 41380 654968
rect 104532 654916 104584 654968
rect 106188 654916 106240 654968
rect 155592 654916 155644 654968
rect 24768 654848 24820 654900
rect 87512 654848 87564 654900
rect 89628 654848 89680 654900
rect 138572 654848 138624 654900
rect 171048 654848 171100 654900
rect 206744 654848 206796 654900
rect 219072 654848 219124 654900
rect 240784 654848 240836 654900
rect 8024 654780 8076 654832
rect 70492 654780 70544 654832
rect 72792 654780 72844 654832
rect 121552 654780 121604 654832
rect 137744 654780 137796 654832
rect 172704 654780 172756 654832
rect 202788 654780 202840 654832
rect 223764 654780 223816 654832
rect 235908 654780 235960 654832
rect 257896 654780 257948 654832
rect 267648 654780 267700 654832
rect 274916 654780 274968 654832
rect 284024 654780 284076 654832
rect 291936 654780 291988 654832
rect 300768 654100 300820 654152
rect 308956 654100 309008 654152
rect 3516 645804 3568 645856
rect 59360 645804 59412 645856
rect 523776 638936 523828 638988
rect 580172 638936 580224 638988
rect 3424 630572 3476 630624
rect 59360 630572 59412 630624
rect 524328 619556 524380 619608
rect 580264 619556 580316 619608
rect 3608 616768 3660 616820
rect 59360 616768 59412 616820
rect 523132 605752 523184 605804
rect 580448 605752 580500 605804
rect 3516 603032 3568 603084
rect 59360 603032 59412 603084
rect 523684 592016 523736 592068
rect 579804 592016 579856 592068
rect 3424 587800 3476 587852
rect 59360 587800 59412 587852
rect 524328 579572 524380 579624
rect 580356 579572 580408 579624
rect 3516 573996 3568 574048
rect 59360 573996 59412 574048
rect 523132 565768 523184 565820
rect 580448 565768 580500 565820
rect 3424 560192 3476 560244
rect 59360 560192 59412 560244
rect 523776 556180 523828 556232
rect 580172 556180 580224 556232
rect 523500 545096 523552 545148
rect 580172 545096 580224 545148
rect 3424 545028 3476 545080
rect 59360 545028 59412 545080
rect 523684 539520 523736 539572
rect 580264 539520 580316 539572
rect 3424 531224 3476 531276
rect 59360 531224 59412 531276
rect 3148 510552 3200 510604
rect 59360 510552 59412 510604
rect 523776 509260 523828 509312
rect 580172 509260 580224 509312
rect 523684 499468 523736 499520
rect 580264 499468 580316 499520
rect 523684 498176 523736 498228
rect 580172 498176 580224 498228
rect 3424 496748 3476 496800
rect 60004 496748 60056 496800
rect 3516 481584 3568 481636
rect 59360 481584 59412 481636
rect 523684 462340 523736 462392
rect 580172 462340 580224 462392
rect 524328 459484 524380 459536
rect 580264 459484 580316 459536
rect 3424 452548 3476 452600
rect 60004 452548 60056 452600
rect 523776 451256 523828 451308
rect 580172 451256 580224 451308
rect 523684 438880 523736 438932
rect 580172 438880 580224 438932
rect 3148 438812 3200 438864
rect 60096 438812 60148 438864
rect 3240 425008 3292 425060
rect 60004 425008 60056 425060
rect 523684 415420 523736 415472
rect 580172 415420 580224 415472
rect 523776 404336 523828 404388
rect 580172 404336 580224 404388
rect 3148 395972 3200 396024
rect 60096 395972 60148 396024
rect 523684 391960 523736 392012
rect 580172 391960 580224 392012
rect 3240 380808 3292 380860
rect 60188 380808 60240 380860
rect 524236 368500 524288 368552
rect 580172 368500 580224 368552
rect 3148 367004 3200 367056
rect 60004 367004 60056 367056
rect 523684 357416 523736 357468
rect 580172 357416 580224 357468
rect 523776 345040 523828 345092
rect 580172 345040 580224 345092
rect 3424 338036 3476 338088
rect 60096 338036 60148 338088
rect 3240 324232 3292 324284
rect 60188 324232 60240 324284
rect 524328 322872 524380 322924
rect 580172 322872 580224 322924
rect 524328 311788 524380 311840
rect 580172 311788 580224 311840
rect 3332 309068 3384 309120
rect 60004 309068 60056 309120
rect 524328 298732 524380 298784
rect 580172 298732 580224 298784
rect 3424 295264 3476 295316
rect 60372 295264 60424 295316
rect 3424 280100 3476 280152
rect 60096 280100 60148 280152
rect 523684 275952 523736 276004
rect 580172 275952 580224 276004
rect 3148 266296 3200 266348
rect 60280 266296 60332 266348
rect 523684 264868 523736 264920
rect 580172 264868 580224 264920
rect 3424 252492 3476 252544
rect 60464 252492 60516 252544
rect 523684 252492 523736 252544
rect 579804 252492 579856 252544
rect 3424 237328 3476 237380
rect 60004 237328 60056 237380
rect 523684 229032 523736 229084
rect 580172 229032 580224 229084
rect 3148 223524 3200 223576
rect 60188 223524 60240 223576
rect 523776 217948 523828 218000
rect 580172 217948 580224 218000
rect 3424 208292 3476 208344
rect 60096 208292 60148 208344
rect 523868 205572 523920 205624
rect 579804 205572 579856 205624
rect 3148 194488 3200 194540
rect 60280 194488 60332 194540
rect 523684 182112 523736 182164
rect 580172 182112 580224 182164
rect 3240 180752 3292 180804
rect 60372 180752 60424 180804
rect 523776 171028 523828 171080
rect 580172 171028 580224 171080
rect 3516 165520 3568 165572
rect 60188 165520 60240 165572
rect 523868 158652 523920 158704
rect 579804 158652 579856 158704
rect 3148 151716 3200 151768
rect 60096 151716 60148 151768
rect 3240 136552 3292 136604
rect 60004 136552 60056 136604
rect 523684 135192 523736 135244
rect 580172 135192 580224 135244
rect 523776 124108 523828 124160
rect 580172 124108 580224 124160
rect 3424 122748 3476 122800
rect 60372 122748 60424 122800
rect 523868 111732 523920 111784
rect 579804 111732 579856 111784
rect 3240 108944 3292 108996
rect 60280 108944 60332 108996
rect 3424 93780 3476 93832
rect 60188 93780 60240 93832
rect 523684 88272 523736 88324
rect 580172 88272 580224 88324
rect 3424 79976 3476 80028
rect 60004 79976 60056 80028
rect 523776 77188 523828 77240
rect 580172 77188 580224 77240
rect 3332 64812 3384 64864
rect 60096 64812 60148 64864
rect 523868 64812 523920 64864
rect 579804 64812 579856 64864
rect 3424 51008 3476 51060
rect 60280 51008 60332 51060
rect 82820 49648 82872 49700
rect 84844 49648 84896 49700
rect 169760 49648 169812 49700
rect 172336 49648 172388 49700
rect 354496 49648 354548 49700
rect 355324 49648 355376 49700
rect 383108 49648 383160 49700
rect 384304 49648 384356 49700
rect 400956 49648 401008 49700
rect 403624 49648 403676 49700
rect 440332 49648 440384 49700
rect 442264 49648 442316 49700
rect 477224 49648 477276 49700
rect 482284 49648 482336 49700
rect 81624 49308 81676 49360
rect 142252 49308 142304 49360
rect 74448 49240 74500 49292
rect 135444 49240 135496 49292
rect 396172 49240 396224 49292
rect 456892 49240 456944 49292
rect 88708 49172 88760 49224
rect 150624 49172 150676 49224
rect 210332 49172 210384 49224
rect 270500 49172 270552 49224
rect 281816 49172 281868 49224
rect 308404 49172 308456 49224
rect 309232 49172 309284 49224
rect 319444 49172 319496 49224
rect 403348 49172 403400 49224
rect 463792 49172 463844 49224
rect 489184 49172 489236 49224
rect 549260 49172 549312 49224
rect 95884 49104 95936 49156
rect 157432 49104 157484 49156
rect 167368 49104 167420 49156
rect 227904 49104 227956 49156
rect 253204 49104 253256 49156
rect 313464 49104 313516 49156
rect 367652 49104 367704 49156
rect 474832 49104 474884 49156
rect 535460 49104 535512 49156
rect 103060 49036 103112 49088
rect 164332 49036 164384 49088
rect 217416 49036 217468 49088
rect 296076 49036 296128 49088
rect 333244 49036 333296 49088
rect 374736 49036 374788 49088
rect 451004 49036 451056 49088
rect 451924 49036 451976 49088
rect 482008 49036 482060 49088
rect 542360 49036 542412 49088
rect 67272 48968 67324 49020
rect 128452 48968 128504 49020
rect 145932 48968 145984 49020
rect 207112 48968 207164 49020
rect 224592 48968 224644 49020
rect 285772 48968 285824 49020
rect 318708 48968 318760 49020
rect 374644 48968 374696 49020
rect 389088 48968 389140 49020
rect 449900 48968 449952 49020
rect 467748 48968 467800 49020
rect 528560 48968 528612 49020
rect 66076 48764 66128 48816
rect 66904 48764 66956 48816
rect 70860 48764 70912 48816
rect 71688 48764 71740 48816
rect 72056 48764 72108 48816
rect 73068 48764 73120 48816
rect 73252 48764 73304 48816
rect 74448 48764 74500 48816
rect 76840 48764 76892 48816
rect 77944 48764 77996 48816
rect 80428 48764 80480 48816
rect 82084 48764 82136 48816
rect 89904 48764 89956 48816
rect 91008 48764 91060 48816
rect 91100 48764 91152 48816
rect 92296 48764 92348 48816
rect 97080 48764 97132 48816
rect 97908 48764 97960 48816
rect 98276 48764 98328 48816
rect 99288 48764 99340 48816
rect 99472 48764 99524 48816
rect 100668 48764 100720 48816
rect 105452 48764 105504 48816
rect 106188 48764 106240 48816
rect 106648 48764 106700 48816
rect 107568 48764 107620 48816
rect 107844 48764 107896 48816
rect 108948 48764 109000 48816
rect 109040 48764 109092 48816
rect 110236 48764 110288 48816
rect 113732 48764 113784 48816
rect 114468 48764 114520 48816
rect 114928 48764 114980 48816
rect 115848 48764 115900 48816
rect 116124 48764 116176 48816
rect 117228 48764 117280 48816
rect 117320 48764 117372 48816
rect 118608 48764 118660 48816
rect 124496 48764 124548 48816
rect 125508 48764 125560 48816
rect 132868 48764 132920 48816
rect 133788 48764 133840 48816
rect 134064 48764 134116 48816
rect 135168 48764 135220 48816
rect 135260 48764 135312 48816
rect 136456 48764 136508 48816
rect 141148 48764 141200 48816
rect 142068 48764 142120 48816
rect 142344 48764 142396 48816
rect 143448 48764 143500 48816
rect 143540 48764 143592 48816
rect 144828 48764 144880 48816
rect 149520 48764 149572 48816
rect 150348 48764 150400 48816
rect 150716 48764 150768 48816
rect 151728 48764 151780 48816
rect 151912 48764 151964 48816
rect 153844 48764 153896 48816
rect 157892 48764 157944 48816
rect 158628 48764 158680 48816
rect 159088 48764 159140 48816
rect 160008 48764 160060 48816
rect 160284 48764 160336 48816
rect 161388 48764 161440 48816
rect 166172 48764 166224 48816
rect 167736 48764 167788 48816
rect 168564 48764 168616 48816
rect 169668 48764 169720 48816
rect 176936 48764 176988 48816
rect 177948 48764 178000 48816
rect 178132 48764 178184 48816
rect 179328 48764 179380 48816
rect 185308 48764 185360 48816
rect 186228 48764 186280 48816
rect 186504 48764 186556 48816
rect 187608 48764 187660 48816
rect 187700 48764 187752 48816
rect 189724 48764 189776 48816
rect 193588 48764 193640 48816
rect 194508 48764 194560 48816
rect 201960 48764 202012 48816
rect 202788 48764 202840 48816
rect 203156 48764 203208 48816
rect 204168 48764 204220 48816
rect 204352 48764 204404 48816
rect 205548 48764 205600 48816
rect 212724 48764 212776 48816
rect 213828 48764 213880 48816
rect 213920 48764 213972 48816
rect 215208 48764 215260 48816
rect 218612 48764 218664 48816
rect 219348 48764 219400 48816
rect 219808 48764 219860 48816
rect 220728 48764 220780 48816
rect 221004 48764 221056 48816
rect 222108 48764 222160 48816
rect 222200 48764 222252 48816
rect 223488 48764 223540 48816
rect 228180 48764 228232 48816
rect 229008 48764 229060 48816
rect 229376 48764 229428 48816
rect 230388 48764 230440 48816
rect 235356 48764 235408 48816
rect 236644 48764 236696 48816
rect 237748 48764 237800 48816
rect 238668 48764 238720 48816
rect 238944 48764 238996 48816
rect 240048 48764 240100 48816
rect 240140 48764 240192 48816
rect 241428 48764 241480 48816
rect 246028 48764 246080 48816
rect 246948 48764 247000 48816
rect 247224 48764 247276 48816
rect 248328 48764 248380 48816
rect 254400 48764 254452 48816
rect 255228 48764 255280 48816
rect 255596 48764 255648 48816
rect 256608 48764 256660 48816
rect 256792 48764 256844 48816
rect 257988 48764 258040 48816
rect 260380 48764 260432 48816
rect 261484 48764 261536 48816
rect 265164 48764 265216 48816
rect 266268 48764 266320 48816
rect 266360 48764 266412 48816
rect 267556 48764 267608 48816
rect 272248 48764 272300 48816
rect 273168 48764 273220 48816
rect 273444 48764 273496 48816
rect 274548 48764 274600 48816
rect 274640 48764 274692 48816
rect 276664 48764 276716 48816
rect 280620 48764 280672 48816
rect 281448 48764 281500 48816
rect 283012 48764 283064 48816
rect 284208 48764 284260 48816
rect 290188 48764 290240 48816
rect 291108 48764 291160 48816
rect 298468 48764 298520 48816
rect 299388 48764 299440 48816
rect 299664 48764 299716 48816
rect 301504 48764 301556 48816
rect 308036 48764 308088 48816
rect 309048 48764 309100 48816
rect 316408 48764 316460 48816
rect 317328 48764 317380 48816
rect 323492 48764 323544 48816
rect 324228 48764 324280 48816
rect 324688 48764 324740 48816
rect 325608 48764 325660 48816
rect 325884 48764 325936 48816
rect 326988 48764 327040 48816
rect 327080 48764 327132 48816
rect 328276 48764 328328 48816
rect 329472 48764 329524 48816
rect 330484 48764 330536 48816
rect 333060 48764 333112 48816
rect 333888 48764 333940 48816
rect 335452 48764 335504 48816
rect 336648 48764 336700 48816
rect 343732 48764 343784 48816
rect 344928 48764 344980 48816
rect 347320 48764 347372 48816
rect 348424 48764 348476 48816
rect 350908 48764 350960 48816
rect 351828 48764 351880 48816
rect 353300 48764 353352 48816
rect 354588 48764 354640 48816
rect 359280 48764 359332 48816
rect 360108 48764 360160 48816
rect 361672 48764 361724 48816
rect 362868 48764 362920 48816
rect 369952 48764 370004 48816
rect 371056 48764 371108 48816
rect 375932 48764 375984 48816
rect 376668 48764 376720 48816
rect 378324 48764 378376 48816
rect 379428 48764 379480 48816
rect 379520 48764 379572 48816
rect 380808 48764 380860 48816
rect 385500 48764 385552 48816
rect 386328 48764 386380 48816
rect 386696 48764 386748 48816
rect 387708 48764 387760 48816
rect 387892 48764 387944 48816
rect 389088 48764 389140 48816
rect 394976 48764 395028 48816
rect 395988 48764 396040 48816
rect 404544 48764 404596 48816
rect 405648 48764 405700 48816
rect 412916 48764 412968 48816
rect 413928 48764 413980 48816
rect 414112 48764 414164 48816
rect 415308 48764 415360 48816
rect 420092 48764 420144 48816
rect 420828 48764 420880 48816
rect 421196 48764 421248 48816
rect 422208 48764 422260 48816
rect 422392 48764 422444 48816
rect 423588 48764 423640 48816
rect 428372 48764 428424 48816
rect 429108 48764 429160 48816
rect 429568 48764 429620 48816
rect 430488 48764 430540 48816
rect 430764 48764 430816 48816
rect 431868 48764 431920 48816
rect 433156 48764 433208 48816
rect 433984 48764 434036 48816
rect 437940 48764 437992 48816
rect 438768 48764 438820 48816
rect 439136 48764 439188 48816
rect 440148 48764 440200 48816
rect 446220 48764 446272 48816
rect 447048 48764 447100 48816
rect 447416 48764 447468 48816
rect 448428 48764 448480 48816
rect 448612 48764 448664 48816
rect 449716 48764 449768 48816
rect 455788 48764 455840 48816
rect 456708 48764 456760 48816
rect 456984 48764 457036 48816
rect 458088 48764 458140 48816
rect 459376 48764 459428 48816
rect 460204 48764 460256 48816
rect 464160 48764 464212 48816
rect 464988 48764 465040 48816
rect 465356 48764 465408 48816
rect 466368 48764 466420 48816
rect 466552 48764 466604 48816
rect 467748 48764 467800 48816
rect 473636 48764 473688 48816
rect 474648 48764 474700 48816
rect 480812 48764 480864 48816
rect 481548 48764 481600 48816
rect 483204 48764 483256 48816
rect 484308 48764 484360 48816
rect 484400 48764 484452 48816
rect 485596 48764 485648 48816
rect 491576 48764 491628 48816
rect 492588 48764 492640 48816
rect 492772 48764 492824 48816
rect 493968 48764 494020 48816
rect 495164 48764 495216 48816
rect 496084 48764 496136 48816
rect 498660 48764 498712 48816
rect 499488 48764 499540 48816
rect 499856 48764 499908 48816
rect 500868 48764 500920 48816
rect 501052 48764 501104 48816
rect 502248 48764 502300 48816
rect 508228 48764 508280 48816
rect 509148 48764 509200 48816
rect 509424 48764 509476 48816
rect 510528 48764 510580 48816
rect 516600 48764 516652 48816
rect 517428 48764 517480 48816
rect 517796 48764 517848 48816
rect 518808 48764 518860 48816
rect 518992 48764 519044 48816
rect 520096 48764 520148 48816
rect 64880 48696 64932 48748
rect 66168 48696 66220 48748
rect 123300 48696 123352 48748
rect 124128 48696 124180 48748
rect 161480 48696 161532 48748
rect 167644 48696 167696 48748
rect 262772 48696 262824 48748
rect 263508 48696 263560 48748
rect 263968 48696 264020 48748
rect 265624 48696 265676 48748
rect 271052 48696 271104 48748
rect 272524 48696 272576 48748
rect 288992 48696 289044 48748
rect 290464 48696 290516 48748
rect 306840 48696 306892 48748
rect 312544 48696 312596 48748
rect 334256 48696 334308 48748
rect 335268 48696 335320 48748
rect 360476 48696 360528 48748
rect 361488 48696 361540 48748
rect 431960 48696 432012 48748
rect 433248 48696 433300 48748
rect 436744 48696 436796 48748
rect 438124 48696 438176 48748
rect 458180 48696 458232 48748
rect 459468 48696 459520 48748
rect 472440 48696 472492 48748
rect 474004 48696 474056 48748
rect 487988 48696 488040 48748
rect 489184 48696 489236 48748
rect 125692 48628 125744 48680
rect 126796 48628 126848 48680
rect 195980 48628 196032 48680
rect 197268 48628 197320 48680
rect 278228 48628 278280 48680
rect 280804 48628 280856 48680
rect 292580 48628 292632 48680
rect 293868 48628 293920 48680
rect 365260 48628 365312 48680
rect 367744 48628 367796 48680
rect 175740 48560 175792 48612
rect 176568 48560 176620 48612
rect 315212 48560 315264 48612
rect 315948 48560 316000 48612
rect 248420 48492 248472 48544
rect 249616 48492 249668 48544
rect 300860 48492 300912 48544
rect 302148 48492 302200 48544
rect 342628 48492 342680 48544
rect 343548 48492 343600 48544
rect 510620 48492 510672 48544
rect 511908 48492 511960 48544
rect 352104 48424 352156 48476
rect 353208 48424 353260 48476
rect 411720 48424 411772 48476
rect 412548 48424 412600 48476
rect 293684 48356 293736 48408
rect 294604 48356 294656 48408
rect 211528 48288 211580 48340
rect 212448 48288 212500 48340
rect 278964 48331 279016 48340
rect 278964 48297 278973 48331
rect 278973 48297 279007 48331
rect 279007 48297 279016 48331
rect 278964 48288 279016 48297
rect 317604 48288 317656 48340
rect 318708 48288 318760 48340
rect 368848 48288 368900 48340
rect 369768 48288 369820 48340
rect 377128 48288 377180 48340
rect 378048 48288 378100 48340
rect 427912 48331 427964 48340
rect 427912 48297 427921 48331
rect 427921 48297 427955 48331
rect 427955 48297 427964 48331
rect 427912 48288 427964 48297
rect 434812 48331 434864 48340
rect 434812 48297 434821 48331
rect 434821 48297 434855 48331
rect 434855 48297 434864 48331
rect 434812 48288 434864 48297
rect 194784 47676 194836 47728
rect 255320 47676 255372 47728
rect 136548 47608 136600 47660
rect 197360 47608 197412 47660
rect 275836 47608 275888 47660
rect 336740 47608 336792 47660
rect 94688 47540 94740 47592
rect 155960 47540 156012 47592
rect 242440 47540 242492 47592
rect 303620 47540 303672 47592
rect 336832 47540 336884 47592
rect 397460 47540 397512 47592
rect 425980 47540 426032 47592
rect 485780 47540 485832 47592
rect 490380 47540 490432 47592
rect 550640 47540 550692 47592
rect 285772 46903 285824 46912
rect 285772 46869 285781 46903
rect 285781 46869 285815 46903
rect 285815 46869 285824 46903
rect 285772 46860 285824 46869
rect 172336 46248 172388 46300
rect 230480 46248 230532 46300
rect 291384 46248 291436 46300
rect 351920 46248 351972 46300
rect 443920 46248 443972 46300
rect 503720 46248 503772 46300
rect 112628 46180 112680 46232
rect 173900 46180 173952 46232
rect 230572 46180 230624 46232
rect 291200 46180 291252 46232
rect 344836 46180 344888 46232
rect 405740 46180 405792 46232
rect 406016 46180 406068 46232
rect 466460 46180 466512 46232
rect 504640 46180 504692 46232
rect 564440 46180 564492 46232
rect 238668 44888 238720 44940
rect 298100 44888 298152 44940
rect 349068 44888 349120 44940
rect 408500 44888 408552 44940
rect 117228 44820 117280 44872
rect 176660 44820 176712 44872
rect 177948 44820 178000 44872
rect 237380 44820 237432 44872
rect 295248 44820 295300 44872
rect 356060 44820 356112 44872
rect 415216 44820 415268 44872
rect 476120 44820 476172 44872
rect 480168 44820 480220 44872
rect 539600 44820 539652 44872
rect 135168 43460 135220 43512
rect 194600 43460 194652 43512
rect 249616 43460 249668 43512
rect 309140 43460 309192 43512
rect 355968 43460 356020 43512
rect 416872 43460 416924 43512
rect 191748 43392 191800 43444
rect 252652 43392 252704 43444
rect 302056 43392 302108 43444
rect 362960 43392 363012 43444
rect 402888 43392 402940 43444
rect 462320 43392 462372 43444
rect 493876 43392 493928 43444
rect 554780 43392 554832 43444
rect 202788 42100 202840 42152
rect 262220 42100 262272 42152
rect 263508 42100 263560 42152
rect 322940 42100 322992 42152
rect 84108 42032 84160 42084
rect 144920 42032 144972 42084
rect 148968 42032 149020 42084
rect 209872 42032 209924 42084
rect 320088 42032 320140 42084
rect 380900 42032 380952 42084
rect 419448 42032 419500 42084
rect 478880 42032 478932 42084
rect 498108 42032 498160 42084
rect 557540 42032 557592 42084
rect 523684 41352 523736 41404
rect 580172 41352 580224 41404
rect 220728 40740 220780 40792
rect 280160 40740 280212 40792
rect 331128 40740 331180 40792
rect 390560 40740 390612 40792
rect 88248 40672 88300 40724
rect 149060 40672 149112 40724
rect 162768 40672 162820 40724
rect 223580 40672 223632 40724
rect 277308 40672 277360 40724
rect 338120 40672 338172 40724
rect 391848 40672 391900 40724
rect 451280 40672 451332 40724
rect 274548 39380 274600 39432
rect 333980 39380 334032 39432
rect 384948 39380 385000 39432
rect 444380 39380 444432 39432
rect 82084 39312 82136 39364
rect 140780 39312 140832 39364
rect 153844 39312 153896 39364
rect 212540 39312 212592 39364
rect 213828 39312 213880 39364
rect 273260 39312 273312 39364
rect 328276 39312 328328 39364
rect 387800 39312 387852 39364
rect 420828 39312 420880 39364
rect 480260 39312 480312 39364
rect 509148 39312 509200 39364
rect 568580 39312 568632 39364
rect 427912 38607 427964 38616
rect 427912 38573 427921 38607
rect 427921 38573 427955 38607
rect 427955 38573 427964 38607
rect 427912 38564 427964 38573
rect 434812 38607 434864 38616
rect 434812 38573 434821 38607
rect 434821 38573 434855 38607
rect 434855 38573 434864 38607
rect 434812 38564 434864 38573
rect 142068 37952 142120 38004
rect 201500 37952 201552 38004
rect 256608 37952 256660 38004
rect 316040 37952 316092 38004
rect 413928 37952 413980 38004
rect 473360 37952 473412 38004
rect 77944 37884 77996 37936
rect 138020 37884 138072 37936
rect 198648 37884 198700 37936
rect 259460 37884 259512 37936
rect 313188 37884 313240 37936
rect 374092 37884 374144 37936
rect 380716 37884 380768 37936
rect 441620 37884 441672 37936
rect 511816 37884 511868 37936
rect 571432 37884 571484 37936
rect 285772 37315 285824 37324
rect 285772 37281 285781 37315
rect 285781 37281 285815 37315
rect 285815 37281 285824 37315
rect 285772 37272 285824 37281
rect 353208 36660 353260 36712
rect 412640 36660 412692 36712
rect 189724 36592 189776 36644
rect 248420 36592 248472 36644
rect 299388 36592 299440 36644
rect 358820 36592 358872 36644
rect 137928 36524 137980 36576
rect 198740 36524 198792 36576
rect 245568 36524 245620 36576
rect 305000 36524 305052 36576
rect 398748 36524 398800 36576
rect 459652 36524 459704 36576
rect 516048 36524 516100 36576
rect 574744 36524 574796 36576
rect 3424 35844 3476 35896
rect 60188 35844 60240 35896
rect 184848 35232 184900 35284
rect 244280 35232 244332 35284
rect 288348 35232 288400 35284
rect 347780 35232 347832 35284
rect 395988 35232 396040 35284
rect 455420 35232 455472 35284
rect 131028 35164 131080 35216
rect 191840 35164 191892 35216
rect 241336 35164 241388 35216
rect 302240 35164 302292 35216
rect 342168 35164 342220 35216
rect 401600 35164 401652 35216
rect 460204 35164 460256 35216
rect 520372 35164 520424 35216
rect 124128 33804 124180 33856
rect 183560 33804 183612 33856
rect 227628 33804 227680 33856
rect 287060 33804 287112 33856
rect 338028 33804 338080 33856
rect 398840 33804 398892 33856
rect 441528 33804 441580 33856
rect 502432 33804 502484 33856
rect 173808 33736 173860 33788
rect 234620 33736 234672 33788
rect 284116 33736 284168 33788
rect 345020 33736 345072 33788
rect 409788 33736 409840 33788
rect 469220 33736 469272 33788
rect 502156 33736 502208 33788
rect 563152 33736 563204 33788
rect 167736 32444 167788 32496
rect 227812 32444 227864 32496
rect 281448 32444 281500 32496
rect 340880 32444 340932 32496
rect 389088 32444 389140 32496
rect 448520 32444 448572 32496
rect 119988 32376 120040 32428
rect 180800 32376 180852 32428
rect 223396 32376 223448 32428
rect 284300 32376 284352 32428
rect 335268 32376 335320 32428
rect 394700 32376 394752 32428
rect 467748 32376 467800 32428
rect 527180 32376 527232 32428
rect 160008 31084 160060 31136
rect 219440 31084 219492 31136
rect 267556 31084 267608 31136
rect 327080 31084 327132 31136
rect 378048 31084 378100 31136
rect 437480 31084 437532 31136
rect 106188 31016 106240 31068
rect 167092 31016 167144 31068
rect 216588 31016 216640 31068
rect 277400 31016 277452 31068
rect 324228 31016 324280 31068
rect 383660 31016 383712 31068
rect 449716 31016 449768 31068
rect 509240 31016 509292 31068
rect 510528 31016 510580 31068
rect 569960 31016 570012 31068
rect 523776 30268 523828 30320
rect 580172 30268 580224 30320
rect 155868 29656 155920 29708
rect 216680 29656 216732 29708
rect 259368 29656 259420 29708
rect 320180 29656 320232 29708
rect 373908 29656 373960 29708
rect 433340 29656 433392 29708
rect 102048 29588 102100 29640
rect 162860 29588 162912 29640
rect 205456 29588 205508 29640
rect 266360 29588 266412 29640
rect 317328 29588 317380 29640
rect 376760 29588 376812 29640
rect 438768 29588 438820 29640
rect 498200 29588 498252 29640
rect 427912 29019 427964 29028
rect 427912 28985 427921 29019
rect 427921 28985 427955 29019
rect 427955 28985 427964 29019
rect 427912 28976 427964 28985
rect 434812 29019 434864 29028
rect 434812 28985 434821 29019
rect 434821 28985 434855 29019
rect 434855 28985 434864 29019
rect 434812 28976 434864 28985
rect 248420 28908 248472 28960
rect 248512 28908 248564 28960
rect 280804 28364 280856 28416
rect 339500 28364 339552 28416
rect 97908 28296 97960 28348
rect 158812 28296 158864 28348
rect 236644 28296 236696 28348
rect 296720 28296 296772 28348
rect 371056 28296 371108 28348
rect 430580 28296 430632 28348
rect 144736 28228 144788 28280
rect 205640 28228 205692 28280
rect 208308 28228 208360 28280
rect 269120 28228 269172 28280
rect 311808 28228 311860 28280
rect 372620 28228 372672 28280
rect 445668 28228 445720 28280
rect 505100 28228 505152 28280
rect 285772 27591 285824 27600
rect 285772 27557 285781 27591
rect 285781 27557 285815 27591
rect 285815 27557 285824 27591
rect 285772 27548 285824 27557
rect 319444 26936 319496 26988
rect 369860 26936 369912 26988
rect 492588 26936 492640 26988
rect 552020 26936 552072 26988
rect 93768 26868 93820 26920
rect 154580 26868 154632 26920
rect 165528 26868 165580 26920
rect 226340 26868 226392 26920
rect 257896 26868 257948 26920
rect 318800 26868 318852 26920
rect 367008 26868 367060 26920
rect 426440 26868 426492 26920
rect 434628 26868 434680 26920
rect 494060 26868 494112 26920
rect 306288 25576 306340 25628
rect 365720 25576 365772 25628
rect 431868 25576 431920 25628
rect 491300 25576 491352 25628
rect 91008 25508 91060 25560
rect 150532 25508 150584 25560
rect 158628 25508 158680 25560
rect 218060 25508 218112 25560
rect 251088 25508 251140 25560
rect 311900 25508 311952 25560
rect 360108 25508 360160 25560
rect 419540 25508 419592 25560
rect 485596 25508 485648 25560
rect 545120 25508 545172 25560
rect 309048 24216 309100 24268
rect 368480 24216 368532 24268
rect 249708 24148 249760 24200
rect 310520 24148 310572 24200
rect 481548 24148 481600 24200
rect 540980 24148 541032 24200
rect 86868 24080 86920 24132
rect 147680 24080 147732 24132
rect 154488 24080 154540 24132
rect 215300 24080 215352 24132
rect 226248 24080 226300 24132
rect 287152 24080 287204 24132
rect 362776 24080 362828 24132
rect 423680 24080 423732 24132
rect 427728 24080 427780 24132
rect 487160 24080 487212 24132
rect 261484 22788 261536 22840
rect 321560 22788 321612 22840
rect 482284 22788 482336 22840
rect 536840 22788 536892 22840
rect 84844 22720 84896 22772
rect 143540 22720 143592 22772
rect 151728 22720 151780 22772
rect 211160 22720 211212 22772
rect 215116 22720 215168 22772
rect 276020 22720 276072 22772
rect 286968 22720 287020 22772
rect 347872 22720 347924 22772
rect 348424 22720 348476 22772
rect 408592 22720 408644 22772
rect 423496 22720 423548 22772
rect 484400 22720 484452 22772
rect 3148 22040 3200 22092
rect 60004 22040 60056 22092
rect 79968 21360 80020 21412
rect 140872 21360 140924 21412
rect 147588 21360 147640 21412
rect 208400 21360 208452 21412
rect 212448 21360 212500 21412
rect 271880 21360 271932 21412
rect 273168 21360 273220 21412
rect 332600 21360 332652 21412
rect 333888 21360 333940 21412
rect 393320 21360 393372 21412
rect 412548 21360 412600 21412
rect 471980 21360 472032 21412
rect 474648 21360 474700 21412
rect 534080 21360 534132 21412
rect 312544 20000 312596 20052
rect 367100 20000 367152 20052
rect 75828 19932 75880 19984
rect 136640 19932 136692 19984
rect 144828 19932 144880 19984
rect 204260 19932 204312 19984
rect 205548 19932 205600 19984
rect 264980 19932 265032 19984
rect 269028 19932 269080 19984
rect 329840 19932 329892 19984
rect 330484 19932 330536 19984
rect 390652 19932 390704 19984
rect 408408 19932 408460 19984
rect 467840 19932 467892 19984
rect 470508 19932 470560 19984
rect 529940 19932 529992 19984
rect 248420 19295 248472 19304
rect 248420 19261 248429 19295
rect 248429 19261 248463 19295
rect 248463 19261 248472 19295
rect 248420 19252 248472 19261
rect 259460 19295 259512 19304
rect 259460 19261 259469 19295
rect 259469 19261 259503 19295
rect 259503 19261 259512 19295
rect 259460 19252 259512 19261
rect 269120 19295 269172 19304
rect 269120 19261 269129 19295
rect 269129 19261 269163 19295
rect 269163 19261 269172 19295
rect 269120 19252 269172 19261
rect 277400 19252 277452 19304
rect 277768 19252 277820 19304
rect 278964 19295 279016 19304
rect 278964 19261 278973 19295
rect 278973 19261 279007 19295
rect 279007 19261 279016 19295
rect 278964 19252 279016 19261
rect 284300 19295 284352 19304
rect 284300 19261 284309 19295
rect 284309 19261 284343 19295
rect 284343 19261 284352 19295
rect 284300 19252 284352 19261
rect 427912 19295 427964 19304
rect 427912 19261 427921 19295
rect 427921 19261 427955 19295
rect 427955 19261 427964 19295
rect 427912 19252 427964 19261
rect 434812 19295 434864 19304
rect 434812 19261 434821 19295
rect 434821 19261 434855 19295
rect 434855 19261 434864 19295
rect 434812 19252 434864 19261
rect 201408 18640 201460 18692
rect 262312 18640 262364 18692
rect 266268 18640 266320 18692
rect 325700 18640 325752 18692
rect 326988 18640 327040 18692
rect 386420 18640 386472 18692
rect 73068 18572 73120 18624
rect 132592 18572 132644 18624
rect 140688 18572 140740 18624
rect 201592 18572 201644 18624
rect 303528 18572 303580 18624
rect 364340 18572 364392 18624
rect 405648 18572 405700 18624
rect 465080 18572 465132 18624
rect 474004 18572 474056 18624
rect 532700 18572 532752 18624
rect 523868 17892 523920 17944
rect 579804 17892 579856 17944
rect 129648 17280 129700 17332
rect 190460 17280 190512 17332
rect 290464 17280 290516 17332
rect 349160 17280 349212 17332
rect 403624 17280 403676 17332
rect 460940 17280 460992 17332
rect 70308 17212 70360 17264
rect 131120 17212 131172 17264
rect 197176 17212 197228 17264
rect 258080 17212 258132 17264
rect 262128 17212 262180 17264
rect 321652 17212 321704 17264
rect 322848 17212 322900 17264
rect 382372 17212 382424 17264
rect 456708 17212 456760 17264
rect 516140 17212 516192 17264
rect 126796 15920 126848 15972
rect 186320 15920 186372 15972
rect 255228 15920 255280 15972
rect 314660 15920 314712 15972
rect 315948 15920 316000 15972
rect 375380 15920 375432 15972
rect 66904 15852 66956 15904
rect 126980 15852 127032 15904
rect 194508 15852 194560 15904
rect 253940 15852 253992 15904
rect 285588 15852 285640 15904
rect 346400 15852 346452 15904
rect 397368 15852 397420 15904
rect 458180 15852 458232 15904
rect 469128 15852 469180 15904
rect 528652 15852 528704 15904
rect 276664 14560 276716 14612
rect 335360 14560 335412 14612
rect 74448 14492 74500 14544
rect 133880 14492 133932 14544
rect 187608 14492 187660 14544
rect 247040 14492 247092 14544
rect 304908 14492 304960 14544
rect 365812 14492 365864 14544
rect 122748 14424 122800 14476
rect 183652 14424 183704 14476
rect 244188 14424 244240 14476
rect 305092 14424 305144 14476
rect 384304 14424 384356 14476
rect 443092 14424 443144 14476
rect 451924 14424 451976 14476
rect 512000 14424 512052 14476
rect 272524 13200 272576 13252
rect 331220 13200 331272 13252
rect 92296 13132 92348 13184
rect 151820 13132 151872 13184
rect 241428 13132 241480 13184
rect 506388 13132 506440 13184
rect 565820 13132 565872 13184
rect 118516 13064 118568 13116
rect 179420 13064 179472 13116
rect 183468 13064 183520 13116
rect 244372 13064 244424 13116
rect 302148 13064 302200 13116
rect 361580 13064 361632 13116
rect 376668 13064 376720 13116
rect 436100 13064 436152 13116
rect 448428 13064 448480 13116
rect 507860 13064 507912 13116
rect 276020 12452 276072 12504
rect 247040 12384 247092 12436
rect 247960 12384 248012 12436
rect 253940 12384 253992 12436
rect 255044 12384 255096 12436
rect 255320 12384 255372 12436
rect 256240 12384 256292 12436
rect 258080 12384 258132 12436
rect 258632 12384 258684 12436
rect 264980 12384 265032 12436
rect 265808 12384 265860 12436
rect 266360 12384 266412 12436
rect 267004 12384 267056 12436
rect 271880 12384 271932 12436
rect 272892 12384 272944 12436
rect 273260 12384 273312 12436
rect 274088 12384 274140 12436
rect 280160 12384 280212 12436
rect 281264 12384 281316 12436
rect 291200 12384 291252 12436
rect 291936 12384 291988 12436
rect 298100 12384 298152 12436
rect 299112 12384 299164 12436
rect 276480 12316 276532 12368
rect 237288 11772 237340 11824
rect 297916 11772 297968 11824
rect 298008 11772 298060 11824
rect 357440 11772 357492 11824
rect 367744 11772 367796 11824
rect 425060 11772 425112 11824
rect 442264 11772 442316 11824
rect 500960 11772 501012 11824
rect 115848 11704 115900 11756
rect 175372 11704 175424 11756
rect 179236 11704 179288 11756
rect 240140 11704 240192 11756
rect 267648 11704 267700 11756
rect 328460 11704 328512 11756
rect 424968 11704 425020 11756
rect 485872 11704 485924 11756
rect 499488 11704 499540 11756
rect 558920 11704 558972 11756
rect 176568 10344 176620 10396
rect 236092 10344 236144 10396
rect 265624 10344 265676 10396
rect 324320 10344 324372 10396
rect 438124 10344 438176 10396
rect 496820 10344 496872 10396
rect 111708 10276 111760 10328
rect 172520 10276 172572 10328
rect 233148 10276 233200 10328
rect 294328 10276 294380 10328
rect 294604 10276 294656 10328
rect 354680 10276 354732 10328
rect 355324 10276 355376 10328
rect 415400 10276 415452 10328
rect 416688 10276 416740 10328
rect 477592 10276 477644 10328
rect 496084 10276 496136 10328
rect 554872 10276 554924 10328
rect 249156 9664 249208 9716
rect 259828 9664 259880 9716
rect 269304 9664 269356 9716
rect 278964 9707 279016 9716
rect 278964 9673 278973 9707
rect 278973 9673 279007 9707
rect 279007 9673 279016 9707
rect 278964 9664 279016 9673
rect 284760 9664 284812 9716
rect 285956 9664 286008 9716
rect 301412 9707 301464 9716
rect 301412 9673 301421 9707
rect 301421 9673 301455 9707
rect 301455 9673 301464 9707
rect 301412 9664 301464 9673
rect 427912 9707 427964 9716
rect 427912 9673 427921 9707
rect 427921 9673 427955 9707
rect 427955 9673 427964 9707
rect 427912 9664 427964 9673
rect 434812 9707 434864 9716
rect 434812 9673 434821 9707
rect 434821 9673 434855 9707
rect 434855 9673 434864 9707
rect 434812 9664 434864 9673
rect 276480 9596 276532 9648
rect 430580 9596 430632 9648
rect 436100 9596 436152 9648
rect 276480 9460 276532 9512
rect 230388 9052 230440 9104
rect 290740 9052 290792 9104
rect 291108 9052 291160 9104
rect 351368 9052 351420 9104
rect 257988 8984 258040 9036
rect 318064 8984 318116 9036
rect 351828 8984 351880 9036
rect 412088 8984 412140 9036
rect 489184 8984 489236 9036
rect 548892 8984 548944 9036
rect 108948 8916 109000 8968
rect 169392 8916 169444 8968
rect 172428 8916 172480 8968
rect 233700 8916 233752 8968
rect 310428 8916 310480 8968
rect 371608 8916 371660 8968
rect 433984 8916 434036 8968
rect 494152 8916 494204 8968
rect 3424 8236 3476 8288
rect 60096 8236 60148 8288
rect 284208 7760 284260 7812
rect 223488 7624 223540 7676
rect 283656 7624 283708 7676
rect 287060 7624 287112 7676
rect 288348 7624 288400 7676
rect 293868 7692 293920 7744
rect 353760 7692 353812 7744
rect 344284 7624 344336 7676
rect 423588 7624 423640 7676
rect 483480 7624 483532 7676
rect 104808 7556 104860 7608
rect 165896 7556 165948 7608
rect 169668 7556 169720 7608
rect 230112 7556 230164 7608
rect 234528 7556 234580 7608
rect 295524 7556 295576 7608
rect 344928 7556 344980 7608
rect 404912 7556 404964 7608
rect 433340 7556 433392 7608
rect 434628 7556 434680 7608
rect 452568 7556 452620 7608
rect 513196 7556 513248 7608
rect 520096 7556 520148 7608
rect 579804 7556 579856 7608
rect 244280 7488 244332 7540
rect 245568 7488 245620 7540
rect 262220 7488 262272 7540
rect 263416 7488 263468 7540
rect 270500 7488 270552 7540
rect 271696 7488 271748 7540
rect 167644 6264 167696 6316
rect 222936 6264 222988 6316
rect 301504 6264 301556 6316
rect 360936 6264 360988 6316
rect 110236 6196 110288 6248
rect 170588 6196 170640 6248
rect 219348 6196 219400 6248
rect 279976 6196 280028 6248
rect 280068 6196 280120 6248
rect 340696 6196 340748 6248
rect 100576 6128 100628 6180
rect 162308 6128 162360 6180
rect 180708 6128 180760 6180
rect 241980 6128 242032 6180
rect 252468 6128 252520 6180
rect 313372 6128 313424 6180
rect 340788 6128 340840 6180
rect 401324 6128 401376 6180
rect 430488 6128 430540 6180
rect 490564 6128 490616 6180
rect 502248 6128 502300 6180
rect 561956 6128 562008 6180
rect 374644 5516 374696 5568
rect 379980 5516 380032 5568
rect 362868 5244 362920 5296
rect 422760 5244 422812 5296
rect 463608 5244 463660 5296
rect 523868 5244 523920 5296
rect 380808 5176 380860 5228
rect 440608 5176 440660 5228
rect 462228 5176 462280 5228
rect 522672 5176 522724 5228
rect 248328 5040 248380 5092
rect 394608 5108 394660 5160
rect 454868 5108 454920 5160
rect 487068 5108 487120 5160
rect 547696 5108 547748 5160
rect 387708 5040 387760 5092
rect 447784 5040 447836 5092
rect 484308 5040 484360 5092
rect 544108 5040 544160 5092
rect 358728 4972 358780 5024
rect 308588 4904 308640 4956
rect 369768 4972 369820 5024
rect 429936 4972 429988 5024
rect 466368 4972 466420 5024
rect 526260 4972 526312 5024
rect 419172 4904 419224 4956
rect 68928 4836 68980 4888
rect 130200 4836 130252 4888
rect 133788 4836 133840 4888
rect 194416 4836 194468 4888
rect 209688 4836 209740 4888
rect 270592 4836 270644 4888
rect 308404 4836 308456 4888
rect 343088 4836 343140 4888
rect 455328 4904 455380 4956
rect 515588 4904 515640 4956
rect 459468 4836 459520 4888
rect 519084 4836 519136 4888
rect 66168 4768 66220 4820
rect 126612 4768 126664 4820
rect 126888 4768 126940 4820
rect 188436 4768 188488 4820
rect 190368 4768 190420 4820
rect 251456 4768 251508 4820
rect 270408 4768 270460 4820
rect 331312 4768 331364 4820
rect 333244 4768 333296 4820
rect 357256 4768 357308 4820
rect 372528 4768 372580 4820
rect 433524 4768 433576 4820
rect 476028 4768 476080 4820
rect 536932 4768 536984 4820
rect 390468 4700 390520 4752
rect 143448 4088 143500 4140
rect 203892 4088 203944 4140
rect 222108 4088 222160 4140
rect 282460 4088 282512 4140
rect 336648 4088 336700 4140
rect 396632 4088 396684 4140
rect 433248 4088 433300 4140
rect 492956 4088 493008 4140
rect 496728 4088 496780 4140
rect 557172 4088 557224 4140
rect 125508 4020 125560 4072
rect 186044 4020 186096 4072
rect 193128 4020 193180 4072
rect 253848 4020 253900 4072
rect 357348 4020 357400 4072
rect 417976 4020 418028 4072
rect 464988 4020 465040 4072
rect 525064 4020 525116 4072
rect 78588 3952 78640 4004
rect 139676 3952 139728 4004
rect 161388 3952 161440 4004
rect 221740 3952 221792 4004
rect 229008 3952 229060 4004
rect 289544 3952 289596 4004
rect 343548 3952 343600 4004
rect 403716 3952 403768 4004
rect 442908 3952 442960 4004
rect 503628 3952 503680 4004
rect 514668 3952 514720 4004
rect 575020 3952 575072 4004
rect 85488 3884 85540 3936
rect 146852 3884 146904 3936
rect 150532 3884 150584 3936
rect 151544 3884 151596 3936
rect 171048 3884 171100 3936
rect 232504 3884 232556 3936
rect 361488 3884 361540 3936
rect 421564 3884 421616 3936
rect 429108 3884 429160 3936
rect 489368 3884 489420 3936
rect 500868 3884 500920 3936
rect 560760 3884 560812 3936
rect 128268 3816 128320 3868
rect 189632 3816 189684 3868
rect 201500 3816 201552 3868
rect 202696 3816 202748 3868
rect 215208 3816 215260 3868
rect 275284 3816 275336 3868
rect 332508 3816 332560 3868
rect 393044 3816 393096 3868
rect 393228 3816 393280 3868
rect 453672 3816 453724 3868
rect 493968 3816 494020 3868
rect 553584 3816 553636 3868
rect 110328 3748 110380 3800
rect 171784 3748 171836 3800
rect 175188 3748 175240 3800
rect 236000 3748 236052 3800
rect 240048 3748 240100 3800
rect 300308 3748 300360 3800
rect 350448 3748 350500 3800
rect 410892 3748 410944 3800
rect 411168 3748 411220 3800
rect 471520 3748 471572 3800
rect 478788 3748 478840 3800
rect 539324 3748 539376 3800
rect 114468 3680 114520 3732
rect 175280 3680 175332 3732
rect 175372 3680 175424 3732
rect 176568 3680 176620 3732
rect 182088 3680 182140 3732
rect 243176 3680 243228 3732
rect 328368 3680 328420 3732
rect 389456 3680 389508 3732
rect 400128 3680 400180 3732
rect 460848 3680 460900 3732
rect 460940 3680 460992 3732
rect 521476 3680 521528 3732
rect 521568 3680 521620 3732
rect 582196 3680 582248 3732
rect 121368 3612 121420 3664
rect 182548 3612 182600 3664
rect 183560 3612 183612 3664
rect 184848 3612 184900 3664
rect 188988 3612 189040 3664
rect 250352 3612 250404 3664
rect 321468 3612 321520 3664
rect 382280 3612 382332 3664
rect 382372 3612 382424 3664
rect 383568 3612 383620 3664
rect 390560 3612 390612 3664
rect 391848 3612 391900 3664
rect 408500 3612 408552 3664
rect 409696 3612 409748 3664
rect 418068 3612 418120 3664
rect 478696 3612 478748 3664
rect 485780 3612 485832 3664
rect 486976 3612 487028 3664
rect 503444 3612 503496 3664
rect 564348 3612 564400 3664
rect 132408 3544 132460 3596
rect 193220 3544 193272 3596
rect 200028 3544 200080 3596
rect 261024 3544 261076 3596
rect 321652 3544 321704 3596
rect 322848 3544 322900 3596
rect 1676 3476 1728 3528
rect 63500 3476 63552 3528
rect 132592 3476 132644 3528
rect 133788 3476 133840 3528
rect 139308 3476 139360 3528
rect 200396 3476 200448 3528
rect 206928 3476 206980 3528
rect 268108 3476 268160 3528
rect 305000 3476 305052 3528
rect 306196 3476 306248 3528
rect 318708 3476 318760 3528
rect 378784 3544 378836 3596
rect 382188 3544 382240 3596
rect 443000 3544 443052 3596
rect 451280 3544 451332 3596
rect 452476 3544 452528 3596
rect 467840 3544 467892 3596
rect 469128 3544 469180 3596
rect 471888 3544 471940 3596
rect 528652 3544 528704 3596
rect 529848 3544 529900 3596
rect 536840 3544 536892 3596
rect 538128 3544 538180 3596
rect 331220 3476 331272 3528
rect 332416 3476 332468 3528
rect 347780 3476 347832 3528
rect 349068 3476 349120 3528
rect 572 3408 624 3460
rect 62120 3408 62172 3460
rect 71688 3408 71740 3460
rect 140780 3408 140832 3460
rect 142068 3408 142120 3460
rect 164148 3408 164200 3460
rect 225328 3408 225380 3460
rect 246948 3408 247000 3460
rect 307392 3408 307444 3460
rect 314568 3408 314620 3460
rect 132592 3340 132644 3392
rect 136456 3340 136508 3392
rect 196808 3340 196860 3392
rect 197268 3340 197320 3392
rect 257436 3340 257488 3392
rect 150348 3272 150400 3324
rect 211068 3272 211120 3324
rect 218060 3272 218112 3324
rect 219348 3272 219400 3324
rect 339408 3408 339460 3460
rect 346308 3340 346360 3392
rect 407304 3476 407356 3528
rect 415308 3476 415360 3528
rect 475108 3476 475160 3528
rect 494060 3476 494112 3528
rect 495348 3476 495400 3528
rect 507768 3476 507820 3528
rect 567844 3476 567896 3528
rect 571432 3476 571484 3528
rect 572628 3476 572680 3528
rect 574744 3476 574796 3528
rect 576216 3476 576268 3528
rect 400220 3408 400272 3460
rect 422208 3408 422260 3460
rect 482284 3408 482336 3460
rect 518808 3408 518860 3460
rect 578608 3408 578660 3460
rect 354588 3340 354640 3392
rect 414480 3340 414532 3392
rect 425060 3340 425112 3392
rect 426348 3340 426400 3392
rect 453948 3340 454000 3392
rect 514392 3340 514444 3392
rect 517428 3340 517480 3392
rect 577412 3340 577464 3392
rect 375196 3272 375248 3324
rect 386328 3272 386380 3324
rect 446588 3272 446640 3324
rect 458088 3272 458140 3324
rect 517888 3272 517940 3324
rect 532240 3272 532292 3324
rect 118608 3204 118660 3256
rect 178960 3204 179012 3256
rect 179328 3204 179380 3256
rect 239588 3204 239640 3256
rect 365720 3204 365772 3256
rect 366916 3204 366968 3256
rect 379428 3204 379480 3256
rect 439412 3204 439464 3256
rect 440148 3204 440200 3256
rect 500132 3204 500184 3256
rect 511908 3204 511960 3256
rect 571432 3204 571484 3256
rect 100668 3136 100720 3188
rect 161112 3136 161164 3188
rect 204168 3136 204220 3188
rect 264612 3136 264664 3188
rect 325608 3136 325660 3188
rect 385868 3136 385920 3188
rect 436008 3136 436060 3188
rect 496544 3136 496596 3188
rect 513288 3136 513340 3188
rect 573824 3136 573876 3188
rect 107568 3068 107620 3120
rect 168196 3068 168248 3120
rect 186228 3068 186280 3120
rect 246764 3068 246816 3120
rect 447048 3068 447100 3120
rect 507216 3068 507268 3120
rect 99288 3000 99340 3052
rect 159916 3000 159968 3052
rect 451280 2932 451332 2984
rect 427912 2796 427964 2848
rect 434812 2796 434864 2848
rect 428740 2728 428792 2780
rect 435824 2728 435876 2780
rect 301320 552 301372 604
rect 301412 552 301464 604
rect 354680 552 354732 604
rect 354956 552 355008 604
rect 357440 552 357492 604
rect 358544 552 358596 604
rect 358820 552 358872 604
rect 359740 552 359792 604
rect 361580 552 361632 604
rect 362132 552 362184 604
rect 431132 595 431184 604
rect 431132 561 431141 595
rect 431141 561 431175 595
rect 431175 561 431184 595
rect 431132 552 431184 561
rect 437020 595 437072 604
rect 437020 561 437029 595
rect 437029 561 437063 595
rect 437063 561 437072 595
rect 437020 552 437072 561
rect 461032 552 461084 604
rect 462044 552 462096 604
rect 462320 552 462372 604
rect 463240 552 463292 604
rect 463792 552 463844 604
rect 464436 552 464488 604
rect 465080 552 465132 604
rect 465632 552 465684 604
rect 466460 552 466512 604
rect 466828 552 466880 604
rect 469220 552 469272 604
rect 470324 552 470376 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3436 630630 3464 667927
rect 3528 645862 3556 682207
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654838 8064 663734
rect 24780 654906 24808 699654
rect 41340 654974 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 692782 72740 698278
rect 72700 692776 72752 692782
rect 72700 692718 72752 692724
rect 72516 683256 72568 683262
rect 72516 683198 72568 683204
rect 72528 683126 72556 683198
rect 72516 683120 72568 683126
rect 72516 683062 72568 683068
rect 72700 678904 72752 678910
rect 72700 678846 72752 678852
rect 72712 669322 72740 678846
rect 72700 669316 72752 669322
rect 72700 669258 72752 669264
rect 72884 669316 72936 669322
rect 72884 669258 72936 669264
rect 72896 666534 72924 669258
rect 72884 666528 72936 666534
rect 72884 666470 72936 666476
rect 72792 656940 72844 656946
rect 72792 656882 72844 656888
rect 41328 654968 41380 654974
rect 41328 654910 41380 654916
rect 24768 654900 24820 654906
rect 24768 654842 24820 654848
rect 72804 654838 72832 656882
rect 89640 654906 89668 699654
rect 106200 654974 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 104532 654968 104584 654974
rect 104532 654910 104584 654916
rect 106188 654968 106240 654974
rect 106188 654910 106240 654916
rect 87512 654900 87564 654906
rect 87512 654842 87564 654848
rect 89628 654900 89680 654906
rect 89628 654842 89680 654848
rect 8024 654832 8076 654838
rect 8024 654774 8076 654780
rect 70492 654832 70544 654838
rect 70492 654774 70544 654780
rect 72792 654832 72844 654838
rect 72792 654774 72844 654780
rect 3606 653576 3662 653585
rect 3606 653511 3662 653520
rect 3516 645856 3568 645862
rect 3516 645798 3568 645804
rect 3424 630624 3476 630630
rect 3424 630566 3476 630572
rect 3514 624880 3570 624889
rect 3514 624815 3570 624824
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 587858 3464 610399
rect 3528 603090 3556 624815
rect 3620 616826 3648 653511
rect 70504 651916 70532 654774
rect 87524 651916 87552 654842
rect 104544 651916 104572 654910
rect 137756 654838 137784 663734
rect 154316 655042 154344 663734
rect 154304 655036 154356 655042
rect 154304 654978 154356 654984
rect 155592 654968 155644 654974
rect 155592 654910 155644 654916
rect 138572 654900 138624 654906
rect 138572 654842 138624 654848
rect 121552 654832 121604 654838
rect 121552 654774 121604 654780
rect 137744 654832 137796 654838
rect 137744 654774 137796 654780
rect 121564 651916 121592 654774
rect 138584 651916 138612 654842
rect 155604 651916 155632 654910
rect 171060 654906 171088 700198
rect 189724 655036 189776 655042
rect 189724 654978 189776 654984
rect 171048 654900 171100 654906
rect 171048 654842 171100 654848
rect 172704 654832 172756 654838
rect 172704 654774 172756 654780
rect 172716 651916 172744 654774
rect 189736 651916 189764 654978
rect 202800 654838 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 679046 219112 685850
rect 219072 679040 219124 679046
rect 219072 678982 219124 678988
rect 218980 678972 219032 678978
rect 218980 678914 219032 678920
rect 218992 669322 219020 678914
rect 218980 669316 219032 669322
rect 218980 669258 219032 669264
rect 219164 669316 219216 669322
rect 219164 669258 219216 669264
rect 219176 666534 219204 669258
rect 219164 666528 219216 666534
rect 219164 666470 219216 666476
rect 219072 656940 219124 656946
rect 219072 656882 219124 656888
rect 219084 654906 219112 656882
rect 206744 654900 206796 654906
rect 206744 654842 206796 654848
rect 219072 654900 219124 654906
rect 219072 654842 219124 654848
rect 202788 654832 202840 654838
rect 202788 654774 202840 654780
rect 206756 651916 206784 654842
rect 235920 654838 235948 699654
rect 240784 654900 240836 654906
rect 240784 654842 240836 654848
rect 223764 654832 223816 654838
rect 223764 654774 223816 654780
rect 235908 654832 235960 654838
rect 235908 654774 235960 654780
rect 223776 651916 223804 654774
rect 240796 651916 240824 654842
rect 267660 654838 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 343548 700324 343600 700330
rect 343548 700266 343600 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 326988 699712 327040 699718
rect 326988 699654 327040 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654838 284064 663734
rect 257896 654832 257948 654838
rect 257896 654774 257948 654780
rect 267648 654832 267700 654838
rect 267648 654774 267700 654780
rect 274916 654832 274968 654838
rect 274916 654774 274968 654780
rect 284024 654832 284076 654838
rect 284024 654774 284076 654780
rect 291936 654832 291988 654838
rect 291936 654774 291988 654780
rect 257908 651916 257936 654774
rect 274928 651916 274956 654774
rect 291948 651916 291976 654774
rect 300780 654158 300808 699654
rect 327000 655178 327028 699654
rect 325976 655172 326028 655178
rect 325976 655114 326028 655120
rect 326988 655172 327040 655178
rect 326988 655114 327040 655120
rect 300768 654152 300820 654158
rect 300768 654094 300820 654100
rect 308956 654152 309008 654158
rect 308956 654094 309008 654100
rect 308968 651916 308996 654094
rect 325988 651916 326016 655114
rect 343560 651794 343588 700266
rect 364996 699718 365024 703520
rect 394608 700392 394660 700398
rect 394608 700334 394660 700340
rect 378048 700324 378100 700330
rect 378048 700266 378100 700272
rect 360108 699712 360160 699718
rect 360108 699654 360160 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 360120 651916 360148 699654
rect 378060 655518 378088 700266
rect 377128 655512 377180 655518
rect 377128 655454 377180 655460
rect 378048 655512 378100 655518
rect 378048 655454 378100 655460
rect 377140 651916 377168 655454
rect 394620 651794 394648 700334
rect 397472 700330 397500 703520
rect 411168 700460 411220 700466
rect 411168 700402 411220 700408
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 411180 651916 411208 700402
rect 413664 700398 413692 703520
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 445668 700392 445720 700398
rect 445668 700334 445720 700340
rect 429108 700324 429160 700330
rect 429108 700266 429160 700272
rect 429120 655518 429148 700266
rect 428188 655512 428240 655518
rect 428188 655454 428240 655460
rect 429108 655512 429160 655518
rect 429108 655454 429160 655460
rect 428200 651916 428228 655454
rect 445680 651930 445708 700334
rect 462332 700330 462360 703520
rect 463608 700460 463660 700466
rect 463608 700402 463660 700408
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 463620 655518 463648 700402
rect 478524 700398 478552 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 514668 700460 514720 700466
rect 514668 700402 514720 700408
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 496728 700392 496780 700398
rect 496728 700334 496780 700340
rect 480168 700324 480220 700330
rect 480168 700266 480220 700272
rect 480180 655518 480208 700266
rect 462320 655512 462372 655518
rect 462320 655454 462372 655460
rect 463608 655512 463660 655518
rect 463608 655454 463660 655460
rect 479340 655512 479392 655518
rect 479340 655454 479392 655460
rect 480168 655512 480220 655518
rect 480168 655454 480220 655460
rect 445326 651902 445708 651930
rect 462332 651916 462360 655454
rect 479352 651916 479380 655454
rect 496740 651930 496768 700334
rect 514680 655314 514708 700402
rect 527192 700330 527220 703520
rect 543476 700398 543504 703520
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 523776 696992 523828 696998
rect 523776 696934 523828 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 523684 685908 523736 685914
rect 523684 685850 523736 685856
rect 513380 655308 513432 655314
rect 513380 655250 513432 655256
rect 514668 655308 514720 655314
rect 514668 655250 514720 655256
rect 496386 651902 496768 651930
rect 513392 651916 513420 655250
rect 343022 651766 343588 651794
rect 394174 651766 394648 651794
rect 59360 645856 59412 645862
rect 59360 645798 59412 645804
rect 59372 644745 59400 645798
rect 59358 644736 59414 644745
rect 59358 644671 59414 644680
rect 523696 631961 523724 685850
rect 523788 645289 523816 696934
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 523774 645280 523830 645289
rect 523774 645215 523830 645224
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 523776 638988 523828 638994
rect 523776 638930 523828 638936
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 523682 631952 523738 631961
rect 523682 631887 523738 631896
rect 59360 630624 59412 630630
rect 59360 630566 59412 630572
rect 59372 630465 59400 630566
rect 59358 630456 59414 630465
rect 59358 630391 59414 630400
rect 3608 616820 3660 616826
rect 3608 616762 3660 616768
rect 59360 616820 59412 616826
rect 59360 616762 59412 616768
rect 59372 616185 59400 616762
rect 59358 616176 59414 616185
rect 59358 616111 59414 616120
rect 523132 605804 523184 605810
rect 523132 605746 523184 605752
rect 523144 605305 523172 605746
rect 523130 605296 523186 605305
rect 523130 605231 523186 605240
rect 3516 603084 3568 603090
rect 3516 603026 3568 603032
rect 59360 603084 59412 603090
rect 59360 603026 59412 603032
rect 59372 601905 59400 603026
rect 59358 601896 59414 601905
rect 59358 601831 59414 601840
rect 3514 596048 3570 596057
rect 3514 595983 3570 595992
rect 3424 587852 3476 587858
rect 3424 587794 3476 587800
rect 3528 574054 3556 595983
rect 523684 592068 523736 592074
rect 523684 592010 523736 592016
rect 59360 587852 59412 587858
rect 59360 587794 59412 587800
rect 59372 587625 59400 587794
rect 59358 587616 59414 587625
rect 59358 587551 59414 587560
rect 3516 574048 3568 574054
rect 3516 573990 3568 573996
rect 59360 574048 59412 574054
rect 59360 573990 59412 573996
rect 59372 573345 59400 573990
rect 59358 573336 59414 573345
rect 59358 573271 59414 573280
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 560250 3464 567287
rect 523132 565820 523184 565826
rect 523132 565762 523184 565768
rect 523144 565321 523172 565762
rect 523130 565312 523186 565321
rect 523130 565247 523186 565256
rect 3424 560244 3476 560250
rect 3424 560186 3476 560192
rect 59360 560244 59412 560250
rect 59360 560186 59412 560192
rect 59372 559065 59400 560186
rect 59358 559056 59414 559065
rect 59358 558991 59414 559000
rect 3422 553072 3478 553081
rect 3422 553007 3478 553016
rect 3436 545086 3464 553007
rect 523696 551993 523724 592010
rect 523788 591977 523816 638930
rect 580276 619614 580304 674591
rect 580446 651128 580502 651137
rect 580446 651063 580502 651072
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 524328 619608 524380 619614
rect 524328 619550 524380 619556
rect 580264 619608 580316 619614
rect 580264 619550 580316 619556
rect 524340 618633 524368 619550
rect 524326 618624 524382 618633
rect 524326 618559 524382 618568
rect 579802 592512 579858 592521
rect 579802 592447 579858 592456
rect 579816 592074 579844 592447
rect 579804 592068 579856 592074
rect 579804 592010 579856 592016
rect 523774 591968 523830 591977
rect 523774 591903 523830 591912
rect 580262 580816 580318 580825
rect 580262 580751 580318 580760
rect 524328 579624 524380 579630
rect 524328 579566 524380 579572
rect 524340 578649 524368 579566
rect 524326 578640 524382 578649
rect 524326 578575 524382 578584
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 523776 556232 523828 556238
rect 523776 556174 523828 556180
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 523682 551984 523738 551993
rect 523682 551919 523738 551928
rect 523500 545148 523552 545154
rect 523500 545090 523552 545096
rect 3424 545080 3476 545086
rect 3424 545022 3476 545028
rect 59360 545080 59412 545086
rect 59360 545022 59412 545028
rect 59372 544785 59400 545022
rect 59358 544776 59414 544785
rect 59358 544711 59414 544720
rect 3422 538656 3478 538665
rect 3422 538591 3478 538600
rect 3436 531282 3464 538591
rect 523512 538234 523540 545090
rect 523684 539572 523736 539578
rect 523684 539514 523736 539520
rect 523696 538665 523724 539514
rect 523682 538656 523738 538665
rect 523682 538591 523738 538600
rect 523512 538206 523724 538234
rect 3424 531276 3476 531282
rect 3424 531218 3476 531224
rect 59360 531276 59412 531282
rect 59360 531218 59412 531224
rect 59372 530505 59400 531218
rect 59358 530496 59414 530505
rect 59358 530431 59414 530440
rect 59358 516216 59414 516225
rect 59358 516151 59414 516160
rect 59372 510610 59400 516151
rect 523696 512009 523724 538206
rect 523788 525337 523816 556174
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580276 539578 580304 580751
rect 580368 579630 580396 627671
rect 580460 605810 580488 651063
rect 580448 605804 580500 605810
rect 580448 605746 580500 605752
rect 580446 604208 580502 604217
rect 580446 604143 580502 604152
rect 580356 579624 580408 579630
rect 580356 579566 580408 579572
rect 580460 565826 580488 604143
rect 580448 565820 580500 565826
rect 580448 565762 580500 565768
rect 580264 539572 580316 539578
rect 580264 539514 580316 539520
rect 580262 533896 580318 533905
rect 580262 533831 580318 533840
rect 523774 525328 523830 525337
rect 523774 525263 523830 525272
rect 523682 512000 523738 512009
rect 523682 511935 523738 511944
rect 3148 510604 3200 510610
rect 3148 510546 3200 510552
rect 59360 510604 59412 510610
rect 59360 510546 59412 510552
rect 3160 509969 3188 510546
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 3146 509960 3202 509969
rect 3146 509895 3202 509904
rect 580184 509318 580212 510303
rect 523776 509312 523828 509318
rect 523776 509254 523828 509260
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 60002 501936 60058 501945
rect 60002 501871 60058 501880
rect 60016 496806 60044 501871
rect 523684 499520 523736 499526
rect 523684 499462 523736 499468
rect 523696 498681 523724 499462
rect 523682 498672 523738 498681
rect 523682 498607 523738 498616
rect 523684 498228 523736 498234
rect 523684 498170 523736 498176
rect 3424 496800 3476 496806
rect 3424 496742 3476 496748
rect 60004 496800 60056 496806
rect 60004 496742 60056 496748
rect 3436 495553 3464 496742
rect 3422 495544 3478 495553
rect 3422 495479 3478 495488
rect 59358 487656 59414 487665
rect 59358 487591 59414 487600
rect 59372 481642 59400 487591
rect 3516 481636 3568 481642
rect 3516 481578 3568 481584
rect 59360 481636 59412 481642
rect 59360 481578 59412 481584
rect 3528 481137 3556 481578
rect 3514 481128 3570 481137
rect 3514 481063 3570 481072
rect 60002 473376 60058 473385
rect 60002 473311 60058 473320
rect 60016 452606 60044 473311
rect 523696 472025 523724 498170
rect 523788 485353 523816 509254
rect 580276 499526 580304 533831
rect 580264 499520 580316 499526
rect 580264 499462 580316 499468
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580262 486840 580318 486849
rect 580262 486775 580318 486784
rect 523774 485344 523830 485353
rect 523774 485279 523830 485288
rect 523682 472016 523738 472025
rect 523682 471951 523738 471960
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 523684 462392 523736 462398
rect 523684 462334 523736 462340
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 60094 459096 60150 459105
rect 60094 459031 60150 459040
rect 3424 452600 3476 452606
rect 3424 452542 3476 452548
rect 60004 452600 60056 452606
rect 60004 452542 60056 452548
rect 3436 452441 3464 452542
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 60002 444816 60058 444825
rect 60002 444751 60058 444760
rect 3148 438864 3200 438870
rect 3148 438806 3200 438812
rect 3160 438025 3188 438806
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 60016 425066 60044 444751
rect 60108 438870 60136 459031
rect 523696 445369 523724 462334
rect 580276 459542 580304 486775
rect 524328 459536 524380 459542
rect 524328 459478 524380 459484
rect 580264 459536 580316 459542
rect 580264 459478 580316 459484
rect 524340 458697 524368 459478
rect 524326 458688 524382 458697
rect 524326 458623 524382 458632
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 523776 451308 523828 451314
rect 523776 451250 523828 451256
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 523682 445360 523738 445369
rect 523682 445295 523738 445304
rect 523684 438932 523736 438938
rect 523684 438874 523736 438880
rect 60096 438864 60148 438870
rect 60096 438806 60148 438812
rect 60094 430536 60150 430545
rect 60094 430471 60150 430480
rect 3240 425060 3292 425066
rect 3240 425002 3292 425008
rect 60004 425060 60056 425066
rect 60004 425002 60056 425008
rect 3252 423745 3280 425002
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 60002 401976 60058 401985
rect 60002 401911 60058 401920
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 60016 367062 60044 401911
rect 60108 396030 60136 430471
rect 523696 418713 523724 438874
rect 523788 432041 523816 451250
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 523774 432032 523830 432041
rect 523774 431967 523830 431976
rect 523682 418704 523738 418713
rect 523682 418639 523738 418648
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 60186 416256 60242 416265
rect 60186 416191 60242 416200
rect 60096 396024 60148 396030
rect 60096 395966 60148 395972
rect 60094 387696 60150 387705
rect 60094 387631 60150 387640
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 60004 367056 60056 367062
rect 60004 366998 60056 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 60002 359136 60058 359145
rect 60002 359071 60058 359080
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 60016 309126 60044 359071
rect 60108 338094 60136 387631
rect 60200 380866 60228 416191
rect 580184 415478 580212 416463
rect 523684 415472 523736 415478
rect 523684 415414 523736 415420
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 523696 405385 523724 415414
rect 523682 405376 523738 405385
rect 523682 405311 523738 405320
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 523776 404388 523828 404394
rect 523776 404330 523828 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 523788 392057 523816 404330
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 523774 392048 523830 392057
rect 523684 392012 523736 392018
rect 580184 392018 580212 392935
rect 523774 391983 523830 391992
rect 580172 392012 580224 392018
rect 523684 391954 523736 391960
rect 580172 391954 580224 391960
rect 60188 380860 60240 380866
rect 60188 380802 60240 380808
rect 523696 378729 523724 391954
rect 523682 378720 523738 378729
rect 523682 378655 523738 378664
rect 60186 373416 60242 373425
rect 60186 373351 60242 373360
rect 60096 338088 60148 338094
rect 60096 338030 60148 338036
rect 60094 330440 60150 330449
rect 60094 330375 60150 330384
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 60004 309120 60056 309126
rect 60004 309062 60056 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3424 295316 3476 295322
rect 3424 295258 3476 295264
rect 3436 294409 3464 295258
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 60002 287600 60058 287609
rect 60002 287535 60058 287544
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 3148 266348 3200 266354
rect 3148 266290 3200 266296
rect 3160 265713 3188 266290
rect 3146 265704 3202 265713
rect 3146 265639 3202 265648
rect 3424 252544 3476 252550
rect 3424 252486 3476 252492
rect 3436 251297 3464 252486
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 60016 237386 60044 287535
rect 60108 280158 60136 330375
rect 60200 324290 60228 373351
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 524236 368552 524288 368558
rect 524236 368494 524288 368500
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 524248 365401 524276 368494
rect 524234 365392 524290 365401
rect 524234 365327 524290 365336
rect 580170 357912 580226 357921
rect 580170 357847 580226 357856
rect 580184 357474 580212 357847
rect 523684 357468 523736 357474
rect 523684 357410 523736 357416
rect 580172 357468 580224 357474
rect 580172 357410 580224 357416
rect 523696 351937 523724 357410
rect 523682 351928 523738 351937
rect 523682 351863 523738 351872
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345098 580212 346015
rect 523776 345092 523828 345098
rect 523776 345034 523828 345040
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 60370 344720 60426 344729
rect 60370 344655 60426 344664
rect 60188 324284 60240 324290
rect 60188 324226 60240 324232
rect 60278 316160 60334 316169
rect 60278 316095 60334 316104
rect 60096 280152 60148 280158
rect 60096 280094 60148 280100
rect 60186 273320 60242 273329
rect 60186 273255 60242 273264
rect 60094 259040 60150 259049
rect 60094 258975 60150 258984
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 60004 237380 60056 237386
rect 60004 237322 60056 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 60108 208350 60136 258975
rect 60200 223582 60228 273255
rect 60292 266354 60320 316095
rect 60384 295322 60412 344655
rect 523788 338609 523816 345034
rect 523774 338600 523830 338609
rect 523774 338535 523830 338544
rect 524326 325272 524382 325281
rect 524326 325207 524382 325216
rect 524340 322930 524368 325207
rect 524328 322924 524380 322930
rect 524328 322866 524380 322872
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 524326 311944 524382 311953
rect 524326 311879 524382 311888
rect 524340 311846 524368 311879
rect 524328 311840 524380 311846
rect 524328 311782 524380 311788
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 60462 301880 60518 301889
rect 60462 301815 60518 301824
rect 60372 295316 60424 295322
rect 60372 295258 60424 295264
rect 60280 266348 60332 266354
rect 60280 266290 60332 266296
rect 60476 252550 60504 301815
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580184 298790 580212 299095
rect 524328 298784 524380 298790
rect 524328 298726 524380 298732
rect 580172 298784 580224 298790
rect 580172 298726 580224 298732
rect 524340 298625 524368 298726
rect 524326 298616 524382 298625
rect 524326 298551 524382 298560
rect 523682 285288 523738 285297
rect 523682 285223 523738 285232
rect 523696 276010 523724 285223
rect 523684 276004 523736 276010
rect 523684 275946 523736 275952
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 523682 271960 523738 271969
rect 523682 271895 523738 271904
rect 523696 264926 523724 271895
rect 523684 264920 523736 264926
rect 523684 264862 523736 264868
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 523682 258632 523738 258641
rect 523682 258567 523738 258576
rect 523696 252550 523724 258567
rect 60464 252544 60516 252550
rect 60464 252486 60516 252492
rect 523684 252544 523736 252550
rect 523684 252486 523736 252492
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 523682 245304 523738 245313
rect 523682 245239 523738 245248
rect 60278 244760 60334 244769
rect 60278 244695 60334 244704
rect 60188 223576 60240 223582
rect 60188 223518 60240 223524
rect 60186 216200 60242 216209
rect 60186 216135 60242 216144
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 60096 208344 60148 208350
rect 60096 208286 60148 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 60094 201920 60150 201929
rect 60094 201855 60150 201864
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 60002 187640 60058 187649
rect 60002 187575 60058 187584
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 60016 136610 60044 187575
rect 60108 151774 60136 201855
rect 60200 165578 60228 216135
rect 60292 194546 60320 244695
rect 60370 230480 60426 230489
rect 60370 230415 60426 230424
rect 60280 194540 60332 194546
rect 60280 194482 60332 194488
rect 60384 180810 60412 230415
rect 523696 229090 523724 245239
rect 523774 231976 523830 231985
rect 523774 231911 523830 231920
rect 523684 229084 523736 229090
rect 523684 229026 523736 229032
rect 523788 218006 523816 231911
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 523866 218648 523922 218657
rect 523866 218583 523922 218592
rect 523776 218000 523828 218006
rect 523776 217942 523828 217948
rect 523880 205630 523908 218583
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 523868 205624 523920 205630
rect 523868 205566 523920 205572
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 523682 205320 523738 205329
rect 523682 205255 523738 205264
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 523696 182170 523724 205255
rect 523774 191992 523830 192001
rect 523774 191927 523830 191936
rect 523684 182164 523736 182170
rect 523684 182106 523736 182112
rect 60372 180804 60424 180810
rect 60372 180746 60424 180752
rect 60370 173360 60426 173369
rect 60370 173295 60426 173304
rect 60188 165572 60240 165578
rect 60188 165514 60240 165520
rect 60278 159080 60334 159089
rect 60278 159015 60334 159024
rect 60096 151768 60148 151774
rect 60096 151710 60148 151716
rect 60186 144800 60242 144809
rect 60186 144735 60242 144744
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 60004 136604 60056 136610
rect 60004 136546 60056 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 60002 130520 60058 130529
rect 60002 130455 60058 130464
rect 3424 122800 3476 122806
rect 3424 122742 3476 122748
rect 3436 122097 3464 122742
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 60016 80034 60044 130455
rect 60094 116240 60150 116249
rect 60094 116175 60150 116184
rect 3424 80028 3476 80034
rect 3424 79970 3476 79976
rect 60004 80028 60056 80034
rect 60004 79970 60056 79976
rect 3436 78985 3464 79970
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 60002 73400 60058 73409
rect 60002 73335 60058 73344
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 60016 22098 60044 73335
rect 60108 64870 60136 116175
rect 60200 93838 60228 144735
rect 60292 109002 60320 159015
rect 60384 122806 60412 173295
rect 523788 171086 523816 191927
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 523866 178664 523922 178673
rect 523866 178599 523922 178608
rect 523776 171080 523828 171086
rect 523776 171022 523828 171028
rect 523682 165336 523738 165345
rect 523682 165271 523738 165280
rect 523696 135250 523724 165271
rect 523880 158710 523908 178599
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 523868 158704 523920 158710
rect 523868 158646 523920 158652
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 523774 152008 523830 152017
rect 523774 151943 523830 151952
rect 523684 135244 523736 135250
rect 523684 135186 523736 135192
rect 523682 125352 523738 125361
rect 523682 125287 523738 125296
rect 60372 122800 60424 122806
rect 60372 122742 60424 122748
rect 60280 108996 60332 109002
rect 60280 108938 60332 108944
rect 60278 101960 60334 101969
rect 60278 101895 60334 101904
rect 60188 93832 60240 93838
rect 60188 93774 60240 93780
rect 60186 87680 60242 87689
rect 60186 87615 60242 87624
rect 60096 64864 60148 64870
rect 60096 64806 60148 64812
rect 60094 59120 60150 59129
rect 60094 59055 60150 59064
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 60004 22092 60056 22098
rect 60004 22034 60056 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 60108 8294 60136 59055
rect 60200 35902 60228 87615
rect 60292 51066 60320 101895
rect 523696 88330 523724 125287
rect 523788 124166 523816 151943
rect 523866 138680 523922 138689
rect 523866 138615 523922 138624
rect 523776 124160 523828 124166
rect 523776 124102 523828 124108
rect 523774 112024 523830 112033
rect 523774 111959 523830 111968
rect 523684 88324 523736 88330
rect 523684 88266 523736 88272
rect 523682 85368 523738 85377
rect 523682 85303 523738 85312
rect 62132 52006 62606 52034
rect 63512 52006 63710 52034
rect 60280 51060 60332 51066
rect 60280 51002 60332 51008
rect 60188 35896 60240 35902
rect 60188 35838 60240 35844
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 60096 8288 60148 8294
rect 60096 8230 60148 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 62132 3466 62160 52006
rect 63512 3534 63540 52006
rect 64892 48754 64920 52020
rect 66088 48822 66116 52020
rect 67284 49026 67312 52020
rect 68494 52006 68968 52034
rect 69690 52006 70348 52034
rect 67272 49020 67324 49026
rect 67272 48962 67324 48968
rect 66076 48816 66128 48822
rect 66076 48758 66128 48764
rect 66904 48816 66956 48822
rect 66904 48758 66956 48764
rect 64880 48748 64932 48754
rect 64880 48690 64932 48696
rect 66168 48748 66220 48754
rect 66168 48690 66220 48696
rect 66180 4826 66208 48690
rect 66916 15910 66944 48758
rect 66904 15904 66956 15910
rect 66904 15846 66956 15852
rect 68940 4894 68968 52006
rect 70320 17270 70348 52006
rect 70872 48822 70900 52020
rect 72068 48822 72096 52020
rect 73264 48822 73292 52020
rect 74460 49298 74488 52020
rect 75670 52006 75868 52034
rect 74448 49292 74500 49298
rect 74448 49234 74500 49240
rect 70860 48816 70912 48822
rect 70860 48758 70912 48764
rect 71688 48816 71740 48822
rect 71688 48758 71740 48764
rect 72056 48816 72108 48822
rect 72056 48758 72108 48764
rect 73068 48816 73120 48822
rect 73068 48758 73120 48764
rect 73252 48816 73304 48822
rect 73252 48758 73304 48764
rect 74448 48816 74500 48822
rect 74448 48758 74500 48764
rect 70308 17264 70360 17270
rect 70308 17206 70360 17212
rect 68928 4888 68980 4894
rect 68928 4830 68980 4836
rect 66168 4820 66220 4826
rect 66168 4762 66220 4768
rect 63500 3528 63552 3534
rect 63500 3470 63552 3476
rect 71700 3466 71728 48758
rect 73080 18630 73108 48758
rect 73068 18624 73120 18630
rect 73068 18566 73120 18572
rect 74460 14550 74488 48758
rect 75840 19990 75868 52006
rect 76852 48822 76880 52020
rect 78062 52006 78628 52034
rect 79258 52006 80008 52034
rect 76840 48816 76892 48822
rect 76840 48758 76892 48764
rect 77944 48816 77996 48822
rect 77944 48758 77996 48764
rect 77956 37942 77984 48758
rect 77944 37936 77996 37942
rect 77944 37878 77996 37884
rect 75828 19984 75880 19990
rect 75828 19926 75880 19932
rect 74448 14544 74500 14550
rect 74448 14486 74500 14492
rect 78600 4010 78628 52006
rect 79980 21418 80008 52006
rect 80440 48822 80468 52020
rect 81636 49366 81664 52020
rect 82832 49706 82860 52020
rect 84042 52006 84148 52034
rect 85238 52006 85528 52034
rect 86434 52006 86908 52034
rect 87630 52006 88288 52034
rect 82820 49700 82872 49706
rect 82820 49642 82872 49648
rect 81624 49360 81676 49366
rect 81624 49302 81676 49308
rect 80428 48816 80480 48822
rect 80428 48758 80480 48764
rect 82084 48816 82136 48822
rect 82084 48758 82136 48764
rect 82096 39370 82124 48758
rect 84120 42090 84148 52006
rect 84844 49700 84896 49706
rect 84844 49642 84896 49648
rect 84108 42084 84160 42090
rect 84108 42026 84160 42032
rect 82084 39364 82136 39370
rect 82084 39306 82136 39312
rect 84856 22778 84884 49642
rect 84844 22772 84896 22778
rect 84844 22714 84896 22720
rect 79968 21412 80020 21418
rect 79968 21354 80020 21360
rect 78588 4004 78640 4010
rect 78588 3946 78640 3952
rect 85500 3942 85528 52006
rect 86880 24138 86908 52006
rect 88260 40730 88288 52006
rect 88720 49230 88748 52020
rect 88708 49224 88760 49230
rect 88708 49166 88760 49172
rect 89916 48822 89944 52020
rect 91112 48822 91140 52020
rect 92322 52006 92428 52034
rect 93518 52006 93808 52034
rect 89904 48816 89956 48822
rect 89904 48758 89956 48764
rect 91008 48816 91060 48822
rect 91008 48758 91060 48764
rect 91100 48816 91152 48822
rect 91100 48758 91152 48764
rect 92296 48816 92348 48822
rect 92296 48758 92348 48764
rect 88248 40724 88300 40730
rect 88248 40666 88300 40672
rect 91020 25566 91048 48758
rect 91008 25560 91060 25566
rect 91008 25502 91060 25508
rect 86868 24132 86920 24138
rect 86868 24074 86920 24080
rect 92308 13190 92336 48758
rect 92296 13184 92348 13190
rect 92296 13126 92348 13132
rect 85488 3936 85540 3942
rect 85488 3878 85540 3884
rect 62120 3460 62172 3466
rect 62120 3402 62172 3408
rect 71688 3460 71740 3466
rect 71688 3402 71740 3408
rect 92400 3369 92428 52006
rect 93780 26926 93808 52006
rect 94700 47598 94728 52020
rect 95896 49162 95924 52020
rect 95884 49156 95936 49162
rect 95884 49098 95936 49104
rect 97092 48822 97120 52020
rect 98288 48822 98316 52020
rect 99484 48822 99512 52020
rect 100588 52006 100694 52034
rect 101890 52006 102088 52034
rect 97080 48816 97132 48822
rect 97080 48758 97132 48764
rect 97908 48816 97960 48822
rect 97908 48758 97960 48764
rect 98276 48816 98328 48822
rect 98276 48758 98328 48764
rect 99288 48816 99340 48822
rect 99288 48758 99340 48764
rect 99472 48816 99524 48822
rect 99472 48758 99524 48764
rect 94688 47592 94740 47598
rect 94688 47534 94740 47540
rect 97920 28354 97948 48758
rect 97908 28348 97960 28354
rect 97908 28290 97960 28296
rect 93768 26920 93820 26926
rect 93768 26862 93820 26868
rect 92386 3360 92442 3369
rect 92386 3295 92442 3304
rect 99300 3058 99328 48758
rect 100588 6186 100616 52006
rect 100668 48816 100720 48822
rect 100668 48758 100720 48764
rect 100576 6180 100628 6186
rect 100576 6122 100628 6128
rect 100680 3194 100708 48758
rect 102060 29646 102088 52006
rect 103072 49094 103100 52020
rect 104282 52006 104848 52034
rect 103060 49088 103112 49094
rect 103060 49030 103112 49036
rect 102048 29640 102100 29646
rect 102048 29582 102100 29588
rect 104820 7614 104848 52006
rect 105464 48822 105492 52020
rect 106660 48822 106688 52020
rect 107856 48822 107884 52020
rect 109052 48822 109080 52020
rect 110262 52006 110368 52034
rect 111458 52006 111748 52034
rect 105452 48816 105504 48822
rect 105452 48758 105504 48764
rect 106188 48816 106240 48822
rect 106188 48758 106240 48764
rect 106648 48816 106700 48822
rect 106648 48758 106700 48764
rect 107568 48816 107620 48822
rect 107568 48758 107620 48764
rect 107844 48816 107896 48822
rect 107844 48758 107896 48764
rect 108948 48816 109000 48822
rect 108948 48758 109000 48764
rect 109040 48816 109092 48822
rect 109040 48758 109092 48764
rect 110236 48816 110288 48822
rect 110236 48758 110288 48764
rect 106200 31074 106228 48758
rect 106188 31068 106240 31074
rect 106188 31010 106240 31016
rect 104808 7608 104860 7614
rect 104808 7550 104860 7556
rect 100668 3188 100720 3194
rect 100668 3130 100720 3136
rect 107580 3126 107608 48758
rect 108960 8974 108988 48758
rect 108948 8968 109000 8974
rect 108948 8910 109000 8916
rect 110248 6254 110276 48758
rect 110236 6248 110288 6254
rect 110236 6190 110288 6196
rect 110340 3806 110368 52006
rect 111720 10334 111748 52006
rect 112640 46238 112668 52020
rect 113744 48822 113772 52020
rect 114940 48822 114968 52020
rect 116136 48822 116164 52020
rect 117332 48822 117360 52020
rect 113732 48816 113784 48822
rect 113732 48758 113784 48764
rect 114468 48816 114520 48822
rect 114468 48758 114520 48764
rect 114928 48816 114980 48822
rect 114928 48758 114980 48764
rect 115848 48816 115900 48822
rect 115848 48758 115900 48764
rect 116124 48816 116176 48822
rect 116124 48758 116176 48764
rect 117228 48816 117280 48822
rect 117228 48758 117280 48764
rect 117320 48816 117372 48822
rect 117320 48758 117372 48764
rect 112628 46232 112680 46238
rect 112628 46174 112680 46180
rect 111708 10328 111760 10334
rect 111708 10270 111760 10276
rect 110328 3800 110380 3806
rect 110328 3742 110380 3748
rect 114480 3738 114508 48758
rect 115860 11762 115888 48758
rect 117240 44878 117268 48758
rect 117228 44872 117280 44878
rect 117228 44814 117280 44820
rect 118528 13122 118556 52020
rect 119738 52006 120028 52034
rect 120934 52006 121408 52034
rect 122130 52006 122788 52034
rect 118608 48816 118660 48822
rect 118608 48758 118660 48764
rect 118516 13116 118568 13122
rect 118516 13058 118568 13064
rect 115848 11756 115900 11762
rect 115848 11698 115900 11704
rect 114468 3732 114520 3738
rect 114468 3674 114520 3680
rect 118620 3262 118648 48758
rect 120000 32434 120028 52006
rect 119988 32428 120040 32434
rect 119988 32370 120040 32376
rect 121380 3670 121408 52006
rect 122760 14482 122788 52006
rect 123312 48754 123340 52020
rect 124508 48822 124536 52020
rect 124496 48816 124548 48822
rect 124496 48758 124548 48764
rect 125508 48816 125560 48822
rect 125508 48758 125560 48764
rect 123300 48748 123352 48754
rect 123300 48690 123352 48696
rect 124128 48748 124180 48754
rect 124128 48690 124180 48696
rect 124140 33862 124168 48690
rect 124128 33856 124180 33862
rect 124128 33798 124180 33804
rect 122748 14476 122800 14482
rect 122748 14418 122800 14424
rect 125520 4078 125548 48758
rect 125704 48686 125732 52020
rect 125692 48680 125744 48686
rect 125692 48622 125744 48628
rect 126796 48680 126848 48686
rect 126796 48622 126848 48628
rect 126808 15978 126836 48622
rect 126796 15972 126848 15978
rect 126796 15914 126848 15920
rect 126900 4826 126928 52020
rect 128110 52006 128308 52034
rect 129306 52006 129688 52034
rect 130502 52006 131068 52034
rect 131698 52006 132448 52034
rect 126980 15904 127032 15910
rect 126980 15846 127032 15852
rect 126612 4820 126664 4826
rect 126612 4762 126664 4768
rect 126888 4820 126940 4826
rect 126888 4762 126940 4768
rect 125508 4072 125560 4078
rect 125508 4014 125560 4020
rect 121368 3664 121420 3670
rect 121368 3606 121420 3612
rect 118608 3256 118660 3262
rect 118608 3198 118660 3204
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 99288 3052 99340 3058
rect 99288 2994 99340 3000
rect 126624 480 126652 4762
rect 126992 3482 127020 15846
rect 128280 3874 128308 52006
rect 128452 49020 128504 49026
rect 128452 48962 128504 48968
rect 128268 3868 128320 3874
rect 128268 3810 128320 3816
rect 128464 3482 128492 48962
rect 129660 17338 129688 52006
rect 131040 35222 131068 52006
rect 131028 35216 131080 35222
rect 131028 35158 131080 35164
rect 129648 17332 129700 17338
rect 129648 17274 129700 17280
rect 131120 17264 131172 17270
rect 131120 17206 131172 17212
rect 130200 4888 130252 4894
rect 130200 4830 130252 4836
rect 126992 3454 127848 3482
rect 128464 3454 129044 3482
rect 127820 480 127848 3454
rect 129016 480 129044 3454
rect 130212 480 130240 4830
rect 131132 3482 131160 17206
rect 132420 3602 132448 52006
rect 132880 48822 132908 52020
rect 134076 48822 134104 52020
rect 135272 48822 135300 52020
rect 136482 52006 136588 52034
rect 137678 52006 137968 52034
rect 138874 52006 139348 52034
rect 139978 52006 140728 52034
rect 135444 49292 135496 49298
rect 135444 49234 135496 49240
rect 132868 48816 132920 48822
rect 132868 48758 132920 48764
rect 133788 48816 133840 48822
rect 133788 48758 133840 48764
rect 134064 48816 134116 48822
rect 134064 48758 134116 48764
rect 135168 48816 135220 48822
rect 135168 48758 135220 48764
rect 135260 48816 135312 48822
rect 135260 48758 135312 48764
rect 132592 18624 132644 18630
rect 132592 18566 132644 18572
rect 132408 3596 132460 3602
rect 132408 3538 132460 3544
rect 132604 3534 132632 18566
rect 133800 4894 133828 48758
rect 135180 43518 135208 48758
rect 135168 43512 135220 43518
rect 135168 43454 135220 43460
rect 133880 14544 133932 14550
rect 133880 14486 133932 14492
rect 133788 4888 133840 4894
rect 133788 4830 133840 4836
rect 132592 3528 132644 3534
rect 131132 3454 131436 3482
rect 132592 3470 132644 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 131408 480 131436 3454
rect 132592 3392 132644 3398
rect 132592 3334 132644 3340
rect 132604 480 132632 3334
rect 133800 480 133828 3470
rect 133892 3346 133920 14486
rect 135456 3346 135484 49234
rect 136456 48816 136508 48822
rect 136456 48758 136508 48764
rect 136468 3398 136496 48758
rect 136560 47666 136588 52006
rect 136548 47660 136600 47666
rect 136548 47602 136600 47608
rect 137940 36582 137968 52006
rect 138020 37936 138072 37942
rect 138020 37878 138072 37884
rect 137928 36576 137980 36582
rect 137928 36518 137980 36524
rect 136640 19984 136692 19990
rect 136640 19926 136692 19932
rect 136456 3392 136508 3398
rect 133892 3318 134932 3346
rect 135456 3318 136128 3346
rect 136456 3334 136508 3340
rect 136652 3346 136680 19926
rect 138032 3346 138060 37878
rect 139320 3534 139348 52006
rect 140700 18630 140728 52006
rect 141160 48822 141188 52020
rect 142252 49360 142304 49366
rect 142252 49302 142304 49308
rect 141148 48816 141200 48822
rect 141148 48758 141200 48764
rect 142068 48816 142120 48822
rect 142068 48758 142120 48764
rect 140780 39364 140832 39370
rect 140780 39306 140832 39312
rect 140688 18624 140740 18630
rect 140688 18566 140740 18572
rect 139676 4004 139728 4010
rect 139676 3946 139728 3952
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 136652 3318 137324 3346
rect 138032 3318 138520 3346
rect 134904 480 134932 3318
rect 136100 480 136128 3318
rect 137296 480 137324 3318
rect 138492 480 138520 3318
rect 139688 480 139716 3946
rect 140792 3466 140820 39306
rect 142080 38010 142108 48758
rect 142068 38004 142120 38010
rect 142068 37946 142120 37952
rect 140872 21412 140924 21418
rect 140872 21354 140924 21360
rect 140780 3460 140832 3466
rect 140780 3402 140832 3408
rect 140884 480 140912 21354
rect 142068 3460 142120 3466
rect 142068 3402 142120 3408
rect 142080 480 142108 3402
rect 142264 3346 142292 49302
rect 142356 48822 142384 52020
rect 143552 48822 143580 52020
rect 142344 48816 142396 48822
rect 142344 48758 142396 48764
rect 143448 48816 143500 48822
rect 143448 48758 143500 48764
rect 143540 48816 143592 48822
rect 143540 48758 143592 48764
rect 143460 4146 143488 48758
rect 144748 28286 144776 52020
rect 145944 49026 145972 52020
rect 147154 52006 147628 52034
rect 148350 52006 149008 52034
rect 145932 49020 145984 49026
rect 145932 48962 145984 48968
rect 144828 48816 144880 48822
rect 144828 48758 144880 48764
rect 144736 28280 144788 28286
rect 144736 28222 144788 28228
rect 143540 22772 143592 22778
rect 143540 22714 143592 22720
rect 143448 4140 143500 4146
rect 143448 4082 143500 4088
rect 143552 3346 143580 22714
rect 144840 19990 144868 48758
rect 144920 42084 144972 42090
rect 144920 42026 144972 42032
rect 144828 19984 144880 19990
rect 144828 19926 144880 19932
rect 144932 3346 144960 42026
rect 147600 21418 147628 52006
rect 148980 42090 149008 52006
rect 149532 48822 149560 52020
rect 150624 49224 150676 49230
rect 150624 49166 150676 49172
rect 149520 48816 149572 48822
rect 149520 48758 149572 48764
rect 150348 48816 150400 48822
rect 150348 48758 150400 48764
rect 148968 42084 149020 42090
rect 148968 42026 149020 42032
rect 149060 40724 149112 40730
rect 149060 40666 149112 40672
rect 147680 24132 147732 24138
rect 147680 24074 147732 24080
rect 147588 21412 147640 21418
rect 147588 21354 147640 21360
rect 146852 3936 146904 3942
rect 146852 3878 146904 3884
rect 142264 3318 143304 3346
rect 143552 3318 144500 3346
rect 144932 3318 145696 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3318
rect 146864 480 146892 3878
rect 147692 3346 147720 24074
rect 149072 3448 149100 40666
rect 149072 3420 149284 3448
rect 147692 3318 148088 3346
rect 148060 480 148088 3318
rect 149256 480 149284 3420
rect 150360 3330 150388 48758
rect 150532 25560 150584 25566
rect 150532 25502 150584 25508
rect 150544 3942 150572 25502
rect 150532 3936 150584 3942
rect 150532 3878 150584 3884
rect 150636 3482 150664 49166
rect 150728 48822 150756 52020
rect 151924 48822 151952 52020
rect 150716 48816 150768 48822
rect 150716 48758 150768 48764
rect 151728 48816 151780 48822
rect 151728 48758 151780 48764
rect 151912 48816 151964 48822
rect 151912 48758 151964 48764
rect 151740 22778 151768 48758
rect 151728 22772 151780 22778
rect 151728 22714 151780 22720
rect 151820 13184 151872 13190
rect 151820 13126 151872 13132
rect 151544 3936 151596 3942
rect 151544 3878 151596 3884
rect 150452 3454 150664 3482
rect 150348 3324 150400 3330
rect 150348 3266 150400 3272
rect 150452 480 150480 3454
rect 151556 480 151584 3878
rect 151832 3346 151860 13126
rect 153120 3505 153148 52020
rect 154330 52006 154528 52034
rect 155526 52006 155908 52034
rect 156722 52006 157288 52034
rect 153844 48816 153896 48822
rect 153844 48758 153896 48764
rect 153856 39370 153884 48758
rect 153844 39364 153896 39370
rect 153844 39306 153896 39312
rect 154500 24138 154528 52006
rect 155880 29714 155908 52006
rect 155960 47592 156012 47598
rect 155960 47534 156012 47540
rect 155868 29708 155920 29714
rect 155868 29650 155920 29656
rect 154580 26920 154632 26926
rect 154580 26862 154632 26868
rect 154488 24132 154540 24138
rect 154488 24074 154540 24080
rect 153106 3496 153162 3505
rect 153106 3431 153162 3440
rect 153934 3360 153990 3369
rect 151832 3318 152780 3346
rect 152752 480 152780 3318
rect 154592 3346 154620 26862
rect 155972 3346 156000 47534
rect 157260 3369 157288 52006
rect 157432 49156 157484 49162
rect 157432 49098 157484 49104
rect 157246 3360 157302 3369
rect 154592 3318 155172 3346
rect 155972 3318 156368 3346
rect 153934 3295 153990 3304
rect 153948 480 153976 3295
rect 155144 480 155172 3318
rect 156340 480 156368 3318
rect 157246 3295 157302 3304
rect 157444 1578 157472 49098
rect 157904 48822 157932 52020
rect 159100 48822 159128 52020
rect 160296 48822 160324 52020
rect 157892 48816 157944 48822
rect 157892 48758 157944 48764
rect 158628 48816 158680 48822
rect 158628 48758 158680 48764
rect 159088 48816 159140 48822
rect 159088 48758 159140 48764
rect 160008 48816 160060 48822
rect 160008 48758 160060 48764
rect 160284 48816 160336 48822
rect 160284 48758 160336 48764
rect 161388 48816 161440 48822
rect 161388 48758 161440 48764
rect 158640 25566 158668 48758
rect 160020 31142 160048 48758
rect 160008 31136 160060 31142
rect 160008 31078 160060 31084
rect 158812 28348 158864 28354
rect 158812 28290 158864 28296
rect 158628 25560 158680 25566
rect 158628 25502 158680 25508
rect 158824 3482 158852 28290
rect 161400 4010 161428 48758
rect 161492 48754 161520 52020
rect 162702 52006 162808 52034
rect 163898 52006 164188 52034
rect 165002 52006 165568 52034
rect 161480 48748 161532 48754
rect 161480 48690 161532 48696
rect 162780 40730 162808 52006
rect 162768 40724 162820 40730
rect 162768 40666 162820 40672
rect 162860 29640 162912 29646
rect 162860 29582 162912 29588
rect 162308 6180 162360 6186
rect 162308 6122 162360 6128
rect 161388 4004 161440 4010
rect 161388 3946 161440 3952
rect 158732 3454 158852 3482
rect 157444 1550 157564 1578
rect 157536 480 157564 1550
rect 158732 480 158760 3454
rect 161112 3188 161164 3194
rect 161112 3130 161164 3136
rect 159916 3052 159968 3058
rect 159916 2994 159968 3000
rect 159928 480 159956 2994
rect 161124 480 161152 3130
rect 162320 480 162348 6122
rect 162872 3482 162900 29582
rect 162872 3454 163544 3482
rect 164160 3466 164188 52006
rect 164332 49088 164384 49094
rect 164332 49030 164384 49036
rect 164344 3482 164372 49030
rect 165540 26926 165568 52006
rect 166184 48822 166212 52020
rect 167380 49162 167408 52020
rect 167368 49156 167420 49162
rect 167368 49098 167420 49104
rect 168576 48822 168604 52020
rect 169772 49706 169800 52020
rect 170982 52006 171088 52034
rect 172178 52006 172468 52034
rect 173374 52006 173848 52034
rect 174570 52006 175228 52034
rect 169760 49700 169812 49706
rect 169760 49642 169812 49648
rect 166172 48816 166224 48822
rect 166172 48758 166224 48764
rect 167736 48816 167788 48822
rect 167736 48758 167788 48764
rect 168564 48816 168616 48822
rect 168564 48758 168616 48764
rect 169668 48816 169720 48822
rect 169668 48758 169720 48764
rect 167644 48748 167696 48754
rect 167644 48690 167696 48696
rect 167092 31068 167144 31074
rect 167092 31010 167144 31016
rect 165528 26920 165580 26926
rect 165528 26862 165580 26868
rect 165896 7608 165948 7614
rect 165896 7550 165948 7556
rect 163516 480 163544 3454
rect 164148 3460 164200 3466
rect 164344 3454 164740 3482
rect 164148 3402 164200 3408
rect 164712 480 164740 3454
rect 165908 480 165936 7550
rect 167104 480 167132 31010
rect 167656 6322 167684 48690
rect 167748 32502 167776 48758
rect 167736 32496 167788 32502
rect 167736 32438 167788 32444
rect 169392 8968 169444 8974
rect 169392 8910 169444 8916
rect 167644 6316 167696 6322
rect 167644 6258 167696 6264
rect 168196 3120 168248 3126
rect 168196 3062 168248 3068
rect 168208 480 168236 3062
rect 169404 480 169432 8910
rect 169680 7614 169708 48758
rect 169668 7608 169720 7614
rect 169668 7550 169720 7556
rect 170588 6248 170640 6254
rect 170588 6190 170640 6196
rect 170600 480 170628 6190
rect 171060 3942 171088 52006
rect 172336 49700 172388 49706
rect 172336 49642 172388 49648
rect 172348 46306 172376 49642
rect 172336 46300 172388 46306
rect 172336 46242 172388 46248
rect 172440 8974 172468 52006
rect 173820 33794 173848 52006
rect 173900 46232 173952 46238
rect 173900 46174 173952 46180
rect 173808 33788 173860 33794
rect 173808 33730 173860 33736
rect 172520 10328 172572 10334
rect 172520 10270 172572 10276
rect 172428 8968 172480 8974
rect 172428 8910 172480 8916
rect 171048 3936 171100 3942
rect 171048 3878 171100 3884
rect 171784 3800 171836 3806
rect 171784 3742 171836 3748
rect 171796 480 171824 3742
rect 172532 3346 172560 10270
rect 173912 3346 173940 46174
rect 175200 3806 175228 52006
rect 175752 48618 175780 52020
rect 176948 48822 176976 52020
rect 178144 48822 178172 52020
rect 179248 52006 179354 52034
rect 180550 52006 180748 52034
rect 181746 52006 182128 52034
rect 182942 52006 183508 52034
rect 184138 52006 184888 52034
rect 176936 48816 176988 48822
rect 176936 48758 176988 48764
rect 177948 48816 178000 48822
rect 177948 48758 178000 48764
rect 178132 48816 178184 48822
rect 178132 48758 178184 48764
rect 175740 48612 175792 48618
rect 175740 48554 175792 48560
rect 176568 48612 176620 48618
rect 176568 48554 176620 48560
rect 175372 11756 175424 11762
rect 175372 11698 175424 11704
rect 175188 3800 175240 3806
rect 175188 3742 175240 3748
rect 175384 3738 175412 11698
rect 176580 10402 176608 48554
rect 177960 44878 177988 48758
rect 176660 44872 176712 44878
rect 176660 44814 176712 44820
rect 177948 44872 178000 44878
rect 177948 44814 178000 44820
rect 176568 10396 176620 10402
rect 176568 10338 176620 10344
rect 175280 3732 175332 3738
rect 175280 3674 175332 3680
rect 175372 3732 175424 3738
rect 175372 3674 175424 3680
rect 176568 3732 176620 3738
rect 176568 3674 176620 3680
rect 175292 3618 175320 3674
rect 175292 3590 175412 3618
rect 172532 3318 173020 3346
rect 173912 3318 174216 3346
rect 172992 480 173020 3318
rect 174188 480 174216 3318
rect 175384 480 175412 3590
rect 176580 480 176608 3674
rect 176672 3346 176700 44814
rect 179248 11762 179276 52006
rect 179328 48816 179380 48822
rect 179328 48758 179380 48764
rect 179236 11756 179288 11762
rect 179236 11698 179288 11704
rect 176672 3318 177804 3346
rect 177776 480 177804 3318
rect 179340 3262 179368 48758
rect 179420 13116 179472 13122
rect 179420 13058 179472 13064
rect 179432 3346 179460 13058
rect 180720 6186 180748 52006
rect 180800 32428 180852 32434
rect 180800 32370 180852 32376
rect 180708 6180 180760 6186
rect 180708 6122 180760 6128
rect 180812 3346 180840 32370
rect 182100 3738 182128 52006
rect 183480 13122 183508 52006
rect 184860 35290 184888 52006
rect 185320 48822 185348 52020
rect 186516 48822 186544 52020
rect 187712 48822 187740 52020
rect 188922 52006 189028 52034
rect 190118 52006 190408 52034
rect 191222 52006 191788 52034
rect 192418 52006 193168 52034
rect 185308 48816 185360 48822
rect 185308 48758 185360 48764
rect 186228 48816 186280 48822
rect 186228 48758 186280 48764
rect 186504 48816 186556 48822
rect 186504 48758 186556 48764
rect 187608 48816 187660 48822
rect 187608 48758 187660 48764
rect 187700 48816 187752 48822
rect 187700 48758 187752 48764
rect 184848 35284 184900 35290
rect 184848 35226 184900 35232
rect 183560 33856 183612 33862
rect 183560 33798 183612 33804
rect 183468 13116 183520 13122
rect 183468 13058 183520 13064
rect 182088 3732 182140 3738
rect 182088 3674 182140 3680
rect 183572 3670 183600 33798
rect 183652 14476 183704 14482
rect 183652 14418 183704 14424
rect 182548 3664 182600 3670
rect 182548 3606 182600 3612
rect 183560 3664 183612 3670
rect 183560 3606 183612 3612
rect 179432 3318 180196 3346
rect 180812 3318 181392 3346
rect 178960 3256 179012 3262
rect 178960 3198 179012 3204
rect 179328 3256 179380 3262
rect 179328 3198 179380 3204
rect 178972 480 179000 3198
rect 180168 480 180196 3318
rect 181364 480 181392 3318
rect 182560 480 182588 3606
rect 183664 3482 183692 14418
rect 186044 4072 186096 4078
rect 186044 4014 186096 4020
rect 184848 3664 184900 3670
rect 184848 3606 184900 3612
rect 183664 3454 183784 3482
rect 183756 480 183784 3454
rect 184860 480 184888 3606
rect 186056 480 186084 4014
rect 186240 3126 186268 48758
rect 186320 15972 186372 15978
rect 186320 15914 186372 15920
rect 186332 3346 186360 15914
rect 187620 14550 187648 48758
rect 187608 14544 187660 14550
rect 187608 14486 187660 14492
rect 188436 4820 188488 4826
rect 188436 4762 188488 4768
rect 186332 3318 187280 3346
rect 186228 3120 186280 3126
rect 186228 3062 186280 3068
rect 187252 480 187280 3318
rect 188448 480 188476 4762
rect 189000 3670 189028 52006
rect 189724 48816 189776 48822
rect 189724 48758 189776 48764
rect 189736 36650 189764 48758
rect 189724 36644 189776 36650
rect 189724 36586 189776 36592
rect 190380 4826 190408 52006
rect 191760 43450 191788 52006
rect 191748 43444 191800 43450
rect 191748 43386 191800 43392
rect 191840 35216 191892 35222
rect 191840 35158 191892 35164
rect 190460 17332 190512 17338
rect 190460 17274 190512 17280
rect 190368 4820 190420 4826
rect 190368 4762 190420 4768
rect 189632 3868 189684 3874
rect 189632 3810 189684 3816
rect 188988 3664 189040 3670
rect 188988 3606 189040 3612
rect 189644 480 189672 3810
rect 190472 3346 190500 17274
rect 191852 3346 191880 35158
rect 193140 4078 193168 52006
rect 193600 48822 193628 52020
rect 193588 48816 193640 48822
rect 193588 48758 193640 48764
rect 194508 48816 194560 48822
rect 194508 48758 194560 48764
rect 194520 15910 194548 48758
rect 194796 47734 194824 52020
rect 195992 48686 196020 52020
rect 195980 48680 196032 48686
rect 195980 48622 196032 48628
rect 194784 47728 194836 47734
rect 194784 47670 194836 47676
rect 194600 43512 194652 43518
rect 194600 43454 194652 43460
rect 194508 15904 194560 15910
rect 194508 15846 194560 15852
rect 194416 4888 194468 4894
rect 194416 4830 194468 4836
rect 193128 4072 193180 4078
rect 193128 4014 193180 4020
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 190472 3318 190868 3346
rect 191852 3318 192064 3346
rect 190840 480 190868 3318
rect 192036 480 192064 3318
rect 193232 480 193260 3538
rect 194428 480 194456 4830
rect 194612 3346 194640 43454
rect 197188 17270 197216 52020
rect 198398 52006 198688 52034
rect 199594 52006 200068 52034
rect 200790 52006 201448 52034
rect 197268 48680 197320 48686
rect 197268 48622 197320 48628
rect 197176 17264 197228 17270
rect 197176 17206 197228 17212
rect 197280 3398 197308 48622
rect 197360 47660 197412 47666
rect 197360 47602 197412 47608
rect 196808 3392 196860 3398
rect 194612 3318 195652 3346
rect 196808 3334 196860 3340
rect 197268 3392 197320 3398
rect 197268 3334 197320 3340
rect 197372 3346 197400 47602
rect 198660 37942 198688 52006
rect 198648 37936 198700 37942
rect 198648 37878 198700 37884
rect 198740 36576 198792 36582
rect 198740 36518 198792 36524
rect 198752 3346 198780 36518
rect 200040 3602 200068 52006
rect 201420 18698 201448 52006
rect 201972 48822 202000 52020
rect 203168 48822 203196 52020
rect 204364 48822 204392 52020
rect 205468 52006 205574 52034
rect 206770 52006 206968 52034
rect 207966 52006 208348 52034
rect 209162 52006 209728 52034
rect 201960 48816 202012 48822
rect 201960 48758 202012 48764
rect 202788 48816 202840 48822
rect 202788 48758 202840 48764
rect 203156 48816 203208 48822
rect 203156 48758 203208 48764
rect 204168 48816 204220 48822
rect 204168 48758 204220 48764
rect 204352 48816 204404 48822
rect 204352 48758 204404 48764
rect 202800 42158 202828 48758
rect 202788 42152 202840 42158
rect 202788 42094 202840 42100
rect 201500 38004 201552 38010
rect 201500 37946 201552 37952
rect 201408 18692 201460 18698
rect 201408 18634 201460 18640
rect 201512 3874 201540 37946
rect 201592 18624 201644 18630
rect 201592 18566 201644 18572
rect 201500 3868 201552 3874
rect 201500 3810 201552 3816
rect 200028 3596 200080 3602
rect 200028 3538 200080 3544
rect 200396 3528 200448 3534
rect 201604 3482 201632 18566
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 202696 3868 202748 3874
rect 202696 3810 202748 3816
rect 200396 3470 200448 3476
rect 195624 480 195652 3318
rect 196820 480 196848 3334
rect 197372 3318 198044 3346
rect 198752 3318 199240 3346
rect 198016 480 198044 3318
rect 199212 480 199240 3318
rect 200408 480 200436 3470
rect 201512 3454 201632 3482
rect 201512 480 201540 3454
rect 202708 480 202736 3810
rect 203904 480 203932 4082
rect 204180 3194 204208 48758
rect 205468 29646 205496 52006
rect 205548 48816 205600 48822
rect 205548 48758 205600 48764
rect 205456 29640 205508 29646
rect 205456 29582 205508 29588
rect 205560 19990 205588 48758
rect 205640 28280 205692 28286
rect 205640 28222 205692 28228
rect 204260 19984 204312 19990
rect 204260 19926 204312 19932
rect 205548 19984 205600 19990
rect 205548 19926 205600 19932
rect 204272 3346 204300 19926
rect 205652 3346 205680 28222
rect 206940 3534 206968 52006
rect 207112 49020 207164 49026
rect 207112 48962 207164 48968
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 207124 3346 207152 48962
rect 208320 28286 208348 52006
rect 208308 28280 208360 28286
rect 208308 28222 208360 28228
rect 208400 21412 208452 21418
rect 208400 21354 208452 21360
rect 208412 3346 208440 21354
rect 209700 4894 209728 52006
rect 210344 49230 210372 52020
rect 210332 49224 210384 49230
rect 210332 49166 210384 49172
rect 211540 48346 211568 52020
rect 212736 48822 212764 52020
rect 213932 48822 213960 52020
rect 212724 48816 212776 48822
rect 212724 48758 212776 48764
rect 213828 48816 213880 48822
rect 213828 48758 213880 48764
rect 213920 48816 213972 48822
rect 213920 48758 213972 48764
rect 211528 48340 211580 48346
rect 211528 48282 211580 48288
rect 212448 48340 212500 48346
rect 212448 48282 212500 48288
rect 209872 42084 209924 42090
rect 209872 42026 209924 42032
rect 209688 4888 209740 4894
rect 209688 4830 209740 4836
rect 204272 3318 205128 3346
rect 205652 3318 206324 3346
rect 207124 3318 207520 3346
rect 208412 3318 208716 3346
rect 204168 3188 204220 3194
rect 204168 3130 204220 3136
rect 205100 480 205128 3318
rect 206296 480 206324 3318
rect 207492 480 207520 3318
rect 208688 480 208716 3318
rect 209884 480 209912 42026
rect 211160 22772 211212 22778
rect 211160 22714 211212 22720
rect 211172 3346 211200 22714
rect 212460 21418 212488 48282
rect 213840 39370 213868 48758
rect 212540 39364 212592 39370
rect 212540 39306 212592 39312
rect 213828 39364 213880 39370
rect 213828 39306 213880 39312
rect 212448 21412 212500 21418
rect 212448 21354 212500 21360
rect 212552 3346 212580 39306
rect 215128 22778 215156 52020
rect 216246 52006 216628 52034
rect 215208 48816 215260 48822
rect 215208 48758 215260 48764
rect 215116 22772 215168 22778
rect 215116 22714 215168 22720
rect 215220 3874 215248 48758
rect 216600 31074 216628 52006
rect 217428 49094 217456 52020
rect 217416 49088 217468 49094
rect 217416 49030 217468 49036
rect 218624 48822 218652 52020
rect 219820 48822 219848 52020
rect 221016 48822 221044 52020
rect 222212 48822 222240 52020
rect 218612 48816 218664 48822
rect 218612 48758 218664 48764
rect 219348 48816 219400 48822
rect 219348 48758 219400 48764
rect 219808 48816 219860 48822
rect 219808 48758 219860 48764
rect 220728 48816 220780 48822
rect 220728 48758 220780 48764
rect 221004 48816 221056 48822
rect 221004 48758 221056 48764
rect 222108 48816 222160 48822
rect 222108 48758 222160 48764
rect 222200 48816 222252 48822
rect 222200 48758 222252 48764
rect 216588 31068 216640 31074
rect 216588 31010 216640 31016
rect 216680 29708 216732 29714
rect 216680 29650 216732 29656
rect 215300 24132 215352 24138
rect 215300 24074 215352 24080
rect 215208 3868 215260 3874
rect 215208 3810 215260 3816
rect 214654 3496 214710 3505
rect 214654 3431 214710 3440
rect 211068 3324 211120 3330
rect 211172 3318 212304 3346
rect 212552 3318 213500 3346
rect 211068 3266 211120 3272
rect 211080 480 211108 3266
rect 212276 480 212304 3318
rect 213472 480 213500 3318
rect 214668 480 214696 3431
rect 215312 3346 215340 24074
rect 216692 3346 216720 29650
rect 218060 25560 218112 25566
rect 218060 25502 218112 25508
rect 215312 3318 215892 3346
rect 216692 3318 217088 3346
rect 218072 3330 218100 25502
rect 219360 6254 219388 48758
rect 220740 40798 220768 48758
rect 220728 40792 220780 40798
rect 220728 40734 220780 40740
rect 219440 31136 219492 31142
rect 219440 31078 219492 31084
rect 219348 6248 219400 6254
rect 219348 6190 219400 6196
rect 218150 3360 218206 3369
rect 215864 480 215892 3318
rect 217060 480 217088 3318
rect 218060 3324 218112 3330
rect 219452 3346 219480 31078
rect 222120 4146 222148 48758
rect 223408 32434 223436 52020
rect 224604 49026 224632 52020
rect 225814 52006 226288 52034
rect 227010 52006 227668 52034
rect 224592 49020 224644 49026
rect 224592 48962 224644 48968
rect 223488 48816 223540 48822
rect 223488 48758 223540 48764
rect 223396 32428 223448 32434
rect 223396 32370 223448 32376
rect 223500 7682 223528 48758
rect 223580 40724 223632 40730
rect 223580 40666 223632 40672
rect 223488 7676 223540 7682
rect 223488 7618 223540 7624
rect 222936 6316 222988 6322
rect 222936 6258 222988 6264
rect 222108 4140 222160 4146
rect 222108 4082 222160 4088
rect 221740 4004 221792 4010
rect 221740 3946 221792 3952
rect 218150 3295 218206 3304
rect 219348 3324 219400 3330
rect 218060 3266 218112 3272
rect 218164 480 218192 3295
rect 219452 3318 220584 3346
rect 219348 3266 219400 3272
rect 219360 480 219388 3266
rect 220556 480 220584 3318
rect 221752 480 221780 3946
rect 222948 480 222976 6258
rect 223592 3346 223620 40666
rect 226260 24138 226288 52006
rect 227640 33862 227668 52006
rect 227904 49156 227956 49162
rect 227904 49098 227956 49104
rect 227628 33856 227680 33862
rect 227628 33798 227680 33804
rect 227812 32496 227864 32502
rect 227812 32438 227864 32444
rect 226340 26920 226392 26926
rect 226340 26862 226392 26868
rect 226248 24132 226300 24138
rect 226248 24074 226300 24080
rect 225328 3460 225380 3466
rect 225328 3402 225380 3408
rect 223592 3318 224172 3346
rect 224144 480 224172 3318
rect 225340 480 225368 3402
rect 226352 3346 226380 26862
rect 227824 3482 227852 32438
rect 227732 3454 227852 3482
rect 226352 3318 226564 3346
rect 226536 480 226564 3318
rect 227732 480 227760 3454
rect 227916 3346 227944 49098
rect 228192 48822 228220 52020
rect 229388 48822 229416 52020
rect 228180 48816 228232 48822
rect 228180 48758 228232 48764
rect 229008 48816 229060 48822
rect 229008 48758 229060 48764
rect 229376 48816 229428 48822
rect 229376 48758 229428 48764
rect 230388 48816 230440 48822
rect 230388 48758 230440 48764
rect 229020 4010 229048 48758
rect 230400 9110 230428 48758
rect 230480 46300 230532 46306
rect 230480 46242 230532 46248
rect 230388 9104 230440 9110
rect 230388 9046 230440 9052
rect 230112 7608 230164 7614
rect 230112 7550 230164 7556
rect 229008 4004 229060 4010
rect 229008 3946 229060 3952
rect 227916 3318 228956 3346
rect 228928 480 228956 3318
rect 230124 480 230152 7550
rect 230492 3482 230520 46242
rect 230584 46238 230612 52020
rect 230572 46232 230624 46238
rect 230572 46174 230624 46180
rect 230492 3454 231348 3482
rect 231320 480 231348 3454
rect 231780 3369 231808 52020
rect 232990 52006 233188 52034
rect 234186 52006 234568 52034
rect 233160 10334 233188 52006
rect 233148 10328 233200 10334
rect 233148 10270 233200 10276
rect 233700 8968 233752 8974
rect 233700 8910 233752 8916
rect 232504 3936 232556 3942
rect 232504 3878 232556 3884
rect 231766 3360 231822 3369
rect 231766 3295 231822 3304
rect 232516 480 232544 3878
rect 233712 480 233740 8910
rect 234540 7614 234568 52006
rect 235368 48822 235396 52020
rect 236578 52006 237328 52034
rect 235356 48816 235408 48822
rect 235356 48758 235408 48764
rect 236644 48816 236696 48822
rect 236644 48758 236696 48764
rect 234620 33788 234672 33794
rect 234620 33730 234672 33736
rect 234528 7608 234580 7614
rect 234528 7550 234580 7556
rect 234632 3482 234660 33730
rect 236656 28354 236684 48758
rect 236644 28348 236696 28354
rect 236644 28290 236696 28296
rect 237300 11830 237328 52006
rect 237760 48822 237788 52020
rect 238956 48822 238984 52020
rect 240152 48822 240180 52020
rect 237748 48816 237800 48822
rect 237748 48758 237800 48764
rect 238668 48816 238720 48822
rect 238668 48758 238720 48764
rect 238944 48816 238996 48822
rect 238944 48758 238996 48764
rect 240048 48816 240100 48822
rect 240048 48758 240100 48764
rect 240140 48816 240192 48822
rect 240140 48758 240192 48764
rect 238680 44946 238708 48758
rect 238668 44940 238720 44946
rect 238668 44882 238720 44888
rect 237380 44872 237432 44878
rect 237380 44814 237432 44820
rect 237288 11824 237340 11830
rect 237288 11766 237340 11772
rect 236092 10396 236144 10402
rect 236092 10338 236144 10344
rect 236000 3800 236052 3806
rect 236000 3742 236052 3748
rect 234632 3454 234844 3482
rect 234816 480 234844 3454
rect 236012 480 236040 3742
rect 236104 3482 236132 10338
rect 237392 3482 237420 44814
rect 240060 3806 240088 48758
rect 241348 35222 241376 52020
rect 241428 48816 241480 48822
rect 241428 48758 241480 48764
rect 241336 35216 241388 35222
rect 241336 35158 241388 35164
rect 241440 13190 241468 48758
rect 242452 47598 242480 52020
rect 243662 52006 244228 52034
rect 244858 52006 245608 52034
rect 242440 47592 242492 47598
rect 242440 47534 242492 47540
rect 244200 14482 244228 52006
rect 245580 36582 245608 52006
rect 246040 48822 246068 52020
rect 247236 48822 247264 52020
rect 246028 48816 246080 48822
rect 246028 48758 246080 48764
rect 246948 48816 247000 48822
rect 246948 48758 247000 48764
rect 247224 48816 247276 48822
rect 247224 48758 247276 48764
rect 248328 48816 248380 48822
rect 248328 48758 248380 48764
rect 245568 36576 245620 36582
rect 245568 36518 245620 36524
rect 244280 35284 244332 35290
rect 244280 35226 244332 35232
rect 244188 14476 244240 14482
rect 244188 14418 244240 14424
rect 241428 13184 241480 13190
rect 241428 13126 241480 13132
rect 240140 11756 240192 11762
rect 240140 11698 240192 11704
rect 240048 3800 240100 3806
rect 240048 3742 240100 3748
rect 236104 3454 237236 3482
rect 237392 3454 238432 3482
rect 237208 480 237236 3454
rect 238404 480 238432 3454
rect 240152 3346 240180 11698
rect 244292 7546 244320 35226
rect 244372 13116 244424 13122
rect 244372 13058 244424 13064
rect 244280 7540 244332 7546
rect 244280 7482 244332 7488
rect 241980 6180 242032 6186
rect 241980 6122 242032 6128
rect 240152 3318 240824 3346
rect 239588 3256 239640 3262
rect 239588 3198 239640 3204
rect 239600 480 239628 3198
rect 240796 480 240824 3318
rect 241992 480 242020 6122
rect 243176 3732 243228 3738
rect 243176 3674 243228 3680
rect 243188 480 243216 3674
rect 244384 480 244412 13058
rect 245568 7540 245620 7546
rect 245568 7482 245620 7488
rect 245580 480 245608 7482
rect 246960 3466 246988 48758
rect 247040 14544 247092 14550
rect 247040 14486 247092 14492
rect 247052 12442 247080 14486
rect 247040 12436 247092 12442
rect 247040 12378 247092 12384
rect 247960 12436 248012 12442
rect 247960 12378 248012 12384
rect 246948 3460 247000 3466
rect 246948 3402 247000 3408
rect 246764 3120 246816 3126
rect 246764 3062 246816 3068
rect 246776 480 246804 3062
rect 247972 480 248000 12378
rect 248340 5098 248368 48758
rect 248432 48550 248460 52020
rect 249642 52006 249748 52034
rect 250838 52006 251128 52034
rect 252034 52006 252508 52034
rect 248420 48544 248472 48550
rect 248420 48486 248472 48492
rect 249616 48544 249668 48550
rect 249616 48486 249668 48492
rect 249628 43518 249656 48486
rect 249616 43512 249668 43518
rect 249616 43454 249668 43460
rect 248420 36644 248472 36650
rect 248420 36586 248472 36592
rect 248432 28966 248460 36586
rect 248420 28960 248472 28966
rect 248420 28902 248472 28908
rect 248512 28960 248564 28966
rect 248512 28902 248564 28908
rect 248524 19394 248552 28902
rect 249720 24206 249748 52006
rect 251100 25566 251128 52006
rect 251088 25560 251140 25566
rect 251088 25502 251140 25508
rect 249708 24200 249760 24206
rect 249708 24142 249760 24148
rect 248432 19366 248552 19394
rect 248432 19310 248460 19366
rect 248420 19304 248472 19310
rect 248420 19246 248472 19252
rect 249156 9716 249208 9722
rect 249156 9658 249208 9664
rect 248328 5092 248380 5098
rect 248328 5034 248380 5040
rect 249168 480 249196 9658
rect 252480 6186 252508 52006
rect 253216 49162 253244 52020
rect 253204 49156 253256 49162
rect 253204 49098 253256 49104
rect 254412 48822 254440 52020
rect 255608 48822 255636 52020
rect 256804 48822 256832 52020
rect 257908 52006 258014 52034
rect 259210 52006 259408 52034
rect 254400 48816 254452 48822
rect 254400 48758 254452 48764
rect 255228 48816 255280 48822
rect 255228 48758 255280 48764
rect 255596 48816 255648 48822
rect 255596 48758 255648 48764
rect 256608 48816 256660 48822
rect 256608 48758 256660 48764
rect 256792 48816 256844 48822
rect 256792 48758 256844 48764
rect 252652 43444 252704 43450
rect 252652 43386 252704 43392
rect 252468 6180 252520 6186
rect 252468 6122 252520 6128
rect 251456 4820 251508 4826
rect 251456 4762 251508 4768
rect 250352 3664 250404 3670
rect 250352 3606 250404 3612
rect 250364 480 250392 3606
rect 251468 480 251496 4762
rect 252664 480 252692 43386
rect 255240 15978 255268 48758
rect 255320 47728 255372 47734
rect 255320 47670 255372 47676
rect 255228 15972 255280 15978
rect 255228 15914 255280 15920
rect 253940 15904 253992 15910
rect 253940 15846 253992 15852
rect 253952 12442 253980 15846
rect 255332 12442 255360 47670
rect 256620 38010 256648 48758
rect 256608 38004 256660 38010
rect 256608 37946 256660 37952
rect 257908 26926 257936 52006
rect 257988 48816 258040 48822
rect 257988 48758 258040 48764
rect 257896 26920 257948 26926
rect 257896 26862 257948 26868
rect 253940 12436 253992 12442
rect 253940 12378 253992 12384
rect 255044 12436 255096 12442
rect 255044 12378 255096 12384
rect 255320 12436 255372 12442
rect 255320 12378 255372 12384
rect 256240 12436 256292 12442
rect 256240 12378 256292 12384
rect 253848 4072 253900 4078
rect 253848 4014 253900 4020
rect 253860 480 253888 4014
rect 255056 480 255084 12378
rect 256252 480 256280 12378
rect 258000 9042 258028 48758
rect 259380 29714 259408 52006
rect 260392 48822 260420 52020
rect 261602 52006 262168 52034
rect 260380 48816 260432 48822
rect 260380 48758 260432 48764
rect 261484 48816 261536 48822
rect 261484 48758 261536 48764
rect 259460 37936 259512 37942
rect 259460 37878 259512 37884
rect 259368 29708 259420 29714
rect 259368 29650 259420 29656
rect 259472 19310 259500 37878
rect 261496 22846 261524 48758
rect 261484 22840 261536 22846
rect 261484 22782 261536 22788
rect 259460 19304 259512 19310
rect 259460 19246 259512 19252
rect 262140 17270 262168 52006
rect 262784 48754 262812 52020
rect 263980 48754 264008 52020
rect 265176 48822 265204 52020
rect 266372 48822 266400 52020
rect 267490 52006 267688 52034
rect 268686 52006 269068 52034
rect 269882 52006 270448 52034
rect 265164 48816 265216 48822
rect 265164 48758 265216 48764
rect 266268 48816 266320 48822
rect 266268 48758 266320 48764
rect 266360 48816 266412 48822
rect 266360 48758 266412 48764
rect 267556 48816 267608 48822
rect 267556 48758 267608 48764
rect 262772 48748 262824 48754
rect 262772 48690 262824 48696
rect 263508 48748 263560 48754
rect 263508 48690 263560 48696
rect 263968 48748 264020 48754
rect 263968 48690 264020 48696
rect 265624 48748 265676 48754
rect 265624 48690 265676 48696
rect 263520 42158 263548 48690
rect 262220 42152 262272 42158
rect 262220 42094 262272 42100
rect 263508 42152 263560 42158
rect 263508 42094 263560 42100
rect 258080 17264 258132 17270
rect 258080 17206 258132 17212
rect 262128 17264 262180 17270
rect 262128 17206 262180 17212
rect 258092 12442 258120 17206
rect 258080 12436 258132 12442
rect 258080 12378 258132 12384
rect 258632 12436 258684 12442
rect 258632 12378 258684 12384
rect 257988 9036 258040 9042
rect 257988 8978 258040 8984
rect 257436 3392 257488 3398
rect 257436 3334 257488 3340
rect 257448 480 257476 3334
rect 258644 480 258672 12378
rect 259828 9716 259880 9722
rect 259828 9658 259880 9664
rect 259840 480 259868 9658
rect 262232 7546 262260 42094
rect 264980 19984 265032 19990
rect 264980 19926 265032 19932
rect 262312 18692 262364 18698
rect 262312 18634 262364 18640
rect 262220 7540 262272 7546
rect 262220 7482 262272 7488
rect 262324 7426 262352 18634
rect 264992 12442 265020 19926
rect 264980 12436 265032 12442
rect 264980 12378 265032 12384
rect 265636 10402 265664 48690
rect 266280 18698 266308 48758
rect 267568 31142 267596 48758
rect 267556 31136 267608 31142
rect 267556 31078 267608 31084
rect 266360 29640 266412 29646
rect 266360 29582 266412 29588
rect 266268 18692 266320 18698
rect 266268 18634 266320 18640
rect 266372 12442 266400 29582
rect 265808 12436 265860 12442
rect 265808 12378 265860 12384
rect 266360 12436 266412 12442
rect 266360 12378 266412 12384
rect 267004 12436 267056 12442
rect 267004 12378 267056 12384
rect 265624 10396 265676 10402
rect 265624 10338 265676 10344
rect 263416 7540 263468 7546
rect 263416 7482 263468 7488
rect 262232 7398 262352 7426
rect 261024 3596 261076 3602
rect 261024 3538 261076 3544
rect 261036 480 261064 3538
rect 262232 480 262260 7398
rect 263428 480 263456 7482
rect 264612 3188 264664 3194
rect 264612 3130 264664 3136
rect 264624 480 264652 3130
rect 265820 480 265848 12378
rect 267016 480 267044 12378
rect 267660 11762 267688 52006
rect 269040 19990 269068 52006
rect 269120 28280 269172 28286
rect 269120 28222 269172 28228
rect 269028 19984 269080 19990
rect 269028 19926 269080 19932
rect 269132 19310 269160 28222
rect 269120 19304 269172 19310
rect 269120 19246 269172 19252
rect 267648 11756 267700 11762
rect 267648 11698 267700 11704
rect 269304 9716 269356 9722
rect 269304 9658 269356 9664
rect 268108 3528 268160 3534
rect 268108 3470 268160 3476
rect 268120 480 268148 3470
rect 269316 480 269344 9658
rect 270420 4826 270448 52006
rect 270500 49224 270552 49230
rect 270500 49166 270552 49172
rect 270512 7546 270540 49166
rect 271064 48754 271092 52020
rect 272260 48822 272288 52020
rect 273456 48822 273484 52020
rect 274652 48822 274680 52020
rect 272248 48816 272300 48822
rect 272248 48758 272300 48764
rect 273168 48816 273220 48822
rect 273168 48758 273220 48764
rect 273444 48816 273496 48822
rect 273444 48758 273496 48764
rect 274548 48816 274600 48822
rect 274548 48758 274600 48764
rect 274640 48816 274692 48822
rect 274640 48758 274692 48764
rect 271052 48748 271104 48754
rect 271052 48690 271104 48696
rect 272524 48748 272576 48754
rect 272524 48690 272576 48696
rect 271880 21412 271932 21418
rect 271880 21354 271932 21360
rect 271892 12442 271920 21354
rect 272536 13258 272564 48690
rect 273180 21418 273208 48758
rect 274560 39438 274588 48758
rect 275848 47666 275876 52020
rect 277058 52006 277348 52034
rect 276664 48816 276716 48822
rect 276664 48758 276716 48764
rect 275836 47660 275888 47666
rect 275836 47602 275888 47608
rect 274548 39432 274600 39438
rect 274548 39374 274600 39380
rect 273260 39364 273312 39370
rect 273260 39306 273312 39312
rect 273168 21412 273220 21418
rect 273168 21354 273220 21360
rect 272524 13252 272576 13258
rect 272524 13194 272576 13200
rect 273272 12442 273300 39306
rect 276020 22772 276072 22778
rect 276020 22714 276072 22720
rect 276032 12510 276060 22714
rect 276676 14618 276704 48758
rect 277320 40730 277348 52006
rect 278240 48686 278268 52020
rect 279450 52006 280108 52034
rect 278228 48680 278280 48686
rect 278228 48622 278280 48628
rect 278964 48340 279016 48346
rect 278964 48282 279016 48288
rect 277308 40724 277360 40730
rect 277308 40666 277360 40672
rect 277400 31068 277452 31074
rect 277400 31010 277452 31016
rect 277412 19310 277440 31010
rect 278976 19310 279004 48282
rect 277400 19304 277452 19310
rect 277400 19246 277452 19252
rect 277768 19304 277820 19310
rect 277768 19246 277820 19252
rect 278964 19304 279016 19310
rect 278964 19246 279016 19252
rect 276664 14612 276716 14618
rect 276664 14554 276716 14560
rect 276020 12504 276072 12510
rect 276020 12446 276072 12452
rect 271880 12436 271932 12442
rect 271880 12378 271932 12384
rect 272892 12436 272944 12442
rect 272892 12378 272944 12384
rect 273260 12436 273312 12442
rect 273260 12378 273312 12384
rect 274088 12436 274140 12442
rect 274088 12378 274140 12384
rect 270500 7540 270552 7546
rect 270500 7482 270552 7488
rect 271696 7540 271748 7546
rect 271696 7482 271748 7488
rect 270592 4888 270644 4894
rect 270592 4830 270644 4836
rect 270408 4820 270460 4826
rect 270408 4762 270460 4768
rect 270604 2666 270632 4830
rect 270512 2638 270632 2666
rect 270512 480 270540 2638
rect 271708 480 271736 7482
rect 272904 480 272932 12378
rect 274100 480 274128 12378
rect 276480 12368 276532 12374
rect 276480 12310 276532 12316
rect 276492 9654 276520 12310
rect 276480 9648 276532 9654
rect 276480 9590 276532 9596
rect 276480 9512 276532 9518
rect 276480 9454 276532 9460
rect 275284 3868 275336 3874
rect 275284 3810 275336 3816
rect 275296 480 275324 3810
rect 276492 480 276520 9454
rect 277780 4876 277808 19246
rect 278964 9716 279016 9722
rect 278964 9658 279016 9664
rect 277688 4848 277808 4876
rect 277688 480 277716 4848
rect 278976 2938 279004 9658
rect 280080 6254 280108 52006
rect 280632 48822 280660 52020
rect 281828 49230 281856 52020
rect 281816 49224 281868 49230
rect 281816 49166 281868 49172
rect 283024 48822 283052 52020
rect 284128 52006 284234 52034
rect 285430 52006 285628 52034
rect 286626 52006 287008 52034
rect 287822 52006 288388 52034
rect 280620 48816 280672 48822
rect 280620 48758 280672 48764
rect 281448 48816 281500 48822
rect 281448 48758 281500 48764
rect 283012 48816 283064 48822
rect 283012 48758 283064 48764
rect 280804 48680 280856 48686
rect 280804 48622 280856 48628
rect 280160 40792 280212 40798
rect 280160 40734 280212 40740
rect 280172 12442 280200 40734
rect 280816 28422 280844 48622
rect 281460 32502 281488 48758
rect 284128 33794 284156 52006
rect 284208 48816 284260 48822
rect 284208 48758 284260 48764
rect 284116 33788 284168 33794
rect 284116 33730 284168 33736
rect 281448 32496 281500 32502
rect 281448 32438 281500 32444
rect 280804 28416 280856 28422
rect 280804 28358 280856 28364
rect 280160 12436 280212 12442
rect 280160 12378 280212 12384
rect 281264 12436 281316 12442
rect 281264 12378 281316 12384
rect 279976 6248 280028 6254
rect 279976 6190 280028 6196
rect 280068 6248 280120 6254
rect 280068 6190 280120 6196
rect 279988 6066 280016 6190
rect 279988 6038 280108 6066
rect 278976 2910 279096 2938
rect 279068 2666 279096 2910
rect 278884 2638 279096 2666
rect 278884 480 278912 2638
rect 280080 480 280108 6038
rect 281276 480 281304 12378
rect 284220 7818 284248 48758
rect 284300 32428 284352 32434
rect 284300 32370 284352 32376
rect 284312 19310 284340 32370
rect 284300 19304 284352 19310
rect 284300 19246 284352 19252
rect 285600 15910 285628 52006
rect 285772 49020 285824 49026
rect 285772 48962 285824 48968
rect 285784 46918 285812 48962
rect 285772 46912 285824 46918
rect 285772 46854 285824 46860
rect 285772 37324 285824 37330
rect 285772 37266 285824 37272
rect 285784 27606 285812 37266
rect 285772 27600 285824 27606
rect 285772 27542 285824 27548
rect 286980 22778 287008 52006
rect 288360 35290 288388 52006
rect 289004 48754 289032 52020
rect 290200 48822 290228 52020
rect 290188 48816 290240 48822
rect 290188 48758 290240 48764
rect 291108 48816 291160 48822
rect 291108 48758 291160 48764
rect 288992 48748 289044 48754
rect 288992 48690 289044 48696
rect 290464 48748 290516 48754
rect 290464 48690 290516 48696
rect 288348 35284 288400 35290
rect 288348 35226 288400 35232
rect 287060 33856 287112 33862
rect 287060 33798 287112 33804
rect 286968 22772 287020 22778
rect 286968 22714 287020 22720
rect 285588 15904 285640 15910
rect 285588 15846 285640 15852
rect 284760 9716 284812 9722
rect 284760 9658 284812 9664
rect 285956 9716 286008 9722
rect 285956 9658 286008 9664
rect 284208 7812 284260 7818
rect 284208 7754 284260 7760
rect 283656 7676 283708 7682
rect 283656 7618 283708 7624
rect 282460 4140 282512 4146
rect 282460 4082 282512 4088
rect 282472 480 282500 4082
rect 283668 480 283696 7618
rect 284772 480 284800 9658
rect 285968 480 285996 9658
rect 287072 7682 287100 33798
rect 287152 24132 287204 24138
rect 287152 24074 287204 24080
rect 287060 7676 287112 7682
rect 287060 7618 287112 7624
rect 287164 480 287192 24074
rect 290476 17338 290504 48690
rect 290464 17332 290516 17338
rect 290464 17274 290516 17280
rect 291120 9110 291148 48758
rect 291396 46306 291424 52020
rect 292592 48686 292620 52020
rect 292580 48680 292632 48686
rect 292580 48622 292632 48628
rect 293696 48414 293724 52020
rect 294906 52006 295288 52034
rect 293868 48680 293920 48686
rect 293868 48622 293920 48628
rect 293684 48408 293736 48414
rect 293684 48350 293736 48356
rect 291384 46300 291436 46306
rect 291384 46242 291436 46248
rect 291200 46232 291252 46238
rect 291200 46174 291252 46180
rect 291212 12442 291240 46174
rect 291200 12436 291252 12442
rect 291200 12378 291252 12384
rect 291936 12436 291988 12442
rect 291936 12378 291988 12384
rect 290740 9104 290792 9110
rect 290740 9046 290792 9052
rect 291108 9104 291160 9110
rect 291108 9046 291160 9052
rect 288348 7676 288400 7682
rect 288348 7618 288400 7624
rect 288360 480 288388 7618
rect 289544 4004 289596 4010
rect 289544 3946 289596 3952
rect 289556 480 289584 3946
rect 290752 480 290780 9046
rect 291948 480 291976 12378
rect 293880 7750 293908 48622
rect 294604 48408 294656 48414
rect 294604 48350 294656 48356
rect 294616 10334 294644 48350
rect 295260 44878 295288 52006
rect 296088 49094 296116 52020
rect 297298 52006 298048 52034
rect 296076 49088 296128 49094
rect 296076 49030 296128 49036
rect 295248 44872 295300 44878
rect 295248 44814 295300 44820
rect 296720 28348 296772 28354
rect 296720 28290 296772 28296
rect 294328 10328 294380 10334
rect 294328 10270 294380 10276
rect 294604 10328 294656 10334
rect 294604 10270 294656 10276
rect 293868 7744 293920 7750
rect 293868 7686 293920 7692
rect 293130 3360 293186 3369
rect 293130 3295 293186 3304
rect 293144 480 293172 3295
rect 294340 480 294368 10270
rect 295524 7608 295576 7614
rect 295524 7550 295576 7556
rect 295536 480 295564 7550
rect 296732 480 296760 28290
rect 298020 11830 298048 52006
rect 298480 48822 298508 52020
rect 299676 48822 299704 52020
rect 298468 48816 298520 48822
rect 298468 48758 298520 48764
rect 299388 48816 299440 48822
rect 299388 48758 299440 48764
rect 299664 48816 299716 48822
rect 299664 48758 299716 48764
rect 298100 44940 298152 44946
rect 298100 44882 298152 44888
rect 298112 12442 298140 44882
rect 299400 36650 299428 48758
rect 300872 48550 300900 52020
rect 301504 48816 301556 48822
rect 301504 48758 301556 48764
rect 300860 48544 300912 48550
rect 300860 48486 300912 48492
rect 299388 36644 299440 36650
rect 299388 36586 299440 36592
rect 298100 12436 298152 12442
rect 298100 12378 298152 12384
rect 299112 12436 299164 12442
rect 299112 12378 299164 12384
rect 297916 11824 297968 11830
rect 297916 11766 297968 11772
rect 298008 11824 298060 11830
rect 298008 11766 298060 11772
rect 297928 480 297956 11766
rect 299124 480 299152 12378
rect 301412 9716 301464 9722
rect 301412 9658 301464 9664
rect 301424 9602 301452 9658
rect 301332 9574 301452 9602
rect 300308 3800 300360 3806
rect 300308 3742 300360 3748
rect 300320 480 300348 3742
rect 301332 610 301360 9574
rect 301516 6322 301544 48758
rect 302068 43450 302096 52020
rect 303278 52006 303568 52034
rect 304474 52006 304948 52034
rect 305670 52006 306328 52034
rect 302148 48544 302200 48550
rect 302148 48486 302200 48492
rect 302056 43444 302108 43450
rect 302056 43386 302108 43392
rect 302160 13122 302188 48486
rect 302240 35216 302292 35222
rect 302240 35158 302292 35164
rect 302148 13116 302200 13122
rect 302148 13058 302200 13064
rect 301504 6316 301556 6322
rect 301504 6258 301556 6264
rect 302252 3482 302280 35158
rect 303540 18630 303568 52006
rect 303620 47592 303672 47598
rect 303620 47534 303672 47540
rect 303528 18624 303580 18630
rect 303528 18566 303580 18572
rect 303632 3482 303660 47534
rect 304920 14550 304948 52006
rect 305000 36576 305052 36582
rect 305000 36518 305052 36524
rect 304908 14544 304960 14550
rect 304908 14486 304960 14492
rect 305012 3534 305040 36518
rect 306300 25634 306328 52006
rect 306852 48754 306880 52020
rect 308048 48822 308076 52020
rect 309244 49230 309272 52020
rect 308404 49224 308456 49230
rect 308404 49166 308456 49172
rect 309232 49224 309284 49230
rect 309232 49166 309284 49172
rect 308036 48816 308088 48822
rect 308036 48758 308088 48764
rect 306840 48748 306892 48754
rect 306840 48690 306892 48696
rect 306288 25628 306340 25634
rect 306288 25570 306340 25576
rect 305092 14476 305144 14482
rect 305092 14418 305144 14424
rect 305000 3528 305052 3534
rect 302252 3454 302648 3482
rect 303632 3454 303844 3482
rect 305000 3470 305052 3476
rect 301320 604 301372 610
rect 301320 546 301372 552
rect 301412 604 301464 610
rect 301412 546 301464 552
rect 301424 480 301452 546
rect 302620 480 302648 3454
rect 303816 480 303844 3454
rect 305104 1442 305132 14418
rect 308416 4894 308444 49166
rect 309048 48816 309100 48822
rect 309048 48758 309100 48764
rect 309060 24274 309088 48758
rect 309140 43512 309192 43518
rect 309140 43454 309192 43460
rect 309048 24268 309100 24274
rect 309048 24210 309100 24216
rect 308588 4956 308640 4962
rect 308588 4898 308640 4904
rect 308404 4888 308456 4894
rect 308404 4830 308456 4836
rect 306196 3528 306248 3534
rect 306196 3470 306248 3476
rect 305012 1414 305132 1442
rect 305012 480 305040 1414
rect 306208 480 306236 3470
rect 307392 3460 307444 3466
rect 307392 3402 307444 3408
rect 307404 480 307432 3402
rect 308600 480 308628 4898
rect 309152 3346 309180 43454
rect 310440 8974 310468 52020
rect 311650 52006 311848 52034
rect 312846 52006 313228 52034
rect 314042 52006 314608 52034
rect 311820 28286 311848 52006
rect 312544 48748 312596 48754
rect 312544 48690 312596 48696
rect 311808 28280 311860 28286
rect 311808 28222 311860 28228
rect 311900 25560 311952 25566
rect 311900 25502 311952 25508
rect 310520 24200 310572 24206
rect 310520 24142 310572 24148
rect 310428 8968 310480 8974
rect 310428 8910 310480 8916
rect 310532 3346 310560 24142
rect 311912 3346 311940 25502
rect 312556 20058 312584 48690
rect 313200 37942 313228 52006
rect 313464 49156 313516 49162
rect 313464 49098 313516 49104
rect 313188 37936 313240 37942
rect 313188 37878 313240 37884
rect 312544 20052 312596 20058
rect 312544 19994 312596 20000
rect 313372 6180 313424 6186
rect 313372 6122 313424 6128
rect 309152 3318 309824 3346
rect 310532 3318 311020 3346
rect 311912 3318 312216 3346
rect 309796 480 309824 3318
rect 310992 480 311020 3318
rect 312188 480 312216 3318
rect 313384 480 313412 6122
rect 313476 3346 313504 49098
rect 314580 3466 314608 52006
rect 315224 48618 315252 52020
rect 316420 48822 316448 52020
rect 316408 48816 316460 48822
rect 316408 48758 316460 48764
rect 317328 48816 317380 48822
rect 317328 48758 317380 48764
rect 315212 48612 315264 48618
rect 315212 48554 315264 48560
rect 315948 48612 316000 48618
rect 315948 48554 316000 48560
rect 315960 15978 315988 48554
rect 316040 38004 316092 38010
rect 316040 37946 316092 37952
rect 314660 15972 314712 15978
rect 314660 15914 314712 15920
rect 315948 15972 316000 15978
rect 315948 15914 316000 15920
rect 314568 3460 314620 3466
rect 314568 3402 314620 3408
rect 314672 3346 314700 15914
rect 316052 3346 316080 37946
rect 317340 29646 317368 48758
rect 317616 48346 317644 52020
rect 318720 49026 318748 52020
rect 319930 52006 320128 52034
rect 321126 52006 321508 52034
rect 322322 52006 322888 52034
rect 319444 49224 319496 49230
rect 319444 49166 319496 49172
rect 318708 49020 318760 49026
rect 318708 48962 318760 48968
rect 317604 48340 317656 48346
rect 317604 48282 317656 48288
rect 318708 48340 318760 48346
rect 318708 48282 318760 48288
rect 317328 29640 317380 29646
rect 317328 29582 317380 29588
rect 318064 9036 318116 9042
rect 318064 8978 318116 8984
rect 313476 3318 314608 3346
rect 314672 3318 315804 3346
rect 316052 3318 317000 3346
rect 314580 480 314608 3318
rect 315776 480 315804 3318
rect 316972 480 317000 3318
rect 318076 480 318104 8978
rect 318720 3534 318748 48282
rect 319456 26994 319484 49166
rect 320100 42090 320128 52006
rect 320088 42084 320140 42090
rect 320088 42026 320140 42032
rect 320180 29708 320232 29714
rect 320180 29650 320232 29656
rect 319444 26988 319496 26994
rect 319444 26930 319496 26936
rect 318800 26920 318852 26926
rect 318800 26862 318852 26868
rect 318708 3528 318760 3534
rect 318708 3470 318760 3476
rect 318812 3346 318840 26862
rect 320192 3346 320220 29650
rect 321480 3670 321508 52006
rect 321560 22840 321612 22846
rect 321560 22782 321612 22788
rect 321468 3664 321520 3670
rect 321468 3606 321520 3612
rect 321572 3482 321600 22782
rect 322860 17270 322888 52006
rect 323504 48822 323532 52020
rect 324700 48822 324728 52020
rect 325896 48822 325924 52020
rect 327092 48822 327120 52020
rect 328302 52006 328408 52034
rect 323492 48816 323544 48822
rect 323492 48758 323544 48764
rect 324228 48816 324280 48822
rect 324228 48758 324280 48764
rect 324688 48816 324740 48822
rect 324688 48758 324740 48764
rect 325608 48816 325660 48822
rect 325608 48758 325660 48764
rect 325884 48816 325936 48822
rect 325884 48758 325936 48764
rect 326988 48816 327040 48822
rect 326988 48758 327040 48764
rect 327080 48816 327132 48822
rect 327080 48758 327132 48764
rect 328276 48816 328328 48822
rect 328276 48758 328328 48764
rect 322940 42152 322992 42158
rect 322940 42094 322992 42100
rect 321652 17264 321704 17270
rect 321652 17206 321704 17212
rect 322848 17264 322900 17270
rect 322848 17206 322900 17212
rect 321664 3602 321692 17206
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 321572 3454 321692 3482
rect 318812 3318 319300 3346
rect 320192 3318 320496 3346
rect 319272 480 319300 3318
rect 320468 480 320496 3318
rect 321664 480 321692 3454
rect 322860 480 322888 3538
rect 322952 3346 322980 42094
rect 324240 31074 324268 48758
rect 324228 31068 324280 31074
rect 324228 31010 324280 31016
rect 324320 10396 324372 10402
rect 324320 10338 324372 10344
rect 324332 3346 324360 10338
rect 322952 3318 324084 3346
rect 324332 3318 325280 3346
rect 324056 480 324084 3318
rect 325252 480 325280 3318
rect 325620 3194 325648 48758
rect 327000 18698 327028 48758
rect 328288 39370 328316 48758
rect 328276 39364 328328 39370
rect 328276 39306 328328 39312
rect 327080 31136 327132 31142
rect 327080 31078 327132 31084
rect 325700 18692 325752 18698
rect 325700 18634 325752 18640
rect 326988 18692 327040 18698
rect 326988 18634 327040 18640
rect 325712 3346 325740 18634
rect 327092 3346 327120 31078
rect 328380 3738 328408 52006
rect 329484 48822 329512 52020
rect 330694 52006 331168 52034
rect 331890 52006 332548 52034
rect 329472 48816 329524 48822
rect 329472 48758 329524 48764
rect 330484 48816 330536 48822
rect 330484 48758 330536 48764
rect 330496 19990 330524 48758
rect 331140 40798 331168 52006
rect 331128 40792 331180 40798
rect 331128 40734 331180 40740
rect 329840 19984 329892 19990
rect 329840 19926 329892 19932
rect 330484 19984 330536 19990
rect 330484 19926 330536 19932
rect 328460 11756 328512 11762
rect 328460 11698 328512 11704
rect 328368 3732 328420 3738
rect 328368 3674 328420 3680
rect 328472 3346 328500 11698
rect 329852 3346 329880 19926
rect 331220 13252 331272 13258
rect 331220 13194 331272 13200
rect 331232 3534 331260 13194
rect 331312 4820 331364 4826
rect 331312 4762 331364 4768
rect 331220 3528 331272 3534
rect 331220 3470 331272 3476
rect 331324 3346 331352 4762
rect 332520 3874 332548 52006
rect 333072 48822 333100 52020
rect 333244 49088 333296 49094
rect 333244 49030 333296 49036
rect 333060 48816 333112 48822
rect 333060 48758 333112 48764
rect 332600 21412 332652 21418
rect 332600 21354 332652 21360
rect 332508 3868 332560 3874
rect 332508 3810 332560 3816
rect 332416 3528 332468 3534
rect 332416 3470 332468 3476
rect 325712 3318 326476 3346
rect 327092 3318 327672 3346
rect 328472 3318 328868 3346
rect 329852 3318 330064 3346
rect 325608 3188 325660 3194
rect 325608 3130 325660 3136
rect 326448 480 326476 3318
rect 327644 480 327672 3318
rect 328840 480 328868 3318
rect 330036 480 330064 3318
rect 331232 3318 331352 3346
rect 331232 480 331260 3318
rect 332428 480 332456 3470
rect 332612 3346 332640 21354
rect 333256 4826 333284 49030
rect 333888 48816 333940 48822
rect 333888 48758 333940 48764
rect 333900 21418 333928 48758
rect 334268 48754 334296 52020
rect 335464 48822 335492 52020
rect 336660 48906 336688 52020
rect 337870 52006 338068 52034
rect 339066 52006 339448 52034
rect 340262 52006 340828 52034
rect 341458 52006 342208 52034
rect 336660 48878 336872 48906
rect 335452 48816 335504 48822
rect 335452 48758 335504 48764
rect 336648 48816 336700 48822
rect 336648 48758 336700 48764
rect 334256 48748 334308 48754
rect 334256 48690 334308 48696
rect 335268 48748 335320 48754
rect 335268 48690 335320 48696
rect 333980 39432 334032 39438
rect 333980 39374 334032 39380
rect 333888 21412 333940 21418
rect 333888 21354 333940 21360
rect 333244 4820 333296 4826
rect 333244 4762 333296 4768
rect 333992 3346 334020 39374
rect 335280 32434 335308 48690
rect 335268 32428 335320 32434
rect 335268 32370 335320 32376
rect 335360 14612 335412 14618
rect 335360 14554 335412 14560
rect 335372 3346 335400 14554
rect 336660 4146 336688 48758
rect 336740 47660 336792 47666
rect 336740 47602 336792 47608
rect 336648 4140 336700 4146
rect 336648 4082 336700 4088
rect 336752 3346 336780 47602
rect 336844 47598 336872 48878
rect 336832 47592 336884 47598
rect 336832 47534 336884 47540
rect 338040 33862 338068 52006
rect 338120 40724 338172 40730
rect 338120 40666 338172 40672
rect 338028 33856 338080 33862
rect 338028 33798 338080 33804
rect 338132 3346 338160 40666
rect 339420 3466 339448 52006
rect 339500 28416 339552 28422
rect 339500 28358 339552 28364
rect 339408 3460 339460 3466
rect 339408 3402 339460 3408
rect 332612 3318 333652 3346
rect 333992 3318 334756 3346
rect 335372 3318 335952 3346
rect 336752 3318 337148 3346
rect 338132 3318 338344 3346
rect 333624 480 333652 3318
rect 334728 480 334756 3318
rect 335924 480 335952 3318
rect 337120 480 337148 3318
rect 338316 480 338344 3318
rect 339512 480 339540 28358
rect 340696 6248 340748 6254
rect 340696 6190 340748 6196
rect 340708 480 340736 6190
rect 340800 6186 340828 52006
rect 342180 35222 342208 52006
rect 342640 48550 342668 52020
rect 343744 48822 343772 52020
rect 344848 52006 344954 52034
rect 346150 52006 346348 52034
rect 343732 48816 343784 48822
rect 343732 48758 343784 48764
rect 342628 48544 342680 48550
rect 342628 48486 342680 48492
rect 343548 48544 343600 48550
rect 343548 48486 343600 48492
rect 342168 35216 342220 35222
rect 342168 35158 342220 35164
rect 340880 32496 340932 32502
rect 340880 32438 340932 32444
rect 340788 6180 340840 6186
rect 340788 6122 340840 6128
rect 340892 3346 340920 32438
rect 343088 4888 343140 4894
rect 343088 4830 343140 4836
rect 340892 3318 341932 3346
rect 341904 480 341932 3318
rect 343100 480 343128 4830
rect 343560 4010 343588 48486
rect 344848 46238 344876 52006
rect 344928 48816 344980 48822
rect 344928 48758 344980 48764
rect 344836 46232 344888 46238
rect 344836 46174 344888 46180
rect 344284 7676 344336 7682
rect 344284 7618 344336 7624
rect 343548 4004 343600 4010
rect 343548 3946 343600 3952
rect 344296 480 344324 7618
rect 344940 7614 344968 48758
rect 345020 33788 345072 33794
rect 345020 33730 345072 33736
rect 344928 7608 344980 7614
rect 344928 7550 344980 7556
rect 345032 3482 345060 33730
rect 345032 3454 345520 3482
rect 345492 480 345520 3454
rect 346320 3398 346348 52006
rect 347332 48822 347360 52020
rect 348542 52006 349108 52034
rect 349738 52006 350488 52034
rect 347320 48816 347372 48822
rect 347320 48758 347372 48764
rect 348424 48816 348476 48822
rect 348424 48758 348476 48764
rect 347780 35284 347832 35290
rect 347780 35226 347832 35232
rect 346400 15904 346452 15910
rect 346400 15846 346452 15852
rect 346412 3482 346440 15846
rect 347792 3534 347820 35226
rect 348436 22778 348464 48758
rect 349080 44946 349108 52006
rect 349068 44940 349120 44946
rect 349068 44882 349120 44888
rect 347872 22772 347924 22778
rect 347872 22714 347924 22720
rect 348424 22772 348476 22778
rect 348424 22714 348476 22720
rect 347780 3528 347832 3534
rect 346412 3454 346716 3482
rect 347780 3470 347832 3476
rect 346308 3392 346360 3398
rect 346308 3334 346360 3340
rect 346688 480 346716 3454
rect 347884 480 347912 22714
rect 349160 17332 349212 17338
rect 349160 17274 349212 17280
rect 349068 3528 349120 3534
rect 349068 3470 349120 3476
rect 349172 3482 349200 17274
rect 350460 3806 350488 52006
rect 350920 48822 350948 52020
rect 350908 48816 350960 48822
rect 350908 48758 350960 48764
rect 351828 48816 351880 48822
rect 351828 48758 351880 48764
rect 351368 9104 351420 9110
rect 351368 9046 351420 9052
rect 350448 3800 350500 3806
rect 350448 3742 350500 3748
rect 349080 480 349108 3470
rect 349172 3454 350304 3482
rect 350276 480 350304 3454
rect 351380 480 351408 9046
rect 351840 9042 351868 48758
rect 352116 48482 352144 52020
rect 353312 48822 353340 52020
rect 354508 49706 354536 52020
rect 355718 52006 356008 52034
rect 356914 52006 357388 52034
rect 358110 52006 358768 52034
rect 354496 49700 354548 49706
rect 354496 49642 354548 49648
rect 355324 49700 355376 49706
rect 355324 49642 355376 49648
rect 353300 48816 353352 48822
rect 353300 48758 353352 48764
rect 354588 48816 354640 48822
rect 354588 48758 354640 48764
rect 352104 48476 352156 48482
rect 352104 48418 352156 48424
rect 353208 48476 353260 48482
rect 353208 48418 353260 48424
rect 351920 46300 351972 46306
rect 351920 46242 351972 46248
rect 351828 9036 351880 9042
rect 351828 8978 351880 8984
rect 351932 3482 351960 46242
rect 353220 36718 353248 48418
rect 353208 36712 353260 36718
rect 353208 36654 353260 36660
rect 353760 7744 353812 7750
rect 353760 7686 353812 7692
rect 351932 3454 352604 3482
rect 352576 480 352604 3454
rect 353772 480 353800 7686
rect 354600 3398 354628 48758
rect 355336 10334 355364 49642
rect 355980 43518 356008 52006
rect 356060 44872 356112 44878
rect 356060 44814 356112 44820
rect 355968 43512 356020 43518
rect 355968 43454 356020 43460
rect 354680 10328 354732 10334
rect 354680 10270 354732 10276
rect 355324 10328 355376 10334
rect 355324 10270 355376 10276
rect 354588 3392 354640 3398
rect 354588 3334 354640 3340
rect 354692 610 354720 10270
rect 356072 626 356100 44814
rect 357256 4820 357308 4826
rect 357256 4762 357308 4768
rect 357268 3890 357296 4762
rect 357360 4078 357388 52006
rect 357440 11824 357492 11830
rect 357440 11766 357492 11772
rect 357348 4072 357400 4078
rect 357348 4014 357400 4020
rect 357268 3862 357388 3890
rect 354680 604 354732 610
rect 354680 546 354732 552
rect 354956 604 355008 610
rect 356072 598 356192 626
rect 354956 546 355008 552
rect 354968 480 354996 546
rect 356164 480 356192 598
rect 357360 480 357388 3862
rect 357452 610 357480 11766
rect 358740 5030 358768 52006
rect 359292 48822 359320 52020
rect 359280 48816 359332 48822
rect 359280 48758 359332 48764
rect 360108 48816 360160 48822
rect 360108 48758 360160 48764
rect 358820 36644 358872 36650
rect 358820 36586 358872 36592
rect 358728 5024 358780 5030
rect 358728 4966 358780 4972
rect 358832 610 358860 36586
rect 360120 25566 360148 48758
rect 360488 48754 360516 52020
rect 361684 48822 361712 52020
rect 362788 52006 362894 52034
rect 364090 52006 364288 52034
rect 361672 48816 361724 48822
rect 361672 48758 361724 48764
rect 360476 48748 360528 48754
rect 360476 48690 360528 48696
rect 361488 48748 361540 48754
rect 361488 48690 361540 48696
rect 360108 25560 360160 25566
rect 360108 25502 360160 25508
rect 360936 6316 360988 6322
rect 360936 6258 360988 6264
rect 357440 604 357492 610
rect 357440 546 357492 552
rect 358544 604 358596 610
rect 358544 546 358596 552
rect 358820 604 358872 610
rect 358820 546 358872 552
rect 359740 604 359792 610
rect 359740 546 359792 552
rect 358556 480 358584 546
rect 359752 480 359780 546
rect 360948 480 360976 6258
rect 361500 3942 361528 48690
rect 362788 24138 362816 52006
rect 362868 48816 362920 48822
rect 362868 48758 362920 48764
rect 362776 24132 362828 24138
rect 362776 24074 362828 24080
rect 361580 13116 361632 13122
rect 361580 13058 361632 13064
rect 361488 3936 361540 3942
rect 361488 3878 361540 3884
rect 361592 610 361620 13058
rect 362880 5302 362908 48758
rect 362960 43444 363012 43450
rect 362960 43386 363012 43392
rect 362868 5296 362920 5302
rect 362868 5238 362920 5244
rect 362972 626 363000 43386
rect 364260 3369 364288 52006
rect 365272 48686 365300 52020
rect 366482 52006 367048 52034
rect 365260 48680 365312 48686
rect 365260 48622 365312 48628
rect 367020 26926 367048 52006
rect 367664 49162 367692 52020
rect 367652 49156 367704 49162
rect 367652 49098 367704 49104
rect 367744 48680 367796 48686
rect 367744 48622 367796 48628
rect 367008 26920 367060 26926
rect 367008 26862 367060 26868
rect 365720 25628 365772 25634
rect 365720 25570 365772 25576
rect 364340 18624 364392 18630
rect 364340 18566 364392 18572
rect 364246 3360 364302 3369
rect 364352 3346 364380 18566
rect 364352 3318 364564 3346
rect 364246 3295 364302 3304
rect 361580 604 361632 610
rect 361580 546 361632 552
rect 362132 604 362184 610
rect 362972 598 363368 626
rect 362132 546 362184 552
rect 362144 480 362172 546
rect 363340 480 363368 598
rect 364536 480 364564 3318
rect 365732 3262 365760 25570
rect 367100 20052 367152 20058
rect 367100 19994 367152 20000
rect 365812 14544 365864 14550
rect 365812 14486 365864 14492
rect 365720 3256 365772 3262
rect 365720 3198 365772 3204
rect 365824 1442 365852 14486
rect 367112 3346 367140 19994
rect 367756 11830 367784 48622
rect 368860 48346 368888 52020
rect 369964 48822 369992 52020
rect 369952 48816 370004 48822
rect 369952 48758 370004 48764
rect 371056 48816 371108 48822
rect 371056 48758 371108 48764
rect 368848 48340 368900 48346
rect 368848 48282 368900 48288
rect 369768 48340 369820 48346
rect 369768 48282 369820 48288
rect 368480 24268 368532 24274
rect 368480 24210 368532 24216
rect 367744 11824 367796 11830
rect 367744 11766 367796 11772
rect 368492 3346 368520 24210
rect 369780 5030 369808 48282
rect 371068 28354 371096 48758
rect 371056 28348 371108 28354
rect 371056 28290 371108 28296
rect 369860 26988 369912 26994
rect 369860 26930 369912 26936
rect 369768 5024 369820 5030
rect 369768 4966 369820 4972
rect 367112 3318 368060 3346
rect 368492 3318 369256 3346
rect 366916 3256 366968 3262
rect 366916 3198 366968 3204
rect 365732 1414 365852 1442
rect 365732 480 365760 1414
rect 366928 480 366956 3198
rect 368032 480 368060 3318
rect 369228 480 369256 3318
rect 369872 2258 369900 26930
rect 371160 3641 371188 52020
rect 372370 52006 372568 52034
rect 373566 52006 373948 52034
rect 371608 8968 371660 8974
rect 371608 8910 371660 8916
rect 371146 3632 371202 3641
rect 371146 3567 371202 3576
rect 369872 2230 370452 2258
rect 370424 480 370452 2230
rect 371620 480 371648 8910
rect 372540 4826 372568 52006
rect 373920 29714 373948 52006
rect 374748 49094 374776 52020
rect 374736 49088 374788 49094
rect 374736 49030 374788 49036
rect 374644 49020 374696 49026
rect 374644 48962 374696 48968
rect 374092 37936 374144 37942
rect 374092 37878 374144 37884
rect 373908 29708 373960 29714
rect 373908 29650 373960 29656
rect 372620 28280 372672 28286
rect 372620 28222 372672 28228
rect 372528 4820 372580 4826
rect 372528 4762 372580 4768
rect 372632 3346 372660 28222
rect 372632 3318 372844 3346
rect 372816 480 372844 3318
rect 374104 1442 374132 37878
rect 374656 5574 374684 48962
rect 375944 48822 375972 52020
rect 375932 48816 375984 48822
rect 375932 48758 375984 48764
rect 376668 48816 376720 48822
rect 376668 48758 376720 48764
rect 375380 15972 375432 15978
rect 375380 15914 375432 15920
rect 374644 5568 374696 5574
rect 374644 5510 374696 5516
rect 375392 3346 375420 15914
rect 376680 13122 376708 48758
rect 377140 48346 377168 52020
rect 378336 48822 378364 52020
rect 379532 48822 379560 52020
rect 378324 48816 378376 48822
rect 378324 48758 378376 48764
rect 379428 48816 379480 48822
rect 379428 48758 379480 48764
rect 379520 48816 379572 48822
rect 379520 48758 379572 48764
rect 377128 48340 377180 48346
rect 377128 48282 377180 48288
rect 378048 48340 378100 48346
rect 378048 48282 378100 48288
rect 378060 31142 378088 48282
rect 378048 31136 378100 31142
rect 378048 31078 378100 31084
rect 376760 29640 376812 29646
rect 376760 29582 376812 29588
rect 376668 13116 376720 13122
rect 376668 13058 376720 13064
rect 376772 3346 376800 29582
rect 378784 3596 378836 3602
rect 378784 3538 378836 3544
rect 375196 3324 375248 3330
rect 375392 3318 376432 3346
rect 376772 3318 377628 3346
rect 375196 3266 375248 3272
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 3266
rect 376404 480 376432 3318
rect 377600 480 377628 3318
rect 378796 480 378824 3538
rect 379440 3262 379468 48758
rect 380728 37942 380756 52020
rect 381938 52006 382228 52034
rect 380808 48816 380860 48822
rect 380808 48758 380860 48764
rect 380716 37936 380768 37942
rect 380716 37878 380768 37884
rect 379980 5568 380032 5574
rect 379980 5510 380032 5516
rect 379428 3256 379480 3262
rect 379428 3198 379480 3204
rect 379992 480 380020 5510
rect 380820 5234 380848 48758
rect 380900 42084 380952 42090
rect 380900 42026 380952 42032
rect 380808 5228 380860 5234
rect 380808 5170 380860 5176
rect 380912 3346 380940 42026
rect 382200 3602 382228 52006
rect 383120 49706 383148 52020
rect 384330 52006 384988 52034
rect 383108 49700 383160 49706
rect 383108 49642 383160 49648
rect 384304 49700 384356 49706
rect 384304 49642 384356 49648
rect 383660 31068 383712 31074
rect 383660 31010 383712 31016
rect 382372 17264 382424 17270
rect 382372 17206 382424 17212
rect 382384 3670 382412 17206
rect 382280 3664 382332 3670
rect 382280 3606 382332 3612
rect 382372 3664 382424 3670
rect 382372 3606 382424 3612
rect 383568 3664 383620 3670
rect 383568 3606 383620 3612
rect 382188 3596 382240 3602
rect 382188 3538 382240 3544
rect 382292 3482 382320 3606
rect 382292 3454 382412 3482
rect 380912 3318 381216 3346
rect 381188 480 381216 3318
rect 382384 480 382412 3454
rect 383580 480 383608 3606
rect 383672 3346 383700 31010
rect 384316 14482 384344 49642
rect 384960 39438 384988 52006
rect 385512 48822 385540 52020
rect 386708 48822 386736 52020
rect 387904 48822 387932 52020
rect 389100 49026 389128 52020
rect 390310 52006 390508 52034
rect 391506 52006 391888 52034
rect 392702 52006 393268 52034
rect 393898 52006 394648 52034
rect 389088 49020 389140 49026
rect 389088 48962 389140 48968
rect 385500 48816 385552 48822
rect 385500 48758 385552 48764
rect 386328 48816 386380 48822
rect 386328 48758 386380 48764
rect 386696 48816 386748 48822
rect 386696 48758 386748 48764
rect 387708 48816 387760 48822
rect 387708 48758 387760 48764
rect 387892 48816 387944 48822
rect 387892 48758 387944 48764
rect 389088 48816 389140 48822
rect 389088 48758 389140 48764
rect 384948 39432 385000 39438
rect 384948 39374 385000 39380
rect 384304 14476 384356 14482
rect 384304 14418 384356 14424
rect 383672 3318 384712 3346
rect 386340 3330 386368 48758
rect 386420 18692 386472 18698
rect 386420 18634 386472 18640
rect 386432 3346 386460 18634
rect 387720 5098 387748 48758
rect 387800 39364 387852 39370
rect 387800 39306 387852 39312
rect 387708 5092 387760 5098
rect 387708 5034 387760 5040
rect 387812 3346 387840 39306
rect 389100 32502 389128 48758
rect 389088 32496 389140 32502
rect 389088 32438 389140 32444
rect 390480 4758 390508 52006
rect 390560 40792 390612 40798
rect 390560 40734 390612 40740
rect 390468 4752 390520 4758
rect 390468 4694 390520 4700
rect 389456 3732 389508 3738
rect 389456 3674 389508 3680
rect 384684 480 384712 3318
rect 386328 3324 386380 3330
rect 386432 3318 387104 3346
rect 387812 3318 388300 3346
rect 386328 3266 386380 3272
rect 385868 3188 385920 3194
rect 385868 3130 385920 3136
rect 385880 480 385908 3130
rect 387076 480 387104 3318
rect 388272 480 388300 3318
rect 389468 480 389496 3674
rect 390572 3670 390600 40734
rect 391860 40730 391888 52006
rect 391848 40724 391900 40730
rect 391848 40666 391900 40672
rect 390652 19984 390704 19990
rect 390652 19926 390704 19932
rect 390560 3664 390612 3670
rect 390560 3606 390612 3612
rect 390664 480 390692 19926
rect 393240 3874 393268 52006
rect 393320 21412 393372 21418
rect 393320 21354 393372 21360
rect 393044 3868 393096 3874
rect 393044 3810 393096 3816
rect 393228 3868 393280 3874
rect 393228 3810 393280 3816
rect 391848 3664 391900 3670
rect 391848 3606 391900 3612
rect 391860 480 391888 3606
rect 393056 480 393084 3810
rect 393332 3346 393360 21354
rect 394620 5166 394648 52006
rect 394988 48822 395016 52020
rect 396184 49298 396212 52020
rect 396172 49292 396224 49298
rect 396172 49234 396224 49240
rect 394976 48816 395028 48822
rect 394976 48758 395028 48764
rect 395988 48816 396040 48822
rect 395988 48758 396040 48764
rect 396000 35290 396028 48758
rect 395988 35284 396040 35290
rect 395988 35226 396040 35232
rect 394700 32428 394752 32434
rect 394700 32370 394752 32376
rect 394608 5160 394660 5166
rect 394608 5102 394660 5108
rect 394712 3346 394740 32370
rect 397380 15910 397408 52020
rect 398590 52006 398788 52034
rect 399786 52006 400168 52034
rect 397460 47592 397512 47598
rect 397460 47534 397512 47540
rect 397368 15904 397420 15910
rect 397368 15846 397420 15852
rect 396632 4140 396684 4146
rect 396632 4082 396684 4088
rect 393332 3318 394280 3346
rect 394712 3318 395476 3346
rect 394252 480 394280 3318
rect 395448 480 395476 3318
rect 396644 480 396672 4082
rect 397472 3346 397500 47534
rect 398760 36582 398788 52006
rect 398748 36576 398800 36582
rect 398748 36518 398800 36524
rect 398840 33856 398892 33862
rect 398840 33798 398892 33804
rect 398852 3346 398880 33798
rect 400140 3738 400168 52006
rect 400968 49706 400996 52020
rect 402178 52006 402928 52034
rect 400956 49700 401008 49706
rect 400956 49642 401008 49648
rect 402900 43450 402928 52006
rect 403360 49230 403388 52020
rect 403624 49700 403676 49706
rect 403624 49642 403676 49648
rect 403348 49224 403400 49230
rect 403348 49166 403400 49172
rect 402888 43444 402940 43450
rect 402888 43386 402940 43392
rect 401600 35216 401652 35222
rect 401600 35158 401652 35164
rect 401324 6180 401376 6186
rect 401324 6122 401376 6128
rect 400128 3732 400180 3738
rect 400128 3674 400180 3680
rect 400220 3460 400272 3466
rect 400220 3402 400272 3408
rect 397472 3318 397868 3346
rect 398852 3318 399064 3346
rect 397840 480 397868 3318
rect 399036 480 399064 3318
rect 400232 480 400260 3402
rect 401336 480 401364 6122
rect 401612 3346 401640 35158
rect 403636 17338 403664 49642
rect 404556 48822 404584 52020
rect 405766 52006 406056 52034
rect 406962 52006 407068 52034
rect 408158 52006 408448 52034
rect 409354 52006 409828 52034
rect 410550 52006 411208 52034
rect 404544 48816 404596 48822
rect 404544 48758 404596 48764
rect 405648 48816 405700 48822
rect 405648 48758 405700 48764
rect 405660 18630 405688 48758
rect 406028 46238 406056 52006
rect 405740 46232 405792 46238
rect 405740 46174 405792 46180
rect 406016 46232 406068 46238
rect 406016 46174 406068 46180
rect 405648 18624 405700 18630
rect 405648 18566 405700 18572
rect 403624 17332 403676 17338
rect 403624 17274 403676 17280
rect 404912 7608 404964 7614
rect 404912 7550 404964 7556
rect 403716 4004 403768 4010
rect 403716 3946 403768 3952
rect 401612 3318 402560 3346
rect 402532 480 402560 3318
rect 403728 480 403756 3946
rect 404924 480 404952 7550
rect 405752 3346 405780 46174
rect 407040 3505 407068 52006
rect 408420 19990 408448 52006
rect 408500 44940 408552 44946
rect 408500 44882 408552 44888
rect 408408 19984 408460 19990
rect 408408 19926 408460 19932
rect 408512 3670 408540 44882
rect 409800 33794 409828 52006
rect 409788 33788 409840 33794
rect 409788 33730 409840 33736
rect 408592 22772 408644 22778
rect 408592 22714 408644 22720
rect 408500 3664 408552 3670
rect 408500 3606 408552 3612
rect 407304 3528 407356 3534
rect 407026 3496 407082 3505
rect 408604 3482 408632 22714
rect 411180 3806 411208 52006
rect 411732 48482 411760 52020
rect 412928 48822 412956 52020
rect 414124 48822 414152 52020
rect 415228 52006 415334 52034
rect 416530 52006 416728 52034
rect 417726 52006 418108 52034
rect 418922 52006 419488 52034
rect 412916 48816 412968 48822
rect 412916 48758 412968 48764
rect 413928 48816 413980 48822
rect 413928 48758 413980 48764
rect 414112 48816 414164 48822
rect 414112 48758 414164 48764
rect 411720 48476 411772 48482
rect 411720 48418 411772 48424
rect 412548 48476 412600 48482
rect 412548 48418 412600 48424
rect 412560 21418 412588 48418
rect 413940 38010 413968 48758
rect 415228 44878 415256 52006
rect 415308 48816 415360 48822
rect 415308 48758 415360 48764
rect 415216 44872 415268 44878
rect 415216 44814 415268 44820
rect 413928 38004 413980 38010
rect 413928 37946 413980 37952
rect 412640 36712 412692 36718
rect 412640 36654 412692 36660
rect 412548 21412 412600 21418
rect 412548 21354 412600 21360
rect 412088 9036 412140 9042
rect 412088 8978 412140 8984
rect 410892 3800 410944 3806
rect 410892 3742 410944 3748
rect 411168 3800 411220 3806
rect 411168 3742 411220 3748
rect 409696 3664 409748 3670
rect 409696 3606 409748 3612
rect 407304 3470 407356 3476
rect 407026 3431 407082 3440
rect 405752 3318 406148 3346
rect 406120 480 406148 3318
rect 407316 480 407344 3470
rect 408512 3454 408632 3482
rect 408512 480 408540 3454
rect 409708 480 409736 3606
rect 410904 480 410932 3742
rect 412100 480 412128 8978
rect 412652 3346 412680 36654
rect 415320 3534 415348 48758
rect 416700 10334 416728 52006
rect 416872 43512 416924 43518
rect 416872 43454 416924 43460
rect 415400 10328 415452 10334
rect 415400 10270 415452 10276
rect 416688 10328 416740 10334
rect 416688 10270 416740 10276
rect 415308 3528 415360 3534
rect 415308 3470 415360 3476
rect 414480 3392 414532 3398
rect 412652 3318 413324 3346
rect 414480 3334 414532 3340
rect 413296 480 413324 3318
rect 414492 480 414520 3334
rect 415412 626 415440 10270
rect 415412 598 415716 626
rect 415688 480 415716 598
rect 416884 480 416912 43454
rect 417976 4072 418028 4078
rect 417976 4014 418028 4020
rect 417988 480 418016 4014
rect 418080 3670 418108 52006
rect 419460 42090 419488 52006
rect 420104 48822 420132 52020
rect 421208 48822 421236 52020
rect 422404 48822 422432 52020
rect 423508 52006 423614 52034
rect 424810 52006 425008 52034
rect 420092 48816 420144 48822
rect 420092 48758 420144 48764
rect 420828 48816 420880 48822
rect 420828 48758 420880 48764
rect 421196 48816 421248 48822
rect 421196 48758 421248 48764
rect 422208 48816 422260 48822
rect 422208 48758 422260 48764
rect 422392 48816 422444 48822
rect 422392 48758 422444 48764
rect 419448 42084 419500 42090
rect 419448 42026 419500 42032
rect 420840 39370 420868 48758
rect 420828 39364 420880 39370
rect 420828 39306 420880 39312
rect 419540 25560 419592 25566
rect 419540 25502 419592 25508
rect 419172 4956 419224 4962
rect 419172 4898 419224 4904
rect 418068 3664 418120 3670
rect 418068 3606 418120 3612
rect 419184 480 419212 4898
rect 419552 3346 419580 25502
rect 421564 3936 421616 3942
rect 421564 3878 421616 3884
rect 419552 3318 420408 3346
rect 420380 480 420408 3318
rect 421576 480 421604 3878
rect 422220 3466 422248 48758
rect 423508 22778 423536 52006
rect 423588 48816 423640 48822
rect 423588 48758 423640 48764
rect 423496 22772 423548 22778
rect 423496 22714 423548 22720
rect 423600 7682 423628 48758
rect 423680 24132 423732 24138
rect 423680 24074 423732 24080
rect 423588 7676 423640 7682
rect 423588 7618 423640 7624
rect 422760 5296 422812 5302
rect 422760 5238 422812 5244
rect 422208 3460 422260 3466
rect 422208 3402 422260 3408
rect 422772 480 422800 5238
rect 423692 3346 423720 24074
rect 424980 11762 425008 52006
rect 425992 47598 426020 52020
rect 427202 52006 427768 52034
rect 425980 47592 426032 47598
rect 425980 47534 426032 47540
rect 426440 26920 426492 26926
rect 426440 26862 426492 26868
rect 425060 11824 425112 11830
rect 425060 11766 425112 11772
rect 424968 11756 425020 11762
rect 424968 11698 425020 11704
rect 425072 3398 425100 11766
rect 425060 3392 425112 3398
rect 423692 3318 423996 3346
rect 426348 3392 426400 3398
rect 425060 3334 425112 3340
rect 425150 3360 425206 3369
rect 423968 480 423996 3318
rect 426348 3334 426400 3340
rect 426452 3346 426480 26862
rect 427740 24138 427768 52006
rect 428384 48822 428412 52020
rect 429580 48822 429608 52020
rect 430776 48822 430804 52020
rect 428372 48816 428424 48822
rect 428372 48758 428424 48764
rect 429108 48816 429160 48822
rect 429108 48758 429160 48764
rect 429568 48816 429620 48822
rect 429568 48758 429620 48764
rect 430488 48816 430540 48822
rect 430488 48758 430540 48764
rect 430764 48816 430816 48822
rect 430764 48758 430816 48764
rect 431868 48816 431920 48822
rect 431868 48758 431920 48764
rect 427912 48340 427964 48346
rect 427912 48282 427964 48288
rect 427924 38622 427952 48282
rect 427912 38616 427964 38622
rect 427912 38558 427964 38564
rect 427912 29028 427964 29034
rect 427912 28970 427964 28976
rect 427728 24132 427780 24138
rect 427728 24074 427780 24080
rect 427924 19310 427952 28970
rect 427912 19304 427964 19310
rect 427912 19246 427964 19252
rect 427912 9716 427964 9722
rect 427912 9658 427964 9664
rect 425150 3295 425206 3304
rect 425164 480 425192 3295
rect 426360 480 426388 3334
rect 426452 3318 427584 3346
rect 427556 480 427584 3318
rect 427924 2854 427952 9658
rect 429120 3942 429148 48758
rect 430500 6186 430528 48758
rect 430580 28348 430632 28354
rect 430580 28290 430632 28296
rect 430592 9654 430620 28290
rect 431880 25634 431908 48758
rect 431972 48754 432000 52020
rect 433168 48822 433196 52020
rect 434378 52006 434668 52034
rect 435574 52006 436048 52034
rect 433156 48816 433208 48822
rect 433156 48758 433208 48764
rect 433984 48816 434036 48822
rect 433984 48758 434036 48764
rect 431960 48748 432012 48754
rect 431960 48690 432012 48696
rect 433248 48748 433300 48754
rect 433248 48690 433300 48696
rect 431868 25628 431920 25634
rect 431868 25570 431920 25576
rect 430580 9648 430632 9654
rect 430580 9590 430632 9596
rect 430488 6180 430540 6186
rect 430488 6122 430540 6128
rect 429936 5024 429988 5030
rect 429936 4966 429988 4972
rect 429108 3936 429160 3942
rect 429108 3878 429160 3884
rect 427912 2848 427964 2854
rect 427912 2790 427964 2796
rect 428740 2780 428792 2786
rect 428740 2722 428792 2728
rect 428752 480 428780 2722
rect 429948 480 429976 4966
rect 433260 4146 433288 48690
rect 433340 29708 433392 29714
rect 433340 29650 433392 29656
rect 433352 7614 433380 29650
rect 433996 8974 434024 48758
rect 434640 26926 434668 52006
rect 434812 48340 434864 48346
rect 434812 48282 434864 48288
rect 434824 38622 434852 48282
rect 434812 38616 434864 38622
rect 434812 38558 434864 38564
rect 434812 29028 434864 29034
rect 434812 28970 434864 28976
rect 434628 26920 434680 26926
rect 434628 26862 434680 26868
rect 434824 19310 434852 28970
rect 434812 19304 434864 19310
rect 434812 19246 434864 19252
rect 434812 9716 434864 9722
rect 434812 9658 434864 9664
rect 433984 8968 434036 8974
rect 433984 8910 434036 8916
rect 433340 7608 433392 7614
rect 433340 7550 433392 7556
rect 434628 7608 434680 7614
rect 434628 7550 434680 7556
rect 433524 4820 433576 4826
rect 433524 4762 433576 4768
rect 433248 4140 433300 4146
rect 433248 4082 433300 4088
rect 432326 3632 432382 3641
rect 432326 3567 432382 3576
rect 431132 604 431184 610
rect 431132 546 431184 552
rect 431144 480 431172 546
rect 432340 480 432368 3567
rect 433536 480 433564 4762
rect 434640 480 434668 7550
rect 434824 2854 434852 9658
rect 436020 3194 436048 52006
rect 436756 48754 436784 52020
rect 437952 48822 437980 52020
rect 439148 48822 439176 52020
rect 440344 49706 440372 52020
rect 440332 49700 440384 49706
rect 440332 49642 440384 49648
rect 437940 48816 437992 48822
rect 437940 48758 437992 48764
rect 438768 48816 438820 48822
rect 438768 48758 438820 48764
rect 439136 48816 439188 48822
rect 439136 48758 439188 48764
rect 440148 48816 440200 48822
rect 440148 48758 440200 48764
rect 436744 48748 436796 48754
rect 436744 48690 436796 48696
rect 438124 48748 438176 48754
rect 438124 48690 438176 48696
rect 437480 31136 437532 31142
rect 437480 31078 437532 31084
rect 436100 13116 436152 13122
rect 436100 13058 436152 13064
rect 436112 9654 436140 13058
rect 436100 9648 436152 9654
rect 436100 9590 436152 9596
rect 437492 3346 437520 31078
rect 438136 10402 438164 48690
rect 438780 29646 438808 48758
rect 438768 29640 438820 29646
rect 438768 29582 438820 29588
rect 438124 10396 438176 10402
rect 438124 10338 438176 10344
rect 437492 3318 438256 3346
rect 436008 3188 436060 3194
rect 436008 3130 436060 3136
rect 434812 2848 434864 2854
rect 434812 2790 434864 2796
rect 435824 2780 435876 2786
rect 435824 2722 435876 2728
rect 435836 480 435864 2722
rect 437020 604 437072 610
rect 437020 546 437072 552
rect 437032 480 437060 546
rect 438228 480 438256 3318
rect 440160 3262 440188 48758
rect 441540 33862 441568 52020
rect 442750 52006 442948 52034
rect 442264 49700 442316 49706
rect 442264 49642 442316 49648
rect 441620 37936 441672 37942
rect 441620 37878 441672 37884
rect 441528 33856 441580 33862
rect 441528 33798 441580 33804
rect 440608 5228 440660 5234
rect 440608 5170 440660 5176
rect 439412 3256 439464 3262
rect 439412 3198 439464 3204
rect 440148 3256 440200 3262
rect 440148 3198 440200 3204
rect 439424 480 439452 3198
rect 440620 480 440648 5170
rect 441632 3346 441660 37878
rect 442276 11830 442304 49642
rect 442264 11824 442316 11830
rect 442264 11766 442316 11772
rect 442920 4010 442948 52006
rect 443932 46306 443960 52020
rect 445142 52006 445708 52034
rect 443920 46300 443972 46306
rect 443920 46242 443972 46248
rect 444380 39432 444432 39438
rect 444380 39374 444432 39380
rect 443092 14476 443144 14482
rect 443092 14418 443144 14424
rect 442908 4004 442960 4010
rect 442908 3946 442960 3952
rect 443000 3596 443052 3602
rect 443000 3538 443052 3544
rect 441632 3318 441844 3346
rect 441816 480 441844 3318
rect 443012 480 443040 3538
rect 443104 3346 443132 14418
rect 444392 3346 444420 39374
rect 445680 28286 445708 52006
rect 446232 48822 446260 52020
rect 447428 48822 447456 52020
rect 448624 48822 448652 52020
rect 446220 48816 446272 48822
rect 446220 48758 446272 48764
rect 447048 48816 447100 48822
rect 447048 48758 447100 48764
rect 447416 48816 447468 48822
rect 447416 48758 447468 48764
rect 448428 48816 448480 48822
rect 448428 48758 448480 48764
rect 448612 48816 448664 48822
rect 448612 48758 448664 48764
rect 449716 48816 449768 48822
rect 449716 48758 449768 48764
rect 445668 28280 445720 28286
rect 445668 28222 445720 28228
rect 443104 3318 444236 3346
rect 444392 3318 445432 3346
rect 444208 480 444236 3318
rect 445404 480 445432 3318
rect 446588 3324 446640 3330
rect 446588 3266 446640 3272
rect 446600 480 446628 3266
rect 447060 3126 447088 48758
rect 448440 13122 448468 48758
rect 448520 32496 448572 32502
rect 448520 32438 448572 32444
rect 448428 13116 448480 13122
rect 448428 13058 448480 13064
rect 447784 5092 447836 5098
rect 447784 5034 447836 5040
rect 447048 3120 447100 3126
rect 447048 3062 447100 3068
rect 447796 480 447824 5034
rect 448532 3346 448560 32438
rect 449728 31074 449756 48758
rect 449716 31068 449768 31074
rect 449716 31010 449768 31016
rect 449820 3369 449848 52020
rect 451016 49094 451044 52020
rect 452226 52006 452608 52034
rect 453422 52006 453988 52034
rect 454618 52006 455368 52034
rect 451004 49088 451056 49094
rect 451004 49030 451056 49036
rect 451924 49088 451976 49094
rect 451924 49030 451976 49036
rect 449900 49020 449952 49026
rect 449900 48962 449952 48968
rect 449806 3360 449862 3369
rect 448532 3318 449020 3346
rect 448992 480 449020 3318
rect 449912 3346 449940 48962
rect 451280 40724 451332 40730
rect 451280 40666 451332 40672
rect 451292 3602 451320 40666
rect 451936 14482 451964 49030
rect 451924 14476 451976 14482
rect 451924 14418 451976 14424
rect 452580 7614 452608 52006
rect 452568 7608 452620 7614
rect 452568 7550 452620 7556
rect 453672 3868 453724 3874
rect 453672 3810 453724 3816
rect 451280 3596 451332 3602
rect 451280 3538 451332 3544
rect 452476 3596 452528 3602
rect 452476 3538 452528 3544
rect 449912 3318 450216 3346
rect 449806 3295 449862 3304
rect 450188 480 450216 3318
rect 451280 2984 451332 2990
rect 451280 2926 451332 2932
rect 451292 480 451320 2926
rect 452488 480 452516 3538
rect 453684 480 453712 3810
rect 453960 3398 453988 52006
rect 454868 5160 454920 5166
rect 454868 5102 454920 5108
rect 453948 3392 454000 3398
rect 453948 3334 454000 3340
rect 454880 480 454908 5102
rect 455340 4962 455368 52006
rect 455800 48822 455828 52020
rect 456892 49292 456944 49298
rect 456892 49234 456944 49240
rect 455788 48816 455840 48822
rect 455788 48758 455840 48764
rect 456708 48816 456760 48822
rect 456708 48758 456760 48764
rect 455420 35284 455472 35290
rect 455420 35226 455472 35232
rect 455328 4956 455380 4962
rect 455328 4898 455380 4904
rect 455432 626 455460 35226
rect 456720 17270 456748 48758
rect 456708 17264 456760 17270
rect 456708 17206 456760 17212
rect 456904 626 456932 49234
rect 456996 48822 457024 52020
rect 456984 48816 457036 48822
rect 456984 48758 457036 48764
rect 458088 48816 458140 48822
rect 458088 48758 458140 48764
rect 458100 3330 458128 48758
rect 458192 48754 458220 52020
rect 459388 48822 459416 52020
rect 460598 52006 460888 52034
rect 461794 52006 462268 52034
rect 462990 52006 463648 52034
rect 459376 48816 459428 48822
rect 459376 48758 459428 48764
rect 460204 48816 460256 48822
rect 460204 48758 460256 48764
rect 458180 48748 458232 48754
rect 458180 48690 458232 48696
rect 459468 48748 459520 48754
rect 459468 48690 459520 48696
rect 458180 15904 458232 15910
rect 458180 15846 458232 15852
rect 458088 3324 458140 3330
rect 458088 3266 458140 3272
rect 458192 626 458220 15846
rect 459480 4894 459508 48690
rect 459652 36576 459704 36582
rect 459652 36518 459704 36524
rect 459468 4888 459520 4894
rect 459468 4830 459520 4836
rect 455432 598 456012 626
rect 456904 598 457208 626
rect 458192 598 458404 626
rect 455984 592 456012 598
rect 457180 592 457208 598
rect 458376 592 458404 598
rect 455984 564 456104 592
rect 457180 564 457300 592
rect 458376 564 458496 592
rect 456076 480 456104 564
rect 457272 480 457300 564
rect 458468 480 458496 564
rect 459664 480 459692 36518
rect 460216 35222 460244 48758
rect 460204 35216 460256 35222
rect 460204 35158 460256 35164
rect 460860 3856 460888 52006
rect 460940 17332 460992 17338
rect 460940 17274 460992 17280
rect 460952 4026 460980 17274
rect 462240 5234 462268 52006
rect 462320 43444 462372 43450
rect 462320 43386 462372 43392
rect 462228 5228 462280 5234
rect 462228 5170 462280 5176
rect 460952 3998 461072 4026
rect 460860 3828 460980 3856
rect 460952 3738 460980 3828
rect 460848 3732 460900 3738
rect 460848 3674 460900 3680
rect 460940 3732 460992 3738
rect 460940 3674 460992 3680
rect 460860 480 460888 3674
rect 461044 610 461072 3998
rect 462332 610 462360 43386
rect 463620 5302 463648 52006
rect 463792 49224 463844 49230
rect 463792 49166 463844 49172
rect 463608 5296 463660 5302
rect 463608 5238 463660 5244
rect 463804 610 463832 49166
rect 464172 48822 464200 52020
rect 465368 48822 465396 52020
rect 466564 48822 466592 52020
rect 467760 49026 467788 52020
rect 468970 52006 469168 52034
rect 470166 52006 470548 52034
rect 471362 52006 471928 52034
rect 467748 49020 467800 49026
rect 467748 48962 467800 48968
rect 464160 48816 464212 48822
rect 464160 48758 464212 48764
rect 464988 48816 465040 48822
rect 464988 48758 465040 48764
rect 465356 48816 465408 48822
rect 465356 48758 465408 48764
rect 466368 48816 466420 48822
rect 466368 48758 466420 48764
rect 466552 48816 466604 48822
rect 466552 48758 466604 48764
rect 467748 48816 467800 48822
rect 467748 48758 467800 48764
rect 465000 4078 465028 48758
rect 465080 18624 465132 18630
rect 465080 18566 465132 18572
rect 464988 4072 465040 4078
rect 464988 4014 465040 4020
rect 465092 610 465120 18566
rect 466380 5030 466408 48758
rect 466460 46232 466512 46238
rect 466460 46174 466512 46180
rect 466368 5024 466420 5030
rect 466368 4966 466420 4972
rect 466472 610 466500 46174
rect 467760 32434 467788 48758
rect 467748 32428 467800 32434
rect 467748 32370 467800 32376
rect 467840 19984 467892 19990
rect 467840 19926 467892 19932
rect 467852 3602 467880 19926
rect 469140 15910 469168 52006
rect 469220 33788 469272 33794
rect 469220 33730 469272 33736
rect 469128 15904 469180 15910
rect 469128 15846 469180 15852
rect 467840 3596 467892 3602
rect 467840 3538 467892 3544
rect 469128 3596 469180 3602
rect 469128 3538 469180 3544
rect 467930 3496 467986 3505
rect 467930 3431 467986 3440
rect 461032 604 461084 610
rect 461032 546 461084 552
rect 462044 604 462096 610
rect 462044 546 462096 552
rect 462320 604 462372 610
rect 462320 546 462372 552
rect 463240 604 463292 610
rect 463240 546 463292 552
rect 463792 604 463844 610
rect 463792 546 463844 552
rect 464436 604 464488 610
rect 464436 546 464488 552
rect 465080 604 465132 610
rect 465080 546 465132 552
rect 465632 604 465684 610
rect 465632 546 465684 552
rect 466460 604 466512 610
rect 466460 546 466512 552
rect 466828 604 466880 610
rect 466828 546 466880 552
rect 462056 480 462084 546
rect 463252 480 463280 546
rect 464448 480 464476 546
rect 465644 480 465672 546
rect 466840 480 466868 546
rect 467944 480 467972 3431
rect 469140 480 469168 3538
rect 469232 610 469260 33730
rect 470520 19990 470548 52006
rect 470508 19984 470560 19990
rect 470508 19926 470560 19932
rect 471520 3800 471572 3806
rect 471520 3742 471572 3748
rect 469220 604 469272 610
rect 469220 546 469272 552
rect 470324 604 470376 610
rect 470324 546 470376 552
rect 470336 480 470364 546
rect 471532 480 471560 3742
rect 471900 3602 471928 52006
rect 472452 48754 472480 52020
rect 473648 48822 473676 52020
rect 474844 49162 474872 52020
rect 474832 49156 474884 49162
rect 474832 49098 474884 49104
rect 473636 48816 473688 48822
rect 473636 48758 473688 48764
rect 474648 48816 474700 48822
rect 474648 48758 474700 48764
rect 472440 48748 472492 48754
rect 472440 48690 472492 48696
rect 474004 48748 474056 48754
rect 474004 48690 474056 48696
rect 473360 38004 473412 38010
rect 473360 37946 473412 37952
rect 471980 21412 472032 21418
rect 471980 21354 472032 21360
rect 471888 3596 471940 3602
rect 471888 3538 471940 3544
rect 471992 3346 472020 21354
rect 473372 3346 473400 37946
rect 474016 18630 474044 48690
rect 474660 21418 474688 48758
rect 474648 21412 474700 21418
rect 474648 21354 474700 21360
rect 474004 18624 474056 18630
rect 474004 18566 474056 18572
rect 476040 4826 476068 52020
rect 477236 49706 477264 52020
rect 478446 52006 478828 52034
rect 479642 52006 480208 52034
rect 477224 49700 477276 49706
rect 477224 49642 477276 49648
rect 476120 44872 476172 44878
rect 476120 44814 476172 44820
rect 476028 4820 476080 4826
rect 476028 4762 476080 4768
rect 475108 3528 475160 3534
rect 475108 3470 475160 3476
rect 471992 3318 472756 3346
rect 473372 3318 473952 3346
rect 472728 480 472756 3318
rect 473924 480 473952 3318
rect 475120 480 475148 3470
rect 476132 3346 476160 44814
rect 477592 10328 477644 10334
rect 477592 10270 477644 10276
rect 477604 3482 477632 10270
rect 478800 3806 478828 52006
rect 480180 44878 480208 52006
rect 480824 48822 480852 52020
rect 482020 49094 482048 52020
rect 482284 49700 482336 49706
rect 482284 49642 482336 49648
rect 482008 49088 482060 49094
rect 482008 49030 482060 49036
rect 480812 48816 480864 48822
rect 480812 48758 480864 48764
rect 481548 48816 481600 48822
rect 481548 48758 481600 48764
rect 480168 44872 480220 44878
rect 480168 44814 480220 44820
rect 478880 42084 478932 42090
rect 478880 42026 478932 42032
rect 478788 3800 478840 3806
rect 478788 3742 478840 3748
rect 478696 3664 478748 3670
rect 478696 3606 478748 3612
rect 477512 3454 477632 3482
rect 476132 3318 476344 3346
rect 476316 480 476344 3318
rect 477512 480 477540 3454
rect 478708 480 478736 3606
rect 478892 3346 478920 42026
rect 480260 39364 480312 39370
rect 480260 39306 480312 39312
rect 480272 3346 480300 39306
rect 481560 24206 481588 48758
rect 481548 24200 481600 24206
rect 481548 24142 481600 24148
rect 482296 22846 482324 49642
rect 483216 48822 483244 52020
rect 484412 48822 484440 52020
rect 485622 52006 485728 52034
rect 486818 52006 487108 52034
rect 483204 48816 483256 48822
rect 483204 48758 483256 48764
rect 484308 48816 484360 48822
rect 484308 48758 484360 48764
rect 484400 48816 484452 48822
rect 484400 48758 484452 48764
rect 485596 48816 485648 48822
rect 485596 48758 485648 48764
rect 482284 22840 482336 22846
rect 482284 22782 482336 22788
rect 483480 7676 483532 7682
rect 483480 7618 483532 7624
rect 482284 3460 482336 3466
rect 482284 3402 482336 3408
rect 478892 3318 479932 3346
rect 480272 3318 481128 3346
rect 479904 480 479932 3318
rect 481100 480 481128 3318
rect 482296 480 482324 3402
rect 483492 480 483520 7618
rect 484320 5098 484348 48758
rect 485608 25566 485636 48758
rect 485596 25560 485648 25566
rect 485596 25502 485648 25508
rect 484400 22772 484452 22778
rect 484400 22714 484452 22720
rect 484308 5092 484360 5098
rect 484308 5034 484360 5040
rect 484412 3346 484440 22714
rect 485700 3505 485728 52006
rect 485780 47592 485832 47598
rect 485780 47534 485832 47540
rect 485792 3670 485820 47534
rect 485872 11756 485924 11762
rect 485872 11698 485924 11704
rect 485780 3664 485832 3670
rect 485780 3606 485832 3612
rect 485686 3496 485742 3505
rect 485884 3482 485912 11698
rect 487080 5166 487108 52006
rect 488000 48754 488028 52020
rect 489196 49230 489224 52020
rect 489184 49224 489236 49230
rect 489184 49166 489236 49172
rect 487988 48748 488040 48754
rect 487988 48690 488040 48696
rect 489184 48748 489236 48754
rect 489184 48690 489236 48696
rect 487160 24132 487212 24138
rect 487160 24074 487212 24080
rect 487068 5160 487120 5166
rect 487068 5102 487120 5108
rect 486976 3664 487028 3670
rect 486976 3606 487028 3612
rect 485686 3431 485742 3440
rect 485792 3454 485912 3482
rect 484412 3318 484624 3346
rect 484596 480 484624 3318
rect 485792 480 485820 3454
rect 486988 480 487016 3606
rect 487172 3346 487200 24074
rect 489196 9042 489224 48690
rect 490392 47598 490420 52020
rect 491588 48822 491616 52020
rect 492784 48822 492812 52020
rect 493888 52006 493994 52034
rect 491576 48816 491628 48822
rect 491576 48758 491628 48764
rect 492588 48816 492640 48822
rect 492588 48758 492640 48764
rect 492772 48816 492824 48822
rect 492772 48758 492824 48764
rect 490380 47592 490432 47598
rect 490380 47534 490432 47540
rect 492600 26994 492628 48758
rect 493888 43450 493916 52006
rect 495176 48822 495204 52020
rect 496386 52006 496768 52034
rect 497490 52006 498148 52034
rect 493968 48816 494020 48822
rect 493968 48758 494020 48764
rect 495164 48816 495216 48822
rect 495164 48758 495216 48764
rect 496084 48816 496136 48822
rect 496084 48758 496136 48764
rect 493876 43444 493928 43450
rect 493876 43386 493928 43392
rect 492588 26988 492640 26994
rect 492588 26930 492640 26936
rect 491300 25628 491352 25634
rect 491300 25570 491352 25576
rect 489184 9036 489236 9042
rect 489184 8978 489236 8984
rect 490564 6180 490616 6186
rect 490564 6122 490616 6128
rect 489368 3936 489420 3942
rect 489368 3878 489420 3884
rect 487172 3318 488212 3346
rect 488184 480 488212 3318
rect 489380 480 489408 3878
rect 490576 480 490604 6122
rect 491312 3482 491340 25570
rect 492956 4140 493008 4146
rect 492956 4082 493008 4088
rect 491312 3454 491800 3482
rect 491772 480 491800 3454
rect 492968 480 492996 4082
rect 493980 3874 494008 48758
rect 494060 26920 494112 26926
rect 494060 26862 494112 26868
rect 493968 3868 494020 3874
rect 493968 3810 494020 3816
rect 494072 3534 494100 26862
rect 496096 10334 496124 48758
rect 496084 10328 496136 10334
rect 496084 10270 496136 10276
rect 494152 8968 494204 8974
rect 494152 8910 494204 8916
rect 494060 3528 494112 3534
rect 494060 3470 494112 3476
rect 494164 480 494192 8910
rect 496740 4146 496768 52006
rect 498120 42090 498148 52006
rect 498672 48822 498700 52020
rect 499868 48822 499896 52020
rect 501064 48822 501092 52020
rect 502168 52006 502274 52034
rect 503470 52006 503668 52034
rect 498660 48816 498712 48822
rect 498660 48758 498712 48764
rect 499488 48816 499540 48822
rect 499488 48758 499540 48764
rect 499856 48816 499908 48822
rect 499856 48758 499908 48764
rect 500868 48816 500920 48822
rect 500868 48758 500920 48764
rect 501052 48816 501104 48822
rect 501052 48758 501104 48764
rect 498108 42084 498160 42090
rect 498108 42026 498160 42032
rect 498200 29640 498252 29646
rect 498200 29582 498252 29588
rect 496820 10396 496872 10402
rect 496820 10338 496872 10344
rect 496728 4140 496780 4146
rect 496728 4082 496780 4088
rect 495348 3528 495400 3534
rect 495348 3470 495400 3476
rect 496832 3482 496860 10338
rect 498212 3482 498240 29582
rect 499500 11762 499528 48758
rect 499488 11756 499540 11762
rect 499488 11698 499540 11704
rect 500880 3942 500908 48758
rect 502168 33794 502196 52006
rect 502248 48816 502300 48822
rect 502248 48758 502300 48764
rect 502156 33788 502208 33794
rect 502156 33730 502208 33736
rect 500960 11824 501012 11830
rect 500960 11766 501012 11772
rect 500868 3936 500920 3942
rect 500868 3878 500920 3884
rect 495360 480 495388 3470
rect 496832 3454 497780 3482
rect 498212 3454 498976 3482
rect 496544 3188 496596 3194
rect 496544 3130 496596 3136
rect 496556 480 496584 3130
rect 497752 480 497780 3454
rect 498948 480 498976 3454
rect 500972 3346 501000 11766
rect 502260 6186 502288 48758
rect 502432 33856 502484 33862
rect 502432 33798 502484 33804
rect 502248 6180 502300 6186
rect 502248 6122 502300 6128
rect 500972 3318 501276 3346
rect 500132 3256 500184 3262
rect 500132 3198 500184 3204
rect 500144 480 500172 3198
rect 501248 480 501276 3318
rect 502444 480 502472 33798
rect 503640 6882 503668 52006
rect 503720 46300 503772 46306
rect 503720 46242 503772 46248
rect 503456 6854 503668 6882
rect 503456 3670 503484 6854
rect 503628 4004 503680 4010
rect 503628 3946 503680 3952
rect 503444 3664 503496 3670
rect 503444 3606 503496 3612
rect 503640 480 503668 3946
rect 503732 3346 503760 46242
rect 504652 46238 504680 52020
rect 505862 52006 506428 52034
rect 507058 52006 507808 52034
rect 504640 46232 504692 46238
rect 504640 46174 504692 46180
rect 505100 28280 505152 28286
rect 505100 28222 505152 28228
rect 505112 3346 505140 28222
rect 506400 13190 506428 52006
rect 506388 13184 506440 13190
rect 506388 13126 506440 13132
rect 507780 3534 507808 52006
rect 508240 48822 508268 52020
rect 509436 48822 509464 52020
rect 508228 48816 508280 48822
rect 508228 48758 508280 48764
rect 509148 48816 509200 48822
rect 509148 48758 509200 48764
rect 509424 48816 509476 48822
rect 509424 48758 509476 48764
rect 510528 48816 510580 48822
rect 510528 48758 510580 48764
rect 509160 39370 509188 48758
rect 509148 39364 509200 39370
rect 509148 39306 509200 39312
rect 510540 31074 510568 48758
rect 510632 48550 510660 52020
rect 510620 48544 510672 48550
rect 510620 48486 510672 48492
rect 511828 37942 511856 52020
rect 513038 52006 513328 52034
rect 514234 52006 514708 52034
rect 515430 52006 516088 52034
rect 511908 48544 511960 48550
rect 511908 48486 511960 48492
rect 511816 37936 511868 37942
rect 511816 37878 511868 37884
rect 509240 31068 509292 31074
rect 509240 31010 509292 31016
rect 510528 31068 510580 31074
rect 510528 31010 510580 31016
rect 507860 13116 507912 13122
rect 507860 13058 507912 13064
rect 507768 3528 507820 3534
rect 507768 3470 507820 3476
rect 507872 3346 507900 13058
rect 509252 3346 509280 31010
rect 510802 3360 510858 3369
rect 503732 3318 504864 3346
rect 505112 3318 506060 3346
rect 507872 3318 508452 3346
rect 509252 3318 509648 3346
rect 504836 480 504864 3318
rect 506032 480 506060 3318
rect 507216 3120 507268 3126
rect 507216 3062 507268 3068
rect 507228 480 507256 3062
rect 508424 480 508452 3318
rect 509620 480 509648 3318
rect 510802 3295 510858 3304
rect 510816 480 510844 3295
rect 511920 3262 511948 48486
rect 512000 14476 512052 14482
rect 512000 14418 512052 14424
rect 511908 3256 511960 3262
rect 511908 3198 511960 3204
rect 512012 480 512040 14418
rect 513196 7608 513248 7614
rect 513196 7550 513248 7556
rect 513208 480 513236 7550
rect 513300 3194 513328 52006
rect 514680 4010 514708 52006
rect 516060 36582 516088 52006
rect 516612 48822 516640 52020
rect 517808 48822 517836 52020
rect 519004 48822 519032 52020
rect 516600 48816 516652 48822
rect 516600 48758 516652 48764
rect 517428 48816 517480 48822
rect 517428 48758 517480 48764
rect 517796 48816 517848 48822
rect 517796 48758 517848 48764
rect 518808 48816 518860 48822
rect 518808 48758 518860 48764
rect 518992 48816 519044 48822
rect 518992 48758 519044 48764
rect 520096 48816 520148 48822
rect 520096 48758 520148 48764
rect 516048 36576 516100 36582
rect 516048 36518 516100 36524
rect 516140 17264 516192 17270
rect 516140 17206 516192 17212
rect 515588 4956 515640 4962
rect 515588 4898 515640 4904
rect 514668 4004 514720 4010
rect 514668 3946 514720 3952
rect 514392 3392 514444 3398
rect 514392 3334 514444 3340
rect 513288 3188 513340 3194
rect 513288 3130 513340 3136
rect 514404 480 514432 3334
rect 515600 480 515628 4898
rect 516152 3346 516180 17206
rect 517440 3398 517468 48758
rect 518820 3466 518848 48758
rect 520108 7614 520136 48758
rect 520096 7608 520148 7614
rect 520096 7550 520148 7556
rect 519084 4888 519136 4894
rect 519084 4830 519136 4836
rect 518808 3460 518860 3466
rect 518808 3402 518860 3408
rect 517428 3392 517480 3398
rect 516152 3318 516824 3346
rect 517428 3334 517480 3340
rect 516796 480 516824 3318
rect 517888 3324 517940 3330
rect 517888 3266 517940 3272
rect 517900 480 517928 3266
rect 519096 480 519124 4830
rect 520200 3369 520228 52020
rect 521410 52006 521608 52034
rect 520372 35216 520424 35222
rect 520372 35158 520424 35164
rect 520384 3482 520412 35158
rect 521580 3738 521608 52006
rect 523696 41410 523724 85303
rect 523788 77246 523816 111959
rect 523880 111790 523908 138615
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 523868 111784 523920 111790
rect 523868 111726 523920 111732
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 523866 98696 523922 98705
rect 523866 98631 523922 98640
rect 523776 77240 523828 77246
rect 523776 77182 523828 77188
rect 523774 72040 523830 72049
rect 523774 71975 523830 71984
rect 523684 41404 523736 41410
rect 523684 41346 523736 41352
rect 523788 30326 523816 71975
rect 523880 64870 523908 98631
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 523868 64864 523920 64870
rect 523868 64806 523920 64812
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 523866 58712 523922 58721
rect 523866 58647 523922 58656
rect 523776 30320 523828 30326
rect 523776 30262 523828 30268
rect 523880 17950 523908 58647
rect 549260 49224 549312 49230
rect 549260 49166 549312 49172
rect 535460 49156 535512 49162
rect 535460 49098 535512 49104
rect 528560 49020 528612 49026
rect 528560 48962 528612 48968
rect 527180 32428 527232 32434
rect 527180 32370 527232 32376
rect 523868 17944 523920 17950
rect 523868 17886 523920 17892
rect 523868 5296 523920 5302
rect 523868 5238 523920 5244
rect 522672 5228 522724 5234
rect 522672 5170 522724 5176
rect 521476 3732 521528 3738
rect 521476 3674 521528 3680
rect 521568 3732 521620 3738
rect 521568 3674 521620 3680
rect 520292 3454 520412 3482
rect 520186 3360 520242 3369
rect 520186 3295 520242 3304
rect 520292 480 520320 3454
rect 521488 480 521516 3674
rect 522684 480 522712 5170
rect 523880 480 523908 5238
rect 526260 5024 526312 5030
rect 526260 4966 526312 4972
rect 525064 4072 525116 4078
rect 525064 4014 525116 4020
rect 525076 480 525104 4014
rect 526272 480 526300 4966
rect 527192 3346 527220 32370
rect 528572 3482 528600 48962
rect 534080 21412 534132 21418
rect 534080 21354 534132 21360
rect 529940 19984 529992 19990
rect 529940 19926 529992 19932
rect 528652 15904 528704 15910
rect 528652 15846 528704 15852
rect 528664 3602 528692 15846
rect 528652 3596 528704 3602
rect 528652 3538 528704 3544
rect 529848 3596 529900 3602
rect 529848 3538 529900 3544
rect 528572 3454 528692 3482
rect 527192 3318 527496 3346
rect 527468 480 527496 3318
rect 528664 480 528692 3454
rect 529860 480 529888 3538
rect 529952 3482 529980 19926
rect 532700 18624 532752 18630
rect 532700 18566 532752 18572
rect 532712 3482 532740 18566
rect 534092 3482 534120 21354
rect 535472 3482 535500 49098
rect 542360 49088 542412 49094
rect 542360 49030 542412 49036
rect 539600 44872 539652 44878
rect 539600 44814 539652 44820
rect 536840 22840 536892 22846
rect 536840 22782 536892 22788
rect 536852 3602 536880 22782
rect 536932 4820 536984 4826
rect 536932 4762 536984 4768
rect 536840 3596 536892 3602
rect 536840 3538 536892 3544
rect 529952 3454 531084 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 531056 480 531084 3454
rect 532240 3324 532292 3330
rect 532240 3266 532292 3272
rect 532252 480 532280 3266
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 4762
rect 539324 3800 539376 3806
rect 539324 3742 539376 3748
rect 538128 3596 538180 3602
rect 538128 3538 538180 3544
rect 538140 480 538168 3538
rect 539336 480 539364 3742
rect 539612 3482 539640 44814
rect 540980 24200 541032 24206
rect 540980 24142 541032 24148
rect 540992 3482 541020 24142
rect 542372 3482 542400 49030
rect 545120 25560 545172 25566
rect 545120 25502 545172 25508
rect 544108 5092 544160 5098
rect 544108 5034 544160 5040
rect 539612 3454 540560 3482
rect 540992 3454 541756 3482
rect 542372 3454 542952 3482
rect 540532 480 540560 3454
rect 541728 480 541756 3454
rect 542924 480 542952 3454
rect 544120 480 544148 5034
rect 545132 3482 545160 25502
rect 548892 9036 548944 9042
rect 548892 8978 548944 8984
rect 547696 5160 547748 5166
rect 547696 5102 547748 5108
rect 546498 3496 546554 3505
rect 545132 3454 545344 3482
rect 545316 480 545344 3454
rect 546498 3431 546554 3440
rect 546512 480 546540 3431
rect 547708 480 547736 5102
rect 548904 480 548932 8978
rect 549272 3482 549300 49166
rect 550640 47592 550692 47598
rect 550640 47534 550692 47540
rect 550652 3482 550680 47534
rect 564440 46232 564492 46238
rect 564440 46174 564492 46180
rect 554780 43444 554832 43450
rect 554780 43386 554832 43392
rect 552020 26988 552072 26994
rect 552020 26930 552072 26936
rect 552032 3482 552060 26930
rect 553584 3868 553636 3874
rect 553584 3810 553636 3816
rect 549272 3454 550128 3482
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 550100 480 550128 3454
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3810
rect 554792 480 554820 43386
rect 557540 42084 557592 42090
rect 557540 42026 557592 42032
rect 554872 10328 554924 10334
rect 554872 10270 554924 10276
rect 554884 3482 554912 10270
rect 557172 4140 557224 4146
rect 557172 4082 557224 4088
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 4082
rect 557552 3482 557580 42026
rect 563152 33788 563204 33794
rect 563152 33730 563204 33736
rect 558920 11756 558972 11762
rect 558920 11698 558972 11704
rect 558932 3482 558960 11698
rect 561956 6180 562008 6186
rect 561956 6122 562008 6128
rect 560760 3936 560812 3942
rect 560760 3878 560812 3884
rect 557552 3454 558408 3482
rect 558932 3454 559604 3482
rect 558380 480 558408 3454
rect 559576 480 559604 3454
rect 560772 480 560800 3878
rect 561968 480 561996 6122
rect 563164 480 563192 33730
rect 564348 3664 564400 3670
rect 564348 3606 564400 3612
rect 564360 480 564388 3606
rect 564452 3482 564480 46174
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 568580 39364 568632 39370
rect 568580 39306 568632 39312
rect 565820 13184 565872 13190
rect 565820 13126 565872 13132
rect 565832 3482 565860 13126
rect 567844 3528 567896 3534
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 567844 3470 567896 3476
rect 568592 3482 568620 39306
rect 571432 37936 571484 37942
rect 571432 37878 571484 37884
rect 569960 31068 570012 31074
rect 569960 31010 570012 31016
rect 569972 3482 570000 31010
rect 571444 3534 571472 37878
rect 574744 36576 574796 36582
rect 574744 36518 574796 36524
rect 574756 3534 574784 36518
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 579804 7608 579856 7614
rect 579804 7550 579856 7556
rect 575020 4004 575072 4010
rect 575020 3946 575072 3952
rect 571432 3528 571484 3534
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3470
rect 568592 3454 569080 3482
rect 569972 3454 570276 3482
rect 571432 3470 571484 3476
rect 572628 3528 572680 3534
rect 572628 3470 572680 3476
rect 574744 3528 574796 3534
rect 574744 3470 574796 3476
rect 569052 480 569080 3454
rect 570248 480 570276 3454
rect 571432 3256 571484 3262
rect 571432 3198 571484 3204
rect 571444 480 571472 3198
rect 572640 480 572668 3470
rect 573824 3188 573876 3194
rect 573824 3130 573876 3136
rect 573836 480 573864 3130
rect 575032 480 575060 3946
rect 576216 3528 576268 3534
rect 576216 3470 576268 3476
rect 576228 480 576256 3470
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 577412 3392 577464 3398
rect 577412 3334 577464 3340
rect 577424 480 577452 3334
rect 578620 480 578648 3402
rect 579816 480 579844 7550
rect 582196 3732 582248 3738
rect 582196 3674 582248 3680
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 3674
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667936 3478 667992
rect 3606 653520 3662 653576
rect 3514 624824 3570 624880
rect 3422 610408 3478 610464
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 580170 697992 580226 698048
rect 59358 644680 59414 644736
rect 580170 686296 580226 686352
rect 580262 674600 580318 674656
rect 523774 645224 523830 645280
rect 580170 639376 580226 639432
rect 523682 631896 523738 631952
rect 59358 630400 59414 630456
rect 59358 616120 59414 616176
rect 523130 605240 523186 605296
rect 59358 601840 59414 601896
rect 3514 595992 3570 596048
rect 59358 587560 59414 587616
rect 59358 573280 59414 573336
rect 3422 567296 3478 567352
rect 523130 565256 523186 565312
rect 59358 559000 59414 559056
rect 3422 553016 3478 553072
rect 580446 651072 580502 651128
rect 580354 627680 580410 627736
rect 524326 618568 524382 618624
rect 579802 592456 579858 592512
rect 523774 591912 523830 591968
rect 580262 580760 580318 580816
rect 524326 578584 524382 578640
rect 580170 557232 580226 557288
rect 523682 551928 523738 551984
rect 59358 544720 59414 544776
rect 3422 538600 3478 538656
rect 523682 538600 523738 538656
rect 59358 530440 59414 530496
rect 59358 516160 59414 516216
rect 580170 545536 580226 545592
rect 580446 604152 580502 604208
rect 580262 533840 580318 533896
rect 523774 525272 523830 525328
rect 523682 511944 523738 512000
rect 580170 510312 580226 510368
rect 3146 509904 3202 509960
rect 60002 501880 60058 501936
rect 523682 498616 523738 498672
rect 3422 495488 3478 495544
rect 59358 487600 59414 487656
rect 3514 481072 3570 481128
rect 60002 473320 60058 473376
rect 580170 498616 580226 498672
rect 580262 486784 580318 486840
rect 523774 485288 523830 485344
rect 523682 471960 523738 472016
rect 580170 463392 580226 463448
rect 60094 459040 60150 459096
rect 3422 452376 3478 452432
rect 60002 444760 60058 444816
rect 3146 437960 3202 438016
rect 524326 458632 524382 458688
rect 580170 451696 580226 451752
rect 523682 445304 523738 445360
rect 60094 430480 60150 430536
rect 3238 423680 3294 423736
rect 60002 401920 60058 401976
rect 3146 394984 3202 395040
rect 3238 380568 3294 380624
rect 580170 439864 580226 439920
rect 523774 431976 523830 432032
rect 523682 418648 523738 418704
rect 580170 416472 580226 416528
rect 60186 416200 60242 416256
rect 60094 387640 60150 387696
rect 3146 366152 3202 366208
rect 60002 359080 60058 359136
rect 3422 337456 3478 337512
rect 3238 323040 3294 323096
rect 523682 405320 523738 405376
rect 580170 404776 580226 404832
rect 580170 392944 580226 393000
rect 523774 391992 523830 392048
rect 523682 378664 523738 378720
rect 60186 373360 60242 373416
rect 60094 330384 60150 330440
rect 3330 308760 3386 308816
rect 3422 294344 3478 294400
rect 60002 287544 60058 287600
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 3146 265648 3202 265704
rect 3422 251232 3478 251288
rect 580170 369552 580226 369608
rect 524234 365336 524290 365392
rect 580170 357856 580226 357912
rect 523682 351872 523738 351928
rect 580170 346024 580226 346080
rect 60370 344664 60426 344720
rect 60278 316104 60334 316160
rect 60186 273264 60242 273320
rect 60094 258984 60150 259040
rect 3422 236952 3478 237008
rect 3146 222536 3202 222592
rect 523774 338544 523830 338600
rect 524326 325216 524382 325272
rect 580170 322632 580226 322688
rect 524326 311888 524382 311944
rect 580170 310800 580226 310856
rect 60462 301824 60518 301880
rect 580170 299104 580226 299160
rect 524326 298560 524382 298616
rect 523682 285232 523738 285288
rect 580170 275712 580226 275768
rect 523682 271904 523738 271960
rect 580170 263880 580226 263936
rect 523682 258576 523738 258632
rect 579802 252184 579858 252240
rect 523682 245248 523738 245304
rect 60278 244704 60334 244760
rect 60186 216144 60242 216200
rect 3422 208120 3478 208176
rect 60094 201864 60150 201920
rect 3146 193840 3202 193896
rect 60002 187584 60058 187640
rect 3238 179424 3294 179480
rect 3514 165008 3570 165064
rect 3146 150728 3202 150784
rect 60370 230424 60426 230480
rect 523774 231920 523830 231976
rect 580170 228792 580226 228848
rect 523866 218592 523922 218648
rect 580170 216960 580226 217016
rect 523682 205264 523738 205320
rect 579802 205264 579858 205320
rect 523774 191936 523830 191992
rect 60370 173304 60426 173360
rect 60278 159024 60334 159080
rect 60186 144744 60242 144800
rect 3238 136312 3294 136368
rect 60002 130464 60058 130520
rect 3422 122032 3478 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 60094 116184 60150 116240
rect 3422 78920 3478 78976
rect 60002 73344 60058 73400
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 580170 181872 580226 181928
rect 523866 178608 523922 178664
rect 523682 165280 523738 165336
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 523774 151952 523830 152008
rect 523682 125296 523738 125352
rect 60278 101904 60334 101960
rect 60186 87624 60242 87680
rect 60094 59064 60150 59120
rect 3146 21392 3202 21448
rect 523866 138624 523922 138680
rect 523774 111968 523830 112024
rect 523682 85312 523738 85368
rect 3422 7112 3478 7168
rect 92386 3304 92442 3360
rect 153106 3440 153162 3496
rect 153934 3304 153990 3360
rect 157246 3304 157302 3360
rect 214654 3440 214710 3496
rect 218150 3304 218206 3360
rect 231766 3304 231822 3360
rect 293130 3304 293186 3360
rect 364246 3304 364302 3360
rect 371146 3576 371202 3632
rect 407026 3440 407082 3496
rect 425150 3304 425206 3360
rect 432326 3576 432382 3632
rect 449806 3304 449862 3360
rect 467930 3440 467986 3496
rect 485686 3440 485742 3496
rect 510802 3304 510858 3360
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 523866 98640 523922 98696
rect 523774 71984 523830 72040
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 523866 58656 523922 58712
rect 520186 3304 520242 3360
rect 546498 3440 546554 3496
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
rect 580998 3304 581054 3360
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3601 653578 3667 653581
rect -960 653576 3667 653578
rect -960 653520 3606 653576
rect 3662 653520 3667 653576
rect -960 653518 3667 653520
rect -960 653428 480 653518
rect 3601 653515 3667 653518
rect 580441 651130 580507 651133
rect 583520 651130 584960 651220
rect 580441 651128 584960 651130
rect 580441 651072 580446 651128
rect 580502 651072 584960 651128
rect 580441 651070 584960 651072
rect 580441 651067 580507 651070
rect 583520 650980 584960 651070
rect 523769 645282 523835 645285
rect 521916 645280 523835 645282
rect 521916 645224 523774 645280
rect 523830 645224 523835 645280
rect 521916 645222 523835 645224
rect 523769 645219 523835 645222
rect 59353 644738 59419 644741
rect 59353 644736 62100 644738
rect 59353 644680 59358 644736
rect 59414 644680 62100 644736
rect 59353 644678 62100 644680
rect 59353 644675 59419 644678
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 523677 631954 523743 631957
rect 521916 631952 523743 631954
rect 521916 631896 523682 631952
rect 523738 631896 523743 631952
rect 521916 631894 523743 631896
rect 523677 631891 523743 631894
rect 59353 630458 59419 630461
rect 59353 630456 62100 630458
rect 59353 630400 59358 630456
rect 59414 630400 62100 630456
rect 59353 630398 62100 630400
rect 59353 630395 59419 630398
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3509 624882 3575 624885
rect -960 624880 3575 624882
rect -960 624824 3514 624880
rect 3570 624824 3575 624880
rect -960 624822 3575 624824
rect -960 624732 480 624822
rect 3509 624819 3575 624822
rect 524321 618626 524387 618629
rect 521916 618624 524387 618626
rect 521916 618568 524326 618624
rect 524382 618568 524387 618624
rect 521916 618566 524387 618568
rect 524321 618563 524387 618566
rect 59353 616178 59419 616181
rect 59353 616176 62100 616178
rect 59353 616120 59358 616176
rect 59414 616120 62100 616176
rect 59353 616118 62100 616120
rect 59353 616115 59419 616118
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 523125 605298 523191 605301
rect 521916 605296 523191 605298
rect 521916 605240 523130 605296
rect 523186 605240 523191 605296
rect 521916 605238 523191 605240
rect 523125 605235 523191 605238
rect 580441 604210 580507 604213
rect 583520 604210 584960 604300
rect 580441 604208 584960 604210
rect 580441 604152 580446 604208
rect 580502 604152 584960 604208
rect 580441 604150 584960 604152
rect 580441 604147 580507 604150
rect 583520 604060 584960 604150
rect 59353 601898 59419 601901
rect 59353 601896 62100 601898
rect 59353 601840 59358 601896
rect 59414 601840 62100 601896
rect 59353 601838 62100 601840
rect 59353 601835 59419 601838
rect -960 596050 480 596140
rect 3509 596050 3575 596053
rect -960 596048 3575 596050
rect -960 595992 3514 596048
rect 3570 595992 3575 596048
rect -960 595990 3575 595992
rect -960 595900 480 595990
rect 3509 595987 3575 595990
rect 579797 592514 579863 592517
rect 583520 592514 584960 592604
rect 579797 592512 584960 592514
rect 579797 592456 579802 592512
rect 579858 592456 584960 592512
rect 579797 592454 584960 592456
rect 579797 592451 579863 592454
rect 583520 592364 584960 592454
rect 523769 591970 523835 591973
rect 521916 591968 523835 591970
rect 521916 591912 523774 591968
rect 523830 591912 523835 591968
rect 521916 591910 523835 591912
rect 523769 591907 523835 591910
rect 59353 587618 59419 587621
rect 59353 587616 62100 587618
rect 59353 587560 59358 587616
rect 59414 587560 62100 587616
rect 59353 587558 62100 587560
rect 59353 587555 59419 587558
rect -960 581620 480 581860
rect 580257 580818 580323 580821
rect 583520 580818 584960 580908
rect 580257 580816 584960 580818
rect 580257 580760 580262 580816
rect 580318 580760 584960 580816
rect 580257 580758 584960 580760
rect 580257 580755 580323 580758
rect 583520 580668 584960 580758
rect 524321 578642 524387 578645
rect 521916 578640 524387 578642
rect 521916 578584 524326 578640
rect 524382 578584 524387 578640
rect 521916 578582 524387 578584
rect 524321 578579 524387 578582
rect 59353 573338 59419 573341
rect 59353 573336 62100 573338
rect 59353 573280 59358 573336
rect 59414 573280 62100 573336
rect 59353 573278 62100 573280
rect 59353 573275 59419 573278
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 523125 565314 523191 565317
rect 521916 565312 523191 565314
rect 521916 565256 523130 565312
rect 523186 565256 523191 565312
rect 521916 565254 523191 565256
rect 523125 565251 523191 565254
rect 59353 559058 59419 559061
rect 59353 559056 62100 559058
rect 59353 559000 59358 559056
rect 59414 559000 62100 559056
rect 59353 558998 62100 559000
rect 59353 558995 59419 558998
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3417 553074 3483 553077
rect -960 553072 3483 553074
rect -960 553016 3422 553072
rect 3478 553016 3483 553072
rect -960 553014 3483 553016
rect -960 552924 480 553014
rect 3417 553011 3483 553014
rect 523677 551986 523743 551989
rect 521916 551984 523743 551986
rect 521916 551928 523682 551984
rect 523738 551928 523743 551984
rect 521916 551926 523743 551928
rect 523677 551923 523743 551926
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 59353 544778 59419 544781
rect 59353 544776 62100 544778
rect 59353 544720 59358 544776
rect 59414 544720 62100 544776
rect 59353 544718 62100 544720
rect 59353 544715 59419 544718
rect -960 538658 480 538748
rect 3417 538658 3483 538661
rect 523677 538658 523743 538661
rect -960 538656 3483 538658
rect -960 538600 3422 538656
rect 3478 538600 3483 538656
rect -960 538598 3483 538600
rect 521916 538656 523743 538658
rect 521916 538600 523682 538656
rect 523738 538600 523743 538656
rect 521916 538598 523743 538600
rect -960 538508 480 538598
rect 3417 538595 3483 538598
rect 523677 538595 523743 538598
rect 580257 533898 580323 533901
rect 583520 533898 584960 533988
rect 580257 533896 584960 533898
rect 580257 533840 580262 533896
rect 580318 533840 584960 533896
rect 580257 533838 584960 533840
rect 580257 533835 580323 533838
rect 583520 533748 584960 533838
rect 59353 530498 59419 530501
rect 59353 530496 62100 530498
rect 59353 530440 59358 530496
rect 59414 530440 62100 530496
rect 59353 530438 62100 530440
rect 59353 530435 59419 530438
rect 523769 525330 523835 525333
rect 521916 525328 523835 525330
rect 521916 525272 523774 525328
rect 523830 525272 523835 525328
rect 521916 525270 523835 525272
rect 523769 525267 523835 525270
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 59353 516218 59419 516221
rect 59353 516216 62100 516218
rect 59353 516160 59358 516216
rect 59414 516160 62100 516216
rect 59353 516158 62100 516160
rect 59353 516155 59419 516158
rect 523677 512002 523743 512005
rect 521916 512000 523743 512002
rect 521916 511944 523682 512000
rect 523738 511944 523743 512000
rect 521916 511942 523743 511944
rect 523677 511939 523743 511942
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3141 509962 3207 509965
rect -960 509960 3207 509962
rect -960 509904 3146 509960
rect 3202 509904 3207 509960
rect -960 509902 3207 509904
rect -960 509812 480 509902
rect 3141 509899 3207 509902
rect 59997 501938 60063 501941
rect 59997 501936 62100 501938
rect 59997 501880 60002 501936
rect 60058 501880 62100 501936
rect 59997 501878 62100 501880
rect 59997 501875 60063 501878
rect 523677 498674 523743 498677
rect 521916 498672 523743 498674
rect 521916 498616 523682 498672
rect 523738 498616 523743 498672
rect 521916 498614 523743 498616
rect 523677 498611 523743 498614
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3417 495546 3483 495549
rect -960 495544 3483 495546
rect -960 495488 3422 495544
rect 3478 495488 3483 495544
rect -960 495486 3483 495488
rect -960 495396 480 495486
rect 3417 495483 3483 495486
rect 59353 487658 59419 487661
rect 59353 487656 62100 487658
rect 59353 487600 59358 487656
rect 59414 487600 62100 487656
rect 59353 487598 62100 487600
rect 59353 487595 59419 487598
rect 580257 486842 580323 486845
rect 583520 486842 584960 486932
rect 580257 486840 584960 486842
rect 580257 486784 580262 486840
rect 580318 486784 584960 486840
rect 580257 486782 584960 486784
rect 580257 486779 580323 486782
rect 583520 486692 584960 486782
rect 523769 485346 523835 485349
rect 521916 485344 523835 485346
rect 521916 485288 523774 485344
rect 523830 485288 523835 485344
rect 521916 485286 523835 485288
rect 523769 485283 523835 485286
rect -960 481130 480 481220
rect 3509 481130 3575 481133
rect -960 481128 3575 481130
rect -960 481072 3514 481128
rect 3570 481072 3575 481128
rect -960 481070 3575 481072
rect -960 480980 480 481070
rect 3509 481067 3575 481070
rect 583520 474996 584960 475236
rect 59997 473378 60063 473381
rect 59997 473376 62100 473378
rect 59997 473320 60002 473376
rect 60058 473320 62100 473376
rect 59997 473318 62100 473320
rect 59997 473315 60063 473318
rect 523677 472018 523743 472021
rect 521916 472016 523743 472018
rect 521916 471960 523682 472016
rect 523738 471960 523743 472016
rect 521916 471958 523743 471960
rect 523677 471955 523743 471958
rect -960 466700 480 466940
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 60089 459098 60155 459101
rect 60089 459096 62100 459098
rect 60089 459040 60094 459096
rect 60150 459040 62100 459096
rect 60089 459038 62100 459040
rect 60089 459035 60155 459038
rect 524321 458690 524387 458693
rect 521916 458688 524387 458690
rect 521916 458632 524326 458688
rect 524382 458632 524387 458688
rect 521916 458630 524387 458632
rect 524321 458627 524387 458630
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 523677 445362 523743 445365
rect 521916 445360 523743 445362
rect 521916 445304 523682 445360
rect 523738 445304 523743 445360
rect 521916 445302 523743 445304
rect 523677 445299 523743 445302
rect 59997 444818 60063 444821
rect 59997 444816 62100 444818
rect 59997 444760 60002 444816
rect 60058 444760 62100 444816
rect 59997 444758 62100 444760
rect 59997 444755 60063 444758
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 523769 432034 523835 432037
rect 521916 432032 523835 432034
rect 521916 431976 523774 432032
rect 523830 431976 523835 432032
rect 521916 431974 523835 431976
rect 523769 431971 523835 431974
rect 60089 430538 60155 430541
rect 60089 430536 62100 430538
rect 60089 430480 60094 430536
rect 60150 430480 62100 430536
rect 60089 430478 62100 430480
rect 60089 430475 60155 430478
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 523677 418706 523743 418709
rect 521916 418704 523743 418706
rect 521916 418648 523682 418704
rect 523738 418648 523743 418704
rect 521916 418646 523743 418648
rect 523677 418643 523743 418646
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 60181 416258 60247 416261
rect 60181 416256 62100 416258
rect 60181 416200 60186 416256
rect 60242 416200 62100 416256
rect 60181 416198 62100 416200
rect 60181 416195 60247 416198
rect -960 409172 480 409412
rect 523677 405378 523743 405381
rect 521916 405376 523743 405378
rect 521916 405320 523682 405376
rect 523738 405320 523743 405376
rect 521916 405318 523743 405320
rect 523677 405315 523743 405318
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 59997 401978 60063 401981
rect 59997 401976 62100 401978
rect 59997 401920 60002 401976
rect 60058 401920 62100 401976
rect 59997 401918 62100 401920
rect 59997 401915 60063 401918
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 523769 392050 523835 392053
rect 521916 392048 523835 392050
rect 521916 391992 523774 392048
rect 523830 391992 523835 392048
rect 521916 391990 523835 391992
rect 523769 391987 523835 391990
rect 60089 387698 60155 387701
rect 60089 387696 62100 387698
rect 60089 387640 60094 387696
rect 60150 387640 62100 387696
rect 60089 387638 62100 387640
rect 60089 387635 60155 387638
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 523677 378722 523743 378725
rect 521916 378720 523743 378722
rect 521916 378664 523682 378720
rect 523738 378664 523743 378720
rect 521916 378662 523743 378664
rect 523677 378659 523743 378662
rect 60181 373418 60247 373421
rect 60181 373416 62100 373418
rect 60181 373360 60186 373416
rect 60242 373360 62100 373416
rect 60181 373358 62100 373360
rect 60181 373355 60247 373358
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 524229 365394 524295 365397
rect 521916 365392 524295 365394
rect 521916 365336 524234 365392
rect 524290 365336 524295 365392
rect 521916 365334 524295 365336
rect 524229 365331 524295 365334
rect 59997 359138 60063 359141
rect 59997 359136 62100 359138
rect 59997 359080 60002 359136
rect 60058 359080 62100 359136
rect 59997 359078 62100 359080
rect 59997 359075 60063 359078
rect 580165 357914 580231 357917
rect 583520 357914 584960 358004
rect 580165 357912 584960 357914
rect 580165 357856 580170 357912
rect 580226 357856 584960 357912
rect 580165 357854 584960 357856
rect 580165 357851 580231 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 523677 351930 523743 351933
rect 521916 351928 523743 351930
rect 521916 351872 523682 351928
rect 523738 351872 523743 351928
rect 521916 351870 523743 351872
rect 523677 351867 523743 351870
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 60365 344722 60431 344725
rect 60365 344720 62100 344722
rect 60365 344664 60370 344720
rect 60426 344664 62100 344720
rect 60365 344662 62100 344664
rect 60365 344659 60431 344662
rect 523769 338602 523835 338605
rect 521916 338600 523835 338602
rect 521916 338544 523774 338600
rect 523830 338544 523835 338600
rect 521916 338542 523835 338544
rect 523769 338539 523835 338542
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 583520 334236 584960 334476
rect 60089 330442 60155 330445
rect 60089 330440 62100 330442
rect 60089 330384 60094 330440
rect 60150 330384 62100 330440
rect 60089 330382 62100 330384
rect 60089 330379 60155 330382
rect 524321 325274 524387 325277
rect 521916 325272 524387 325274
rect 521916 325216 524326 325272
rect 524382 325216 524387 325272
rect 521916 325214 524387 325216
rect 524321 325211 524387 325214
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 60273 316162 60339 316165
rect 60273 316160 62100 316162
rect 60273 316104 60278 316160
rect 60334 316104 62100 316160
rect 60273 316102 62100 316104
rect 60273 316099 60339 316102
rect 524321 311946 524387 311949
rect 521916 311944 524387 311946
rect 521916 311888 524326 311944
rect 524382 311888 524387 311944
rect 521916 311886 524387 311888
rect 524321 311883 524387 311886
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 60457 301882 60523 301885
rect 60457 301880 62100 301882
rect 60457 301824 60462 301880
rect 60518 301824 62100 301880
rect 60457 301822 62100 301824
rect 60457 301819 60523 301822
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect 524321 298618 524387 298621
rect 521916 298616 524387 298618
rect 521916 298560 524326 298616
rect 524382 298560 524387 298616
rect 521916 298558 524387 298560
rect 524321 298555 524387 298558
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 59997 287602 60063 287605
rect 59997 287600 62100 287602
rect 59997 287544 60002 287600
rect 60058 287544 62100 287600
rect 59997 287542 62100 287544
rect 59997 287539 60063 287542
rect 583520 287316 584960 287556
rect 523677 285290 523743 285293
rect 521916 285288 523743 285290
rect 521916 285232 523682 285288
rect 523738 285232 523743 285288
rect 521916 285230 523743 285232
rect 523677 285227 523743 285230
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 60181 273322 60247 273325
rect 60181 273320 62100 273322
rect 60181 273264 60186 273320
rect 60242 273264 62100 273320
rect 60181 273262 62100 273264
rect 60181 273259 60247 273262
rect 523677 271962 523743 271965
rect 521916 271960 523743 271962
rect 521916 271904 523682 271960
rect 523738 271904 523743 271960
rect 521916 271902 523743 271904
rect 523677 271899 523743 271902
rect -960 265706 480 265796
rect 3141 265706 3207 265709
rect -960 265704 3207 265706
rect -960 265648 3146 265704
rect 3202 265648 3207 265704
rect -960 265646 3207 265648
rect -960 265556 480 265646
rect 3141 265643 3207 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 60089 259042 60155 259045
rect 60089 259040 62100 259042
rect 60089 258984 60094 259040
rect 60150 258984 62100 259040
rect 60089 258982 62100 258984
rect 60089 258979 60155 258982
rect 523677 258634 523743 258637
rect 521916 258632 523743 258634
rect 521916 258576 523682 258632
rect 523738 258576 523743 258632
rect 521916 258574 523743 258576
rect 523677 258571 523743 258574
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 523677 245306 523743 245309
rect 521916 245304 523743 245306
rect 521916 245248 523682 245304
rect 523738 245248 523743 245304
rect 521916 245246 523743 245248
rect 523677 245243 523743 245246
rect 60273 244762 60339 244765
rect 60273 244760 62100 244762
rect 60273 244704 60278 244760
rect 60334 244704 62100 244760
rect 60273 244702 62100 244704
rect 60273 244699 60339 244702
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 523769 231978 523835 231981
rect 521916 231976 523835 231978
rect 521916 231920 523774 231976
rect 523830 231920 523835 231976
rect 521916 231918 523835 231920
rect 523769 231915 523835 231918
rect 60365 230482 60431 230485
rect 60365 230480 62100 230482
rect 60365 230424 60370 230480
rect 60426 230424 62100 230480
rect 60365 230422 62100 230424
rect 60365 230419 60431 230422
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 523861 218650 523927 218653
rect 521916 218648 523927 218650
rect 521916 218592 523866 218648
rect 523922 218592 523927 218648
rect 521916 218590 523927 218592
rect 523861 218587 523927 218590
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 60181 216202 60247 216205
rect 60181 216200 62100 216202
rect 60181 216144 60186 216200
rect 60242 216144 62100 216200
rect 60181 216142 62100 216144
rect 60181 216139 60247 216142
rect -960 208178 480 208268
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 523677 205322 523743 205325
rect 521916 205320 523743 205322
rect 521916 205264 523682 205320
rect 523738 205264 523743 205320
rect 521916 205262 523743 205264
rect 523677 205259 523743 205262
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 60089 201922 60155 201925
rect 60089 201920 62100 201922
rect 60089 201864 60094 201920
rect 60150 201864 62100 201920
rect 60089 201862 62100 201864
rect 60089 201859 60155 201862
rect -960 193898 480 193988
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 523769 191994 523835 191997
rect 521916 191992 523835 191994
rect 521916 191936 523774 191992
rect 523830 191936 523835 191992
rect 521916 191934 523835 191936
rect 523769 191931 523835 191934
rect 59997 187642 60063 187645
rect 59997 187640 62100 187642
rect 59997 187584 60002 187640
rect 60058 187584 62100 187640
rect 59997 187582 62100 187584
rect 59997 187579 60063 187582
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 523861 178666 523927 178669
rect 521916 178664 523927 178666
rect 521916 178608 523866 178664
rect 523922 178608 523927 178664
rect 521916 178606 523927 178608
rect 523861 178603 523927 178606
rect 60365 173362 60431 173365
rect 60365 173360 62100 173362
rect 60365 173304 60370 173360
rect 60426 173304 62100 173360
rect 60365 173302 62100 173304
rect 60365 173299 60431 173302
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 523677 165338 523743 165341
rect 521916 165336 523743 165338
rect 521916 165280 523682 165336
rect 523738 165280 523743 165336
rect 521916 165278 523743 165280
rect 523677 165275 523743 165278
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 60273 159082 60339 159085
rect 60273 159080 62100 159082
rect 60273 159024 60278 159080
rect 60334 159024 62100 159080
rect 60273 159022 62100 159024
rect 60273 159019 60339 159022
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 523769 152010 523835 152013
rect 521916 152008 523835 152010
rect 521916 151952 523774 152008
rect 523830 151952 523835 152008
rect 521916 151950 523835 151952
rect 523769 151947 523835 151950
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect 60181 144802 60247 144805
rect 60181 144800 62100 144802
rect 60181 144744 60186 144800
rect 60242 144744 62100 144800
rect 60181 144742 62100 144744
rect 60181 144739 60247 144742
rect 523861 138682 523927 138685
rect 521916 138680 523927 138682
rect 521916 138624 523866 138680
rect 523922 138624 523927 138680
rect 521916 138622 523927 138624
rect 523861 138619 523927 138622
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 59997 130522 60063 130525
rect 59997 130520 62100 130522
rect 59997 130464 60002 130520
rect 60058 130464 62100 130520
rect 59997 130462 62100 130464
rect 59997 130459 60063 130462
rect 523677 125354 523743 125357
rect 521916 125352 523743 125354
rect 521916 125296 523682 125352
rect 523738 125296 523743 125352
rect 521916 125294 523743 125296
rect 523677 125291 523743 125294
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 60089 116242 60155 116245
rect 60089 116240 62100 116242
rect 60089 116184 60094 116240
rect 60150 116184 62100 116240
rect 60089 116182 62100 116184
rect 60089 116179 60155 116182
rect 523769 112026 523835 112029
rect 521916 112024 523835 112026
rect 521916 111968 523774 112024
rect 523830 111968 523835 112024
rect 521916 111966 523835 111968
rect 523769 111963 523835 111966
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 60273 101962 60339 101965
rect 60273 101960 62100 101962
rect 60273 101904 60278 101960
rect 60334 101904 62100 101960
rect 60273 101902 62100 101904
rect 60273 101899 60339 101902
rect 583520 99636 584960 99876
rect 523861 98698 523927 98701
rect 521916 98696 523927 98698
rect 521916 98640 523866 98696
rect 523922 98640 523927 98696
rect 521916 98638 523927 98640
rect 523861 98635 523927 98638
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 60181 87682 60247 87685
rect 60181 87680 62100 87682
rect 60181 87624 60186 87680
rect 60242 87624 62100 87680
rect 60181 87622 62100 87624
rect 60181 87619 60247 87622
rect 523677 85370 523743 85373
rect 521916 85368 523743 85370
rect 521916 85312 523682 85368
rect 523738 85312 523743 85368
rect 521916 85310 523743 85312
rect 523677 85307 523743 85310
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 59997 73402 60063 73405
rect 59997 73400 62100 73402
rect 59997 73344 60002 73400
rect 60058 73344 62100 73400
rect 59997 73342 62100 73344
rect 59997 73339 60063 73342
rect 523769 72042 523835 72045
rect 521916 72040 523835 72042
rect 521916 71984 523774 72040
rect 523830 71984 523835 72040
rect 521916 71982 523835 71984
rect 523769 71979 523835 71982
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 60089 59122 60155 59125
rect 60089 59120 62100 59122
rect 60089 59064 60094 59120
rect 60150 59064 62100 59120
rect 60089 59062 62100 59064
rect 60089 59059 60155 59062
rect 523861 58714 523927 58717
rect 521916 58712 523927 58714
rect 521916 58656 523866 58712
rect 523922 58656 523927 58712
rect 521916 58654 523927 58656
rect 523861 58651 523927 58654
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 371141 3634 371207 3637
rect 432321 3634 432387 3637
rect 371141 3632 432387 3634
rect 371141 3576 371146 3632
rect 371202 3576 432326 3632
rect 432382 3576 432387 3632
rect 371141 3574 432387 3576
rect 371141 3571 371207 3574
rect 432321 3571 432387 3574
rect 153101 3498 153167 3501
rect 214649 3498 214715 3501
rect 153101 3496 214715 3498
rect 153101 3440 153106 3496
rect 153162 3440 214654 3496
rect 214710 3440 214715 3496
rect 153101 3438 214715 3440
rect 153101 3435 153167 3438
rect 214649 3435 214715 3438
rect 407021 3498 407087 3501
rect 467925 3498 467991 3501
rect 407021 3496 467991 3498
rect 407021 3440 407026 3496
rect 407082 3440 467930 3496
rect 467986 3440 467991 3496
rect 407021 3438 467991 3440
rect 407021 3435 407087 3438
rect 467925 3435 467991 3438
rect 485681 3498 485747 3501
rect 546493 3498 546559 3501
rect 485681 3496 546559 3498
rect 485681 3440 485686 3496
rect 485742 3440 546498 3496
rect 546554 3440 546559 3496
rect 485681 3438 546559 3440
rect 485681 3435 485747 3438
rect 546493 3435 546559 3438
rect 92381 3362 92447 3365
rect 153929 3362 153995 3365
rect 92381 3360 153995 3362
rect 92381 3304 92386 3360
rect 92442 3304 153934 3360
rect 153990 3304 153995 3360
rect 92381 3302 153995 3304
rect 92381 3299 92447 3302
rect 153929 3299 153995 3302
rect 157241 3362 157307 3365
rect 218145 3362 218211 3365
rect 157241 3360 218211 3362
rect 157241 3304 157246 3360
rect 157302 3304 218150 3360
rect 218206 3304 218211 3360
rect 157241 3302 218211 3304
rect 157241 3299 157307 3302
rect 218145 3299 218211 3302
rect 231761 3362 231827 3365
rect 293125 3362 293191 3365
rect 231761 3360 293191 3362
rect 231761 3304 231766 3360
rect 231822 3304 293130 3360
rect 293186 3304 293191 3360
rect 231761 3302 293191 3304
rect 231761 3299 231827 3302
rect 293125 3299 293191 3302
rect 364241 3362 364307 3365
rect 425145 3362 425211 3365
rect 364241 3360 425211 3362
rect 364241 3304 364246 3360
rect 364302 3304 425150 3360
rect 425206 3304 425211 3360
rect 364241 3302 425211 3304
rect 364241 3299 364307 3302
rect 425145 3299 425211 3302
rect 449801 3362 449867 3365
rect 510797 3362 510863 3365
rect 449801 3360 510863 3362
rect 449801 3304 449806 3360
rect 449862 3304 510802 3360
rect 510858 3304 510863 3360
rect 449801 3302 510863 3304
rect 449801 3299 449867 3302
rect 510797 3299 510863 3302
rect 520181 3362 520247 3365
rect 580993 3362 581059 3365
rect 520181 3360 581059 3362
rect 520181 3304 520186 3360
rect 520242 3304 580998 3360
rect 581054 3304 581059 3360
rect 520181 3302 581059 3304
rect 520181 3299 520247 3302
rect 580993 3299 581059 3302
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 652000 62604 675098
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 652000 66204 678698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 652000 73404 685898
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 652000 77004 653498
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 652000 80604 657098
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 652000 84204 660698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 652000 91404 667898
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 652000 95004 671498
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 652000 98604 675098
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 652000 102204 678698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 652000 109404 685898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 652000 113004 653498
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 652000 116604 657098
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 652000 120204 660698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 652000 127404 667898
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 652000 131004 671498
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 652000 134604 675098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 652000 138204 678698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 652000 145404 685898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 652000 149004 653498
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 652000 152604 657098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 652000 156204 660698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 652000 163404 667898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 652000 167004 671498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 652000 170604 675098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 652000 174204 678698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 652000 181404 685898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 652000 185004 653498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 652000 188604 657098
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 652000 192204 660698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 652000 199404 667898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 652000 203004 671498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 652000 206604 675098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 652000 210204 678698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 652000 217404 685898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 652000 221004 653498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 652000 224604 657098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 652000 228204 660698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 652000 235404 667898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 652000 239004 671498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 652000 242604 675098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 652000 246204 678698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 652000 253404 685898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 652000 257004 653498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 652000 260604 657098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 652000 264204 660698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 652000 271404 667898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 652000 275004 671498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 652000 278604 675098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 652000 282204 678698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 652000 289404 685898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 652000 293004 653498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 652000 296604 657098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 652000 300204 660698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 652000 307404 667898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 652000 311004 671498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 652000 314604 675098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 652000 318204 678698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 652000 325404 685898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 652000 329004 653498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 652000 332604 657098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 652000 336204 660698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 652000 343404 667898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 652000 347004 671498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 652000 350604 675098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 652000 354204 678698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 652000 361404 685898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 652000 365004 653498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 652000 368604 657098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 652000 372204 660698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 652000 379404 667898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 652000 383004 671498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 652000 386604 675098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 652000 390204 678698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 652000 397404 685898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 652000 401004 653498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 652000 404604 657098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 652000 408204 660698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 652000 415404 667898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 652000 419004 671498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 652000 422604 675098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 652000 426204 678698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 652000 433404 685898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 652000 437004 653498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 652000 440604 657098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 652000 444204 660698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 652000 451404 667898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 652000 455004 671498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 652000 458604 675098
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 652000 462204 678698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 652000 469404 685898
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 652000 473004 653498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 652000 476604 657098
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 652000 480204 660698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 652000 487404 667898
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 652000 491004 671498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 652000 494604 675098
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 652000 498204 678698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 652000 505404 685898
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 652000 509004 653498
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 652000 512604 657098
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 652000 516204 660698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 27654 62604 52000
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 31254 66204 52000
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 38454 73404 52000
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 42054 77004 52000
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 45654 80604 52000
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 49254 84204 52000
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 20454 91404 52000
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 24054 95004 52000
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 27654 98604 52000
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 31254 102204 52000
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 38454 109404 52000
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 42054 113004 52000
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 45654 116604 52000
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 49254 120204 52000
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 20454 127404 52000
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 24054 131004 52000
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 27654 134604 52000
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 31254 138204 52000
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 38454 145404 52000
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 42054 149004 52000
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 45654 152604 52000
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 49254 156204 52000
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 20454 163404 52000
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 24054 167004 52000
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 27654 170604 52000
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 31254 174204 52000
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 38454 181404 52000
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 42054 185004 52000
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 45654 188604 52000
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 49254 192204 52000
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 20454 199404 52000
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 24054 203004 52000
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 27654 206604 52000
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 31254 210204 52000
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 38454 217404 52000
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 42054 221004 52000
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 45654 224604 52000
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 49254 228204 52000
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 20454 235404 52000
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 24054 239004 52000
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 27654 242604 52000
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 31254 246204 52000
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 38454 253404 52000
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 42054 257004 52000
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 45654 260604 52000
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 49254 264204 52000
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 20454 271404 52000
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 24054 275004 52000
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 27654 278604 52000
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 31254 282204 52000
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 38454 289404 52000
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 42054 293004 52000
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 45654 296604 52000
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 49254 300204 52000
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 20454 307404 52000
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 24054 311004 52000
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 27654 314604 52000
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 31254 318204 52000
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 38454 325404 52000
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 42054 329004 52000
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 45654 332604 52000
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 49254 336204 52000
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 20454 343404 52000
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 24054 347004 52000
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 27654 350604 52000
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 31254 354204 52000
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 38454 361404 52000
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 42054 365004 52000
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 45654 368604 52000
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 49254 372204 52000
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 20454 379404 52000
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 24054 383004 52000
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 27654 386604 52000
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 31254 390204 52000
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 38454 397404 52000
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 42054 401004 52000
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 45654 404604 52000
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 49254 408204 52000
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 20454 415404 52000
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 24054 419004 52000
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 27654 422604 52000
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 31254 426204 52000
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 38454 433404 52000
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 42054 437004 52000
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 45654 440604 52000
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 49254 444204 52000
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 20454 451404 52000
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 24054 455004 52000
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 27654 458604 52000
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 31254 462204 52000
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 38454 469404 52000
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 42054 473004 52000
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 45654 476604 52000
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 49254 480204 52000
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 20454 487404 52000
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 24054 491004 52000
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 27654 494604 52000
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 31254 498204 52000
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 38454 505404 52000
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 42054 509004 52000
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 45654 512604 52000
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 49254 516204 52000
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use ghazi_top_dffram_csv  mprj
timestamp 1607663363
transform 1 0 62000 0 1 52000
box 0 0 460000 600000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
