VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3519.700 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3519.700 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3519.700 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3519.700 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3519.700 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3519.700 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3519.700 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3519.700 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3519.700 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 0.300 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 0.300 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 0.300 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 0.300 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 0.300 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 0.300 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 0.300 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2619.310 89.660 2619.630 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2619.310 89.520 2899.310 89.660 ;
        RECT 2619.310 89.460 2619.630 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2619.340 89.460 2619.600 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2619.330 293.235 2619.610 293.605 ;
        RECT 2619.400 89.750 2619.540 293.235 ;
        RECT 2619.340 89.430 2619.600 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2619.330 293.280 2619.610 293.560 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 293.570 2610.000 293.960 ;
        RECT 2619.305 293.570 2619.635 293.585 ;
        RECT 2606.000 293.360 2619.635 293.570 ;
        RECT 2609.580 293.270 2619.635 293.360 ;
        RECT 2619.305 293.255 2619.635 293.270 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
=======
        RECT 2919.700 87.460 2924.800 88.660 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2621.610 2297.620 2621.930 2297.680 ;
        RECT 2901.290 2297.620 2901.610 2297.680 ;
        RECT 2621.610 2297.480 2901.610 2297.620 ;
        RECT 2621.610 2297.420 2621.930 2297.480 ;
        RECT 2901.290 2297.420 2901.610 2297.480 ;
      LAYER via ;
        RECT 2621.640 2297.420 2621.900 2297.680 ;
        RECT 2901.320 2297.420 2901.580 2297.680 ;
      LAYER met2 ;
        RECT 2901.310 2433.875 2901.590 2434.245 ;
        RECT 2901.380 2297.710 2901.520 2433.875 ;
        RECT 2621.640 2297.390 2621.900 2297.710 ;
        RECT 2901.320 2297.390 2901.580 2297.710 ;
        RECT 2621.700 2293.485 2621.840 2297.390 ;
        RECT 2621.630 2293.115 2621.910 2293.485 ;
      LAYER via2 ;
        RECT 2901.310 2433.920 2901.590 2434.200 ;
        RECT 2621.630 2293.160 2621.910 2293.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2901.285 2434.210 2901.615 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2901.285 2433.910 2924.800 2434.210 ;
        RECT 2901.285 2433.895 2901.615 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2606.000 2293.450 2610.000 2293.840 ;
        RECT 2621.605 2293.450 2621.935 2293.465 ;
        RECT 2606.000 2293.240 2621.935 2293.450 ;
        RECT 2609.580 2293.150 2621.935 2293.240 ;
        RECT 2621.605 2293.135 2621.935 2293.150 ;
=======
        RECT 2919.700 2433.460 2924.800 2434.660 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2497.540 2618.710 2497.600 ;
        RECT 2901.290 2497.540 2901.610 2497.600 ;
        RECT 2618.390 2497.400 2901.610 2497.540 ;
        RECT 2618.390 2497.340 2618.710 2497.400 ;
        RECT 2901.290 2497.340 2901.610 2497.400 ;
      LAYER via ;
        RECT 2618.420 2497.340 2618.680 2497.600 ;
        RECT 2901.320 2497.340 2901.580 2497.600 ;
      LAYER met2 ;
        RECT 2901.310 2669.155 2901.590 2669.525 ;
        RECT 2901.380 2497.630 2901.520 2669.155 ;
        RECT 2618.420 2497.310 2618.680 2497.630 ;
        RECT 2901.320 2497.310 2901.580 2497.630 ;
        RECT 2618.480 2493.405 2618.620 2497.310 ;
        RECT 2618.410 2493.035 2618.690 2493.405 ;
      LAYER via2 ;
        RECT 2901.310 2669.200 2901.590 2669.480 ;
        RECT 2618.410 2493.080 2618.690 2493.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2901.285 2669.490 2901.615 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2901.285 2669.190 2924.800 2669.490 ;
        RECT 2901.285 2669.175 2901.615 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2606.000 2493.370 2610.000 2493.760 ;
        RECT 2618.385 2493.370 2618.715 2493.385 ;
        RECT 2606.000 2493.160 2618.715 2493.370 ;
        RECT 2609.580 2493.070 2618.715 2493.160 ;
        RECT 2618.385 2493.055 2618.715 2493.070 ;
=======
        RECT 2919.700 2668.740 2924.800 2669.940 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2697.800 2618.710 2697.860 ;
        RECT 2901.290 2697.800 2901.610 2697.860 ;
        RECT 2618.390 2697.660 2901.610 2697.800 ;
        RECT 2618.390 2697.600 2618.710 2697.660 ;
        RECT 2901.290 2697.600 2901.610 2697.660 ;
      LAYER via ;
        RECT 2618.420 2697.600 2618.680 2697.860 ;
        RECT 2901.320 2697.600 2901.580 2697.860 ;
      LAYER met2 ;
        RECT 2901.310 2903.755 2901.590 2904.125 ;
        RECT 2901.380 2697.890 2901.520 2903.755 ;
        RECT 2618.420 2697.570 2618.680 2697.890 ;
        RECT 2901.320 2697.570 2901.580 2697.890 ;
        RECT 2618.480 2693.325 2618.620 2697.570 ;
        RECT 2618.410 2692.955 2618.690 2693.325 ;
      LAYER via2 ;
        RECT 2901.310 2903.800 2901.590 2904.080 ;
        RECT 2618.410 2693.000 2618.690 2693.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2901.285 2904.090 2901.615 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2901.285 2903.790 2924.800 2904.090 ;
        RECT 2901.285 2903.775 2901.615 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2606.000 2693.290 2610.000 2693.680 ;
        RECT 2618.385 2693.290 2618.715 2693.305 ;
        RECT 2606.000 2693.080 2618.715 2693.290 ;
        RECT 2609.580 2692.990 2618.715 2693.080 ;
        RECT 2618.385 2692.975 2618.715 2692.990 ;
=======
        RECT 2919.700 2903.340 2924.800 2904.540 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2621.610 2898.060 2621.930 2898.120 ;
        RECT 2901.750 2898.060 2902.070 2898.120 ;
        RECT 2621.610 2897.920 2902.070 2898.060 ;
        RECT 2621.610 2897.860 2621.930 2897.920 ;
        RECT 2901.750 2897.860 2902.070 2897.920 ;
      LAYER via ;
        RECT 2621.640 2897.860 2621.900 2898.120 ;
        RECT 2901.780 2897.860 2902.040 2898.120 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 2901.840 2898.150 2901.980 3138.355 ;
        RECT 2621.640 2897.830 2621.900 2898.150 ;
        RECT 2901.780 2897.830 2902.040 2898.150 ;
        RECT 2621.700 2893.245 2621.840 2897.830 ;
        RECT 2621.630 2892.875 2621.910 2893.245 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
        RECT 2621.630 2892.920 2621.910 2893.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2606.000 2893.210 2610.000 2893.600 ;
        RECT 2621.605 2893.210 2621.935 2893.225 ;
        RECT 2606.000 2893.000 2621.935 2893.210 ;
        RECT 2609.580 2892.910 2621.935 2893.000 ;
        RECT 2621.605 2892.895 2621.935 2892.910 ;
=======
        RECT 2919.700 3137.940 2924.800 3139.140 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2621.610 3097.980 2621.930 3098.040 ;
        RECT 2901.290 3097.980 2901.610 3098.040 ;
        RECT 2621.610 3097.840 2901.610 3097.980 ;
        RECT 2621.610 3097.780 2621.930 3097.840 ;
        RECT 2901.290 3097.780 2901.610 3097.840 ;
      LAYER via ;
        RECT 2621.640 3097.780 2621.900 3098.040 ;
        RECT 2901.320 3097.780 2901.580 3098.040 ;
      LAYER met2 ;
        RECT 2901.310 3372.955 2901.590 3373.325 ;
        RECT 2901.380 3098.070 2901.520 3372.955 ;
        RECT 2621.640 3097.750 2621.900 3098.070 ;
        RECT 2901.320 3097.750 2901.580 3098.070 ;
        RECT 2621.700 3093.165 2621.840 3097.750 ;
        RECT 2621.630 3092.795 2621.910 3093.165 ;
      LAYER via2 ;
        RECT 2901.310 3373.000 2901.590 3373.280 ;
        RECT 2621.630 3092.840 2621.910 3093.120 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2901.285 3373.290 2901.615 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2901.285 3372.990 2924.800 3373.290 ;
        RECT 2901.285 3372.975 2901.615 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2606.000 3093.130 2610.000 3093.520 ;
        RECT 2621.605 3093.130 2621.935 3093.145 ;
        RECT 2606.000 3092.920 2621.935 3093.130 ;
        RECT 2609.580 3092.830 2621.935 3092.920 ;
        RECT 2621.605 3092.815 2621.935 3092.830 ;
=======
        RECT 2919.700 3372.540 2924.800 3373.740 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2573.310 3502.240 2573.630 3502.300 ;
        RECT 2798.250 3502.240 2798.570 3502.300 ;
        RECT 2573.310 3502.100 2798.570 3502.240 ;
        RECT 2573.310 3502.040 2573.630 3502.100 ;
        RECT 2798.250 3502.040 2798.570 3502.100 ;
        RECT 2566.870 3276.480 2567.190 3276.540 ;
        RECT 2573.310 3276.480 2573.630 3276.540 ;
        RECT 2566.870 3276.340 2573.630 3276.480 ;
        RECT 2566.870 3276.280 2567.190 3276.340 ;
        RECT 2573.310 3276.280 2573.630 3276.340 ;
      LAYER via ;
        RECT 2573.340 3502.040 2573.600 3502.300 ;
        RECT 2798.280 3502.040 2798.540 3502.300 ;
        RECT 2566.900 3276.280 2567.160 3276.540 ;
        RECT 2573.340 3276.280 2573.600 3276.540 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3502.330 2798.480 3517.600 ;
        RECT 2573.340 3502.010 2573.600 3502.330 ;
        RECT 2798.280 3502.010 2798.540 3502.330 ;
        RECT 2573.400 3276.570 2573.540 3502.010 ;
        RECT 2566.900 3276.250 2567.160 3276.570 ;
        RECT 2573.340 3276.250 2573.600 3276.570 ;
        RECT 2566.960 3260.000 2567.100 3276.250 ;
        RECT 2566.850 3256.000 2567.130 3260.000 ;
=======
        RECT 2798.130 3519.700 2798.690 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2318.010 3502.240 2318.330 3502.300 ;
        RECT 2473.950 3502.240 2474.270 3502.300 ;
        RECT 2318.010 3502.100 2474.270 3502.240 ;
        RECT 2318.010 3502.040 2318.330 3502.100 ;
        RECT 2473.950 3502.040 2474.270 3502.100 ;
        RECT 2311.570 3277.500 2311.890 3277.560 ;
        RECT 2318.010 3277.500 2318.330 3277.560 ;
        RECT 2311.570 3277.360 2318.330 3277.500 ;
        RECT 2311.570 3277.300 2311.890 3277.360 ;
        RECT 2318.010 3277.300 2318.330 3277.360 ;
      LAYER via ;
        RECT 2318.040 3502.040 2318.300 3502.300 ;
        RECT 2473.980 3502.040 2474.240 3502.300 ;
        RECT 2311.600 3277.300 2311.860 3277.560 ;
        RECT 2318.040 3277.300 2318.300 3277.560 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3502.330 2474.180 3517.600 ;
        RECT 2318.040 3502.010 2318.300 3502.330 ;
        RECT 2473.980 3502.010 2474.240 3502.330 ;
        RECT 2318.100 3277.590 2318.240 3502.010 ;
        RECT 2311.600 3277.270 2311.860 3277.590 ;
        RECT 2318.040 3277.270 2318.300 3277.590 ;
        RECT 2311.660 3260.000 2311.800 3277.270 ;
        RECT 2311.550 3256.000 2311.830 3260.000 ;
=======
        RECT 2473.830 3519.700 2474.390 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2055.810 3502.240 2056.130 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 2055.810 3502.100 2149.510 3502.240 ;
        RECT 2055.810 3502.040 2056.130 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
      LAYER via ;
        RECT 2055.840 3502.040 2056.100 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 2055.840 3502.010 2056.100 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 2055.900 3260.000 2056.040 3502.010 ;
        RECT 2055.790 3256.000 2056.070 3260.000 ;
=======
        RECT 2149.070 3519.700 2149.630 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1800.510 3498.500 1800.830 3498.560 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1800.510 3498.360 1825.210 3498.500 ;
        RECT 1800.510 3498.300 1800.830 3498.360 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
      LAYER via ;
        RECT 1800.540 3498.300 1800.800 3498.560 ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1800.540 3498.270 1800.800 3498.590 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1800.600 3260.000 1800.740 3498.270 ;
        RECT 1800.490 3256.000 1800.770 3260.000 ;
=======
        RECT 1824.770 3519.700 1825.330 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 3270.700 1504.130 3270.760 ;
        RECT 1544.750 3270.700 1545.070 3270.760 ;
        RECT 1503.810 3270.560 1545.070 3270.700 ;
        RECT 1503.810 3270.500 1504.130 3270.560 ;
        RECT 1544.750 3270.500 1545.070 3270.560 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 3270.500 1504.100 3270.760 ;
        RECT 1544.780 3270.500 1545.040 3270.760 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3270.790 1504.040 3498.270 ;
        RECT 1503.840 3270.470 1504.100 3270.790 ;
        RECT 1544.780 3270.470 1545.040 3270.790 ;
        RECT 1544.840 3260.000 1544.980 3270.470 ;
        RECT 1544.730 3256.000 1545.010 3260.000 ;
=======
        RECT 1500.470 3519.700 1501.030 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2619.310 324.260 2619.630 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2619.310 324.120 2899.310 324.260 ;
        RECT 2619.310 324.060 2619.630 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2619.340 324.060 2619.600 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2619.330 493.155 2619.610 493.525 ;
        RECT 2619.400 324.350 2619.540 493.155 ;
        RECT 2619.340 324.030 2619.600 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2619.330 493.200 2619.610 493.480 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 493.490 2610.000 493.880 ;
        RECT 2619.305 493.490 2619.635 493.505 ;
        RECT 2606.000 493.280 2619.635 493.490 ;
        RECT 2609.580 493.190 2619.635 493.280 ;
        RECT 2619.305 493.175 2619.635 493.190 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
=======
        RECT 2919.700 322.060 2924.800 323.260 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3274.100 1179.830 3274.160 ;
        RECT 1289.450 3274.100 1289.770 3274.160 ;
        RECT 1179.510 3273.960 1289.770 3274.100 ;
        RECT 1179.510 3273.900 1179.830 3273.960 ;
        RECT 1289.450 3273.900 1289.770 3273.960 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3273.900 1179.800 3274.160 ;
        RECT 1289.480 3273.900 1289.740 3274.160 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3274.190 1179.740 3498.270 ;
        RECT 1179.540 3273.870 1179.800 3274.190 ;
        RECT 1289.480 3273.870 1289.740 3274.190 ;
        RECT 1289.540 3260.000 1289.680 3273.870 ;
        RECT 1289.430 3256.000 1289.710 3260.000 ;
=======
        RECT 1175.710 3519.700 1176.270 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 855.210 3501.220 855.530 3501.280 ;
        RECT 851.530 3501.080 855.530 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 855.210 3501.020 855.530 3501.080 ;
        RECT 855.210 3274.440 855.530 3274.500 ;
        RECT 1033.690 3274.440 1034.010 3274.500 ;
        RECT 855.210 3274.300 1034.010 3274.440 ;
        RECT 855.210 3274.240 855.530 3274.300 ;
        RECT 1033.690 3274.240 1034.010 3274.300 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 855.240 3501.020 855.500 3501.280 ;
        RECT 855.240 3274.240 855.500 3274.500 ;
        RECT 1033.720 3274.240 1033.980 3274.500 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 855.240 3500.990 855.500 3501.310 ;
        RECT 855.300 3274.530 855.440 3500.990 ;
        RECT 855.240 3274.210 855.500 3274.530 ;
        RECT 1033.720 3274.210 1033.980 3274.530 ;
        RECT 1033.780 3260.000 1033.920 3274.210 ;
        RECT 1033.670 3256.000 1033.950 3260.000 ;
=======
        RECT 851.410 3519.700 851.970 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 3274.440 531.230 3274.500 ;
        RECT 777.930 3274.440 778.250 3274.500 ;
        RECT 530.910 3274.300 778.250 3274.440 ;
        RECT 530.910 3274.240 531.230 3274.300 ;
        RECT 777.930 3274.240 778.250 3274.300 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 3274.240 531.200 3274.500 ;
        RECT 777.960 3274.240 778.220 3274.500 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 3274.530 531.140 3498.270 ;
        RECT 530.940 3274.210 531.200 3274.530 ;
        RECT 777.960 3274.210 778.220 3274.530 ;
        RECT 778.020 3260.000 778.160 3274.210 ;
        RECT 777.910 3256.000 778.190 3260.000 ;
=======
        RECT 527.110 3519.700 527.670 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 3274.440 206.930 3274.500 ;
        RECT 522.630 3274.440 522.950 3274.500 ;
        RECT 206.610 3274.300 522.950 3274.440 ;
        RECT 206.610 3274.240 206.930 3274.300 ;
        RECT 522.630 3274.240 522.950 3274.300 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 3274.240 206.900 3274.500 ;
        RECT 522.660 3274.240 522.920 3274.500 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 3274.530 206.840 3501.670 ;
        RECT 206.640 3274.210 206.900 3274.530 ;
        RECT 522.660 3274.210 522.920 3274.530 ;
        RECT 522.720 3260.000 522.860 3274.210 ;
        RECT 522.610 3256.000 522.890 3260.000 ;
=======
        RECT 202.350 3519.700 202.910 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 3229.220 18.330 3229.280 ;
        RECT 296.770 3229.220 297.090 3229.280 ;
        RECT 18.010 3229.080 297.090 3229.220 ;
        RECT 18.010 3229.020 18.330 3229.080 ;
        RECT 296.770 3229.020 297.090 3229.080 ;
      LAYER via ;
        RECT 18.040 3229.020 18.300 3229.280 ;
        RECT 296.800 3229.020 297.060 3229.280 ;
      LAYER met2 ;
        RECT 18.030 3411.035 18.310 3411.405 ;
        RECT 18.100 3229.310 18.240 3411.035 ;
        RECT 18.040 3228.990 18.300 3229.310 ;
        RECT 296.800 3228.990 297.060 3229.310 ;
        RECT 296.860 3223.725 297.000 3228.990 ;
        RECT 296.790 3223.355 297.070 3223.725 ;
      LAYER via2 ;
        RECT 18.030 3411.080 18.310 3411.360 ;
        RECT 296.790 3223.400 297.070 3223.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 18.005 3411.370 18.335 3411.385 ;
        RECT -4.800 3411.070 18.335 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 18.005 3411.055 18.335 3411.070 ;
        RECT 296.765 3223.690 297.095 3223.705 ;
        RECT 310.000 3223.690 314.000 3224.080 ;
        RECT 296.765 3223.480 314.000 3223.690 ;
        RECT 296.765 3223.390 310.500 3223.480 ;
        RECT 296.765 3223.375 297.095 3223.390 ;
=======
        RECT -4.800 3410.620 0.300 3411.820 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 3015.360 18.330 3015.420 ;
        RECT 296.770 3015.360 297.090 3015.420 ;
        RECT 18.010 3015.220 297.090 3015.360 ;
        RECT 18.010 3015.160 18.330 3015.220 ;
        RECT 296.770 3015.160 297.090 3015.220 ;
      LAYER via ;
        RECT 18.040 3015.160 18.300 3015.420 ;
        RECT 296.800 3015.160 297.060 3015.420 ;
      LAYER met2 ;
        RECT 18.030 3124.075 18.310 3124.445 ;
        RECT 18.100 3015.450 18.240 3124.075 ;
        RECT 18.040 3015.130 18.300 3015.450 ;
        RECT 296.800 3015.130 297.060 3015.450 ;
        RECT 296.860 3009.525 297.000 3015.130 ;
        RECT 296.790 3009.155 297.070 3009.525 ;
      LAYER via2 ;
        RECT 18.030 3124.120 18.310 3124.400 ;
        RECT 296.790 3009.200 297.070 3009.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 18.005 3124.410 18.335 3124.425 ;
        RECT -4.800 3124.110 18.335 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 18.005 3124.095 18.335 3124.110 ;
        RECT 296.765 3009.490 297.095 3009.505 ;
        RECT 310.000 3009.490 314.000 3009.880 ;
        RECT 296.765 3009.280 314.000 3009.490 ;
        RECT 296.765 3009.190 310.500 3009.280 ;
        RECT 296.765 3009.175 297.095 3009.190 ;
=======
        RECT -4.800 3123.660 0.300 3124.860 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2801.160 17.410 2801.220 ;
        RECT 296.770 2801.160 297.090 2801.220 ;
        RECT 17.090 2801.020 297.090 2801.160 ;
        RECT 17.090 2800.960 17.410 2801.020 ;
        RECT 296.770 2800.960 297.090 2801.020 ;
      LAYER via ;
        RECT 17.120 2800.960 17.380 2801.220 ;
        RECT 296.800 2800.960 297.060 2801.220 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2801.250 17.320 2836.435 ;
        RECT 17.120 2800.930 17.380 2801.250 ;
        RECT 296.800 2800.930 297.060 2801.250 ;
        RECT 296.860 2795.325 297.000 2800.930 ;
        RECT 296.790 2794.955 297.070 2795.325 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
        RECT 296.790 2795.000 297.070 2795.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
        RECT 296.765 2795.290 297.095 2795.305 ;
        RECT 310.000 2795.290 314.000 2795.680 ;
        RECT 296.765 2795.080 314.000 2795.290 ;
        RECT 296.765 2794.990 310.500 2795.080 ;
        RECT 296.765 2794.975 297.095 2794.990 ;
=======
        RECT -4.800 2836.020 0.300 2837.220 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2580.840 17.410 2580.900 ;
        RECT 296.770 2580.840 297.090 2580.900 ;
        RECT 17.090 2580.700 297.090 2580.840 ;
        RECT 17.090 2580.640 17.410 2580.700 ;
        RECT 296.770 2580.640 297.090 2580.700 ;
      LAYER via ;
        RECT 17.120 2580.640 17.380 2580.900 ;
        RECT 296.800 2580.640 297.060 2580.900 ;
      LAYER met2 ;
        RECT 17.120 2580.610 17.380 2580.930 ;
        RECT 296.790 2580.755 297.070 2581.125 ;
        RECT 296.800 2580.610 297.060 2580.755 ;
        RECT 17.180 2549.845 17.320 2580.610 ;
        RECT 17.110 2549.475 17.390 2549.845 ;
      LAYER via2 ;
        RECT 296.790 2580.800 297.070 2581.080 ;
        RECT 17.110 2549.520 17.390 2549.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2581.090 297.095 2581.105 ;
        RECT 310.000 2581.090 314.000 2581.480 ;
        RECT 296.765 2580.880 314.000 2581.090 ;
        RECT 296.765 2580.790 310.500 2580.880 ;
        RECT 296.765 2580.775 297.095 2580.790 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 17.085 2549.810 17.415 2549.825 ;
        RECT -4.800 2549.510 17.415 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 17.085 2549.495 17.415 2549.510 ;
=======
        RECT -4.800 2549.060 0.300 2550.260 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2366.980 17.410 2367.040 ;
        RECT 296.770 2366.980 297.090 2367.040 ;
        RECT 17.090 2366.840 297.090 2366.980 ;
        RECT 17.090 2366.780 17.410 2366.840 ;
        RECT 296.770 2366.780 297.090 2366.840 ;
      LAYER via ;
        RECT 17.120 2366.780 17.380 2367.040 ;
        RECT 296.800 2366.780 297.060 2367.040 ;
      LAYER met2 ;
        RECT 17.120 2366.750 17.380 2367.070 ;
        RECT 296.800 2366.925 297.060 2367.070 ;
        RECT 17.180 2262.205 17.320 2366.750 ;
        RECT 296.790 2366.555 297.070 2366.925 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
      LAYER via2 ;
        RECT 296.790 2366.600 297.070 2366.880 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2366.890 297.095 2366.905 ;
        RECT 310.000 2366.890 314.000 2367.280 ;
        RECT 296.765 2366.680 314.000 2366.890 ;
        RECT 296.765 2366.590 310.500 2366.680 ;
        RECT 296.765 2366.575 297.095 2366.590 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
=======
        RECT -4.800 2261.420 0.300 2262.620 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2145.980 17.870 2146.040 ;
        RECT 296.770 2145.980 297.090 2146.040 ;
        RECT 17.550 2145.840 297.090 2145.980 ;
        RECT 17.550 2145.780 17.870 2145.840 ;
        RECT 296.770 2145.780 297.090 2145.840 ;
      LAYER via ;
        RECT 17.580 2145.780 17.840 2146.040 ;
        RECT 296.800 2145.780 297.060 2146.040 ;
      LAYER met2 ;
        RECT 296.790 2152.355 297.070 2152.725 ;
        RECT 296.860 2146.070 297.000 2152.355 ;
        RECT 17.580 2145.750 17.840 2146.070 ;
        RECT 296.800 2145.750 297.060 2146.070 ;
        RECT 17.640 1975.245 17.780 2145.750 ;
        RECT 17.570 1974.875 17.850 1975.245 ;
      LAYER via2 ;
        RECT 296.790 2152.400 297.070 2152.680 ;
        RECT 17.570 1974.920 17.850 1975.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2152.690 297.095 2152.705 ;
        RECT 310.000 2152.690 314.000 2153.080 ;
        RECT 296.765 2152.480 314.000 2152.690 ;
        RECT 296.765 2152.390 310.500 2152.480 ;
        RECT 296.765 2152.375 297.095 2152.390 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 17.545 1975.210 17.875 1975.225 ;
        RECT -4.800 1974.910 17.875 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 17.545 1974.895 17.875 1974.910 ;
=======
        RECT -4.800 1974.460 0.300 1975.660 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2619.310 558.860 2619.630 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2619.310 558.720 2899.310 558.860 ;
        RECT 2619.310 558.660 2619.630 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2619.340 558.660 2619.600 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2619.330 693.075 2619.610 693.445 ;
        RECT 2619.400 558.950 2619.540 693.075 ;
        RECT 2619.340 558.630 2619.600 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2619.330 693.120 2619.610 693.400 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 693.410 2610.000 693.800 ;
        RECT 2619.305 693.410 2619.635 693.425 ;
        RECT 2606.000 693.200 2619.635 693.410 ;
        RECT 2609.580 693.110 2619.635 693.200 ;
        RECT 2619.305 693.095 2619.635 693.110 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
=======
        RECT 2919.700 556.660 2924.800 557.860 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 1690.380 18.330 1690.440 ;
        RECT 299.990 1690.380 300.310 1690.440 ;
        RECT 18.010 1690.240 300.310 1690.380 ;
        RECT 18.010 1690.180 18.330 1690.240 ;
        RECT 299.990 1690.180 300.310 1690.240 ;
      LAYER via ;
        RECT 18.040 1690.180 18.300 1690.440 ;
        RECT 300.020 1690.180 300.280 1690.440 ;
      LAYER met2 ;
        RECT 300.010 1938.155 300.290 1938.525 ;
        RECT 300.080 1690.470 300.220 1938.155 ;
        RECT 18.040 1690.150 18.300 1690.470 ;
        RECT 300.020 1690.150 300.280 1690.470 ;
        RECT 18.100 1687.605 18.240 1690.150 ;
        RECT 18.030 1687.235 18.310 1687.605 ;
      LAYER via2 ;
        RECT 300.010 1938.200 300.290 1938.480 ;
        RECT 18.030 1687.280 18.310 1687.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 299.985 1938.490 300.315 1938.505 ;
        RECT 310.000 1938.490 314.000 1938.880 ;
        RECT 299.985 1938.280 314.000 1938.490 ;
        RECT 299.985 1938.190 310.500 1938.280 ;
        RECT 299.985 1938.175 300.315 1938.190 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 18.005 1687.570 18.335 1687.585 ;
        RECT -4.800 1687.270 18.335 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 18.005 1687.255 18.335 1687.270 ;
=======
        RECT -4.800 1686.820 0.300 1688.020 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1476.520 15.570 1476.580 ;
        RECT 300.910 1476.520 301.230 1476.580 ;
        RECT 15.250 1476.380 301.230 1476.520 ;
        RECT 15.250 1476.320 15.570 1476.380 ;
        RECT 300.910 1476.320 301.230 1476.380 ;
      LAYER via ;
        RECT 15.280 1476.320 15.540 1476.580 ;
        RECT 300.940 1476.320 301.200 1476.580 ;
      LAYER met2 ;
        RECT 300.930 1723.275 301.210 1723.645 ;
        RECT 301.000 1476.610 301.140 1723.275 ;
        RECT 15.280 1476.290 15.540 1476.610 ;
        RECT 300.940 1476.290 301.200 1476.610 ;
        RECT 15.340 1472.045 15.480 1476.290 ;
        RECT 15.270 1471.675 15.550 1472.045 ;
      LAYER via2 ;
        RECT 300.930 1723.320 301.210 1723.600 ;
        RECT 15.270 1471.720 15.550 1472.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 300.905 1723.610 301.235 1723.625 ;
        RECT 310.000 1723.610 314.000 1724.000 ;
        RECT 300.905 1723.400 314.000 1723.610 ;
        RECT 300.905 1723.310 310.500 1723.400 ;
        RECT 300.905 1723.295 301.235 1723.310 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.245 1472.010 15.575 1472.025 ;
        RECT -4.800 1471.710 15.575 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.245 1471.695 15.575 1471.710 ;
=======
        RECT -4.800 1471.260 0.300 1472.460 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1262.660 16.030 1262.720 ;
        RECT 300.450 1262.660 300.770 1262.720 ;
        RECT 15.710 1262.520 300.770 1262.660 ;
        RECT 15.710 1262.460 16.030 1262.520 ;
        RECT 300.450 1262.460 300.770 1262.520 ;
      LAYER via ;
        RECT 15.740 1262.460 16.000 1262.720 ;
        RECT 300.480 1262.460 300.740 1262.720 ;
      LAYER met2 ;
        RECT 300.470 1509.075 300.750 1509.445 ;
        RECT 300.540 1262.750 300.680 1509.075 ;
        RECT 15.740 1262.430 16.000 1262.750 ;
        RECT 300.480 1262.430 300.740 1262.750 ;
        RECT 15.800 1256.485 15.940 1262.430 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
      LAYER via2 ;
        RECT 300.470 1509.120 300.750 1509.400 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 300.445 1509.410 300.775 1509.425 ;
        RECT 310.000 1509.410 314.000 1509.800 ;
        RECT 300.445 1509.200 314.000 1509.410 ;
        RECT 300.445 1509.110 310.500 1509.200 ;
        RECT 300.445 1509.095 300.775 1509.110 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
=======
        RECT -4.800 1255.700 0.300 1256.900 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1041.660 16.030 1041.720 ;
        RECT 299.990 1041.660 300.310 1041.720 ;
        RECT 15.710 1041.520 300.310 1041.660 ;
        RECT 15.710 1041.460 16.030 1041.520 ;
        RECT 299.990 1041.460 300.310 1041.520 ;
      LAYER via ;
        RECT 15.740 1041.460 16.000 1041.720 ;
        RECT 300.020 1041.460 300.280 1041.720 ;
      LAYER met2 ;
        RECT 300.010 1294.875 300.290 1295.245 ;
        RECT 300.080 1041.750 300.220 1294.875 ;
        RECT 15.740 1041.430 16.000 1041.750 ;
        RECT 300.020 1041.430 300.280 1041.750 ;
        RECT 15.800 1040.925 15.940 1041.430 ;
        RECT 15.730 1040.555 16.010 1040.925 ;
      LAYER via2 ;
        RECT 300.010 1294.920 300.290 1295.200 ;
        RECT 15.730 1040.600 16.010 1040.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 299.985 1295.210 300.315 1295.225 ;
        RECT 310.000 1295.210 314.000 1295.600 ;
        RECT 299.985 1295.000 314.000 1295.210 ;
        RECT 299.985 1294.910 310.500 1295.000 ;
        RECT 299.985 1294.895 300.315 1294.910 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 15.705 1040.890 16.035 1040.905 ;
        RECT -4.800 1040.590 16.035 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 15.705 1040.575 16.035 1040.590 ;
=======
        RECT -4.800 1040.140 0.300 1041.340 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 827.800 17.410 827.860 ;
        RECT 300.450 827.800 300.770 827.860 ;
        RECT 17.090 827.660 300.770 827.800 ;
        RECT 17.090 827.600 17.410 827.660 ;
        RECT 300.450 827.600 300.770 827.660 ;
      LAYER via ;
        RECT 17.120 827.600 17.380 827.860 ;
        RECT 300.480 827.600 300.740 827.860 ;
      LAYER met2 ;
        RECT 300.470 1080.675 300.750 1081.045 ;
        RECT 300.540 827.890 300.680 1080.675 ;
        RECT 17.120 827.570 17.380 827.890 ;
        RECT 300.480 827.570 300.740 827.890 ;
        RECT 17.180 825.365 17.320 827.570 ;
        RECT 17.110 824.995 17.390 825.365 ;
      LAYER via2 ;
        RECT 300.470 1080.720 300.750 1081.000 ;
        RECT 17.110 825.040 17.390 825.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 300.445 1081.010 300.775 1081.025 ;
        RECT 310.000 1081.010 314.000 1081.400 ;
        RECT 300.445 1080.800 314.000 1081.010 ;
        RECT 300.445 1080.710 310.500 1080.800 ;
        RECT 300.445 1080.695 300.775 1080.710 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.085 825.330 17.415 825.345 ;
        RECT -4.800 825.030 17.415 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.085 825.015 17.415 825.030 ;
=======
        RECT -4.800 824.580 0.300 825.780 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 14.790 613.940 15.110 614.000 ;
        RECT 299.990 613.940 300.310 614.000 ;
        RECT 14.790 613.800 300.310 613.940 ;
        RECT 14.790 613.740 15.110 613.800 ;
        RECT 299.990 613.740 300.310 613.800 ;
      LAYER via ;
        RECT 14.820 613.740 15.080 614.000 ;
        RECT 300.020 613.740 300.280 614.000 ;
      LAYER met2 ;
        RECT 300.010 866.475 300.290 866.845 ;
        RECT 300.080 614.030 300.220 866.475 ;
        RECT 14.820 613.710 15.080 614.030 ;
        RECT 300.020 613.710 300.280 614.030 ;
        RECT 14.880 610.485 15.020 613.710 ;
        RECT 14.810 610.115 15.090 610.485 ;
      LAYER via2 ;
        RECT 300.010 866.520 300.290 866.800 ;
        RECT 14.810 610.160 15.090 610.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 299.985 866.810 300.315 866.825 ;
        RECT 310.000 866.810 314.000 867.200 ;
        RECT 299.985 866.600 314.000 866.810 ;
        RECT 299.985 866.510 310.500 866.600 ;
        RECT 299.985 866.495 300.315 866.510 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 14.785 610.450 15.115 610.465 ;
        RECT -4.800 610.150 15.115 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 14.785 610.135 15.115 610.150 ;
=======
        RECT -4.800 609.700 0.300 610.900 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 400.080 15.570 400.140 ;
        RECT 300.450 400.080 300.770 400.140 ;
        RECT 15.250 399.940 300.770 400.080 ;
        RECT 15.250 399.880 15.570 399.940 ;
        RECT 300.450 399.880 300.770 399.940 ;
      LAYER via ;
        RECT 15.280 399.880 15.540 400.140 ;
        RECT 300.480 399.880 300.740 400.140 ;
      LAYER met2 ;
        RECT 300.470 652.275 300.750 652.645 ;
        RECT 300.540 400.170 300.680 652.275 ;
        RECT 15.280 399.850 15.540 400.170 ;
        RECT 300.480 399.850 300.740 400.170 ;
        RECT 15.340 394.925 15.480 399.850 ;
        RECT 15.270 394.555 15.550 394.925 ;
      LAYER via2 ;
        RECT 300.470 652.320 300.750 652.600 ;
        RECT 15.270 394.600 15.550 394.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 300.445 652.610 300.775 652.625 ;
        RECT 310.000 652.610 314.000 653.000 ;
        RECT 300.445 652.400 314.000 652.610 ;
        RECT 300.445 652.310 310.500 652.400 ;
        RECT 300.445 652.295 300.775 652.310 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 15.245 394.890 15.575 394.905 ;
        RECT -4.800 394.590 15.575 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 15.245 394.575 15.575 394.590 ;
=======
        RECT -4.800 394.140 0.300 395.340 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 179.420 16.950 179.480 ;
        RECT 299.990 179.420 300.310 179.480 ;
        RECT 16.630 179.280 300.310 179.420 ;
        RECT 16.630 179.220 16.950 179.280 ;
        RECT 299.990 179.220 300.310 179.280 ;
      LAYER via ;
        RECT 16.660 179.220 16.920 179.480 ;
        RECT 300.020 179.220 300.280 179.480 ;
      LAYER met2 ;
        RECT 300.010 438.075 300.290 438.445 ;
        RECT 300.080 179.510 300.220 438.075 ;
        RECT 16.660 179.365 16.920 179.510 ;
        RECT 16.650 178.995 16.930 179.365 ;
        RECT 300.020 179.190 300.280 179.510 ;
      LAYER via2 ;
        RECT 300.010 438.120 300.290 438.400 ;
        RECT 16.650 179.040 16.930 179.320 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 299.985 438.410 300.315 438.425 ;
        RECT 310.000 438.410 314.000 438.800 ;
        RECT 299.985 438.200 314.000 438.410 ;
        RECT 299.985 438.110 310.500 438.200 ;
        RECT 299.985 438.095 300.315 438.110 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 16.625 179.330 16.955 179.345 ;
        RECT -4.800 179.030 16.955 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 16.625 179.015 16.955 179.030 ;
=======
        RECT -4.800 178.580 0.300 179.780 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2619.310 793.460 2619.630 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2619.310 793.320 2899.310 793.460 ;
        RECT 2619.310 793.260 2619.630 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2619.340 793.260 2619.600 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2619.330 892.995 2619.610 893.365 ;
        RECT 2619.400 793.550 2619.540 892.995 ;
        RECT 2619.340 793.230 2619.600 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2619.330 893.040 2619.610 893.320 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 893.330 2610.000 893.720 ;
        RECT 2619.305 893.330 2619.635 893.345 ;
        RECT 2606.000 893.120 2619.635 893.330 ;
        RECT 2609.580 893.030 2619.635 893.120 ;
        RECT 2619.305 893.015 2619.635 893.030 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
=======
        RECT 2919.700 791.260 2924.800 792.460 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2619.310 1028.060 2619.630 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2619.310 1027.920 2899.310 1028.060 ;
        RECT 2619.310 1027.860 2619.630 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2619.340 1027.860 2619.600 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2619.330 1092.915 2619.610 1093.285 ;
        RECT 2619.400 1028.150 2619.540 1092.915 ;
        RECT 2619.340 1027.830 2619.600 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2619.330 1092.960 2619.610 1093.240 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1093.250 2610.000 1093.640 ;
        RECT 2619.305 1093.250 2619.635 1093.265 ;
        RECT 2606.000 1093.040 2619.635 1093.250 ;
        RECT 2609.580 1092.950 2619.635 1093.040 ;
        RECT 2619.305 1092.935 2619.635 1092.950 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
=======
        RECT 2919.700 1025.860 2924.800 1027.060 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1262.660 2618.710 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 2618.390 1262.520 2899.310 1262.660 ;
        RECT 2618.390 1262.460 2618.710 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 2618.420 1262.460 2618.680 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 2618.410 1292.835 2618.690 1293.205 ;
        RECT 2618.480 1262.750 2618.620 1292.835 ;
        RECT 2618.420 1262.430 2618.680 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2618.410 1292.880 2618.690 1293.160 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1293.170 2610.000 1293.560 ;
        RECT 2618.385 1293.170 2618.715 1293.185 ;
        RECT 2606.000 1292.960 2618.715 1293.170 ;
        RECT 2609.580 1292.870 2618.715 1292.960 ;
        RECT 2618.385 1292.855 2618.715 1292.870 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
=======
        RECT 2919.700 1260.460 2924.800 1261.660 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1493.860 2621.930 1493.920 ;
        RECT 2900.830 1493.860 2901.150 1493.920 ;
        RECT 2621.610 1493.720 2901.150 1493.860 ;
        RECT 2621.610 1493.660 2621.930 1493.720 ;
        RECT 2900.830 1493.660 2901.150 1493.720 ;
      LAYER via ;
        RECT 2621.640 1493.660 2621.900 1493.920 ;
        RECT 2900.860 1493.660 2901.120 1493.920 ;
      LAYER met2 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
        RECT 2900.920 1493.950 2901.060 1495.475 ;
        RECT 2621.640 1493.630 2621.900 1493.950 ;
        RECT 2900.860 1493.630 2901.120 1493.950 ;
        RECT 2621.700 1493.125 2621.840 1493.630 ;
        RECT 2621.630 1492.755 2621.910 1493.125 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
        RECT 2621.630 1492.800 2621.910 1493.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2606.000 1493.090 2610.000 1493.480 ;
        RECT 2621.605 1493.090 2621.935 1493.105 ;
        RECT 2606.000 1492.880 2621.935 1493.090 ;
        RECT 2609.580 1492.790 2621.935 1492.880 ;
        RECT 2621.605 1492.775 2621.935 1492.790 ;
=======
        RECT 2919.700 1495.060 2924.800 1496.260 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1725.400 2619.170 1725.460 ;
        RECT 2900.830 1725.400 2901.150 1725.460 ;
        RECT 2618.850 1725.260 2901.150 1725.400 ;
        RECT 2618.850 1725.200 2619.170 1725.260 ;
        RECT 2900.830 1725.200 2901.150 1725.260 ;
      LAYER via ;
        RECT 2618.880 1725.200 2619.140 1725.460 ;
        RECT 2900.860 1725.200 2901.120 1725.460 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 2900.920 1725.490 2901.060 1730.075 ;
        RECT 2618.880 1725.170 2619.140 1725.490 ;
        RECT 2900.860 1725.170 2901.120 1725.490 ;
        RECT 2618.940 1693.045 2619.080 1725.170 ;
        RECT 2618.870 1692.675 2619.150 1693.045 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
        RECT 2618.870 1692.720 2619.150 1693.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2606.000 1693.010 2610.000 1693.400 ;
        RECT 2618.845 1693.010 2619.175 1693.025 ;
        RECT 2606.000 1692.800 2619.175 1693.010 ;
        RECT 2609.580 1692.710 2619.175 1692.800 ;
        RECT 2618.845 1692.695 2619.175 1692.710 ;
=======
        RECT 2919.700 1729.660 2924.800 1730.860 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1960.000 2618.710 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 2618.390 1959.860 2901.150 1960.000 ;
        RECT 2618.390 1959.800 2618.710 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
      LAYER via ;
        RECT 2618.420 1959.800 2618.680 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 2618.420 1959.770 2618.680 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 2618.480 1893.645 2618.620 1959.770 ;
        RECT 2618.410 1893.275 2618.690 1893.645 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
        RECT 2618.410 1893.320 2618.690 1893.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2606.000 1893.610 2610.000 1894.000 ;
        RECT 2618.385 1893.610 2618.715 1893.625 ;
        RECT 2606.000 1893.400 2618.715 1893.610 ;
        RECT 2609.580 1893.310 2618.715 1893.400 ;
        RECT 2618.385 1893.295 2618.715 1893.310 ;
=======
        RECT 2919.700 1964.260 2924.800 1965.460 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2194.600 2618.710 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2618.390 2194.460 2901.150 2194.600 ;
        RECT 2618.390 2194.400 2618.710 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
      LAYER via ;
        RECT 2618.420 2194.400 2618.680 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2618.420 2194.370 2618.680 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2618.480 2093.565 2618.620 2194.370 ;
        RECT 2618.410 2093.195 2618.690 2093.565 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2618.410 2093.240 2618.690 2093.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2606.000 2093.530 2610.000 2093.920 ;
        RECT 2618.385 2093.530 2618.715 2093.545 ;
        RECT 2606.000 2093.320 2618.715 2093.530 ;
        RECT 2609.580 2093.230 2618.715 2093.320 ;
        RECT 2618.385 2093.215 2618.715 2093.230 ;
=======
        RECT 2919.700 2198.860 2924.800 2200.060 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 206.960 2618.710 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2618.390 206.820 2901.150 206.960 ;
        RECT 2618.390 206.760 2618.710 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2618.420 206.760 2618.680 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2618.410 426.515 2618.690 426.885 ;
        RECT 2618.480 207.050 2618.620 426.515 ;
        RECT 2618.420 206.730 2618.680 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2618.410 426.560 2618.690 426.840 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 426.850 2610.000 427.240 ;
        RECT 2618.385 426.850 2618.715 426.865 ;
        RECT 2606.000 426.640 2618.715 426.850 ;
        RECT 2609.580 426.550 2618.715 426.640 ;
        RECT 2618.385 426.535 2618.715 426.550 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
=======
        RECT 2919.700 204.420 2924.800 205.620 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2546.500 2619.170 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2618.850 2546.360 2901.150 2546.500 ;
        RECT 2618.850 2546.300 2619.170 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
      LAYER via ;
        RECT 2618.880 2546.300 2619.140 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2618.880 2546.270 2619.140 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2618.940 2426.765 2619.080 2546.270 ;
        RECT 2618.870 2426.395 2619.150 2426.765 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2618.870 2426.440 2619.150 2426.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2606.000 2426.730 2610.000 2427.120 ;
        RECT 2618.845 2426.730 2619.175 2426.745 ;
        RECT 2606.000 2426.520 2619.175 2426.730 ;
        RECT 2609.580 2426.430 2619.175 2426.520 ;
        RECT 2618.845 2426.415 2619.175 2426.430 ;
=======
        RECT 2919.700 2551.100 2924.800 2552.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2781.100 2619.170 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2618.850 2780.960 2901.150 2781.100 ;
        RECT 2618.850 2780.900 2619.170 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 2618.880 2780.900 2619.140 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2618.880 2780.870 2619.140 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2618.940 2626.685 2619.080 2780.870 ;
        RECT 2618.870 2626.315 2619.150 2626.685 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2618.870 2626.360 2619.150 2626.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2606.000 2626.650 2610.000 2627.040 ;
        RECT 2618.845 2626.650 2619.175 2626.665 ;
        RECT 2606.000 2626.440 2619.175 2626.650 ;
        RECT 2609.580 2626.350 2619.175 2626.440 ;
        RECT 2618.845 2626.335 2619.175 2626.350 ;
=======
        RECT 2919.700 2785.700 2924.800 2786.900 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2615.630 2829.040 2615.950 2829.100 ;
        RECT 2902.210 2829.040 2902.530 2829.100 ;
        RECT 2615.630 2828.900 2902.530 2829.040 ;
        RECT 2615.630 2828.840 2615.950 2828.900 ;
        RECT 2902.210 2828.840 2902.530 2828.900 ;
      LAYER via ;
        RECT 2615.660 2828.840 2615.920 2829.100 ;
        RECT 2902.240 2828.840 2902.500 2829.100 ;
      LAYER met2 ;
        RECT 2902.230 3020.715 2902.510 3021.085 ;
        RECT 2902.300 2829.130 2902.440 3020.715 ;
        RECT 2615.660 2828.810 2615.920 2829.130 ;
        RECT 2902.240 2828.810 2902.500 2829.130 ;
        RECT 2615.720 2826.605 2615.860 2828.810 ;
        RECT 2615.650 2826.235 2615.930 2826.605 ;
      LAYER via2 ;
        RECT 2902.230 3020.760 2902.510 3021.040 ;
        RECT 2615.650 2826.280 2615.930 2826.560 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2902.205 3021.050 2902.535 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2902.205 3020.750 2924.800 3021.050 ;
        RECT 2902.205 3020.735 2902.535 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2606.000 2826.570 2610.000 2826.960 ;
        RECT 2615.625 2826.570 2615.955 2826.585 ;
        RECT 2606.000 2826.360 2615.955 2826.570 ;
        RECT 2609.580 2826.270 2615.955 2826.360 ;
        RECT 2615.625 2826.255 2615.955 2826.270 ;
=======
        RECT 2919.700 3020.300 2924.800 3021.500 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2615.630 3028.960 2615.950 3029.020 ;
        RECT 2902.210 3028.960 2902.530 3029.020 ;
        RECT 2615.630 3028.820 2902.530 3028.960 ;
        RECT 2615.630 3028.760 2615.950 3028.820 ;
        RECT 2902.210 3028.760 2902.530 3028.820 ;
      LAYER via ;
        RECT 2615.660 3028.760 2615.920 3029.020 ;
        RECT 2902.240 3028.760 2902.500 3029.020 ;
      LAYER met2 ;
        RECT 2902.230 3255.315 2902.510 3255.685 ;
        RECT 2902.300 3029.050 2902.440 3255.315 ;
        RECT 2615.660 3028.730 2615.920 3029.050 ;
        RECT 2902.240 3028.730 2902.500 3029.050 ;
        RECT 2615.720 3026.525 2615.860 3028.730 ;
        RECT 2615.650 3026.155 2615.930 3026.525 ;
      LAYER via2 ;
        RECT 2902.230 3255.360 2902.510 3255.640 ;
        RECT 2615.650 3026.200 2615.930 3026.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2902.205 3255.650 2902.535 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2902.205 3255.350 2924.800 3255.650 ;
        RECT 2902.205 3255.335 2902.535 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2606.000 3026.490 2610.000 3026.880 ;
        RECT 2615.625 3026.490 2615.955 3026.505 ;
        RECT 2606.000 3026.280 2615.955 3026.490 ;
        RECT 2609.580 3026.190 2615.955 3026.280 ;
        RECT 2615.625 3026.175 2615.955 3026.190 ;
=======
        RECT 2919.700 3254.900 2924.800 3256.100 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3484.900 2619.170 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2618.850 3484.760 2901.150 3484.900 ;
        RECT 2618.850 3484.700 2619.170 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 2618.880 3484.700 2619.140 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2618.880 3484.670 2619.140 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2618.940 3226.445 2619.080 3484.670 ;
        RECT 2618.870 3226.075 2619.150 3226.445 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2618.870 3226.120 2619.150 3226.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2606.000 3226.410 2610.000 3226.800 ;
        RECT 2618.845 3226.410 2619.175 3226.425 ;
        RECT 2606.000 3226.200 2619.175 3226.410 ;
        RECT 2609.580 3226.110 2619.175 3226.200 ;
        RECT 2618.845 3226.095 2619.175 3226.110 ;
=======
        RECT 2919.700 3489.500 2924.800 3490.700 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2400.810 3501.560 2401.130 3501.620 ;
        RECT 2635.870 3501.560 2636.190 3501.620 ;
        RECT 2400.810 3501.420 2636.190 3501.560 ;
        RECT 2400.810 3501.360 2401.130 3501.420 ;
        RECT 2635.870 3501.360 2636.190 3501.420 ;
        RECT 2396.670 3277.500 2396.990 3277.560 ;
        RECT 2400.810 3277.500 2401.130 3277.560 ;
        RECT 2396.670 3277.360 2401.130 3277.500 ;
        RECT 2396.670 3277.300 2396.990 3277.360 ;
        RECT 2400.810 3277.300 2401.130 3277.360 ;
      LAYER via ;
        RECT 2400.840 3501.360 2401.100 3501.620 ;
        RECT 2635.900 3501.360 2636.160 3501.620 ;
        RECT 2396.700 3277.300 2396.960 3277.560 ;
        RECT 2400.840 3277.300 2401.100 3277.560 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.650 2636.100 3517.600 ;
        RECT 2400.840 3501.330 2401.100 3501.650 ;
        RECT 2635.900 3501.330 2636.160 3501.650 ;
        RECT 2400.900 3277.590 2401.040 3501.330 ;
        RECT 2396.700 3277.270 2396.960 3277.590 ;
        RECT 2400.840 3277.270 2401.100 3277.590 ;
        RECT 2396.760 3260.000 2396.900 3277.270 ;
        RECT 2396.650 3256.000 2396.930 3260.000 ;
=======
        RECT 2635.750 3519.700 2636.310 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2145.510 3501.560 2145.830 3501.620 ;
        RECT 2311.570 3501.560 2311.890 3501.620 ;
        RECT 2145.510 3501.420 2311.890 3501.560 ;
        RECT 2145.510 3501.360 2145.830 3501.420 ;
        RECT 2311.570 3501.360 2311.890 3501.420 ;
        RECT 2140.910 3277.500 2141.230 3277.560 ;
        RECT 2145.510 3277.500 2145.830 3277.560 ;
        RECT 2140.910 3277.360 2145.830 3277.500 ;
        RECT 2140.910 3277.300 2141.230 3277.360 ;
        RECT 2145.510 3277.300 2145.830 3277.360 ;
      LAYER via ;
        RECT 2145.540 3501.360 2145.800 3501.620 ;
        RECT 2311.600 3501.360 2311.860 3501.620 ;
        RECT 2140.940 3277.300 2141.200 3277.560 ;
        RECT 2145.540 3277.300 2145.800 3277.560 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.650 2311.800 3517.600 ;
        RECT 2145.540 3501.330 2145.800 3501.650 ;
        RECT 2311.600 3501.330 2311.860 3501.650 ;
        RECT 2145.600 3277.590 2145.740 3501.330 ;
        RECT 2140.940 3277.270 2141.200 3277.590 ;
        RECT 2145.540 3277.270 2145.800 3277.590 ;
        RECT 2141.000 3260.000 2141.140 3277.270 ;
        RECT 2140.890 3256.000 2141.170 3260.000 ;
=======
        RECT 2311.450 3519.700 2312.010 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1890.210 3501.560 1890.530 3501.620 ;
        RECT 1987.270 3501.560 1987.590 3501.620 ;
        RECT 1890.210 3501.420 1987.590 3501.560 ;
        RECT 1890.210 3501.360 1890.530 3501.420 ;
        RECT 1987.270 3501.360 1987.590 3501.420 ;
        RECT 1885.610 3277.500 1885.930 3277.560 ;
        RECT 1890.210 3277.500 1890.530 3277.560 ;
        RECT 1885.610 3277.360 1890.530 3277.500 ;
        RECT 1885.610 3277.300 1885.930 3277.360 ;
        RECT 1890.210 3277.300 1890.530 3277.360 ;
      LAYER via ;
        RECT 1890.240 3501.360 1890.500 3501.620 ;
        RECT 1987.300 3501.360 1987.560 3501.620 ;
        RECT 1885.640 3277.300 1885.900 3277.560 ;
        RECT 1890.240 3277.300 1890.500 3277.560 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3501.650 1987.500 3517.600 ;
        RECT 1890.240 3501.330 1890.500 3501.650 ;
        RECT 1987.300 3501.330 1987.560 3501.650 ;
        RECT 1890.300 3277.590 1890.440 3501.330 ;
        RECT 1885.640 3277.270 1885.900 3277.590 ;
        RECT 1890.240 3277.270 1890.500 3277.590 ;
        RECT 1885.700 3260.000 1885.840 3277.270 ;
        RECT 1885.590 3256.000 1885.870 3260.000 ;
=======
        RECT 1987.150 3519.700 1987.710 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1634.910 3498.500 1635.230 3498.560 ;
        RECT 1662.510 3498.500 1662.830 3498.560 ;
        RECT 1634.910 3498.360 1662.830 3498.500 ;
        RECT 1634.910 3498.300 1635.230 3498.360 ;
        RECT 1662.510 3498.300 1662.830 3498.360 ;
        RECT 1629.850 3275.800 1630.170 3275.860 ;
        RECT 1634.910 3275.800 1635.230 3275.860 ;
        RECT 1629.850 3275.660 1635.230 3275.800 ;
        RECT 1629.850 3275.600 1630.170 3275.660 ;
        RECT 1634.910 3275.600 1635.230 3275.660 ;
      LAYER via ;
        RECT 1634.940 3498.300 1635.200 3498.560 ;
        RECT 1662.540 3498.300 1662.800 3498.560 ;
        RECT 1629.880 3275.600 1630.140 3275.860 ;
        RECT 1634.940 3275.600 1635.200 3275.860 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3498.590 1662.740 3517.600 ;
        RECT 1634.940 3498.270 1635.200 3498.590 ;
        RECT 1662.540 3498.270 1662.800 3498.590 ;
        RECT 1635.000 3275.890 1635.140 3498.270 ;
        RECT 1629.880 3275.570 1630.140 3275.890 ;
        RECT 1634.940 3275.570 1635.200 3275.890 ;
        RECT 1629.940 3260.000 1630.080 3275.570 ;
        RECT 1629.830 3256.000 1630.110 3260.000 ;
=======
        RECT 1662.390 3519.700 1662.950 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3274.100 1338.530 3274.160 ;
        RECT 1374.550 3274.100 1374.870 3274.160 ;
        RECT 1338.210 3273.960 1374.870 3274.100 ;
        RECT 1338.210 3273.900 1338.530 3273.960 ;
        RECT 1374.550 3273.900 1374.870 3273.960 ;
      LAYER via ;
        RECT 1338.240 3273.900 1338.500 3274.160 ;
        RECT 1374.580 3273.900 1374.840 3274.160 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3274.190 1338.440 3517.600 ;
        RECT 1338.240 3273.870 1338.500 3274.190 ;
        RECT 1374.580 3273.870 1374.840 3274.190 ;
        RECT 1374.640 3260.000 1374.780 3273.870 ;
        RECT 1374.530 3256.000 1374.810 3260.000 ;
=======
        RECT 1338.090 3519.700 1338.650 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 441.560 2618.710 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2618.390 441.420 2901.150 441.560 ;
        RECT 2618.390 441.360 2618.710 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2618.420 441.360 2618.680 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2618.410 626.435 2618.690 626.805 ;
        RECT 2618.480 441.650 2618.620 626.435 ;
        RECT 2618.420 441.330 2618.680 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2618.410 626.480 2618.690 626.760 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 626.770 2610.000 627.160 ;
        RECT 2618.385 626.770 2618.715 626.785 ;
        RECT 2606.000 626.560 2618.715 626.770 ;
        RECT 2609.580 626.470 2618.715 626.560 ;
        RECT 2618.385 626.455 2618.715 626.470 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
=======
        RECT 2919.700 439.020 2924.800 440.220 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3274.100 1014.230 3274.160 ;
        RECT 1118.790 3274.100 1119.110 3274.160 ;
        RECT 1013.910 3273.960 1119.110 3274.100 ;
        RECT 1013.910 3273.900 1014.230 3273.960 ;
        RECT 1118.790 3273.900 1119.110 3273.960 ;
      LAYER via ;
        RECT 1013.940 3273.900 1014.200 3274.160 ;
        RECT 1118.820 3273.900 1119.080 3274.160 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3274.190 1014.140 3517.600 ;
        RECT 1013.940 3273.870 1014.200 3274.190 ;
        RECT 1118.820 3273.870 1119.080 3274.190 ;
        RECT 1118.880 3260.000 1119.020 3273.870 ;
        RECT 1118.770 3256.000 1119.050 3260.000 ;
=======
        RECT 1013.790 3519.700 1014.350 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 689.225 3429.325 689.395 3477.435 ;
      LAYER mcon ;
        RECT 689.225 3477.265 689.395 3477.435 ;
      LAYER met1 ;
        RECT 688.690 3491.360 689.010 3491.420 ;
        RECT 689.610 3491.360 689.930 3491.420 ;
        RECT 688.690 3491.220 689.930 3491.360 ;
        RECT 688.690 3491.160 689.010 3491.220 ;
        RECT 689.610 3491.160 689.930 3491.220 ;
        RECT 689.165 3477.420 689.455 3477.465 ;
        RECT 689.610 3477.420 689.930 3477.480 ;
        RECT 689.165 3477.280 689.930 3477.420 ;
        RECT 689.165 3477.235 689.455 3477.280 ;
        RECT 689.610 3477.220 689.930 3477.280 ;
        RECT 689.150 3429.480 689.470 3429.540 ;
        RECT 688.955 3429.340 689.470 3429.480 ;
        RECT 689.150 3429.280 689.470 3429.340 ;
        RECT 689.150 3395.140 689.470 3395.200 ;
        RECT 688.780 3395.000 689.470 3395.140 ;
        RECT 688.780 3394.860 688.920 3395.000 ;
        RECT 689.150 3394.940 689.470 3395.000 ;
        RECT 688.690 3394.600 689.010 3394.860 ;
        RECT 688.690 3367.600 689.010 3367.660 ;
        RECT 689.610 3367.600 689.930 3367.660 ;
        RECT 688.690 3367.460 689.930 3367.600 ;
        RECT 688.690 3367.400 689.010 3367.460 ;
        RECT 689.610 3367.400 689.930 3367.460 ;
        RECT 688.690 3274.780 689.010 3274.840 ;
        RECT 863.490 3274.780 863.810 3274.840 ;
        RECT 688.690 3274.640 863.810 3274.780 ;
        RECT 688.690 3274.580 689.010 3274.640 ;
        RECT 863.490 3274.580 863.810 3274.640 ;
      LAYER via ;
        RECT 688.720 3491.160 688.980 3491.420 ;
        RECT 689.640 3491.160 689.900 3491.420 ;
        RECT 689.640 3477.220 689.900 3477.480 ;
        RECT 689.180 3429.280 689.440 3429.540 ;
        RECT 689.180 3394.940 689.440 3395.200 ;
        RECT 688.720 3394.600 688.980 3394.860 ;
        RECT 688.720 3367.400 688.980 3367.660 ;
        RECT 689.640 3367.400 689.900 3367.660 ;
        RECT 688.720 3274.580 688.980 3274.840 ;
        RECT 863.520 3274.580 863.780 3274.840 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.780 3517.230 689.380 3517.370 ;
        RECT 688.780 3491.450 688.920 3517.230 ;
        RECT 688.720 3491.130 688.980 3491.450 ;
        RECT 689.640 3491.130 689.900 3491.450 ;
        RECT 689.700 3477.510 689.840 3491.130 ;
        RECT 689.640 3477.190 689.900 3477.510 ;
        RECT 689.180 3429.250 689.440 3429.570 ;
        RECT 689.240 3395.230 689.380 3429.250 ;
        RECT 689.180 3394.910 689.440 3395.230 ;
        RECT 688.720 3394.570 688.980 3394.890 ;
        RECT 688.780 3367.690 688.920 3394.570 ;
        RECT 688.720 3367.370 688.980 3367.690 ;
        RECT 689.640 3367.370 689.900 3367.690 ;
        RECT 689.700 3318.810 689.840 3367.370 ;
        RECT 688.780 3318.670 689.840 3318.810 ;
        RECT 688.780 3274.870 688.920 3318.670 ;
        RECT 688.720 3274.550 688.980 3274.870 ;
        RECT 863.520 3274.550 863.780 3274.870 ;
        RECT 863.580 3260.000 863.720 3274.550 ;
        RECT 863.470 3256.000 863.750 3260.000 ;
=======
        RECT 689.030 3519.700 689.590 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 362.625 3416.065 362.795 3463.835 ;
        RECT 363.545 3394.305 363.715 3415.555 ;
        RECT 364.005 3284.485 364.175 3332.595 ;
      LAYER mcon ;
        RECT 362.625 3463.665 362.795 3463.835 ;
        RECT 363.545 3415.385 363.715 3415.555 ;
        RECT 364.005 3332.425 364.175 3332.595 ;
      LAYER met1 ;
        RECT 362.565 3463.820 362.855 3463.865 ;
        RECT 363.470 3463.820 363.790 3463.880 ;
        RECT 362.565 3463.680 363.790 3463.820 ;
        RECT 362.565 3463.635 362.855 3463.680 ;
        RECT 363.470 3463.620 363.790 3463.680 ;
        RECT 362.550 3416.220 362.870 3416.280 ;
        RECT 362.355 3416.080 362.870 3416.220 ;
        RECT 362.550 3416.020 362.870 3416.080 ;
        RECT 362.550 3415.540 362.870 3415.600 ;
        RECT 363.485 3415.540 363.775 3415.585 ;
        RECT 362.550 3415.400 363.775 3415.540 ;
        RECT 362.550 3415.340 362.870 3415.400 ;
        RECT 363.485 3415.355 363.775 3415.400 ;
        RECT 363.470 3394.460 363.790 3394.520 ;
        RECT 363.275 3394.320 363.790 3394.460 ;
        RECT 363.470 3394.260 363.790 3394.320 ;
        RECT 363.470 3346.520 363.790 3346.580 ;
        RECT 364.390 3346.520 364.710 3346.580 ;
        RECT 363.470 3346.380 364.710 3346.520 ;
        RECT 363.470 3346.320 363.790 3346.380 ;
        RECT 364.390 3346.320 364.710 3346.380 ;
        RECT 363.945 3332.580 364.235 3332.625 ;
        RECT 364.390 3332.580 364.710 3332.640 ;
        RECT 363.945 3332.440 364.710 3332.580 ;
        RECT 363.945 3332.395 364.235 3332.440 ;
        RECT 364.390 3332.380 364.710 3332.440 ;
        RECT 363.930 3284.640 364.250 3284.700 ;
        RECT 363.735 3284.500 364.250 3284.640 ;
        RECT 363.930 3284.440 364.250 3284.500 ;
        RECT 363.930 3274.780 364.250 3274.840 ;
        RECT 607.730 3274.780 608.050 3274.840 ;
        RECT 363.930 3274.640 608.050 3274.780 ;
        RECT 363.930 3274.580 364.250 3274.640 ;
        RECT 607.730 3274.580 608.050 3274.640 ;
      LAYER via ;
        RECT 363.500 3463.620 363.760 3463.880 ;
        RECT 362.580 3416.020 362.840 3416.280 ;
        RECT 362.580 3415.340 362.840 3415.600 ;
        RECT 363.500 3394.260 363.760 3394.520 ;
        RECT 363.500 3346.320 363.760 3346.580 ;
        RECT 364.420 3346.320 364.680 3346.580 ;
        RECT 364.420 3332.380 364.680 3332.640 ;
        RECT 363.960 3284.440 364.220 3284.700 ;
        RECT 363.960 3274.580 364.220 3274.840 ;
        RECT 607.760 3274.580 608.020 3274.840 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3463.910 363.700 3491.390 ;
        RECT 363.500 3463.590 363.760 3463.910 ;
        RECT 362.580 3415.990 362.840 3416.310 ;
        RECT 362.640 3415.630 362.780 3415.990 ;
        RECT 362.580 3415.310 362.840 3415.630 ;
        RECT 363.500 3394.230 363.760 3394.550 ;
        RECT 363.560 3346.610 363.700 3394.230 ;
        RECT 363.500 3346.290 363.760 3346.610 ;
        RECT 364.420 3346.290 364.680 3346.610 ;
        RECT 364.480 3332.670 364.620 3346.290 ;
        RECT 364.420 3332.350 364.680 3332.670 ;
        RECT 363.960 3284.410 364.220 3284.730 ;
        RECT 364.020 3274.870 364.160 3284.410 ;
        RECT 363.960 3274.550 364.220 3274.870 ;
        RECT 607.760 3274.550 608.020 3274.870 ;
        RECT 607.820 3260.000 607.960 3274.550 ;
        RECT 607.710 3256.000 607.990 3260.000 ;
=======
        RECT 364.730 3519.700 365.290 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3274.780 40.410 3274.840 ;
        RECT 352.430 3274.780 352.750 3274.840 ;
        RECT 40.090 3274.640 352.750 3274.780 ;
        RECT 40.090 3274.580 40.410 3274.640 ;
        RECT 352.430 3274.580 352.750 3274.640 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3274.580 40.380 3274.840 ;
        RECT 352.460 3274.580 352.720 3274.840 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3274.870 40.320 3318.670 ;
        RECT 40.120 3274.550 40.380 3274.870 ;
        RECT 352.460 3274.550 352.720 3274.870 ;
        RECT 352.520 3260.000 352.660 3274.550 ;
        RECT 352.410 3256.000 352.690 3260.000 ;
=======
        RECT 40.430 3519.700 40.990 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 3084.040 17.870 3084.100 ;
        RECT 296.770 3084.040 297.090 3084.100 ;
        RECT 17.550 3083.900 297.090 3084.040 ;
        RECT 17.550 3083.840 17.870 3083.900 ;
        RECT 296.770 3083.840 297.090 3083.900 ;
      LAYER via ;
        RECT 17.580 3083.840 17.840 3084.100 ;
        RECT 296.800 3083.840 297.060 3084.100 ;
      LAYER met2 ;
        RECT 17.570 3267.555 17.850 3267.925 ;
        RECT 17.640 3084.130 17.780 3267.555 ;
        RECT 17.580 3083.810 17.840 3084.130 ;
        RECT 296.800 3083.810 297.060 3084.130 ;
        RECT 296.860 3080.925 297.000 3083.810 ;
        RECT 296.790 3080.555 297.070 3080.925 ;
      LAYER via2 ;
        RECT 17.570 3267.600 17.850 3267.880 ;
        RECT 296.790 3080.600 297.070 3080.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 17.545 3267.890 17.875 3267.905 ;
        RECT -4.800 3267.590 17.875 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 17.545 3267.575 17.875 3267.590 ;
        RECT 296.765 3080.890 297.095 3080.905 ;
        RECT 310.000 3080.890 314.000 3081.280 ;
        RECT 296.765 3080.680 314.000 3080.890 ;
        RECT 296.765 3080.590 310.500 3080.680 ;
        RECT 296.765 3080.575 297.095 3080.590 ;
=======
        RECT -4.800 3267.140 0.300 3268.340 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2870.180 17.870 2870.240 ;
        RECT 296.770 2870.180 297.090 2870.240 ;
        RECT 17.550 2870.040 297.090 2870.180 ;
        RECT 17.550 2869.980 17.870 2870.040 ;
        RECT 296.770 2869.980 297.090 2870.040 ;
      LAYER via ;
        RECT 17.580 2869.980 17.840 2870.240 ;
        RECT 296.800 2869.980 297.060 2870.240 ;
      LAYER met2 ;
        RECT 17.570 2979.915 17.850 2980.285 ;
        RECT 17.640 2870.270 17.780 2979.915 ;
        RECT 17.580 2869.950 17.840 2870.270 ;
        RECT 296.800 2869.950 297.060 2870.270 ;
        RECT 296.860 2866.725 297.000 2869.950 ;
        RECT 296.790 2866.355 297.070 2866.725 ;
      LAYER via2 ;
        RECT 17.570 2979.960 17.850 2980.240 ;
        RECT 296.790 2866.400 297.070 2866.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 17.545 2980.250 17.875 2980.265 ;
        RECT -4.800 2979.950 17.875 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 17.545 2979.935 17.875 2979.950 ;
        RECT 296.765 2866.690 297.095 2866.705 ;
        RECT 310.000 2866.690 314.000 2867.080 ;
        RECT 296.765 2866.480 314.000 2866.690 ;
        RECT 296.765 2866.390 310.500 2866.480 ;
        RECT 296.765 2866.375 297.095 2866.390 ;
=======
        RECT -4.800 2979.500 0.300 2980.700 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2656.320 17.410 2656.380 ;
        RECT 296.770 2656.320 297.090 2656.380 ;
        RECT 17.090 2656.180 297.090 2656.320 ;
        RECT 17.090 2656.120 17.410 2656.180 ;
        RECT 296.770 2656.120 297.090 2656.180 ;
      LAYER via ;
        RECT 17.120 2656.120 17.380 2656.380 ;
        RECT 296.800 2656.120 297.060 2656.380 ;
      LAYER met2 ;
        RECT 17.110 2692.955 17.390 2693.325 ;
        RECT 17.180 2656.410 17.320 2692.955 ;
        RECT 17.120 2656.090 17.380 2656.410 ;
        RECT 296.800 2656.090 297.060 2656.410 ;
        RECT 296.860 2652.525 297.000 2656.090 ;
        RECT 296.790 2652.155 297.070 2652.525 ;
      LAYER via2 ;
        RECT 17.110 2693.000 17.390 2693.280 ;
        RECT 296.790 2652.200 297.070 2652.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.085 2693.290 17.415 2693.305 ;
        RECT -4.800 2692.990 17.415 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.085 2692.975 17.415 2692.990 ;
        RECT 296.765 2652.490 297.095 2652.505 ;
        RECT 310.000 2652.490 314.000 2652.880 ;
        RECT 296.765 2652.280 314.000 2652.490 ;
        RECT 296.765 2652.190 310.500 2652.280 ;
        RECT 296.765 2652.175 297.095 2652.190 ;
=======
        RECT -4.800 2692.540 0.300 2693.740 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2436.000 17.410 2436.060 ;
        RECT 296.770 2436.000 297.090 2436.060 ;
        RECT 17.090 2435.860 297.090 2436.000 ;
        RECT 17.090 2435.800 17.410 2435.860 ;
        RECT 296.770 2435.800 297.090 2435.860 ;
      LAYER via ;
        RECT 17.120 2435.800 17.380 2436.060 ;
        RECT 296.800 2435.800 297.060 2436.060 ;
      LAYER met2 ;
        RECT 296.790 2437.955 297.070 2438.325 ;
        RECT 296.860 2436.090 297.000 2437.955 ;
        RECT 17.120 2435.770 17.380 2436.090 ;
        RECT 296.800 2435.770 297.060 2436.090 ;
        RECT 17.180 2405.685 17.320 2435.770 ;
        RECT 17.110 2405.315 17.390 2405.685 ;
      LAYER via2 ;
        RECT 296.790 2438.000 297.070 2438.280 ;
        RECT 17.110 2405.360 17.390 2405.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2438.290 297.095 2438.305 ;
        RECT 310.000 2438.290 314.000 2438.680 ;
        RECT 296.765 2438.080 314.000 2438.290 ;
        RECT 296.765 2437.990 310.500 2438.080 ;
        RECT 296.765 2437.975 297.095 2437.990 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 17.085 2405.650 17.415 2405.665 ;
        RECT -4.800 2405.350 17.415 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 17.085 2405.335 17.415 2405.350 ;
=======
        RECT -4.800 2404.900 0.300 2406.100 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2222.140 17.410 2222.200 ;
        RECT 296.770 2222.140 297.090 2222.200 ;
        RECT 17.090 2222.000 297.090 2222.140 ;
        RECT 17.090 2221.940 17.410 2222.000 ;
        RECT 296.770 2221.940 297.090 2222.000 ;
      LAYER via ;
        RECT 17.120 2221.940 17.380 2222.200 ;
        RECT 296.800 2221.940 297.060 2222.200 ;
      LAYER met2 ;
        RECT 296.790 2223.755 297.070 2224.125 ;
        RECT 296.860 2222.230 297.000 2223.755 ;
        RECT 17.120 2221.910 17.380 2222.230 ;
        RECT 296.800 2221.910 297.060 2222.230 ;
        RECT 17.180 2118.725 17.320 2221.910 ;
        RECT 17.110 2118.355 17.390 2118.725 ;
      LAYER via2 ;
        RECT 296.790 2223.800 297.070 2224.080 ;
        RECT 17.110 2118.400 17.390 2118.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2224.090 297.095 2224.105 ;
        RECT 310.000 2224.090 314.000 2224.480 ;
        RECT 296.765 2223.880 314.000 2224.090 ;
        RECT 296.765 2223.790 310.500 2223.880 ;
        RECT 296.765 2223.775 297.095 2223.790 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 17.085 2118.690 17.415 2118.705 ;
        RECT -4.800 2118.390 17.415 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 17.085 2118.375 17.415 2118.390 ;
=======
        RECT -4.800 2117.940 0.300 2119.140 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 2008.280 18.330 2008.340 ;
        RECT 296.770 2008.280 297.090 2008.340 ;
        RECT 18.010 2008.140 297.090 2008.280 ;
        RECT 18.010 2008.080 18.330 2008.140 ;
        RECT 296.770 2008.080 297.090 2008.140 ;
      LAYER via ;
        RECT 18.040 2008.080 18.300 2008.340 ;
        RECT 296.800 2008.080 297.060 2008.340 ;
      LAYER met2 ;
        RECT 296.790 2009.555 297.070 2009.925 ;
        RECT 296.860 2008.370 297.000 2009.555 ;
        RECT 18.040 2008.050 18.300 2008.370 ;
        RECT 296.800 2008.050 297.060 2008.370 ;
        RECT 18.100 1831.085 18.240 2008.050 ;
        RECT 18.030 1830.715 18.310 1831.085 ;
      LAYER via2 ;
        RECT 296.790 2009.600 297.070 2009.880 ;
        RECT 18.030 1830.760 18.310 1831.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2009.890 297.095 2009.905 ;
        RECT 310.000 2009.890 314.000 2010.280 ;
        RECT 296.765 2009.680 314.000 2009.890 ;
        RECT 296.765 2009.590 310.500 2009.680 ;
        RECT 296.765 2009.575 297.095 2009.590 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 18.005 1831.050 18.335 1831.065 ;
        RECT -4.800 1830.750 18.335 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 18.005 1830.735 18.335 1830.750 ;
=======
        RECT -4.800 1830.300 0.300 1831.500 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 676.160 2618.710 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2618.390 676.020 2901.150 676.160 ;
        RECT 2618.390 675.960 2618.710 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2618.420 675.960 2618.680 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2618.410 826.355 2618.690 826.725 ;
        RECT 2618.480 676.250 2618.620 826.355 ;
        RECT 2618.420 675.930 2618.680 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2618.410 826.400 2618.690 826.680 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 826.690 2610.000 827.080 ;
        RECT 2618.385 826.690 2618.715 826.705 ;
        RECT 2606.000 826.480 2618.715 826.690 ;
        RECT 2609.580 826.390 2618.715 826.480 ;
        RECT 2618.385 826.375 2618.715 826.390 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
=======
        RECT 2919.700 673.620 2924.800 674.820 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1794.080 17.410 1794.140 ;
        RECT 296.770 1794.080 297.090 1794.140 ;
        RECT 17.090 1793.940 297.090 1794.080 ;
        RECT 17.090 1793.880 17.410 1793.940 ;
        RECT 296.770 1793.880 297.090 1793.940 ;
      LAYER via ;
        RECT 17.120 1793.880 17.380 1794.140 ;
        RECT 296.800 1793.880 297.060 1794.140 ;
      LAYER met2 ;
        RECT 296.790 1795.355 297.070 1795.725 ;
        RECT 296.860 1794.170 297.000 1795.355 ;
        RECT 17.120 1793.850 17.380 1794.170 ;
        RECT 296.800 1793.850 297.060 1794.170 ;
        RECT 17.180 1544.125 17.320 1793.850 ;
        RECT 17.110 1543.755 17.390 1544.125 ;
      LAYER via2 ;
        RECT 296.790 1795.400 297.070 1795.680 ;
        RECT 17.110 1543.800 17.390 1544.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1795.690 297.095 1795.705 ;
        RECT 310.000 1795.690 314.000 1796.080 ;
        RECT 296.765 1795.480 314.000 1795.690 ;
        RECT 296.765 1795.390 310.500 1795.480 ;
        RECT 296.765 1795.375 297.095 1795.390 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 17.085 1544.090 17.415 1544.105 ;
        RECT -4.800 1543.790 17.415 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 17.085 1543.775 17.415 1543.790 ;
=======
        RECT -4.800 1543.340 0.300 1544.540 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 1580.220 18.790 1580.280 ;
        RECT 296.770 1580.220 297.090 1580.280 ;
        RECT 18.470 1580.080 297.090 1580.220 ;
        RECT 18.470 1580.020 18.790 1580.080 ;
        RECT 296.770 1580.020 297.090 1580.080 ;
      LAYER via ;
        RECT 18.500 1580.020 18.760 1580.280 ;
        RECT 296.800 1580.020 297.060 1580.280 ;
      LAYER met2 ;
        RECT 296.790 1580.475 297.070 1580.845 ;
        RECT 296.860 1580.310 297.000 1580.475 ;
        RECT 18.500 1579.990 18.760 1580.310 ;
        RECT 296.800 1579.990 297.060 1580.310 ;
        RECT 18.560 1328.565 18.700 1579.990 ;
        RECT 18.490 1328.195 18.770 1328.565 ;
      LAYER via2 ;
        RECT 296.790 1580.520 297.070 1580.800 ;
        RECT 18.490 1328.240 18.770 1328.520 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1580.810 297.095 1580.825 ;
        RECT 310.000 1580.810 314.000 1581.200 ;
        RECT 296.765 1580.600 314.000 1580.810 ;
        RECT 296.765 1580.510 310.500 1580.600 ;
        RECT 296.765 1580.495 297.095 1580.510 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 18.465 1328.530 18.795 1328.545 ;
        RECT -4.800 1328.230 18.795 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 18.465 1328.215 18.795 1328.230 ;
=======
        RECT -4.800 1327.780 0.300 1328.980 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 1366.360 18.330 1366.420 ;
        RECT 296.770 1366.360 297.090 1366.420 ;
        RECT 18.010 1366.220 297.090 1366.360 ;
        RECT 18.010 1366.160 18.330 1366.220 ;
        RECT 296.770 1366.160 297.090 1366.220 ;
      LAYER via ;
        RECT 18.040 1366.160 18.300 1366.420 ;
        RECT 296.800 1366.160 297.060 1366.420 ;
      LAYER met2 ;
        RECT 18.040 1366.130 18.300 1366.450 ;
        RECT 296.790 1366.275 297.070 1366.645 ;
        RECT 296.800 1366.130 297.060 1366.275 ;
        RECT 18.100 1113.005 18.240 1366.130 ;
        RECT 18.030 1112.635 18.310 1113.005 ;
      LAYER via2 ;
        RECT 296.790 1366.320 297.070 1366.600 ;
        RECT 18.030 1112.680 18.310 1112.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1366.610 297.095 1366.625 ;
        RECT 310.000 1366.610 314.000 1367.000 ;
        RECT 296.765 1366.400 314.000 1366.610 ;
        RECT 296.765 1366.310 310.500 1366.400 ;
        RECT 296.765 1366.295 297.095 1366.310 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 18.005 1112.970 18.335 1112.985 ;
        RECT -4.800 1112.670 18.335 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 18.005 1112.655 18.335 1112.670 ;
=======
        RECT -4.800 1112.220 0.300 1113.420 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 1145.700 18.790 1145.760 ;
        RECT 296.770 1145.700 297.090 1145.760 ;
        RECT 18.470 1145.560 297.090 1145.700 ;
        RECT 18.470 1145.500 18.790 1145.560 ;
        RECT 296.770 1145.500 297.090 1145.560 ;
      LAYER via ;
        RECT 18.500 1145.500 18.760 1145.760 ;
        RECT 296.800 1145.500 297.060 1145.760 ;
      LAYER met2 ;
        RECT 296.790 1152.075 297.070 1152.445 ;
        RECT 296.860 1145.790 297.000 1152.075 ;
        RECT 18.500 1145.470 18.760 1145.790 ;
        RECT 296.800 1145.470 297.060 1145.790 ;
        RECT 18.560 897.445 18.700 1145.470 ;
        RECT 18.490 897.075 18.770 897.445 ;
      LAYER via2 ;
        RECT 296.790 1152.120 297.070 1152.400 ;
        RECT 18.490 897.120 18.770 897.400 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1152.410 297.095 1152.425 ;
        RECT 310.000 1152.410 314.000 1152.800 ;
        RECT 296.765 1152.200 314.000 1152.410 ;
        RECT 296.765 1152.110 310.500 1152.200 ;
        RECT 296.765 1152.095 297.095 1152.110 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 18.465 897.410 18.795 897.425 ;
        RECT -4.800 897.110 18.795 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 18.465 897.095 18.795 897.110 ;
=======
        RECT -4.800 896.660 0.300 897.860 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 931.840 18.330 931.900 ;
        RECT 296.770 931.840 297.090 931.900 ;
        RECT 18.010 931.700 297.090 931.840 ;
        RECT 18.010 931.640 18.330 931.700 ;
        RECT 296.770 931.640 297.090 931.700 ;
      LAYER via ;
        RECT 18.040 931.640 18.300 931.900 ;
        RECT 296.800 931.640 297.060 931.900 ;
      LAYER met2 ;
        RECT 296.790 937.875 297.070 938.245 ;
        RECT 296.860 931.930 297.000 937.875 ;
        RECT 18.040 931.610 18.300 931.930 ;
        RECT 296.800 931.610 297.060 931.930 ;
        RECT 18.100 681.885 18.240 931.610 ;
        RECT 18.030 681.515 18.310 681.885 ;
      LAYER via2 ;
        RECT 296.790 937.920 297.070 938.200 ;
        RECT 18.030 681.560 18.310 681.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 938.210 297.095 938.225 ;
        RECT 310.000 938.210 314.000 938.600 ;
        RECT 296.765 938.000 314.000 938.210 ;
        RECT 296.765 937.910 310.500 938.000 ;
        RECT 296.765 937.895 297.095 937.910 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 18.005 681.850 18.335 681.865 ;
        RECT -4.800 681.550 18.335 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 18.005 681.535 18.335 681.550 ;
=======
        RECT -4.800 681.100 0.300 682.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 717.980 18.790 718.040 ;
        RECT 296.770 717.980 297.090 718.040 ;
        RECT 18.470 717.840 297.090 717.980 ;
        RECT 18.470 717.780 18.790 717.840 ;
        RECT 296.770 717.780 297.090 717.840 ;
      LAYER via ;
        RECT 18.500 717.780 18.760 718.040 ;
        RECT 296.800 717.780 297.060 718.040 ;
      LAYER met2 ;
        RECT 296.790 723.675 297.070 724.045 ;
        RECT 296.860 718.070 297.000 723.675 ;
        RECT 18.500 717.750 18.760 718.070 ;
        RECT 296.800 717.750 297.060 718.070 ;
        RECT 18.560 466.325 18.700 717.750 ;
        RECT 18.490 465.955 18.770 466.325 ;
      LAYER via2 ;
        RECT 296.790 723.720 297.070 724.000 ;
        RECT 18.490 466.000 18.770 466.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 724.010 297.095 724.025 ;
        RECT 310.000 724.010 314.000 724.400 ;
        RECT 296.765 723.800 314.000 724.010 ;
        RECT 296.765 723.710 310.500 723.800 ;
        RECT 296.765 723.695 297.095 723.710 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 18.465 466.290 18.795 466.305 ;
        RECT -4.800 465.990 18.795 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 18.465 465.975 18.795 465.990 ;
=======
        RECT -4.800 465.540 0.300 466.740 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 503.780 18.330 503.840 ;
        RECT 296.770 503.780 297.090 503.840 ;
        RECT 18.010 503.640 297.090 503.780 ;
        RECT 18.010 503.580 18.330 503.640 ;
        RECT 296.770 503.580 297.090 503.640 ;
      LAYER via ;
        RECT 18.040 503.580 18.300 503.840 ;
        RECT 296.800 503.580 297.060 503.840 ;
      LAYER met2 ;
        RECT 296.790 509.475 297.070 509.845 ;
        RECT 296.860 503.870 297.000 509.475 ;
        RECT 18.040 503.550 18.300 503.870 ;
        RECT 296.800 503.550 297.060 503.870 ;
        RECT 18.100 250.765 18.240 503.550 ;
        RECT 18.030 250.395 18.310 250.765 ;
      LAYER via2 ;
        RECT 296.790 509.520 297.070 509.800 ;
        RECT 18.030 250.440 18.310 250.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 509.810 297.095 509.825 ;
        RECT 310.000 509.810 314.000 510.200 ;
        RECT 296.765 509.600 314.000 509.810 ;
        RECT 296.765 509.510 310.500 509.600 ;
        RECT 296.765 509.495 297.095 509.510 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 18.005 250.730 18.335 250.745 ;
        RECT -4.800 250.430 18.335 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 18.005 250.415 18.335 250.430 ;
=======
        RECT -4.800 249.980 0.300 251.180 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 289.920 17.870 289.980 ;
        RECT 296.770 289.920 297.090 289.980 ;
        RECT 17.550 289.780 297.090 289.920 ;
        RECT 17.550 289.720 17.870 289.780 ;
        RECT 296.770 289.720 297.090 289.780 ;
      LAYER via ;
        RECT 17.580 289.720 17.840 289.980 ;
        RECT 296.800 289.720 297.060 289.980 ;
      LAYER met2 ;
        RECT 296.790 295.275 297.070 295.645 ;
        RECT 296.860 290.010 297.000 295.275 ;
        RECT 17.580 289.690 17.840 290.010 ;
        RECT 296.800 289.690 297.060 290.010 ;
        RECT 17.640 35.885 17.780 289.690 ;
        RECT 17.570 35.515 17.850 35.885 ;
      LAYER via2 ;
        RECT 296.790 295.320 297.070 295.600 ;
        RECT 17.570 35.560 17.850 35.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 295.610 297.095 295.625 ;
        RECT 310.000 295.610 314.000 296.000 ;
        RECT 296.765 295.400 314.000 295.610 ;
        RECT 296.765 295.310 310.500 295.400 ;
        RECT 296.765 295.295 297.095 295.310 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.545 35.850 17.875 35.865 ;
        RECT -4.800 35.550 17.875 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.545 35.535 17.875 35.550 ;
=======
        RECT -4.800 35.100 0.300 36.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 910.760 2618.710 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2618.390 910.620 2901.150 910.760 ;
        RECT 2618.390 910.560 2618.710 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2618.420 910.560 2618.680 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2618.410 1026.275 2618.690 1026.645 ;
        RECT 2618.480 910.850 2618.620 1026.275 ;
        RECT 2618.420 910.530 2618.680 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2618.410 1026.320 2618.690 1026.600 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1026.610 2610.000 1027.000 ;
        RECT 2618.385 1026.610 2618.715 1026.625 ;
        RECT 2606.000 1026.400 2618.715 1026.610 ;
        RECT 2609.580 1026.310 2618.715 1026.400 ;
        RECT 2618.385 1026.295 2618.715 1026.310 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
=======
        RECT 2919.700 908.900 2924.800 910.100 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1145.360 2618.710 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2618.390 1145.220 2901.150 1145.360 ;
        RECT 2618.390 1145.160 2618.710 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2618.420 1145.160 2618.680 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2618.410 1226.195 2618.690 1226.565 ;
        RECT 2618.480 1145.450 2618.620 1226.195 ;
        RECT 2618.420 1145.130 2618.680 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2618.410 1226.240 2618.690 1226.520 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1226.530 2610.000 1226.920 ;
        RECT 2618.385 1226.530 2618.715 1226.545 ;
        RECT 2606.000 1226.320 2618.715 1226.530 ;
        RECT 2609.580 1226.230 2618.715 1226.320 ;
        RECT 2618.385 1226.215 2618.715 1226.230 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
=======
        RECT 2919.700 1143.500 2924.800 1144.700 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1379.960 2618.710 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2618.390 1379.820 2901.150 1379.960 ;
        RECT 2618.390 1379.760 2618.710 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 2618.420 1379.760 2618.680 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 2618.410 1426.115 2618.690 1426.485 ;
        RECT 2618.480 1380.050 2618.620 1426.115 ;
        RECT 2618.420 1379.730 2618.680 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2618.410 1426.160 2618.690 1426.440 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1426.450 2610.000 1426.840 ;
        RECT 2618.385 1426.450 2618.715 1426.465 ;
        RECT 2606.000 1426.240 2618.715 1426.450 ;
        RECT 2609.580 1426.150 2618.715 1426.240 ;
        RECT 2618.385 1426.135 2618.715 1426.150 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
=======
        RECT 2919.700 1378.100 2924.800 1379.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1614.560 2621.930 1614.620 ;
        RECT 2900.830 1614.560 2901.150 1614.620 ;
        RECT 2621.610 1614.420 2901.150 1614.560 ;
        RECT 2621.610 1614.360 2621.930 1614.420 ;
        RECT 2900.830 1614.360 2901.150 1614.420 ;
      LAYER via ;
        RECT 2621.640 1614.360 2621.900 1614.620 ;
        RECT 2900.860 1614.360 2901.120 1614.620 ;
      LAYER met2 ;
        RECT 2621.630 1626.035 2621.910 1626.405 ;
        RECT 2621.700 1614.650 2621.840 1626.035 ;
        RECT 2621.640 1614.330 2621.900 1614.650 ;
        RECT 2900.860 1614.330 2901.120 1614.650 ;
        RECT 2900.920 1613.485 2901.060 1614.330 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2621.630 1626.080 2621.910 1626.360 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1626.370 2610.000 1626.760 ;
        RECT 2621.605 1626.370 2621.935 1626.385 ;
        RECT 2606.000 1626.160 2621.935 1626.370 ;
        RECT 2609.580 1626.070 2621.935 1626.160 ;
        RECT 2621.605 1626.055 2621.935 1626.070 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
=======
        RECT 2919.700 1612.700 2924.800 1613.900 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2621.150 1842.700 2621.470 1842.760 ;
        RECT 2900.830 1842.700 2901.150 1842.760 ;
        RECT 2621.150 1842.560 2901.150 1842.700 ;
        RECT 2621.150 1842.500 2621.470 1842.560 ;
        RECT 2900.830 1842.500 2901.150 1842.560 ;
      LAYER via ;
        RECT 2621.180 1842.500 2621.440 1842.760 ;
        RECT 2900.860 1842.500 2901.120 1842.760 ;
      LAYER met2 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
        RECT 2900.920 1842.790 2901.060 1847.715 ;
        RECT 2621.180 1842.470 2621.440 1842.790 ;
        RECT 2900.860 1842.470 2901.120 1842.790 ;
        RECT 2621.240 1827.005 2621.380 1842.470 ;
        RECT 2621.170 1826.635 2621.450 1827.005 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
        RECT 2621.170 1826.680 2621.450 1826.960 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2606.000 1826.970 2610.000 1827.360 ;
        RECT 2621.145 1826.970 2621.475 1826.985 ;
        RECT 2606.000 1826.760 2621.475 1826.970 ;
        RECT 2609.580 1826.670 2621.475 1826.760 ;
        RECT 2621.145 1826.655 2621.475 1826.670 ;
=======
        RECT 2919.700 1847.300 2924.800 1848.500 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2077.300 2618.710 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 2618.390 2077.160 2901.150 2077.300 ;
        RECT 2618.390 2077.100 2618.710 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
      LAYER via ;
        RECT 2618.420 2077.100 2618.680 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 2618.420 2077.070 2618.680 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 2618.480 2026.925 2618.620 2077.070 ;
        RECT 2618.410 2026.555 2618.690 2026.925 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
        RECT 2618.410 2026.600 2618.690 2026.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2606.000 2026.890 2610.000 2027.280 ;
        RECT 2618.385 2026.890 2618.715 2026.905 ;
        RECT 2606.000 2026.680 2618.715 2026.890 ;
        RECT 2609.580 2026.590 2618.715 2026.680 ;
        RECT 2618.385 2026.575 2618.715 2026.590 ;
=======
        RECT 2919.700 2081.900 2924.800 2083.100 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2311.900 2618.710 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2618.390 2311.760 2901.150 2311.900 ;
        RECT 2618.390 2311.700 2618.710 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
      LAYER via ;
        RECT 2618.420 2311.700 2618.680 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2618.420 2311.670 2618.680 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2618.480 2226.845 2618.620 2311.670 ;
        RECT 2618.410 2226.475 2618.690 2226.845 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2618.410 2226.520 2618.690 2226.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2606.000 2226.810 2610.000 2227.200 ;
        RECT 2618.385 2226.810 2618.715 2226.825 ;
        RECT 2606.000 2226.600 2618.715 2226.810 ;
        RECT 2609.580 2226.510 2618.715 2226.600 ;
        RECT 2618.385 2226.495 2618.715 2226.510 ;
=======
        RECT 2919.700 2316.500 2924.800 2317.700 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 151.540 2619.170 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2618.850 151.400 2901.150 151.540 ;
        RECT 2618.850 151.340 2619.170 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2618.880 151.340 2619.140 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2618.870 359.875 2619.150 360.245 ;
        RECT 2618.940 151.630 2619.080 359.875 ;
        RECT 2618.880 151.310 2619.140 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2618.870 359.920 2619.150 360.200 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 360.210 2610.000 360.600 ;
        RECT 2618.845 360.210 2619.175 360.225 ;
        RECT 2606.000 360.000 2619.175 360.210 ;
        RECT 2609.580 359.910 2619.175 360.000 ;
        RECT 2618.845 359.895 2619.175 359.910 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
=======
        RECT 2919.700 145.940 2924.800 147.140 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2491.080 2618.710 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 2618.390 2490.940 2901.150 2491.080 ;
        RECT 2618.390 2490.880 2618.710 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
      LAYER via ;
        RECT 2618.420 2490.880 2618.680 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 2618.420 2490.850 2618.680 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 2618.480 2360.125 2618.620 2490.850 ;
        RECT 2618.410 2359.755 2618.690 2360.125 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 2618.410 2359.800 2618.690 2360.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2606.000 2360.090 2610.000 2360.480 ;
        RECT 2618.385 2360.090 2618.715 2360.105 ;
        RECT 2606.000 2359.880 2618.715 2360.090 ;
        RECT 2609.580 2359.790 2618.715 2359.880 ;
        RECT 2618.385 2359.775 2618.715 2359.790 ;
=======
        RECT 2919.700 2492.620 2924.800 2493.820 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2617.470 2725.680 2617.790 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2617.470 2725.540 2901.150 2725.680 ;
        RECT 2617.470 2725.480 2617.790 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 2617.500 2725.480 2617.760 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2617.500 2725.450 2617.760 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 2617.560 2691.170 2617.700 2725.450 ;
        RECT 2617.560 2691.030 2618.620 2691.170 ;
        RECT 2618.480 2560.045 2618.620 2691.030 ;
        RECT 2618.410 2559.675 2618.690 2560.045 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 2618.410 2559.720 2618.690 2560.000 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2606.000 2560.010 2610.000 2560.400 ;
        RECT 2618.385 2560.010 2618.715 2560.025 ;
        RECT 2606.000 2559.800 2618.715 2560.010 ;
        RECT 2609.580 2559.710 2618.715 2559.800 ;
        RECT 2618.385 2559.695 2618.715 2559.710 ;
=======
        RECT 2919.700 2727.220 2924.800 2728.420 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2960.280 2618.710 2960.340 ;
        RECT 2898.990 2960.280 2899.310 2960.340 ;
        RECT 2618.390 2960.140 2899.310 2960.280 ;
        RECT 2618.390 2960.080 2618.710 2960.140 ;
        RECT 2898.990 2960.080 2899.310 2960.140 ;
      LAYER via ;
        RECT 2618.420 2960.080 2618.680 2960.340 ;
        RECT 2899.020 2960.080 2899.280 2960.340 ;
      LAYER met2 ;
        RECT 2899.010 2962.235 2899.290 2962.605 ;
        RECT 2899.080 2960.370 2899.220 2962.235 ;
        RECT 2618.420 2960.050 2618.680 2960.370 ;
        RECT 2899.020 2960.050 2899.280 2960.370 ;
        RECT 2618.480 2759.965 2618.620 2960.050 ;
        RECT 2618.410 2759.595 2618.690 2759.965 ;
      LAYER via2 ;
        RECT 2899.010 2962.280 2899.290 2962.560 ;
        RECT 2618.410 2759.640 2618.690 2759.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2898.985 2962.570 2899.315 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2898.985 2962.270 2924.800 2962.570 ;
        RECT 2898.985 2962.255 2899.315 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2606.000 2759.930 2610.000 2760.320 ;
        RECT 2618.385 2759.930 2618.715 2759.945 ;
        RECT 2606.000 2759.720 2618.715 2759.930 ;
        RECT 2609.580 2759.630 2618.715 2759.720 ;
        RECT 2618.385 2759.615 2618.715 2759.630 ;
=======
        RECT 2919.700 2961.820 2924.800 2963.020 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 3194.880 2619.170 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2618.850 3194.740 2901.150 3194.880 ;
        RECT 2618.850 3194.680 2619.170 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 2618.880 3194.680 2619.140 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2618.880 3194.650 2619.140 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 2618.940 2959.885 2619.080 3194.650 ;
        RECT 2618.870 2959.515 2619.150 2959.885 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 2618.870 2959.560 2619.150 2959.840 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2606.000 2959.850 2610.000 2960.240 ;
        RECT 2618.845 2959.850 2619.175 2959.865 ;
        RECT 2606.000 2959.640 2619.175 2959.850 ;
        RECT 2609.580 2959.550 2619.175 2959.640 ;
        RECT 2618.845 2959.535 2619.175 2959.550 ;
=======
        RECT 2919.700 3196.420 2924.800 3197.620 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 3429.480 2618.710 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2618.390 3429.340 2901.150 3429.480 ;
        RECT 2618.390 3429.280 2618.710 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 2618.420 3429.280 2618.680 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 2618.420 3429.250 2618.680 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 2618.480 3159.805 2618.620 3429.250 ;
        RECT 2618.410 3159.435 2618.690 3159.805 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 2618.410 3159.480 2618.690 3159.760 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2606.000 3159.770 2610.000 3160.160 ;
        RECT 2618.385 3159.770 2618.715 3159.785 ;
        RECT 2606.000 3159.560 2618.715 3159.770 ;
        RECT 2609.580 3159.470 2618.715 3159.560 ;
        RECT 2618.385 3159.455 2618.715 3159.470 ;
=======
        RECT 2919.700 3431.020 2924.800 3432.220 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2483.610 3501.900 2483.930 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 2483.610 3501.760 2717.610 3501.900 ;
        RECT 2483.610 3501.700 2483.930 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 2483.640 3501.700 2483.900 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 2483.640 3501.670 2483.900 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 2481.750 3259.650 2482.030 3260.000 ;
        RECT 2483.700 3259.650 2483.840 3501.670 ;
        RECT 2481.750 3259.510 2483.840 3259.650 ;
        RECT 2481.750 3256.000 2482.030 3259.510 ;
=======
        RECT 2717.170 3519.700 2717.730 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2228.310 3501.900 2228.630 3501.960 ;
        RECT 2392.530 3501.900 2392.850 3501.960 ;
        RECT 2228.310 3501.760 2392.850 3501.900 ;
        RECT 2228.310 3501.700 2228.630 3501.760 ;
        RECT 2392.530 3501.700 2392.850 3501.760 ;
      LAYER via ;
        RECT 2228.340 3501.700 2228.600 3501.960 ;
        RECT 2392.560 3501.700 2392.820 3501.960 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.990 2392.760 3517.600 ;
        RECT 2228.340 3501.670 2228.600 3501.990 ;
        RECT 2392.560 3501.670 2392.820 3501.990 ;
        RECT 2226.450 3259.650 2226.730 3260.000 ;
        RECT 2228.400 3259.650 2228.540 3501.670 ;
        RECT 2226.450 3259.510 2228.540 3259.650 ;
        RECT 2226.450 3256.000 2226.730 3259.510 ;
=======
        RECT 2392.410 3519.700 2392.970 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1973.010 3501.900 1973.330 3501.960 ;
        RECT 2068.230 3501.900 2068.550 3501.960 ;
        RECT 1973.010 3501.760 2068.550 3501.900 ;
        RECT 1973.010 3501.700 1973.330 3501.760 ;
        RECT 2068.230 3501.700 2068.550 3501.760 ;
      LAYER via ;
        RECT 1973.040 3501.700 1973.300 3501.960 ;
        RECT 2068.260 3501.700 2068.520 3501.960 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.990 2068.460 3517.600 ;
        RECT 1973.040 3501.670 1973.300 3501.990 ;
        RECT 2068.260 3501.670 2068.520 3501.990 ;
        RECT 1970.690 3258.970 1970.970 3260.000 ;
        RECT 1973.100 3258.970 1973.240 3501.670 ;
        RECT 1970.690 3258.830 1973.240 3258.970 ;
        RECT 1970.690 3256.000 1970.970 3258.830 ;
=======
        RECT 2068.110 3519.700 2068.670 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1717.710 3501.560 1718.030 3501.620 ;
        RECT 1743.930 3501.560 1744.250 3501.620 ;
        RECT 1717.710 3501.420 1744.250 3501.560 ;
        RECT 1717.710 3501.360 1718.030 3501.420 ;
        RECT 1743.930 3501.360 1744.250 3501.420 ;
      LAYER via ;
        RECT 1717.740 3501.360 1718.000 3501.620 ;
        RECT 1743.960 3501.360 1744.220 3501.620 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3501.650 1744.160 3517.600 ;
        RECT 1717.740 3501.330 1718.000 3501.650 ;
        RECT 1743.960 3501.330 1744.220 3501.650 ;
        RECT 1714.930 3258.970 1715.210 3260.000 ;
        RECT 1717.800 3258.970 1717.940 3501.330 ;
        RECT 1714.930 3258.830 1717.940 3258.970 ;
        RECT 1714.930 3256.000 1715.210 3258.830 ;
=======
        RECT 1743.810 3519.700 1744.370 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1420.165 3381.045 1420.335 3429.155 ;
      LAYER mcon ;
        RECT 1420.165 3428.985 1420.335 3429.155 ;
      LAYER met1 ;
        RECT 1419.170 3477.760 1419.490 3477.820 ;
        RECT 1419.630 3477.760 1419.950 3477.820 ;
        RECT 1419.170 3477.620 1419.950 3477.760 ;
        RECT 1419.170 3477.560 1419.490 3477.620 ;
        RECT 1419.630 3477.560 1419.950 3477.620 ;
        RECT 1419.630 3443.080 1419.950 3443.140 ;
        RECT 1420.550 3443.080 1420.870 3443.140 ;
        RECT 1419.630 3442.940 1420.870 3443.080 ;
        RECT 1419.630 3442.880 1419.950 3442.940 ;
        RECT 1420.550 3442.880 1420.870 3442.940 ;
        RECT 1420.105 3429.140 1420.395 3429.185 ;
        RECT 1420.550 3429.140 1420.870 3429.200 ;
        RECT 1420.105 3429.000 1420.870 3429.140 ;
        RECT 1420.105 3428.955 1420.395 3429.000 ;
        RECT 1420.550 3428.940 1420.870 3429.000 ;
        RECT 1420.090 3381.200 1420.410 3381.260 ;
        RECT 1419.895 3381.060 1420.410 3381.200 ;
        RECT 1420.090 3381.000 1420.410 3381.060 ;
        RECT 1420.090 3367.600 1420.410 3367.660 ;
        RECT 1421.010 3367.600 1421.330 3367.660 ;
        RECT 1420.090 3367.460 1421.330 3367.600 ;
        RECT 1420.090 3367.400 1420.410 3367.460 ;
        RECT 1421.010 3367.400 1421.330 3367.460 ;
        RECT 1420.090 3274.100 1420.410 3274.160 ;
        RECT 1459.650 3274.100 1459.970 3274.160 ;
        RECT 1420.090 3273.960 1459.970 3274.100 ;
        RECT 1420.090 3273.900 1420.410 3273.960 ;
        RECT 1459.650 3273.900 1459.970 3273.960 ;
      LAYER via ;
        RECT 1419.200 3477.560 1419.460 3477.820 ;
        RECT 1419.660 3477.560 1419.920 3477.820 ;
        RECT 1419.660 3442.880 1419.920 3443.140 ;
        RECT 1420.580 3442.880 1420.840 3443.140 ;
        RECT 1420.580 3428.940 1420.840 3429.200 ;
        RECT 1420.120 3381.000 1420.380 3381.260 ;
        RECT 1420.120 3367.400 1420.380 3367.660 ;
        RECT 1421.040 3367.400 1421.300 3367.660 ;
        RECT 1420.120 3273.900 1420.380 3274.160 ;
        RECT 1459.680 3273.900 1459.940 3274.160 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3477.850 1419.400 3517.600 ;
        RECT 1419.200 3477.530 1419.460 3477.850 ;
        RECT 1419.660 3477.530 1419.920 3477.850 ;
        RECT 1419.720 3443.170 1419.860 3477.530 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3274.190 1420.320 3318.670 ;
        RECT 1420.120 3273.870 1420.380 3274.190 ;
        RECT 1459.680 3273.870 1459.940 3274.190 ;
        RECT 1459.740 3260.000 1459.880 3273.870 ;
        RECT 1459.630 3256.000 1459.910 3260.000 ;
=======
        RECT 1419.050 3519.700 1419.610 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 386.140 2619.170 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2618.850 386.000 2901.150 386.140 ;
        RECT 2618.850 385.940 2619.170 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2618.880 385.940 2619.140 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2618.870 559.795 2619.150 560.165 ;
        RECT 2618.940 386.230 2619.080 559.795 ;
        RECT 2618.880 385.910 2619.140 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2618.870 559.840 2619.150 560.120 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 560.130 2610.000 560.520 ;
        RECT 2618.845 560.130 2619.175 560.145 ;
        RECT 2606.000 559.920 2619.175 560.130 ;
        RECT 2609.580 559.830 2619.175 559.920 ;
        RECT 2618.845 559.815 2619.175 559.830 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
=======
        RECT 2919.700 380.540 2924.800 381.740 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1095.405 3284.485 1095.575 3332.595 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1095.405 3332.425 1095.575 3332.595 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1095.330 3395.140 1095.650 3395.200 ;
        RECT 1094.960 3395.000 1095.650 3395.140 ;
        RECT 1094.960 3394.860 1095.100 3395.000 ;
        RECT 1095.330 3394.940 1095.650 3395.000 ;
        RECT 1094.870 3394.600 1095.190 3394.860 ;
        RECT 1094.870 3346.520 1095.190 3346.580 ;
        RECT 1095.790 3346.520 1096.110 3346.580 ;
        RECT 1094.870 3346.380 1096.110 3346.520 ;
        RECT 1094.870 3346.320 1095.190 3346.380 ;
        RECT 1095.790 3346.320 1096.110 3346.380 ;
        RECT 1095.345 3332.580 1095.635 3332.625 ;
        RECT 1095.790 3332.580 1096.110 3332.640 ;
        RECT 1095.345 3332.440 1096.110 3332.580 ;
        RECT 1095.345 3332.395 1095.635 3332.440 ;
        RECT 1095.790 3332.380 1096.110 3332.440 ;
        RECT 1095.330 3284.640 1095.650 3284.700 ;
        RECT 1095.135 3284.500 1095.650 3284.640 ;
        RECT 1095.330 3284.440 1095.650 3284.500 ;
        RECT 1095.330 3274.440 1095.650 3274.500 ;
        RECT 1203.890 3274.440 1204.210 3274.500 ;
        RECT 1095.330 3274.300 1204.210 3274.440 ;
        RECT 1095.330 3274.240 1095.650 3274.300 ;
        RECT 1203.890 3274.240 1204.210 3274.300 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1095.360 3394.940 1095.620 3395.200 ;
        RECT 1094.900 3394.600 1095.160 3394.860 ;
        RECT 1094.900 3346.320 1095.160 3346.580 ;
        RECT 1095.820 3346.320 1096.080 3346.580 ;
        RECT 1095.820 3332.380 1096.080 3332.640 ;
        RECT 1095.360 3284.440 1095.620 3284.700 ;
        RECT 1095.360 3274.240 1095.620 3274.500 ;
        RECT 1203.920 3274.240 1204.180 3274.500 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3395.230 1095.560 3429.250 ;
        RECT 1095.360 3394.910 1095.620 3395.230 ;
        RECT 1094.900 3394.570 1095.160 3394.890 ;
        RECT 1094.960 3346.610 1095.100 3394.570 ;
        RECT 1094.900 3346.290 1095.160 3346.610 ;
        RECT 1095.820 3346.290 1096.080 3346.610 ;
        RECT 1095.880 3332.670 1096.020 3346.290 ;
        RECT 1095.820 3332.350 1096.080 3332.670 ;
        RECT 1095.360 3284.410 1095.620 3284.730 ;
        RECT 1095.420 3274.530 1095.560 3284.410 ;
        RECT 1095.360 3274.210 1095.620 3274.530 ;
        RECT 1203.920 3274.210 1204.180 3274.530 ;
        RECT 1203.980 3260.000 1204.120 3274.210 ;
        RECT 1203.870 3256.000 1204.150 3260.000 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
=======
        RECT 1094.750 3519.700 1095.310 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3274.100 771.810 3274.160 ;
        RECT 948.590 3274.100 948.910 3274.160 ;
        RECT 771.490 3273.960 948.910 3274.100 ;
        RECT 771.490 3273.900 771.810 3273.960 ;
        RECT 948.590 3273.900 948.910 3273.960 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3273.900 771.780 3274.160 ;
        RECT 948.620 3273.900 948.880 3274.160 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3274.190 771.720 3318.670 ;
        RECT 771.520 3273.870 771.780 3274.190 ;
        RECT 948.620 3273.870 948.880 3274.190 ;
        RECT 948.680 3260.000 948.820 3273.870 ;
        RECT 948.570 3256.000 948.850 3260.000 ;
=======
        RECT 770.450 3519.700 771.010 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 3274.100 448.430 3274.160 ;
        RECT 692.830 3274.100 693.150 3274.160 ;
        RECT 448.110 3273.960 693.150 3274.100 ;
        RECT 448.110 3273.900 448.430 3273.960 ;
        RECT 692.830 3273.900 693.150 3273.960 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 3273.900 448.400 3274.160 ;
        RECT 692.860 3273.900 693.120 3274.160 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 3274.190 448.340 3498.270 ;
        RECT 448.140 3273.870 448.400 3274.190 ;
        RECT 692.860 3273.870 693.120 3274.190 ;
        RECT 692.920 3260.000 693.060 3273.870 ;
        RECT 692.810 3256.000 693.090 3260.000 ;
=======
        RECT 445.690 3519.700 446.250 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 3274.100 124.130 3274.160 ;
        RECT 437.530 3274.100 437.850 3274.160 ;
        RECT 123.810 3273.960 437.850 3274.100 ;
        RECT 123.810 3273.900 124.130 3273.960 ;
        RECT 437.530 3273.900 437.850 3273.960 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 3273.900 124.100 3274.160 ;
        RECT 437.560 3273.900 437.820 3274.160 ;
      LAYER met2 ;
<<<<<<< HEAD
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 3274.190 124.040 3498.270 ;
        RECT 123.840 3273.870 124.100 3274.190 ;
        RECT 437.560 3273.870 437.820 3274.190 ;
        RECT 437.620 3260.000 437.760 3273.870 ;
        RECT 437.510 3256.000 437.790 3260.000 ;
=======
        RECT 121.390 3519.700 121.950 3524.800 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3153.060 17.410 3153.120 ;
        RECT 296.770 3153.060 297.090 3153.120 ;
        RECT 17.090 3152.920 297.090 3153.060 ;
        RECT 17.090 3152.860 17.410 3152.920 ;
        RECT 296.770 3152.860 297.090 3152.920 ;
      LAYER via ;
        RECT 17.120 3152.860 17.380 3153.120 ;
        RECT 296.800 3152.860 297.060 3153.120 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 3153.150 17.320 3339.635 ;
        RECT 17.120 3152.830 17.380 3153.150 ;
        RECT 296.800 3152.830 297.060 3153.150 ;
        RECT 296.860 3152.325 297.000 3152.830 ;
        RECT 296.790 3151.955 297.070 3152.325 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 296.790 3152.000 297.070 3152.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 296.765 3152.290 297.095 3152.305 ;
        RECT 310.000 3152.290 314.000 3152.680 ;
        RECT 296.765 3152.080 314.000 3152.290 ;
        RECT 296.765 3151.990 310.500 3152.080 ;
        RECT 296.765 3151.975 297.095 3151.990 ;
=======
        RECT -4.800 3339.220 0.300 3340.420 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2939.200 17.410 2939.260 ;
        RECT 296.770 2939.200 297.090 2939.260 ;
        RECT 17.090 2939.060 297.090 2939.200 ;
        RECT 17.090 2939.000 17.410 2939.060 ;
        RECT 296.770 2939.000 297.090 2939.060 ;
      LAYER via ;
        RECT 17.120 2939.000 17.380 2939.260 ;
        RECT 296.800 2939.000 297.060 2939.260 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 2939.290 17.320 3051.995 ;
        RECT 17.120 2938.970 17.380 2939.290 ;
        RECT 296.800 2938.970 297.060 2939.290 ;
        RECT 296.860 2938.125 297.000 2938.970 ;
        RECT 296.790 2937.755 297.070 2938.125 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 296.790 2937.800 297.070 2938.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 296.765 2938.090 297.095 2938.105 ;
        RECT 310.000 2938.090 314.000 2938.480 ;
        RECT 296.765 2937.880 314.000 2938.090 ;
        RECT 296.765 2937.790 310.500 2937.880 ;
        RECT 296.765 2937.775 297.095 2937.790 ;
=======
        RECT -4.800 3051.580 0.300 3052.780 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2725.340 17.410 2725.400 ;
        RECT 296.770 2725.340 297.090 2725.400 ;
        RECT 17.090 2725.200 297.090 2725.340 ;
        RECT 17.090 2725.140 17.410 2725.200 ;
        RECT 296.770 2725.140 297.090 2725.200 ;
      LAYER via ;
        RECT 17.120 2725.140 17.380 2725.400 ;
        RECT 296.800 2725.140 297.060 2725.400 ;
      LAYER met2 ;
        RECT 17.110 2765.035 17.390 2765.405 ;
        RECT 17.180 2725.430 17.320 2765.035 ;
        RECT 17.120 2725.110 17.380 2725.430 ;
        RECT 296.800 2725.110 297.060 2725.430 ;
        RECT 296.860 2723.925 297.000 2725.110 ;
        RECT 296.790 2723.555 297.070 2723.925 ;
      LAYER via2 ;
        RECT 17.110 2765.080 17.390 2765.360 ;
        RECT 296.790 2723.600 297.070 2723.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 17.085 2765.370 17.415 2765.385 ;
        RECT -4.800 2765.070 17.415 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 17.085 2765.055 17.415 2765.070 ;
        RECT 296.765 2723.890 297.095 2723.905 ;
        RECT 310.000 2723.890 314.000 2724.280 ;
        RECT 296.765 2723.680 314.000 2723.890 ;
        RECT 296.765 2723.590 310.500 2723.680 ;
        RECT 296.765 2723.575 297.095 2723.590 ;
=======
        RECT -4.800 2764.620 0.300 2765.820 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2505.020 16.950 2505.080 ;
        RECT 296.770 2505.020 297.090 2505.080 ;
        RECT 16.630 2504.880 297.090 2505.020 ;
        RECT 16.630 2504.820 16.950 2504.880 ;
        RECT 296.770 2504.820 297.090 2504.880 ;
      LAYER via ;
        RECT 16.660 2504.820 16.920 2505.080 ;
        RECT 296.800 2504.820 297.060 2505.080 ;
      LAYER met2 ;
        RECT 296.790 2509.355 297.070 2509.725 ;
        RECT 296.860 2505.110 297.000 2509.355 ;
        RECT 16.660 2504.790 16.920 2505.110 ;
        RECT 296.800 2504.790 297.060 2505.110 ;
        RECT 16.720 2477.765 16.860 2504.790 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
      LAYER via2 ;
        RECT 296.790 2509.400 297.070 2509.680 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2509.690 297.095 2509.705 ;
        RECT 310.000 2509.690 314.000 2510.080 ;
        RECT 296.765 2509.480 314.000 2509.690 ;
        RECT 296.765 2509.390 310.500 2509.480 ;
        RECT 296.765 2509.375 297.095 2509.390 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
=======
        RECT -4.800 2476.980 0.300 2478.180 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2291.160 17.870 2291.220 ;
        RECT 296.770 2291.160 297.090 2291.220 ;
        RECT 17.550 2291.020 297.090 2291.160 ;
        RECT 17.550 2290.960 17.870 2291.020 ;
        RECT 296.770 2290.960 297.090 2291.020 ;
      LAYER via ;
        RECT 17.580 2290.960 17.840 2291.220 ;
        RECT 296.800 2290.960 297.060 2291.220 ;
      LAYER met2 ;
        RECT 296.790 2295.155 297.070 2295.525 ;
        RECT 296.860 2291.250 297.000 2295.155 ;
        RECT 17.580 2290.930 17.840 2291.250 ;
        RECT 296.800 2290.930 297.060 2291.250 ;
        RECT 17.640 2190.125 17.780 2290.930 ;
        RECT 17.570 2189.755 17.850 2190.125 ;
      LAYER via2 ;
        RECT 296.790 2295.200 297.070 2295.480 ;
        RECT 17.570 2189.800 17.850 2190.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2295.490 297.095 2295.505 ;
        RECT 310.000 2295.490 314.000 2295.880 ;
        RECT 296.765 2295.280 314.000 2295.490 ;
        RECT 296.765 2295.190 310.500 2295.280 ;
        RECT 296.765 2295.175 297.095 2295.190 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 17.545 2190.090 17.875 2190.105 ;
        RECT -4.800 2189.790 17.875 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 17.545 2189.775 17.875 2189.790 ;
=======
        RECT -4.800 2189.340 0.300 2190.540 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2077.300 17.410 2077.360 ;
        RECT 296.770 2077.300 297.090 2077.360 ;
        RECT 17.090 2077.160 297.090 2077.300 ;
        RECT 17.090 2077.100 17.410 2077.160 ;
        RECT 296.770 2077.100 297.090 2077.160 ;
      LAYER via ;
        RECT 17.120 2077.100 17.380 2077.360 ;
        RECT 296.800 2077.100 297.060 2077.360 ;
      LAYER met2 ;
        RECT 296.790 2080.955 297.070 2081.325 ;
        RECT 296.860 2077.390 297.000 2080.955 ;
        RECT 17.120 2077.070 17.380 2077.390 ;
        RECT 296.800 2077.070 297.060 2077.390 ;
        RECT 17.180 1903.165 17.320 2077.070 ;
        RECT 17.110 1902.795 17.390 1903.165 ;
      LAYER via2 ;
        RECT 296.790 2081.000 297.070 2081.280 ;
        RECT 17.110 1902.840 17.390 1903.120 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 2081.290 297.095 2081.305 ;
        RECT 310.000 2081.290 314.000 2081.680 ;
        RECT 296.765 2081.080 314.000 2081.290 ;
        RECT 296.765 2080.990 310.500 2081.080 ;
        RECT 296.765 2080.975 297.095 2080.990 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 17.085 1903.130 17.415 1903.145 ;
        RECT -4.800 1902.830 17.415 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 17.085 1902.815 17.415 1902.830 ;
=======
        RECT -4.800 1902.380 0.300 1903.580 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 620.740 2619.170 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2618.850 620.600 2901.150 620.740 ;
        RECT 2618.850 620.540 2619.170 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2618.880 620.540 2619.140 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2618.870 759.715 2619.150 760.085 ;
        RECT 2618.940 620.830 2619.080 759.715 ;
        RECT 2618.880 620.510 2619.140 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2618.870 759.760 2619.150 760.040 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 760.050 2610.000 760.440 ;
        RECT 2618.845 760.050 2619.175 760.065 ;
        RECT 2606.000 759.840 2619.175 760.050 ;
        RECT 2609.580 759.750 2619.175 759.840 ;
        RECT 2618.845 759.735 2619.175 759.750 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
=======
        RECT 2919.700 615.140 2924.800 616.340 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1863.100 17.870 1863.160 ;
        RECT 296.770 1863.100 297.090 1863.160 ;
        RECT 17.550 1862.960 297.090 1863.100 ;
        RECT 17.550 1862.900 17.870 1862.960 ;
        RECT 296.770 1862.900 297.090 1862.960 ;
      LAYER via ;
        RECT 17.580 1862.900 17.840 1863.160 ;
        RECT 296.800 1862.900 297.060 1863.160 ;
      LAYER met2 ;
        RECT 296.790 1866.755 297.070 1867.125 ;
        RECT 296.860 1863.190 297.000 1866.755 ;
        RECT 17.580 1862.870 17.840 1863.190 ;
        RECT 296.800 1862.870 297.060 1863.190 ;
        RECT 17.640 1615.525 17.780 1862.870 ;
        RECT 17.570 1615.155 17.850 1615.525 ;
      LAYER via2 ;
        RECT 296.790 1866.800 297.070 1867.080 ;
        RECT 17.570 1615.200 17.850 1615.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1867.090 297.095 1867.105 ;
        RECT 310.000 1867.090 314.000 1867.480 ;
        RECT 296.765 1866.880 314.000 1867.090 ;
        RECT 296.765 1866.790 310.500 1866.880 ;
        RECT 296.765 1866.775 297.095 1866.790 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 17.545 1615.490 17.875 1615.505 ;
        RECT -4.800 1615.190 17.875 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 17.545 1615.175 17.875 1615.190 ;
=======
        RECT -4.800 1614.740 0.300 1615.940 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 1649.240 18.330 1649.300 ;
        RECT 296.770 1649.240 297.090 1649.300 ;
        RECT 18.010 1649.100 297.090 1649.240 ;
        RECT 18.010 1649.040 18.330 1649.100 ;
        RECT 296.770 1649.040 297.090 1649.100 ;
      LAYER via ;
        RECT 18.040 1649.040 18.300 1649.300 ;
        RECT 296.800 1649.040 297.060 1649.300 ;
      LAYER met2 ;
        RECT 296.790 1651.875 297.070 1652.245 ;
        RECT 296.860 1649.330 297.000 1651.875 ;
        RECT 18.040 1649.010 18.300 1649.330 ;
        RECT 296.800 1649.010 297.060 1649.330 ;
        RECT 18.100 1400.645 18.240 1649.010 ;
        RECT 18.030 1400.275 18.310 1400.645 ;
      LAYER via2 ;
        RECT 296.790 1651.920 297.070 1652.200 ;
        RECT 18.030 1400.320 18.310 1400.600 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1652.210 297.095 1652.225 ;
        RECT 310.000 1652.210 314.000 1652.600 ;
        RECT 296.765 1652.000 314.000 1652.210 ;
        RECT 296.765 1651.910 310.500 1652.000 ;
        RECT 296.765 1651.895 297.095 1651.910 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 18.005 1400.610 18.335 1400.625 ;
        RECT -4.800 1400.310 18.335 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 18.005 1400.295 18.335 1400.310 ;
=======
        RECT -4.800 1399.860 0.300 1401.060 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1435.380 17.870 1435.440 ;
        RECT 296.770 1435.380 297.090 1435.440 ;
        RECT 17.550 1435.240 297.090 1435.380 ;
        RECT 17.550 1435.180 17.870 1435.240 ;
        RECT 296.770 1435.180 297.090 1435.240 ;
      LAYER via ;
        RECT 17.580 1435.180 17.840 1435.440 ;
        RECT 296.800 1435.180 297.060 1435.440 ;
      LAYER met2 ;
        RECT 296.790 1437.675 297.070 1438.045 ;
        RECT 296.860 1435.470 297.000 1437.675 ;
        RECT 17.580 1435.150 17.840 1435.470 ;
        RECT 296.800 1435.150 297.060 1435.470 ;
        RECT 17.640 1185.085 17.780 1435.150 ;
        RECT 17.570 1184.715 17.850 1185.085 ;
      LAYER via2 ;
        RECT 296.790 1437.720 297.070 1438.000 ;
        RECT 17.570 1184.760 17.850 1185.040 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1438.010 297.095 1438.025 ;
        RECT 310.000 1438.010 314.000 1438.400 ;
        RECT 296.765 1437.800 314.000 1438.010 ;
        RECT 296.765 1437.710 310.500 1437.800 ;
        RECT 296.765 1437.695 297.095 1437.710 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.545 1185.050 17.875 1185.065 ;
        RECT -4.800 1184.750 17.875 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.545 1184.735 17.875 1184.750 ;
=======
        RECT -4.800 1184.300 0.300 1185.500 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1221.520 17.410 1221.580 ;
        RECT 296.770 1221.520 297.090 1221.580 ;
        RECT 17.090 1221.380 297.090 1221.520 ;
        RECT 17.090 1221.320 17.410 1221.380 ;
        RECT 296.770 1221.320 297.090 1221.380 ;
      LAYER via ;
        RECT 17.120 1221.320 17.380 1221.580 ;
        RECT 296.800 1221.320 297.060 1221.580 ;
      LAYER met2 ;
        RECT 296.790 1223.475 297.070 1223.845 ;
        RECT 296.860 1221.610 297.000 1223.475 ;
        RECT 17.120 1221.290 17.380 1221.610 ;
        RECT 296.800 1221.290 297.060 1221.610 ;
        RECT 17.180 969.525 17.320 1221.290 ;
        RECT 17.110 969.155 17.390 969.525 ;
      LAYER via2 ;
        RECT 296.790 1223.520 297.070 1223.800 ;
        RECT 17.110 969.200 17.390 969.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1223.810 297.095 1223.825 ;
        RECT 310.000 1223.810 314.000 1224.200 ;
        RECT 296.765 1223.600 314.000 1223.810 ;
        RECT 296.765 1223.510 310.500 1223.600 ;
        RECT 296.765 1223.495 297.095 1223.510 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 17.085 969.490 17.415 969.505 ;
        RECT -4.800 969.190 17.415 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 17.085 969.175 17.415 969.190 ;
=======
        RECT -4.800 968.740 0.300 969.940 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1007.660 17.870 1007.720 ;
        RECT 296.770 1007.660 297.090 1007.720 ;
        RECT 17.550 1007.520 297.090 1007.660 ;
        RECT 17.550 1007.460 17.870 1007.520 ;
        RECT 296.770 1007.460 297.090 1007.520 ;
      LAYER via ;
        RECT 17.580 1007.460 17.840 1007.720 ;
        RECT 296.800 1007.460 297.060 1007.720 ;
      LAYER met2 ;
        RECT 296.790 1009.275 297.070 1009.645 ;
        RECT 296.860 1007.750 297.000 1009.275 ;
        RECT 17.580 1007.430 17.840 1007.750 ;
        RECT 296.800 1007.430 297.060 1007.750 ;
        RECT 17.640 753.965 17.780 1007.430 ;
        RECT 17.570 753.595 17.850 753.965 ;
      LAYER via2 ;
        RECT 296.790 1009.320 297.070 1009.600 ;
        RECT 17.570 753.640 17.850 753.920 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 1009.610 297.095 1009.625 ;
        RECT 310.000 1009.610 314.000 1010.000 ;
        RECT 296.765 1009.400 314.000 1009.610 ;
        RECT 296.765 1009.310 310.500 1009.400 ;
        RECT 296.765 1009.295 297.095 1009.310 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 17.545 753.930 17.875 753.945 ;
        RECT -4.800 753.630 17.875 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 17.545 753.615 17.875 753.630 ;
=======
        RECT -4.800 753.180 0.300 754.380 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 793.800 17.410 793.860 ;
        RECT 296.770 793.800 297.090 793.860 ;
        RECT 17.090 793.660 297.090 793.800 ;
        RECT 17.090 793.600 17.410 793.660 ;
        RECT 296.770 793.600 297.090 793.660 ;
      LAYER via ;
        RECT 17.120 793.600 17.380 793.860 ;
        RECT 296.800 793.600 297.060 793.860 ;
      LAYER met2 ;
        RECT 296.790 795.075 297.070 795.445 ;
        RECT 296.860 793.890 297.000 795.075 ;
        RECT 17.120 793.570 17.380 793.890 ;
        RECT 296.800 793.570 297.060 793.890 ;
        RECT 17.180 538.405 17.320 793.570 ;
        RECT 17.110 538.035 17.390 538.405 ;
      LAYER via2 ;
        RECT 296.790 795.120 297.070 795.400 ;
        RECT 17.110 538.080 17.390 538.360 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 795.410 297.095 795.425 ;
        RECT 310.000 795.410 314.000 795.800 ;
        RECT 296.765 795.200 314.000 795.410 ;
        RECT 296.765 795.110 310.500 795.200 ;
        RECT 296.765 795.095 297.095 795.110 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.085 538.370 17.415 538.385 ;
        RECT -4.800 538.070 17.415 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.085 538.055 17.415 538.070 ;
=======
        RECT -4.800 537.620 0.300 538.820 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 579.940 17.870 580.000 ;
        RECT 296.770 579.940 297.090 580.000 ;
        RECT 17.550 579.800 297.090 579.940 ;
        RECT 17.550 579.740 17.870 579.800 ;
        RECT 296.770 579.740 297.090 579.800 ;
      LAYER via ;
        RECT 17.580 579.740 17.840 580.000 ;
        RECT 296.800 579.740 297.060 580.000 ;
      LAYER met2 ;
        RECT 296.790 580.875 297.070 581.245 ;
        RECT 296.860 580.030 297.000 580.875 ;
        RECT 17.580 579.710 17.840 580.030 ;
        RECT 296.800 579.710 297.060 580.030 ;
        RECT 17.640 322.845 17.780 579.710 ;
        RECT 17.570 322.475 17.850 322.845 ;
      LAYER via2 ;
        RECT 296.790 580.920 297.070 581.200 ;
        RECT 17.570 322.520 17.850 322.800 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 581.210 297.095 581.225 ;
        RECT 310.000 581.210 314.000 581.600 ;
        RECT 296.765 581.000 314.000 581.210 ;
        RECT 296.765 580.910 310.500 581.000 ;
        RECT 296.765 580.895 297.095 580.910 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 17.545 322.810 17.875 322.825 ;
        RECT -4.800 322.510 17.875 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 17.545 322.495 17.875 322.510 ;
=======
        RECT -4.800 322.060 0.300 323.260 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 366.080 17.410 366.140 ;
        RECT 296.770 366.080 297.090 366.140 ;
        RECT 17.090 365.940 297.090 366.080 ;
        RECT 17.090 365.880 17.410 365.940 ;
        RECT 296.770 365.880 297.090 365.940 ;
      LAYER via ;
        RECT 17.120 365.880 17.380 366.140 ;
        RECT 296.800 365.880 297.060 366.140 ;
      LAYER met2 ;
        RECT 296.790 366.675 297.070 367.045 ;
        RECT 296.860 366.170 297.000 366.675 ;
        RECT 17.120 365.850 17.380 366.170 ;
        RECT 296.800 365.850 297.060 366.170 ;
        RECT 17.180 107.285 17.320 365.850 ;
        RECT 17.110 106.915 17.390 107.285 ;
      LAYER via2 ;
        RECT 296.790 366.720 297.070 367.000 ;
        RECT 17.110 106.960 17.390 107.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.765 367.010 297.095 367.025 ;
        RECT 310.000 367.010 314.000 367.400 ;
        RECT 296.765 366.800 314.000 367.010 ;
        RECT 296.765 366.710 310.500 366.800 ;
        RECT 296.765 366.695 297.095 366.710 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 17.085 107.250 17.415 107.265 ;
        RECT -4.800 106.950 17.415 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 17.085 106.935 17.415 106.950 ;
=======
        RECT -4.800 106.500 0.300 107.700 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 855.340 2619.170 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2618.850 855.200 2901.150 855.340 ;
        RECT 2618.850 855.140 2619.170 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2618.880 855.140 2619.140 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2618.870 959.635 2619.150 960.005 ;
        RECT 2618.940 855.430 2619.080 959.635 ;
        RECT 2618.880 855.110 2619.140 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2618.870 959.680 2619.150 959.960 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 959.970 2610.000 960.360 ;
        RECT 2618.845 959.970 2619.175 959.985 ;
        RECT 2606.000 959.760 2619.175 959.970 ;
        RECT 2609.580 959.670 2619.175 959.760 ;
        RECT 2618.845 959.655 2619.175 959.670 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
=======
        RECT 2919.700 849.740 2924.800 850.940 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 1089.940 2619.170 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2618.850 1089.800 2901.150 1089.940 ;
        RECT 2618.850 1089.740 2619.170 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2618.880 1089.740 2619.140 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2618.870 1159.555 2619.150 1159.925 ;
        RECT 2618.940 1090.030 2619.080 1159.555 ;
        RECT 2618.880 1089.710 2619.140 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2618.870 1159.600 2619.150 1159.880 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1159.890 2610.000 1160.280 ;
        RECT 2618.845 1159.890 2619.175 1159.905 ;
        RECT 2606.000 1159.680 2619.175 1159.890 ;
        RECT 2609.580 1159.590 2619.175 1159.680 ;
        RECT 2618.845 1159.575 2619.175 1159.590 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
=======
        RECT 2919.700 1084.340 2924.800 1085.540 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1324.540 2618.710 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2618.390 1324.400 2901.150 1324.540 ;
        RECT 2618.390 1324.340 2618.710 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 2618.420 1324.340 2618.680 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 2618.410 1359.475 2618.690 1359.845 ;
        RECT 2618.480 1324.630 2618.620 1359.475 ;
        RECT 2618.420 1324.310 2618.680 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2618.410 1359.520 2618.690 1359.800 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1359.810 2610.000 1360.200 ;
        RECT 2618.385 1359.810 2618.715 1359.825 ;
        RECT 2606.000 1359.600 2618.715 1359.810 ;
        RECT 2609.580 1359.510 2618.715 1359.600 ;
        RECT 2618.385 1359.495 2618.715 1359.510 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
=======
        RECT 2919.700 1318.940 2924.800 1320.140 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2621.610 1559.140 2621.930 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2621.610 1559.000 2901.150 1559.140 ;
        RECT 2621.610 1558.940 2621.930 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 2621.640 1558.940 2621.900 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 2621.630 1559.395 2621.910 1559.765 ;
        RECT 2621.700 1559.230 2621.840 1559.395 ;
        RECT 2621.640 1558.910 2621.900 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2621.630 1559.440 2621.910 1559.720 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2606.000 1559.730 2610.000 1560.120 ;
        RECT 2621.605 1559.730 2621.935 1559.745 ;
        RECT 2606.000 1559.520 2621.935 1559.730 ;
        RECT 2609.580 1559.430 2621.935 1559.520 ;
        RECT 2621.605 1559.415 2621.935 1559.430 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
=======
        RECT 2919.700 1553.540 2924.800 1554.740 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.390 1787.280 2618.710 1787.340 ;
        RECT 2900.830 1787.280 2901.150 1787.340 ;
        RECT 2618.390 1787.140 2901.150 1787.280 ;
        RECT 2618.390 1787.080 2618.710 1787.140 ;
        RECT 2900.830 1787.080 2901.150 1787.140 ;
      LAYER via ;
        RECT 2618.420 1787.080 2618.680 1787.340 ;
        RECT 2900.860 1787.080 2901.120 1787.340 ;
      LAYER met2 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
        RECT 2900.920 1787.370 2901.060 1789.235 ;
        RECT 2618.420 1787.050 2618.680 1787.370 ;
        RECT 2900.860 1787.050 2901.120 1787.370 ;
        RECT 2618.480 1759.685 2618.620 1787.050 ;
        RECT 2618.410 1759.315 2618.690 1759.685 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
        RECT 2618.410 1759.360 2618.690 1759.640 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2606.000 1759.650 2610.000 1760.040 ;
        RECT 2618.385 1759.650 2618.715 1759.665 ;
        RECT 2606.000 1759.440 2618.715 1759.650 ;
        RECT 2609.580 1759.350 2618.715 1759.440 ;
        RECT 2618.385 1759.335 2618.715 1759.350 ;
=======
        RECT 2919.700 1788.820 2924.800 1790.020 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2021.880 2619.170 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 2618.850 2021.740 2901.150 2021.880 ;
        RECT 2618.850 2021.680 2619.170 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 2618.880 2021.680 2619.140 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 2618.880 2021.650 2619.140 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 2618.940 1960.285 2619.080 2021.650 ;
        RECT 2618.870 1959.915 2619.150 1960.285 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
        RECT 2618.870 1959.960 2619.150 1960.240 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2606.000 1960.250 2610.000 1960.640 ;
        RECT 2618.845 1960.250 2619.175 1960.265 ;
        RECT 2606.000 1960.040 2619.175 1960.250 ;
        RECT 2609.580 1959.950 2619.175 1960.040 ;
        RECT 2618.845 1959.935 2619.175 1959.950 ;
=======
        RECT 2919.700 2023.420 2924.800 2024.620 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2256.480 2619.170 2256.540 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 2618.850 2256.340 2901.150 2256.480 ;
        RECT 2618.850 2256.280 2619.170 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
      LAYER via ;
        RECT 2618.880 2256.280 2619.140 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 2618.880 2256.250 2619.140 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 2618.940 2160.205 2619.080 2256.250 ;
        RECT 2618.870 2159.835 2619.150 2160.205 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
        RECT 2618.870 2159.880 2619.150 2160.160 ;
      LAYER met3 ;
<<<<<<< HEAD
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2606.000 2160.170 2610.000 2160.560 ;
        RECT 2618.845 2160.170 2619.175 2160.185 ;
        RECT 2606.000 2159.960 2619.175 2160.170 ;
        RECT 2609.580 2159.870 2619.175 2159.960 ;
        RECT 2618.845 2159.855 2619.175 2159.870 ;
=======
        RECT 2919.700 2258.020 2924.800 2259.220 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 324.370 243.680 324.690 243.740 ;
        RECT 330.810 243.680 331.130 243.740 ;
        RECT 324.370 243.540 331.130 243.680 ;
        RECT 324.370 243.480 324.690 243.540 ;
        RECT 330.810 243.480 331.130 243.540 ;
        RECT 330.810 24.380 331.130 24.440 ;
        RECT 633.030 24.380 633.350 24.440 ;
        RECT 330.810 24.240 633.350 24.380 ;
        RECT 330.810 24.180 331.130 24.240 ;
        RECT 633.030 24.180 633.350 24.240 ;
      LAYER via ;
        RECT 324.400 243.480 324.660 243.740 ;
        RECT 330.840 243.480 331.100 243.740 ;
        RECT 330.840 24.180 331.100 24.440 ;
        RECT 633.060 24.180 633.320 24.440 ;
      LAYER met2 ;
        RECT 324.350 260.000 324.630 264.000 ;
        RECT 324.460 243.770 324.600 260.000 ;
        RECT 324.400 243.450 324.660 243.770 ;
        RECT 330.840 243.450 331.100 243.770 ;
        RECT 330.900 24.470 331.040 243.450 ;
        RECT 330.840 24.150 331.100 24.470 ;
        RECT 633.060 24.150 633.320 24.470 ;
        RECT 633.120 2.400 633.260 24.150 ;
        RECT 632.910 -4.800 633.470 2.400 ;
=======
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2111.930 241.640 2112.250 241.700 ;
        RECT 2117.910 241.640 2118.230 241.700 ;
        RECT 2111.930 241.500 2118.230 241.640 ;
        RECT 2111.930 241.440 2112.250 241.500 ;
        RECT 2117.910 241.440 2118.230 241.500 ;
        RECT 2117.910 37.980 2118.230 38.040 ;
        RECT 2417.370 37.980 2417.690 38.040 ;
        RECT 2117.910 37.840 2417.690 37.980 ;
        RECT 2117.910 37.780 2118.230 37.840 ;
        RECT 2417.370 37.780 2417.690 37.840 ;
      LAYER via ;
        RECT 2111.960 241.440 2112.220 241.700 ;
        RECT 2117.940 241.440 2118.200 241.700 ;
        RECT 2117.940 37.780 2118.200 38.040 ;
        RECT 2417.400 37.780 2417.660 38.040 ;
      LAYER met2 ;
        RECT 2111.910 260.000 2112.190 264.000 ;
        RECT 2112.020 241.730 2112.160 260.000 ;
        RECT 2111.960 241.410 2112.220 241.730 ;
        RECT 2117.940 241.410 2118.200 241.730 ;
        RECT 2118.000 38.070 2118.140 241.410 ;
        RECT 2117.940 37.750 2118.200 38.070 ;
        RECT 2417.400 37.750 2417.660 38.070 ;
        RECT 2417.460 2.400 2417.600 37.750 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
=======
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2131.710 30.840 2132.030 30.900 ;
        RECT 2434.850 30.840 2435.170 30.900 ;
        RECT 2131.710 30.700 2435.170 30.840 ;
        RECT 2131.710 30.640 2132.030 30.700 ;
        RECT 2434.850 30.640 2435.170 30.700 ;
      LAYER via ;
        RECT 2131.740 30.640 2132.000 30.900 ;
        RECT 2434.880 30.640 2435.140 30.900 ;
      LAYER met2 ;
        RECT 2129.850 260.170 2130.130 264.000 ;
        RECT 2129.850 260.030 2131.940 260.170 ;
        RECT 2129.850 260.000 2130.130 260.030 ;
        RECT 2131.800 30.930 2131.940 260.030 ;
        RECT 2131.740 30.610 2132.000 30.930 ;
        RECT 2434.880 30.610 2435.140 30.930 ;
        RECT 2434.940 2.400 2435.080 30.610 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
=======
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2147.810 244.020 2148.130 244.080 ;
        RECT 2152.410 244.020 2152.730 244.080 ;
        RECT 2147.810 243.880 2152.730 244.020 ;
        RECT 2147.810 243.820 2148.130 243.880 ;
        RECT 2152.410 243.820 2152.730 243.880 ;
        RECT 2152.410 44.780 2152.730 44.840 ;
        RECT 2452.790 44.780 2453.110 44.840 ;
        RECT 2152.410 44.640 2453.110 44.780 ;
        RECT 2152.410 44.580 2152.730 44.640 ;
        RECT 2452.790 44.580 2453.110 44.640 ;
      LAYER via ;
        RECT 2147.840 243.820 2148.100 244.080 ;
        RECT 2152.440 243.820 2152.700 244.080 ;
        RECT 2152.440 44.580 2152.700 44.840 ;
        RECT 2452.820 44.580 2453.080 44.840 ;
      LAYER met2 ;
        RECT 2147.790 260.000 2148.070 264.000 ;
        RECT 2147.900 244.110 2148.040 260.000 ;
        RECT 2147.840 243.790 2148.100 244.110 ;
        RECT 2152.440 243.790 2152.700 244.110 ;
        RECT 2152.500 44.870 2152.640 243.790 ;
        RECT 2152.440 44.550 2152.700 44.870 ;
        RECT 2452.820 44.550 2453.080 44.870 ;
        RECT 2452.880 2.400 2453.020 44.550 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
=======
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2166.210 237.900 2166.530 237.960 ;
        RECT 2470.270 237.900 2470.590 237.960 ;
        RECT 2166.210 237.760 2470.590 237.900 ;
        RECT 2166.210 237.700 2166.530 237.760 ;
        RECT 2470.270 237.700 2470.590 237.760 ;
      LAYER via ;
        RECT 2166.240 237.700 2166.500 237.960 ;
        RECT 2470.300 237.700 2470.560 237.960 ;
      LAYER met2 ;
        RECT 2165.730 260.170 2166.010 264.000 ;
        RECT 2165.730 260.030 2166.440 260.170 ;
        RECT 2165.730 260.000 2166.010 260.030 ;
        RECT 2166.300 237.990 2166.440 260.030 ;
        RECT 2166.240 237.670 2166.500 237.990 ;
        RECT 2470.300 237.670 2470.560 237.990 ;
        RECT 2470.360 17.410 2470.500 237.670 ;
        RECT 2470.360 17.270 2470.960 17.410 ;
        RECT 2470.820 2.400 2470.960 17.270 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
=======
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2183.690 231.100 2184.010 231.160 ;
        RECT 2484.070 231.100 2484.390 231.160 ;
        RECT 2183.690 230.960 2484.390 231.100 ;
        RECT 2183.690 230.900 2184.010 230.960 ;
        RECT 2484.070 230.900 2484.390 230.960 ;
      LAYER via ;
        RECT 2183.720 230.900 2183.980 231.160 ;
        RECT 2484.100 230.900 2484.360 231.160 ;
      LAYER met2 ;
        RECT 2183.670 260.000 2183.950 264.000 ;
        RECT 2183.780 231.190 2183.920 260.000 ;
        RECT 2183.720 230.870 2183.980 231.190 ;
        RECT 2484.100 230.870 2484.360 231.190 ;
        RECT 2484.160 17.410 2484.300 230.870 ;
        RECT 2484.160 17.270 2488.900 17.410 ;
        RECT 2488.760 2.400 2488.900 17.270 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
=======
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2201.630 244.020 2201.950 244.080 ;
        RECT 2207.610 244.020 2207.930 244.080 ;
        RECT 2201.630 243.880 2207.930 244.020 ;
        RECT 2201.630 243.820 2201.950 243.880 ;
        RECT 2207.610 243.820 2207.930 243.880 ;
        RECT 2207.610 51.920 2207.930 51.980 ;
        RECT 2504.770 51.920 2505.090 51.980 ;
        RECT 2207.610 51.780 2505.090 51.920 ;
        RECT 2207.610 51.720 2207.930 51.780 ;
        RECT 2504.770 51.720 2505.090 51.780 ;
      LAYER via ;
        RECT 2201.660 243.820 2201.920 244.080 ;
        RECT 2207.640 243.820 2207.900 244.080 ;
        RECT 2207.640 51.720 2207.900 51.980 ;
        RECT 2504.800 51.720 2505.060 51.980 ;
      LAYER met2 ;
        RECT 2201.610 260.000 2201.890 264.000 ;
        RECT 2201.720 244.110 2201.860 260.000 ;
        RECT 2201.660 243.790 2201.920 244.110 ;
        RECT 2207.640 243.790 2207.900 244.110 ;
        RECT 2207.700 52.010 2207.840 243.790 ;
        RECT 2207.640 51.690 2207.900 52.010 ;
        RECT 2504.800 51.690 2505.060 52.010 ;
        RECT 2504.860 4.490 2505.000 51.690 ;
        RECT 2504.860 4.350 2506.380 4.490 ;
        RECT 2506.240 2.400 2506.380 4.350 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
=======
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2221.410 58.720 2221.730 58.780 ;
        RECT 2518.570 58.720 2518.890 58.780 ;
        RECT 2221.410 58.580 2518.890 58.720 ;
        RECT 2221.410 58.520 2221.730 58.580 ;
        RECT 2518.570 58.520 2518.890 58.580 ;
      LAYER via ;
        RECT 2221.440 58.520 2221.700 58.780 ;
        RECT 2518.600 58.520 2518.860 58.780 ;
      LAYER met2 ;
        RECT 2219.550 260.170 2219.830 264.000 ;
        RECT 2219.550 260.030 2221.640 260.170 ;
        RECT 2219.550 260.000 2219.830 260.030 ;
        RECT 2221.500 58.810 2221.640 260.030 ;
        RECT 2221.440 58.490 2221.700 58.810 ;
        RECT 2518.600 58.490 2518.860 58.810 ;
        RECT 2518.660 16.730 2518.800 58.490 ;
        RECT 2518.660 16.590 2524.320 16.730 ;
        RECT 2524.180 2.400 2524.320 16.590 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
=======
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2237.050 244.020 2237.370 244.080 ;
        RECT 2242.110 244.020 2242.430 244.080 ;
        RECT 2237.050 243.880 2242.430 244.020 ;
        RECT 2237.050 243.820 2237.370 243.880 ;
        RECT 2242.110 243.820 2242.430 243.880 ;
        RECT 2242.110 65.520 2242.430 65.580 ;
        RECT 2539.270 65.520 2539.590 65.580 ;
        RECT 2242.110 65.380 2539.590 65.520 ;
        RECT 2242.110 65.320 2242.430 65.380 ;
        RECT 2539.270 65.320 2539.590 65.380 ;
      LAYER via ;
        RECT 2237.080 243.820 2237.340 244.080 ;
        RECT 2242.140 243.820 2242.400 244.080 ;
        RECT 2242.140 65.320 2242.400 65.580 ;
        RECT 2539.300 65.320 2539.560 65.580 ;
      LAYER met2 ;
        RECT 2237.030 260.000 2237.310 264.000 ;
        RECT 2237.140 244.110 2237.280 260.000 ;
        RECT 2237.080 243.790 2237.340 244.110 ;
        RECT 2242.140 243.790 2242.400 244.110 ;
        RECT 2242.200 65.610 2242.340 243.790 ;
        RECT 2242.140 65.290 2242.400 65.610 ;
        RECT 2539.300 65.290 2539.560 65.610 ;
        RECT 2539.360 16.730 2539.500 65.290 ;
        RECT 2539.360 16.590 2542.260 16.730 ;
        RECT 2542.120 2.400 2542.260 16.590 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
=======
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2255.910 224.300 2256.230 224.360 ;
        RECT 2559.970 224.300 2560.290 224.360 ;
        RECT 2255.910 224.160 2560.290 224.300 ;
        RECT 2255.910 224.100 2256.230 224.160 ;
        RECT 2559.970 224.100 2560.290 224.160 ;
      LAYER via ;
        RECT 2255.940 224.100 2256.200 224.360 ;
        RECT 2560.000 224.100 2560.260 224.360 ;
      LAYER met2 ;
        RECT 2254.970 260.170 2255.250 264.000 ;
        RECT 2254.970 260.030 2256.140 260.170 ;
        RECT 2254.970 260.000 2255.250 260.030 ;
        RECT 2256.000 224.390 2256.140 260.030 ;
        RECT 2255.940 224.070 2256.200 224.390 ;
        RECT 2560.000 224.070 2560.260 224.390 ;
        RECT 2560.060 2.400 2560.200 224.070 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
=======
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2276.610 25.400 2276.930 25.460 ;
        RECT 2577.910 25.400 2578.230 25.460 ;
        RECT 2276.610 25.260 2578.230 25.400 ;
        RECT 2276.610 25.200 2276.930 25.260 ;
        RECT 2577.910 25.200 2578.230 25.260 ;
      LAYER via ;
        RECT 2276.640 25.200 2276.900 25.460 ;
        RECT 2577.940 25.200 2578.200 25.460 ;
      LAYER met2 ;
        RECT 2272.910 260.170 2273.190 264.000 ;
        RECT 2272.910 260.030 2276.840 260.170 ;
        RECT 2272.910 260.000 2273.190 260.030 ;
        RECT 2276.700 25.490 2276.840 260.030 ;
        RECT 2276.640 25.170 2276.900 25.490 ;
        RECT 2577.940 25.170 2578.200 25.490 ;
        RECT 2578.000 2.400 2578.140 25.170 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
=======
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 502.850 30.840 503.170 30.900 ;
        RECT 811.510 30.840 811.830 30.900 ;
        RECT 502.850 30.700 811.830 30.840 ;
        RECT 502.850 30.640 503.170 30.700 ;
        RECT 811.510 30.640 811.830 30.700 ;
      LAYER via ;
        RECT 502.880 30.640 503.140 30.900 ;
        RECT 811.540 30.640 811.800 30.900 ;
      LAYER met2 ;
        RECT 503.290 260.170 503.570 264.000 ;
        RECT 502.940 260.030 503.570 260.170 ;
        RECT 502.940 30.930 503.080 260.030 ;
        RECT 503.290 260.000 503.570 260.030 ;
        RECT 502.880 30.610 503.140 30.930 ;
        RECT 811.540 30.610 811.800 30.930 ;
        RECT 811.600 2.400 811.740 30.610 ;
        RECT 811.390 -4.800 811.950 2.400 ;
=======
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2290.870 244.020 2291.190 244.080 ;
        RECT 2297.310 244.020 2297.630 244.080 ;
        RECT 2290.870 243.880 2297.630 244.020 ;
        RECT 2290.870 243.820 2291.190 243.880 ;
        RECT 2297.310 243.820 2297.630 243.880 ;
        RECT 2297.310 24.380 2297.630 24.440 ;
        RECT 2595.390 24.380 2595.710 24.440 ;
        RECT 2297.310 24.240 2595.710 24.380 ;
        RECT 2297.310 24.180 2297.630 24.240 ;
        RECT 2595.390 24.180 2595.710 24.240 ;
      LAYER via ;
        RECT 2290.900 243.820 2291.160 244.080 ;
        RECT 2297.340 243.820 2297.600 244.080 ;
        RECT 2297.340 24.180 2297.600 24.440 ;
        RECT 2595.420 24.180 2595.680 24.440 ;
      LAYER met2 ;
        RECT 2290.850 260.000 2291.130 264.000 ;
        RECT 2290.960 244.110 2291.100 260.000 ;
        RECT 2290.900 243.790 2291.160 244.110 ;
        RECT 2297.340 243.790 2297.600 244.110 ;
        RECT 2297.400 24.470 2297.540 243.790 ;
        RECT 2297.340 24.150 2297.600 24.470 ;
        RECT 2595.420 24.150 2595.680 24.470 ;
        RECT 2595.480 2.400 2595.620 24.150 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
=======
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2311.110 24.720 2311.430 24.780 ;
        RECT 2613.330 24.720 2613.650 24.780 ;
        RECT 2311.110 24.580 2613.650 24.720 ;
        RECT 2311.110 24.520 2311.430 24.580 ;
        RECT 2613.330 24.520 2613.650 24.580 ;
      LAYER via ;
        RECT 2311.140 24.520 2311.400 24.780 ;
        RECT 2613.360 24.520 2613.620 24.780 ;
      LAYER met2 ;
        RECT 2308.790 260.170 2309.070 264.000 ;
        RECT 2308.790 260.030 2311.340 260.170 ;
        RECT 2308.790 260.000 2309.070 260.030 ;
        RECT 2311.200 24.810 2311.340 260.030 ;
        RECT 2311.140 24.490 2311.400 24.810 ;
        RECT 2613.360 24.490 2613.620 24.810 ;
        RECT 2613.420 2.400 2613.560 24.490 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
=======
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2326.750 244.020 2327.070 244.080 ;
        RECT 2331.810 244.020 2332.130 244.080 ;
        RECT 2326.750 243.880 2332.130 244.020 ;
        RECT 2326.750 243.820 2327.070 243.880 ;
        RECT 2331.810 243.820 2332.130 243.880 ;
        RECT 2331.810 25.060 2332.130 25.120 ;
        RECT 2631.270 25.060 2631.590 25.120 ;
        RECT 2331.810 24.920 2631.590 25.060 ;
        RECT 2331.810 24.860 2332.130 24.920 ;
        RECT 2631.270 24.860 2631.590 24.920 ;
      LAYER via ;
        RECT 2326.780 243.820 2327.040 244.080 ;
        RECT 2331.840 243.820 2332.100 244.080 ;
        RECT 2331.840 24.860 2332.100 25.120 ;
        RECT 2631.300 24.860 2631.560 25.120 ;
      LAYER met2 ;
        RECT 2326.730 260.000 2327.010 264.000 ;
        RECT 2326.840 244.110 2326.980 260.000 ;
        RECT 2326.780 243.790 2327.040 244.110 ;
        RECT 2331.840 243.790 2332.100 244.110 ;
        RECT 2331.900 25.150 2332.040 243.790 ;
        RECT 2331.840 24.830 2332.100 25.150 ;
        RECT 2631.300 24.830 2631.560 25.150 ;
        RECT 2631.360 2.400 2631.500 24.830 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
=======
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2345.610 72.320 2345.930 72.380 ;
        RECT 2643.230 72.320 2643.550 72.380 ;
        RECT 2345.610 72.180 2643.550 72.320 ;
        RECT 2345.610 72.120 2345.930 72.180 ;
        RECT 2643.230 72.120 2643.550 72.180 ;
        RECT 2643.230 18.940 2643.550 19.000 ;
        RECT 2649.210 18.940 2649.530 19.000 ;
        RECT 2643.230 18.800 2649.530 18.940 ;
        RECT 2643.230 18.740 2643.550 18.800 ;
        RECT 2649.210 18.740 2649.530 18.800 ;
      LAYER via ;
        RECT 2345.640 72.120 2345.900 72.380 ;
        RECT 2643.260 72.120 2643.520 72.380 ;
        RECT 2643.260 18.740 2643.520 19.000 ;
        RECT 2649.240 18.740 2649.500 19.000 ;
      LAYER met2 ;
        RECT 2344.670 260.170 2344.950 264.000 ;
        RECT 2344.670 260.030 2345.840 260.170 ;
        RECT 2344.670 260.000 2344.950 260.030 ;
        RECT 2345.700 72.410 2345.840 260.030 ;
        RECT 2345.640 72.090 2345.900 72.410 ;
        RECT 2643.260 72.090 2643.520 72.410 ;
        RECT 2643.320 19.030 2643.460 72.090 ;
        RECT 2643.260 18.710 2643.520 19.030 ;
        RECT 2649.240 18.710 2649.500 19.030 ;
        RECT 2649.300 2.400 2649.440 18.710 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
=======
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2362.170 243.680 2362.490 243.740 ;
        RECT 2369.990 243.680 2370.310 243.740 ;
        RECT 2362.170 243.540 2370.310 243.680 ;
        RECT 2362.170 243.480 2362.490 243.540 ;
        RECT 2369.990 243.480 2370.310 243.540 ;
        RECT 2369.990 217.160 2370.310 217.220 ;
        RECT 2663.470 217.160 2663.790 217.220 ;
        RECT 2369.990 217.020 2663.790 217.160 ;
        RECT 2369.990 216.960 2370.310 217.020 ;
        RECT 2663.470 216.960 2663.790 217.020 ;
      LAYER via ;
        RECT 2362.200 243.480 2362.460 243.740 ;
        RECT 2370.020 243.480 2370.280 243.740 ;
        RECT 2370.020 216.960 2370.280 217.220 ;
        RECT 2663.500 216.960 2663.760 217.220 ;
      LAYER met2 ;
        RECT 2362.150 260.000 2362.430 264.000 ;
        RECT 2362.260 243.770 2362.400 260.000 ;
        RECT 2362.200 243.450 2362.460 243.770 ;
        RECT 2370.020 243.450 2370.280 243.770 ;
        RECT 2370.080 217.250 2370.220 243.450 ;
        RECT 2370.020 216.930 2370.280 217.250 ;
        RECT 2663.500 216.930 2663.760 217.250 ;
        RECT 2663.560 17.410 2663.700 216.930 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
=======
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2380.110 24.040 2380.430 24.100 ;
        RECT 2684.630 24.040 2684.950 24.100 ;
        RECT 2380.110 23.900 2684.950 24.040 ;
        RECT 2380.110 23.840 2380.430 23.900 ;
        RECT 2684.630 23.840 2684.950 23.900 ;
      LAYER via ;
        RECT 2380.140 23.840 2380.400 24.100 ;
        RECT 2684.660 23.840 2684.920 24.100 ;
      LAYER met2 ;
        RECT 2380.090 260.000 2380.370 264.000 ;
        RECT 2380.200 24.130 2380.340 260.000 ;
        RECT 2380.140 23.810 2380.400 24.130 ;
        RECT 2684.660 23.810 2684.920 24.130 ;
        RECT 2684.720 2.400 2684.860 23.810 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
=======
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2400.810 26.760 2401.130 26.820 ;
        RECT 2702.570 26.760 2702.890 26.820 ;
        RECT 2400.810 26.620 2702.890 26.760 ;
        RECT 2400.810 26.560 2401.130 26.620 ;
        RECT 2702.570 26.560 2702.890 26.620 ;
      LAYER via ;
        RECT 2400.840 26.560 2401.100 26.820 ;
        RECT 2702.600 26.560 2702.860 26.820 ;
      LAYER met2 ;
        RECT 2398.030 260.170 2398.310 264.000 ;
        RECT 2398.030 260.030 2401.040 260.170 ;
        RECT 2398.030 260.000 2398.310 260.030 ;
        RECT 2400.900 26.850 2401.040 260.030 ;
        RECT 2400.840 26.530 2401.100 26.850 ;
        RECT 2702.600 26.530 2702.860 26.850 ;
        RECT 2702.660 2.400 2702.800 26.530 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
=======
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2415.990 244.020 2416.310 244.080 ;
        RECT 2421.510 244.020 2421.830 244.080 ;
        RECT 2415.990 243.880 2421.830 244.020 ;
        RECT 2415.990 243.820 2416.310 243.880 ;
        RECT 2421.510 243.820 2421.830 243.880 ;
        RECT 2421.510 26.420 2421.830 26.480 ;
        RECT 2720.510 26.420 2720.830 26.480 ;
        RECT 2421.510 26.280 2720.830 26.420 ;
        RECT 2421.510 26.220 2421.830 26.280 ;
        RECT 2720.510 26.220 2720.830 26.280 ;
      LAYER via ;
        RECT 2416.020 243.820 2416.280 244.080 ;
        RECT 2421.540 243.820 2421.800 244.080 ;
        RECT 2421.540 26.220 2421.800 26.480 ;
        RECT 2720.540 26.220 2720.800 26.480 ;
      LAYER met2 ;
        RECT 2415.970 260.000 2416.250 264.000 ;
        RECT 2416.080 244.110 2416.220 260.000 ;
        RECT 2416.020 243.790 2416.280 244.110 ;
        RECT 2421.540 243.790 2421.800 244.110 ;
        RECT 2421.600 26.510 2421.740 243.790 ;
        RECT 2421.540 26.190 2421.800 26.510 ;
        RECT 2720.540 26.190 2720.800 26.510 ;
        RECT 2720.600 2.400 2720.740 26.190 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
=======
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2435.310 26.080 2435.630 26.140 ;
        RECT 2738.450 26.080 2738.770 26.140 ;
        RECT 2435.310 25.940 2738.770 26.080 ;
        RECT 2435.310 25.880 2435.630 25.940 ;
        RECT 2738.450 25.880 2738.770 25.940 ;
      LAYER via ;
        RECT 2435.340 25.880 2435.600 26.140 ;
        RECT 2738.480 25.880 2738.740 26.140 ;
      LAYER met2 ;
        RECT 2433.910 260.170 2434.190 264.000 ;
        RECT 2433.910 260.030 2435.540 260.170 ;
        RECT 2433.910 260.000 2434.190 260.030 ;
        RECT 2435.400 26.170 2435.540 260.030 ;
        RECT 2435.340 25.850 2435.600 26.170 ;
        RECT 2738.480 25.850 2738.740 26.170 ;
        RECT 2738.540 2.400 2738.680 25.850 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
=======
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2451.870 238.240 2452.190 238.300 ;
        RECT 2753.170 238.240 2753.490 238.300 ;
        RECT 2451.870 238.100 2753.490 238.240 ;
        RECT 2451.870 238.040 2452.190 238.100 ;
        RECT 2753.170 238.040 2753.490 238.100 ;
      LAYER via ;
        RECT 2451.900 238.040 2452.160 238.300 ;
        RECT 2753.200 238.040 2753.460 238.300 ;
      LAYER met2 ;
        RECT 2451.850 260.000 2452.130 264.000 ;
        RECT 2451.960 238.330 2452.100 260.000 ;
        RECT 2451.900 238.010 2452.160 238.330 ;
        RECT 2753.200 238.010 2753.460 238.330 ;
        RECT 2753.260 17.410 2753.400 238.010 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
=======
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 524.010 38.320 524.330 38.380 ;
        RECT 829.450 38.320 829.770 38.380 ;
        RECT 524.010 38.180 829.770 38.320 ;
        RECT 524.010 38.120 524.330 38.180 ;
        RECT 829.450 38.120 829.770 38.180 ;
      LAYER via ;
        RECT 524.040 38.120 524.300 38.380 ;
        RECT 829.480 38.120 829.740 38.380 ;
      LAYER met2 ;
        RECT 521.230 260.170 521.510 264.000 ;
        RECT 521.230 260.030 524.240 260.170 ;
        RECT 521.230 260.000 521.510 260.030 ;
        RECT 524.100 38.410 524.240 260.030 ;
        RECT 524.040 38.090 524.300 38.410 ;
        RECT 829.480 38.090 829.740 38.410 ;
        RECT 829.540 2.400 829.680 38.090 ;
        RECT 829.330 -4.800 829.890 2.400 ;
=======
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2469.350 210.360 2469.670 210.420 ;
        RECT 2773.870 210.360 2774.190 210.420 ;
        RECT 2469.350 210.220 2774.190 210.360 ;
        RECT 2469.350 210.160 2469.670 210.220 ;
        RECT 2773.870 210.160 2774.190 210.220 ;
      LAYER via ;
        RECT 2469.380 210.160 2469.640 210.420 ;
        RECT 2773.900 210.160 2774.160 210.420 ;
      LAYER met2 ;
        RECT 2469.790 260.170 2470.070 264.000 ;
        RECT 2469.440 260.030 2470.070 260.170 ;
        RECT 2469.440 210.450 2469.580 260.030 ;
        RECT 2469.790 260.000 2470.070 260.030 ;
        RECT 2469.380 210.130 2469.640 210.450 ;
        RECT 2773.900 210.130 2774.160 210.450 ;
        RECT 2773.960 2.400 2774.100 210.130 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
=======
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2487.290 231.100 2487.610 231.160 ;
        RECT 2787.670 231.100 2787.990 231.160 ;
        RECT 2487.290 230.960 2787.990 231.100 ;
        RECT 2487.290 230.900 2487.610 230.960 ;
        RECT 2787.670 230.900 2787.990 230.960 ;
        RECT 2787.670 2.960 2787.990 3.020 ;
        RECT 2791.810 2.960 2792.130 3.020 ;
        RECT 2787.670 2.820 2792.130 2.960 ;
        RECT 2787.670 2.760 2787.990 2.820 ;
        RECT 2791.810 2.760 2792.130 2.820 ;
      LAYER via ;
        RECT 2487.320 230.900 2487.580 231.160 ;
        RECT 2787.700 230.900 2787.960 231.160 ;
        RECT 2787.700 2.760 2787.960 3.020 ;
        RECT 2791.840 2.760 2792.100 3.020 ;
      LAYER met2 ;
        RECT 2487.270 260.000 2487.550 264.000 ;
        RECT 2487.380 231.190 2487.520 260.000 ;
        RECT 2487.320 230.870 2487.580 231.190 ;
        RECT 2787.700 230.870 2787.960 231.190 ;
        RECT 2787.760 3.050 2787.900 230.870 ;
        RECT 2787.700 2.730 2787.960 3.050 ;
        RECT 2791.840 2.730 2792.100 3.050 ;
        RECT 2791.900 2.400 2792.040 2.730 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
=======
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2505.230 244.020 2505.550 244.080 ;
        RECT 2511.210 244.020 2511.530 244.080 ;
        RECT 2505.230 243.880 2511.530 244.020 ;
        RECT 2505.230 243.820 2505.550 243.880 ;
        RECT 2511.210 243.820 2511.530 243.880 ;
        RECT 2511.210 30.840 2511.530 30.900 ;
        RECT 2809.750 30.840 2810.070 30.900 ;
        RECT 2511.210 30.700 2810.070 30.840 ;
        RECT 2511.210 30.640 2511.530 30.700 ;
        RECT 2809.750 30.640 2810.070 30.700 ;
      LAYER via ;
        RECT 2505.260 243.820 2505.520 244.080 ;
        RECT 2511.240 243.820 2511.500 244.080 ;
        RECT 2511.240 30.640 2511.500 30.900 ;
        RECT 2809.780 30.640 2810.040 30.900 ;
      LAYER met2 ;
        RECT 2505.210 260.000 2505.490 264.000 ;
        RECT 2505.320 244.110 2505.460 260.000 ;
        RECT 2505.260 243.790 2505.520 244.110 ;
        RECT 2511.240 243.790 2511.500 244.110 ;
        RECT 2511.300 30.930 2511.440 243.790 ;
        RECT 2511.240 30.610 2511.500 30.930 ;
        RECT 2809.780 30.610 2810.040 30.930 ;
        RECT 2809.840 2.400 2809.980 30.610 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
=======
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2525.010 79.460 2525.330 79.520 ;
        RECT 2822.170 79.460 2822.490 79.520 ;
        RECT 2525.010 79.320 2822.490 79.460 ;
        RECT 2525.010 79.260 2525.330 79.320 ;
        RECT 2822.170 79.260 2822.490 79.320 ;
        RECT 2822.170 2.960 2822.490 3.020 ;
        RECT 2827.690 2.960 2828.010 3.020 ;
        RECT 2822.170 2.820 2828.010 2.960 ;
        RECT 2822.170 2.760 2822.490 2.820 ;
        RECT 2827.690 2.760 2828.010 2.820 ;
      LAYER via ;
        RECT 2525.040 79.260 2525.300 79.520 ;
        RECT 2822.200 79.260 2822.460 79.520 ;
        RECT 2822.200 2.760 2822.460 3.020 ;
        RECT 2827.720 2.760 2827.980 3.020 ;
      LAYER met2 ;
        RECT 2523.150 260.170 2523.430 264.000 ;
        RECT 2523.150 260.030 2525.240 260.170 ;
        RECT 2523.150 260.000 2523.430 260.030 ;
        RECT 2525.100 79.550 2525.240 260.030 ;
        RECT 2525.040 79.230 2525.300 79.550 ;
        RECT 2822.200 79.230 2822.460 79.550 ;
        RECT 2822.260 3.050 2822.400 79.230 ;
        RECT 2822.200 2.730 2822.460 3.050 ;
        RECT 2827.720 2.730 2827.980 3.050 ;
        RECT 2827.780 2.400 2827.920 2.730 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
=======
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2541.110 244.020 2541.430 244.080 ;
        RECT 2545.710 244.020 2546.030 244.080 ;
        RECT 2541.110 243.880 2546.030 244.020 ;
        RECT 2541.110 243.820 2541.430 243.880 ;
        RECT 2545.710 243.820 2546.030 243.880 ;
        RECT 2545.710 224.640 2546.030 224.700 ;
        RECT 2842.870 224.640 2843.190 224.700 ;
        RECT 2545.710 224.500 2843.190 224.640 ;
        RECT 2545.710 224.440 2546.030 224.500 ;
        RECT 2842.870 224.440 2843.190 224.500 ;
      LAYER via ;
        RECT 2541.140 243.820 2541.400 244.080 ;
        RECT 2545.740 243.820 2546.000 244.080 ;
        RECT 2545.740 224.440 2546.000 224.700 ;
        RECT 2842.900 224.440 2843.160 224.700 ;
      LAYER met2 ;
        RECT 2541.090 260.000 2541.370 264.000 ;
        RECT 2541.200 244.110 2541.340 260.000 ;
        RECT 2541.140 243.790 2541.400 244.110 ;
        RECT 2545.740 243.790 2546.000 244.110 ;
        RECT 2545.800 224.730 2545.940 243.790 ;
        RECT 2545.740 224.410 2546.000 224.730 ;
        RECT 2842.900 224.410 2843.160 224.730 ;
        RECT 2842.960 6.530 2843.100 224.410 ;
        RECT 2842.960 6.390 2845.400 6.530 ;
        RECT 2845.260 2.400 2845.400 6.390 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
=======
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2559.050 196.760 2559.370 196.820 ;
        RECT 2857.130 196.760 2857.450 196.820 ;
        RECT 2559.050 196.620 2857.450 196.760 ;
        RECT 2559.050 196.560 2559.370 196.620 ;
        RECT 2857.130 196.560 2857.450 196.620 ;
        RECT 2857.130 17.580 2857.450 17.640 ;
        RECT 2863.110 17.580 2863.430 17.640 ;
        RECT 2857.130 17.440 2863.430 17.580 ;
        RECT 2857.130 17.380 2857.450 17.440 ;
        RECT 2863.110 17.380 2863.430 17.440 ;
      LAYER via ;
        RECT 2559.080 196.560 2559.340 196.820 ;
        RECT 2857.160 196.560 2857.420 196.820 ;
        RECT 2857.160 17.380 2857.420 17.640 ;
        RECT 2863.140 17.380 2863.400 17.640 ;
      LAYER met2 ;
        RECT 2559.030 260.000 2559.310 264.000 ;
        RECT 2559.140 196.850 2559.280 260.000 ;
        RECT 2559.080 196.530 2559.340 196.850 ;
        RECT 2857.160 196.530 2857.420 196.850 ;
        RECT 2857.220 17.670 2857.360 196.530 ;
        RECT 2857.160 17.350 2857.420 17.670 ;
        RECT 2863.140 17.350 2863.400 17.670 ;
        RECT 2863.200 2.400 2863.340 17.350 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
=======
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2580.210 51.580 2580.530 51.640 ;
        RECT 2877.370 51.580 2877.690 51.640 ;
        RECT 2580.210 51.440 2877.690 51.580 ;
        RECT 2580.210 51.380 2580.530 51.440 ;
        RECT 2877.370 51.380 2877.690 51.440 ;
      LAYER via ;
        RECT 2580.240 51.380 2580.500 51.640 ;
        RECT 2877.400 51.380 2877.660 51.640 ;
      LAYER met2 ;
        RECT 2576.970 260.170 2577.250 264.000 ;
        RECT 2576.970 260.030 2580.440 260.170 ;
        RECT 2576.970 260.000 2577.250 260.030 ;
        RECT 2580.300 51.670 2580.440 260.030 ;
        RECT 2580.240 51.350 2580.500 51.670 ;
        RECT 2877.400 51.350 2877.660 51.670 ;
        RECT 2877.460 17.410 2877.600 51.350 ;
        RECT 2877.460 17.270 2881.280 17.410 ;
        RECT 2881.140 2.400 2881.280 17.270 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
=======
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2594.930 244.020 2595.250 244.080 ;
        RECT 2600.450 244.020 2600.770 244.080 ;
        RECT 2594.930 243.880 2600.770 244.020 ;
        RECT 2594.930 243.820 2595.250 243.880 ;
        RECT 2600.450 243.820 2600.770 243.880 ;
        RECT 2600.450 189.620 2600.770 189.680 ;
        RECT 2894.390 189.620 2894.710 189.680 ;
        RECT 2600.450 189.480 2894.710 189.620 ;
        RECT 2600.450 189.420 2600.770 189.480 ;
        RECT 2894.390 189.420 2894.710 189.480 ;
        RECT 2894.390 17.580 2894.710 17.640 ;
        RECT 2898.990 17.580 2899.310 17.640 ;
        RECT 2894.390 17.440 2899.310 17.580 ;
        RECT 2894.390 17.380 2894.710 17.440 ;
        RECT 2898.990 17.380 2899.310 17.440 ;
      LAYER via ;
        RECT 2594.960 243.820 2595.220 244.080 ;
        RECT 2600.480 243.820 2600.740 244.080 ;
        RECT 2600.480 189.420 2600.740 189.680 ;
        RECT 2894.420 189.420 2894.680 189.680 ;
        RECT 2894.420 17.380 2894.680 17.640 ;
        RECT 2899.020 17.380 2899.280 17.640 ;
      LAYER met2 ;
        RECT 2594.910 260.000 2595.190 264.000 ;
        RECT 2595.020 244.110 2595.160 260.000 ;
        RECT 2594.960 243.790 2595.220 244.110 ;
        RECT 2600.480 243.790 2600.740 244.110 ;
        RECT 2600.540 189.710 2600.680 243.790 ;
        RECT 2600.480 189.390 2600.740 189.710 ;
        RECT 2894.420 189.390 2894.680 189.710 ;
        RECT 2894.480 17.670 2894.620 189.390 ;
        RECT 2894.420 17.350 2894.680 17.670 ;
        RECT 2899.020 17.350 2899.280 17.670 ;
        RECT 2899.080 2.400 2899.220 17.350 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
=======
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 539.190 244.020 539.510 244.080 ;
        RECT 544.710 244.020 545.030 244.080 ;
        RECT 539.190 243.880 545.030 244.020 ;
        RECT 539.190 243.820 539.510 243.880 ;
        RECT 544.710 243.820 545.030 243.880 ;
        RECT 544.710 44.780 545.030 44.840 ;
        RECT 846.930 44.780 847.250 44.840 ;
        RECT 544.710 44.640 847.250 44.780 ;
        RECT 544.710 44.580 545.030 44.640 ;
        RECT 846.930 44.580 847.250 44.640 ;
      LAYER via ;
        RECT 539.220 243.820 539.480 244.080 ;
        RECT 544.740 243.820 545.000 244.080 ;
        RECT 544.740 44.580 545.000 44.840 ;
        RECT 846.960 44.580 847.220 44.840 ;
      LAYER met2 ;
        RECT 539.170 260.000 539.450 264.000 ;
        RECT 539.280 244.110 539.420 260.000 ;
        RECT 539.220 243.790 539.480 244.110 ;
        RECT 544.740 243.790 545.000 244.110 ;
        RECT 544.800 44.870 544.940 243.790 ;
        RECT 544.740 44.550 545.000 44.870 ;
        RECT 846.960 44.550 847.220 44.870 ;
        RECT 847.020 2.400 847.160 44.550 ;
        RECT 846.810 -4.800 847.370 2.400 ;
=======
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 558.510 51.580 558.830 51.640 ;
        RECT 862.570 51.580 862.890 51.640 ;
        RECT 558.510 51.440 862.890 51.580 ;
        RECT 558.510 51.380 558.830 51.440 ;
        RECT 862.570 51.380 862.890 51.440 ;
      LAYER via ;
        RECT 558.540 51.380 558.800 51.640 ;
        RECT 862.600 51.380 862.860 51.640 ;
      LAYER met2 ;
        RECT 557.110 260.170 557.390 264.000 ;
        RECT 557.110 260.030 558.740 260.170 ;
        RECT 557.110 260.000 557.390 260.030 ;
        RECT 558.600 51.670 558.740 260.030 ;
        RECT 558.540 51.350 558.800 51.670 ;
        RECT 862.600 51.350 862.860 51.670 ;
        RECT 862.660 16.730 862.800 51.350 ;
        RECT 862.660 16.590 865.100 16.730 ;
        RECT 864.960 2.400 865.100 16.590 ;
        RECT 864.750 -4.800 865.310 2.400 ;
=======
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 574.610 244.020 574.930 244.080 ;
        RECT 579.210 244.020 579.530 244.080 ;
        RECT 574.610 243.880 579.530 244.020 ;
        RECT 574.610 243.820 574.930 243.880 ;
        RECT 579.210 243.820 579.530 243.880 ;
        RECT 579.210 58.720 579.530 58.780 ;
        RECT 876.830 58.720 877.150 58.780 ;
        RECT 579.210 58.580 877.150 58.720 ;
        RECT 579.210 58.520 579.530 58.580 ;
        RECT 876.830 58.520 877.150 58.580 ;
        RECT 876.830 16.560 877.150 16.620 ;
        RECT 882.810 16.560 883.130 16.620 ;
        RECT 876.830 16.420 883.130 16.560 ;
        RECT 876.830 16.360 877.150 16.420 ;
        RECT 882.810 16.360 883.130 16.420 ;
      LAYER via ;
        RECT 574.640 243.820 574.900 244.080 ;
        RECT 579.240 243.820 579.500 244.080 ;
        RECT 579.240 58.520 579.500 58.780 ;
        RECT 876.860 58.520 877.120 58.780 ;
        RECT 876.860 16.360 877.120 16.620 ;
        RECT 882.840 16.360 883.100 16.620 ;
      LAYER met2 ;
        RECT 574.590 260.000 574.870 264.000 ;
        RECT 574.700 244.110 574.840 260.000 ;
        RECT 574.640 243.790 574.900 244.110 ;
        RECT 579.240 243.790 579.500 244.110 ;
        RECT 579.300 58.810 579.440 243.790 ;
        RECT 579.240 58.490 579.500 58.810 ;
        RECT 876.860 58.490 877.120 58.810 ;
        RECT 876.920 16.650 877.060 58.490 ;
        RECT 876.860 16.330 877.120 16.650 ;
        RECT 882.840 16.330 883.100 16.650 ;
        RECT 882.900 2.400 883.040 16.330 ;
        RECT 882.690 -4.800 883.250 2.400 ;
=======
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 592.550 65.520 592.870 65.580 ;
        RECT 897.070 65.520 897.390 65.580 ;
        RECT 592.550 65.380 897.390 65.520 ;
        RECT 592.550 65.320 592.870 65.380 ;
        RECT 897.070 65.320 897.390 65.380 ;
      LAYER via ;
        RECT 592.580 65.320 592.840 65.580 ;
        RECT 897.100 65.320 897.360 65.580 ;
      LAYER met2 ;
        RECT 592.530 260.000 592.810 264.000 ;
        RECT 592.640 65.610 592.780 260.000 ;
        RECT 592.580 65.290 592.840 65.610 ;
        RECT 897.100 65.290 897.360 65.610 ;
        RECT 897.160 16.730 897.300 65.290 ;
        RECT 897.160 16.590 900.980 16.730 ;
        RECT 900.840 2.400 900.980 16.590 ;
        RECT 900.630 -4.800 901.190 2.400 ;
=======
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 613.710 72.320 614.030 72.380 ;
        RECT 918.230 72.320 918.550 72.380 ;
        RECT 613.710 72.180 918.550 72.320 ;
        RECT 613.710 72.120 614.030 72.180 ;
        RECT 918.230 72.120 918.550 72.180 ;
      LAYER via ;
        RECT 613.740 72.120 614.000 72.380 ;
        RECT 918.260 72.120 918.520 72.380 ;
      LAYER met2 ;
        RECT 610.470 260.170 610.750 264.000 ;
        RECT 610.470 260.030 613.940 260.170 ;
        RECT 610.470 260.000 610.750 260.030 ;
        RECT 613.800 72.410 613.940 260.030 ;
        RECT 613.740 72.090 614.000 72.410 ;
        RECT 918.260 72.090 918.520 72.410 ;
        RECT 918.320 17.410 918.460 72.090 ;
        RECT 918.320 17.270 918.920 17.410 ;
        RECT 918.780 2.400 918.920 17.270 ;
        RECT 918.570 -4.800 919.130 2.400 ;
=======
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 628.430 243.340 628.750 243.400 ;
        RECT 634.410 243.340 634.730 243.400 ;
        RECT 628.430 243.200 634.730 243.340 ;
        RECT 628.430 243.140 628.750 243.200 ;
        RECT 634.410 243.140 634.730 243.200 ;
        RECT 634.410 79.800 634.730 79.860 ;
        RECT 931.570 79.800 931.890 79.860 ;
        RECT 634.410 79.660 931.890 79.800 ;
        RECT 634.410 79.600 634.730 79.660 ;
        RECT 931.570 79.600 931.890 79.660 ;
      LAYER via ;
        RECT 628.460 243.140 628.720 243.400 ;
        RECT 634.440 243.140 634.700 243.400 ;
        RECT 634.440 79.600 634.700 79.860 ;
        RECT 931.600 79.600 931.860 79.860 ;
      LAYER met2 ;
        RECT 628.410 260.000 628.690 264.000 ;
        RECT 628.520 243.430 628.660 260.000 ;
        RECT 628.460 243.110 628.720 243.430 ;
        RECT 634.440 243.110 634.700 243.430 ;
        RECT 634.500 79.890 634.640 243.110 ;
        RECT 634.440 79.570 634.700 79.890 ;
        RECT 931.600 79.570 931.860 79.890 ;
        RECT 931.660 16.730 931.800 79.570 ;
        RECT 931.660 16.590 936.400 16.730 ;
        RECT 936.260 2.400 936.400 16.590 ;
        RECT 936.050 -4.800 936.610 2.400 ;
=======
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 648.210 86.260 648.530 86.320 ;
        RECT 952.270 86.260 952.590 86.320 ;
        RECT 648.210 86.120 952.590 86.260 ;
        RECT 648.210 86.060 648.530 86.120 ;
        RECT 952.270 86.060 952.590 86.120 ;
      LAYER via ;
        RECT 648.240 86.060 648.500 86.320 ;
        RECT 952.300 86.060 952.560 86.320 ;
      LAYER met2 ;
        RECT 646.350 260.170 646.630 264.000 ;
        RECT 646.350 260.030 648.440 260.170 ;
        RECT 646.350 260.000 646.630 260.030 ;
        RECT 648.300 86.350 648.440 260.030 ;
        RECT 648.240 86.030 648.500 86.350 ;
        RECT 952.300 86.030 952.560 86.350 ;
        RECT 952.360 16.730 952.500 86.030 ;
        RECT 952.360 16.590 954.340 16.730 ;
        RECT 954.200 2.400 954.340 16.590 ;
        RECT 953.990 -4.800 954.550 2.400 ;
=======
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 664.310 244.020 664.630 244.080 ;
        RECT 668.910 244.020 669.230 244.080 ;
        RECT 664.310 243.880 669.230 244.020 ;
        RECT 664.310 243.820 664.630 243.880 ;
        RECT 668.910 243.820 669.230 243.880 ;
        RECT 668.910 24.720 669.230 24.780 ;
        RECT 972.050 24.720 972.370 24.780 ;
        RECT 668.910 24.580 972.370 24.720 ;
        RECT 668.910 24.520 669.230 24.580 ;
        RECT 972.050 24.520 972.370 24.580 ;
      LAYER via ;
        RECT 664.340 243.820 664.600 244.080 ;
        RECT 668.940 243.820 669.200 244.080 ;
        RECT 668.940 24.520 669.200 24.780 ;
        RECT 972.080 24.520 972.340 24.780 ;
      LAYER met2 ;
        RECT 664.290 260.000 664.570 264.000 ;
        RECT 664.400 244.110 664.540 260.000 ;
        RECT 664.340 243.790 664.600 244.110 ;
        RECT 668.940 243.790 669.200 244.110 ;
        RECT 669.000 24.810 669.140 243.790 ;
        RECT 668.940 24.490 669.200 24.810 ;
        RECT 972.080 24.490 972.340 24.810 ;
        RECT 972.140 2.400 972.280 24.490 ;
        RECT 971.930 -4.800 972.490 2.400 ;
=======
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 344.610 24.040 344.930 24.100 ;
        RECT 650.970 24.040 651.290 24.100 ;
        RECT 344.610 23.900 651.290 24.040 ;
        RECT 344.610 23.840 344.930 23.900 ;
        RECT 650.970 23.840 651.290 23.900 ;
      LAYER via ;
        RECT 344.640 23.840 344.900 24.100 ;
        RECT 651.000 23.840 651.260 24.100 ;
      LAYER met2 ;
        RECT 342.290 260.170 342.570 264.000 ;
        RECT 342.290 260.030 344.840 260.170 ;
        RECT 342.290 260.000 342.570 260.030 ;
        RECT 344.700 24.130 344.840 260.030 ;
        RECT 344.640 23.810 344.900 24.130 ;
        RECT 651.000 23.810 651.260 24.130 ;
        RECT 651.060 2.400 651.200 23.810 ;
        RECT 650.850 -4.800 651.410 2.400 ;
=======
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 682.710 237.900 683.030 237.960 ;
        RECT 986.770 237.900 987.090 237.960 ;
        RECT 682.710 237.760 987.090 237.900 ;
        RECT 682.710 237.700 683.030 237.760 ;
        RECT 986.770 237.700 987.090 237.760 ;
      LAYER via ;
        RECT 682.740 237.700 683.000 237.960 ;
        RECT 986.800 237.700 987.060 237.960 ;
      LAYER met2 ;
        RECT 682.230 260.170 682.510 264.000 ;
        RECT 682.230 260.030 682.940 260.170 ;
        RECT 682.230 260.000 682.510 260.030 ;
        RECT 682.800 237.990 682.940 260.030 ;
        RECT 682.740 237.670 683.000 237.990 ;
        RECT 986.800 237.670 987.060 237.990 ;
        RECT 986.860 16.730 987.000 237.670 ;
        RECT 986.860 16.590 990.220 16.730 ;
        RECT 990.080 2.400 990.220 16.590 ;
        RECT 989.870 -4.800 990.430 2.400 ;
=======
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 703.410 93.060 703.730 93.120 ;
        RECT 1007.930 93.060 1008.250 93.120 ;
        RECT 703.410 92.920 1008.250 93.060 ;
        RECT 703.410 92.860 703.730 92.920 ;
        RECT 1007.930 92.860 1008.250 92.920 ;
      LAYER via ;
        RECT 703.440 92.860 703.700 93.120 ;
        RECT 1007.960 92.860 1008.220 93.120 ;
      LAYER met2 ;
        RECT 699.710 260.170 699.990 264.000 ;
        RECT 699.710 260.030 703.640 260.170 ;
        RECT 699.710 260.000 699.990 260.030 ;
        RECT 703.500 93.150 703.640 260.030 ;
        RECT 703.440 92.830 703.700 93.150 ;
        RECT 1007.960 92.830 1008.220 93.150 ;
        RECT 1008.020 17.410 1008.160 92.830 ;
        RECT 1007.560 17.270 1008.160 17.410 ;
        RECT 1007.560 2.400 1007.700 17.270 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
=======
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 717.670 242.660 717.990 242.720 ;
        RECT 724.110 242.660 724.430 242.720 ;
        RECT 717.670 242.520 724.430 242.660 ;
        RECT 717.670 242.460 717.990 242.520 ;
        RECT 724.110 242.460 724.430 242.520 ;
        RECT 724.110 99.860 724.430 99.920 ;
        RECT 1021.270 99.860 1021.590 99.920 ;
        RECT 724.110 99.720 1021.590 99.860 ;
        RECT 724.110 99.660 724.430 99.720 ;
        RECT 1021.270 99.660 1021.590 99.720 ;
      LAYER via ;
        RECT 717.700 242.460 717.960 242.720 ;
        RECT 724.140 242.460 724.400 242.720 ;
        RECT 724.140 99.660 724.400 99.920 ;
        RECT 1021.300 99.660 1021.560 99.920 ;
      LAYER met2 ;
        RECT 717.650 260.000 717.930 264.000 ;
        RECT 717.760 242.750 717.900 260.000 ;
        RECT 717.700 242.430 717.960 242.750 ;
        RECT 724.140 242.430 724.400 242.750 ;
        RECT 724.200 99.950 724.340 242.430 ;
        RECT 724.140 99.630 724.400 99.950 ;
        RECT 1021.300 99.630 1021.560 99.950 ;
        RECT 1021.360 16.730 1021.500 99.630 ;
        RECT 1021.360 16.590 1025.640 16.730 ;
        RECT 1025.500 2.400 1025.640 16.590 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
=======
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 737.910 107.000 738.230 107.060 ;
        RECT 1041.970 107.000 1042.290 107.060 ;
        RECT 737.910 106.860 1042.290 107.000 ;
        RECT 737.910 106.800 738.230 106.860 ;
        RECT 1041.970 106.800 1042.290 106.860 ;
      LAYER via ;
        RECT 737.940 106.800 738.200 107.060 ;
        RECT 1042.000 106.800 1042.260 107.060 ;
      LAYER met2 ;
        RECT 735.590 260.170 735.870 264.000 ;
        RECT 735.590 260.030 738.140 260.170 ;
        RECT 735.590 260.000 735.870 260.030 ;
        RECT 738.000 107.090 738.140 260.030 ;
        RECT 737.940 106.770 738.200 107.090 ;
        RECT 1042.000 106.770 1042.260 107.090 ;
        RECT 1042.060 16.730 1042.200 106.770 ;
        RECT 1042.060 16.590 1043.580 16.730 ;
        RECT 1043.440 2.400 1043.580 16.590 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
=======
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 753.550 244.020 753.870 244.080 ;
        RECT 758.610 244.020 758.930 244.080 ;
        RECT 753.550 243.880 758.930 244.020 ;
        RECT 753.550 243.820 753.870 243.880 ;
        RECT 758.610 243.820 758.930 243.880 ;
        RECT 758.610 113.800 758.930 113.860 ;
        RECT 1055.770 113.800 1056.090 113.860 ;
        RECT 758.610 113.660 1056.090 113.800 ;
        RECT 758.610 113.600 758.930 113.660 ;
        RECT 1055.770 113.600 1056.090 113.660 ;
      LAYER via ;
        RECT 753.580 243.820 753.840 244.080 ;
        RECT 758.640 243.820 758.900 244.080 ;
        RECT 758.640 113.600 758.900 113.860 ;
        RECT 1055.800 113.600 1056.060 113.860 ;
      LAYER met2 ;
        RECT 753.530 260.000 753.810 264.000 ;
        RECT 753.640 244.110 753.780 260.000 ;
        RECT 753.580 243.790 753.840 244.110 ;
        RECT 758.640 243.790 758.900 244.110 ;
        RECT 758.700 113.890 758.840 243.790 ;
        RECT 758.640 113.570 758.900 113.890 ;
        RECT 1055.800 113.570 1056.060 113.890 ;
        RECT 1055.860 16.730 1056.000 113.570 ;
        RECT 1055.860 16.590 1061.520 16.730 ;
        RECT 1061.380 2.400 1061.520 16.590 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
=======
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 772.410 120.600 772.730 120.660 ;
        RECT 1076.470 120.600 1076.790 120.660 ;
        RECT 772.410 120.460 1076.790 120.600 ;
        RECT 772.410 120.400 772.730 120.460 ;
        RECT 1076.470 120.400 1076.790 120.460 ;
      LAYER via ;
        RECT 772.440 120.400 772.700 120.660 ;
        RECT 1076.500 120.400 1076.760 120.660 ;
      LAYER met2 ;
        RECT 771.470 260.170 771.750 264.000 ;
        RECT 771.470 260.030 772.640 260.170 ;
        RECT 771.470 260.000 771.750 260.030 ;
        RECT 772.500 120.690 772.640 260.030 ;
        RECT 772.440 120.370 772.700 120.690 ;
        RECT 1076.500 120.370 1076.760 120.690 ;
        RECT 1076.560 16.730 1076.700 120.370 ;
        RECT 1076.560 16.590 1079.460 16.730 ;
        RECT 1079.320 2.400 1079.460 16.590 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
=======
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 789.430 244.020 789.750 244.080 ;
        RECT 793.110 244.020 793.430 244.080 ;
        RECT 789.430 243.880 793.430 244.020 ;
        RECT 789.430 243.820 789.750 243.880 ;
        RECT 793.110 243.820 793.430 243.880 ;
        RECT 793.110 127.740 793.430 127.800 ;
        RECT 1090.730 127.740 1091.050 127.800 ;
        RECT 793.110 127.600 1091.050 127.740 ;
        RECT 793.110 127.540 793.430 127.600 ;
        RECT 1090.730 127.540 1091.050 127.600 ;
        RECT 1090.730 17.920 1091.050 17.980 ;
        RECT 1096.710 17.920 1097.030 17.980 ;
        RECT 1090.730 17.780 1097.030 17.920 ;
        RECT 1090.730 17.720 1091.050 17.780 ;
        RECT 1096.710 17.720 1097.030 17.780 ;
      LAYER via ;
        RECT 789.460 243.820 789.720 244.080 ;
        RECT 793.140 243.820 793.400 244.080 ;
        RECT 793.140 127.540 793.400 127.800 ;
        RECT 1090.760 127.540 1091.020 127.800 ;
        RECT 1090.760 17.720 1091.020 17.980 ;
        RECT 1096.740 17.720 1097.000 17.980 ;
      LAYER met2 ;
        RECT 789.410 260.000 789.690 264.000 ;
        RECT 789.520 244.110 789.660 260.000 ;
        RECT 789.460 243.790 789.720 244.110 ;
        RECT 793.140 243.790 793.400 244.110 ;
        RECT 793.200 127.830 793.340 243.790 ;
        RECT 793.140 127.510 793.400 127.830 ;
        RECT 1090.760 127.510 1091.020 127.830 ;
        RECT 1090.820 18.010 1090.960 127.510 ;
        RECT 1090.760 17.690 1091.020 18.010 ;
        RECT 1096.740 17.690 1097.000 18.010 ;
        RECT 1096.800 2.400 1096.940 17.690 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
=======
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 807.370 244.020 807.690 244.080 ;
        RECT 813.810 244.020 814.130 244.080 ;
        RECT 807.370 243.880 814.130 244.020 ;
        RECT 807.370 243.820 807.690 243.880 ;
        RECT 813.810 243.820 814.130 243.880 ;
        RECT 813.810 31.520 814.130 31.580 ;
        RECT 1114.650 31.520 1114.970 31.580 ;
        RECT 813.810 31.380 1114.970 31.520 ;
        RECT 813.810 31.320 814.130 31.380 ;
        RECT 1114.650 31.320 1114.970 31.380 ;
      LAYER via ;
        RECT 807.400 243.820 807.660 244.080 ;
        RECT 813.840 243.820 814.100 244.080 ;
        RECT 813.840 31.320 814.100 31.580 ;
        RECT 1114.680 31.320 1114.940 31.580 ;
      LAYER met2 ;
        RECT 807.350 260.000 807.630 264.000 ;
        RECT 807.460 244.110 807.600 260.000 ;
        RECT 807.400 243.790 807.660 244.110 ;
        RECT 813.840 243.790 814.100 244.110 ;
        RECT 813.900 31.610 814.040 243.790 ;
        RECT 813.840 31.290 814.100 31.610 ;
        RECT 1114.680 31.290 1114.940 31.610 ;
        RECT 1114.740 2.400 1114.880 31.290 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
=======
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 827.610 134.540 827.930 134.600 ;
        RECT 1131.670 134.540 1131.990 134.600 ;
        RECT 827.610 134.400 1131.990 134.540 ;
        RECT 827.610 134.340 827.930 134.400 ;
        RECT 1131.670 134.340 1131.990 134.400 ;
      LAYER via ;
        RECT 827.640 134.340 827.900 134.600 ;
        RECT 1131.700 134.340 1131.960 134.600 ;
      LAYER met2 ;
        RECT 824.830 260.170 825.110 264.000 ;
        RECT 824.830 260.030 827.840 260.170 ;
        RECT 824.830 260.000 825.110 260.030 ;
        RECT 827.700 134.630 827.840 260.030 ;
        RECT 827.640 134.310 827.900 134.630 ;
        RECT 1131.700 134.310 1131.960 134.630 ;
        RECT 1131.760 16.730 1131.900 134.310 ;
        RECT 1131.760 16.590 1132.820 16.730 ;
        RECT 1132.680 2.400 1132.820 16.590 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
=======
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 842.790 244.020 843.110 244.080 ;
        RECT 848.310 244.020 848.630 244.080 ;
        RECT 842.790 243.880 848.630 244.020 ;
        RECT 842.790 243.820 843.110 243.880 ;
        RECT 848.310 243.820 848.630 243.880 ;
        RECT 848.310 38.320 848.630 38.380 ;
        RECT 1150.530 38.320 1150.850 38.380 ;
        RECT 848.310 38.180 1150.850 38.320 ;
        RECT 848.310 38.120 848.630 38.180 ;
        RECT 1150.530 38.120 1150.850 38.180 ;
      LAYER via ;
        RECT 842.820 243.820 843.080 244.080 ;
        RECT 848.340 243.820 848.600 244.080 ;
        RECT 848.340 38.120 848.600 38.380 ;
        RECT 1150.560 38.120 1150.820 38.380 ;
      LAYER met2 ;
        RECT 842.770 260.000 843.050 264.000 ;
        RECT 842.880 244.110 843.020 260.000 ;
        RECT 842.820 243.790 843.080 244.110 ;
        RECT 848.340 243.790 848.600 244.110 ;
        RECT 848.400 38.410 848.540 243.790 ;
        RECT 848.340 38.090 848.600 38.410 ;
        RECT 1150.560 38.090 1150.820 38.410 ;
        RECT 1150.620 2.400 1150.760 38.090 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
=======
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 360.250 244.020 360.570 244.080 ;
        RECT 365.310 244.020 365.630 244.080 ;
        RECT 360.250 243.880 365.630 244.020 ;
        RECT 360.250 243.820 360.570 243.880 ;
        RECT 365.310 243.820 365.630 243.880 ;
        RECT 365.310 93.060 365.630 93.120 ;
        RECT 662.930 93.060 663.250 93.120 ;
        RECT 365.310 92.920 663.250 93.060 ;
        RECT 365.310 92.860 365.630 92.920 ;
        RECT 662.930 92.860 663.250 92.920 ;
        RECT 662.930 20.300 663.250 20.360 ;
        RECT 668.910 20.300 669.230 20.360 ;
        RECT 662.930 20.160 669.230 20.300 ;
        RECT 662.930 20.100 663.250 20.160 ;
        RECT 668.910 20.100 669.230 20.160 ;
      LAYER via ;
        RECT 360.280 243.820 360.540 244.080 ;
        RECT 365.340 243.820 365.600 244.080 ;
        RECT 365.340 92.860 365.600 93.120 ;
        RECT 662.960 92.860 663.220 93.120 ;
        RECT 662.960 20.100 663.220 20.360 ;
        RECT 668.940 20.100 669.200 20.360 ;
      LAYER met2 ;
        RECT 360.230 260.000 360.510 264.000 ;
        RECT 360.340 244.110 360.480 260.000 ;
        RECT 360.280 243.790 360.540 244.110 ;
        RECT 365.340 243.790 365.600 244.110 ;
        RECT 365.400 93.150 365.540 243.790 ;
        RECT 365.340 92.830 365.600 93.150 ;
        RECT 662.960 92.830 663.220 93.150 ;
        RECT 663.020 20.390 663.160 92.830 ;
        RECT 662.960 20.070 663.220 20.390 ;
        RECT 668.940 20.070 669.200 20.390 ;
        RECT 669.000 2.400 669.140 20.070 ;
        RECT 668.790 -4.800 669.350 2.400 ;
=======
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 862.110 44.780 862.430 44.840 ;
        RECT 1168.470 44.780 1168.790 44.840 ;
        RECT 862.110 44.640 1168.790 44.780 ;
        RECT 862.110 44.580 862.430 44.640 ;
        RECT 1168.470 44.580 1168.790 44.640 ;
      LAYER via ;
        RECT 862.140 44.580 862.400 44.840 ;
        RECT 1168.500 44.580 1168.760 44.840 ;
      LAYER met2 ;
        RECT 860.710 260.170 860.990 264.000 ;
        RECT 860.710 260.030 862.340 260.170 ;
        RECT 860.710 260.000 860.990 260.030 ;
        RECT 862.200 44.870 862.340 260.030 ;
        RECT 862.140 44.550 862.400 44.870 ;
        RECT 1168.500 44.550 1168.760 44.870 ;
        RECT 1168.560 2.400 1168.700 44.550 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
=======
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 878.670 244.020 878.990 244.080 ;
        RECT 882.810 244.020 883.130 244.080 ;
        RECT 878.670 243.880 883.130 244.020 ;
        RECT 878.670 243.820 878.990 243.880 ;
        RECT 882.810 243.820 883.130 243.880 ;
        RECT 882.810 51.920 883.130 51.980 ;
        RECT 1180.430 51.920 1180.750 51.980 ;
        RECT 882.810 51.780 1180.750 51.920 ;
        RECT 882.810 51.720 883.130 51.780 ;
        RECT 1180.430 51.720 1180.750 51.780 ;
        RECT 1180.430 17.920 1180.750 17.980 ;
        RECT 1185.950 17.920 1186.270 17.980 ;
        RECT 1180.430 17.780 1186.270 17.920 ;
        RECT 1180.430 17.720 1180.750 17.780 ;
        RECT 1185.950 17.720 1186.270 17.780 ;
      LAYER via ;
        RECT 878.700 243.820 878.960 244.080 ;
        RECT 882.840 243.820 883.100 244.080 ;
        RECT 882.840 51.720 883.100 51.980 ;
        RECT 1180.460 51.720 1180.720 51.980 ;
        RECT 1180.460 17.720 1180.720 17.980 ;
        RECT 1185.980 17.720 1186.240 17.980 ;
      LAYER met2 ;
        RECT 878.650 260.000 878.930 264.000 ;
        RECT 878.760 244.110 878.900 260.000 ;
        RECT 878.700 243.790 878.960 244.110 ;
        RECT 882.840 243.790 883.100 244.110 ;
        RECT 882.900 52.010 883.040 243.790 ;
        RECT 882.840 51.690 883.100 52.010 ;
        RECT 1180.460 51.690 1180.720 52.010 ;
        RECT 1180.520 18.010 1180.660 51.690 ;
        RECT 1180.460 17.690 1180.720 18.010 ;
        RECT 1185.980 17.690 1186.240 18.010 ;
        RECT 1186.040 2.400 1186.180 17.690 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
=======
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 896.150 58.720 896.470 58.780 ;
        RECT 1200.670 58.720 1200.990 58.780 ;
        RECT 896.150 58.580 1200.990 58.720 ;
        RECT 896.150 58.520 896.470 58.580 ;
        RECT 1200.670 58.520 1200.990 58.580 ;
      LAYER via ;
        RECT 896.180 58.520 896.440 58.780 ;
        RECT 1200.700 58.520 1200.960 58.780 ;
      LAYER met2 ;
        RECT 896.590 260.170 896.870 264.000 ;
        RECT 896.240 260.030 896.870 260.170 ;
        RECT 896.240 58.810 896.380 260.030 ;
        RECT 896.590 260.000 896.870 260.030 ;
        RECT 896.180 58.490 896.440 58.810 ;
        RECT 1200.700 58.490 1200.960 58.810 ;
        RECT 1200.760 16.730 1200.900 58.490 ;
        RECT 1200.760 16.590 1204.120 16.730 ;
        RECT 1203.980 2.400 1204.120 16.590 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
=======
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 917.310 65.520 917.630 65.580 ;
        RECT 1221.830 65.520 1222.150 65.580 ;
        RECT 917.310 65.380 1222.150 65.520 ;
        RECT 917.310 65.320 917.630 65.380 ;
        RECT 1221.830 65.320 1222.150 65.380 ;
      LAYER via ;
        RECT 917.340 65.320 917.600 65.580 ;
        RECT 1221.860 65.320 1222.120 65.580 ;
      LAYER met2 ;
        RECT 914.530 260.170 914.810 264.000 ;
        RECT 914.530 260.030 917.540 260.170 ;
        RECT 914.530 260.000 914.810 260.030 ;
        RECT 917.400 65.610 917.540 260.030 ;
        RECT 917.340 65.290 917.600 65.610 ;
        RECT 1221.860 65.290 1222.120 65.610 ;
        RECT 1221.920 2.400 1222.060 65.290 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
=======
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 932.490 244.020 932.810 244.080 ;
        RECT 938.010 244.020 938.330 244.080 ;
        RECT 932.490 243.880 938.330 244.020 ;
        RECT 932.490 243.820 932.810 243.880 ;
        RECT 938.010 243.820 938.330 243.880 ;
        RECT 938.010 72.320 938.330 72.380 ;
        RECT 1235.170 72.320 1235.490 72.380 ;
        RECT 938.010 72.180 1235.490 72.320 ;
        RECT 938.010 72.120 938.330 72.180 ;
        RECT 1235.170 72.120 1235.490 72.180 ;
      LAYER via ;
        RECT 932.520 243.820 932.780 244.080 ;
        RECT 938.040 243.820 938.300 244.080 ;
        RECT 938.040 72.120 938.300 72.380 ;
        RECT 1235.200 72.120 1235.460 72.380 ;
      LAYER met2 ;
        RECT 932.470 260.000 932.750 264.000 ;
        RECT 932.580 244.110 932.720 260.000 ;
        RECT 932.520 243.790 932.780 244.110 ;
        RECT 938.040 243.790 938.300 244.110 ;
        RECT 938.100 72.410 938.240 243.790 ;
        RECT 938.040 72.090 938.300 72.410 ;
        RECT 1235.200 72.090 1235.460 72.410 ;
        RECT 1235.260 16.730 1235.400 72.090 ;
        RECT 1235.260 16.590 1240.000 16.730 ;
        RECT 1239.860 2.400 1240.000 16.590 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
=======
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 951.810 24.040 952.130 24.100 ;
        RECT 1257.250 24.040 1257.570 24.100 ;
        RECT 951.810 23.900 1257.570 24.040 ;
        RECT 951.810 23.840 952.130 23.900 ;
        RECT 1257.250 23.840 1257.570 23.900 ;
      LAYER via ;
        RECT 951.840 23.840 952.100 24.100 ;
        RECT 1257.280 23.840 1257.540 24.100 ;
      LAYER met2 ;
        RECT 950.410 260.170 950.690 264.000 ;
        RECT 950.410 260.030 952.040 260.170 ;
        RECT 950.410 260.000 950.690 260.030 ;
        RECT 951.900 24.130 952.040 260.030 ;
        RECT 951.840 23.810 952.100 24.130 ;
        RECT 1257.280 23.810 1257.540 24.130 ;
        RECT 1257.340 2.400 1257.480 23.810 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
=======
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 967.910 244.020 968.230 244.080 ;
        RECT 972.510 244.020 972.830 244.080 ;
        RECT 967.910 243.880 972.830 244.020 ;
        RECT 967.910 243.820 968.230 243.880 ;
        RECT 972.510 243.820 972.830 243.880 ;
        RECT 972.510 79.460 972.830 79.520 ;
        RECT 1269.670 79.460 1269.990 79.520 ;
        RECT 972.510 79.320 1269.990 79.460 ;
        RECT 972.510 79.260 972.830 79.320 ;
        RECT 1269.670 79.260 1269.990 79.320 ;
      LAYER via ;
        RECT 967.940 243.820 968.200 244.080 ;
        RECT 972.540 243.820 972.800 244.080 ;
        RECT 972.540 79.260 972.800 79.520 ;
        RECT 1269.700 79.260 1269.960 79.520 ;
      LAYER met2 ;
        RECT 967.890 260.000 968.170 264.000 ;
        RECT 968.000 244.110 968.140 260.000 ;
        RECT 967.940 243.790 968.200 244.110 ;
        RECT 972.540 243.790 972.800 244.110 ;
        RECT 972.600 79.550 972.740 243.790 ;
        RECT 972.540 79.230 972.800 79.550 ;
        RECT 1269.700 79.230 1269.960 79.550 ;
        RECT 1269.760 16.730 1269.900 79.230 ;
        RECT 1269.760 16.590 1275.420 16.730 ;
        RECT 1275.280 2.400 1275.420 16.590 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
=======
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 985.850 86.260 986.170 86.320 ;
        RECT 1290.370 86.260 1290.690 86.320 ;
        RECT 985.850 86.120 1290.690 86.260 ;
        RECT 985.850 86.060 986.170 86.120 ;
        RECT 1290.370 86.060 1290.690 86.120 ;
      LAYER via ;
        RECT 985.880 86.060 986.140 86.320 ;
        RECT 1290.400 86.060 1290.660 86.320 ;
      LAYER met2 ;
        RECT 985.830 260.000 986.110 264.000 ;
        RECT 985.940 86.350 986.080 260.000 ;
        RECT 985.880 86.030 986.140 86.350 ;
        RECT 1290.400 86.030 1290.660 86.350 ;
        RECT 1290.460 17.410 1290.600 86.030 ;
        RECT 1290.460 17.270 1293.360 17.410 ;
        RECT 1293.220 2.400 1293.360 17.270 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
=======
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1007.010 141.340 1007.330 141.400 ;
        RECT 1311.530 141.340 1311.850 141.400 ;
        RECT 1007.010 141.200 1311.850 141.340 ;
        RECT 1007.010 141.140 1007.330 141.200 ;
        RECT 1311.530 141.140 1311.850 141.200 ;
      LAYER via ;
        RECT 1007.040 141.140 1007.300 141.400 ;
        RECT 1311.560 141.140 1311.820 141.400 ;
      LAYER met2 ;
        RECT 1003.770 260.170 1004.050 264.000 ;
        RECT 1003.770 260.030 1007.240 260.170 ;
        RECT 1003.770 260.000 1004.050 260.030 ;
        RECT 1007.100 141.430 1007.240 260.030 ;
        RECT 1007.040 141.110 1007.300 141.430 ;
        RECT 1311.560 141.110 1311.820 141.430 ;
        RECT 1311.620 17.410 1311.760 141.110 ;
        RECT 1311.160 17.270 1311.760 17.410 ;
        RECT 1311.160 2.400 1311.300 17.270 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
=======
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1021.730 244.020 1022.050 244.080 ;
        RECT 1027.710 244.020 1028.030 244.080 ;
        RECT 1021.730 243.880 1028.030 244.020 ;
        RECT 1021.730 243.820 1022.050 243.880 ;
        RECT 1027.710 243.820 1028.030 243.880 ;
        RECT 1027.710 99.860 1028.030 99.920 ;
        RECT 1324.870 99.860 1325.190 99.920 ;
        RECT 1027.710 99.720 1325.190 99.860 ;
        RECT 1027.710 99.660 1028.030 99.720 ;
        RECT 1324.870 99.660 1325.190 99.720 ;
      LAYER via ;
        RECT 1021.760 243.820 1022.020 244.080 ;
        RECT 1027.740 243.820 1028.000 244.080 ;
        RECT 1027.740 99.660 1028.000 99.920 ;
        RECT 1324.900 99.660 1325.160 99.920 ;
      LAYER met2 ;
        RECT 1021.710 260.000 1021.990 264.000 ;
        RECT 1021.820 244.110 1021.960 260.000 ;
        RECT 1021.760 243.790 1022.020 244.110 ;
        RECT 1027.740 243.790 1028.000 244.110 ;
        RECT 1027.800 99.950 1027.940 243.790 ;
        RECT 1027.740 99.630 1028.000 99.950 ;
        RECT 1324.900 99.630 1325.160 99.950 ;
        RECT 1324.960 17.410 1325.100 99.630 ;
        RECT 1324.960 17.270 1329.240 17.410 ;
        RECT 1329.100 2.400 1329.240 17.270 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
=======
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 379.110 99.860 379.430 99.920 ;
        RECT 683.170 99.860 683.490 99.920 ;
        RECT 379.110 99.720 683.490 99.860 ;
        RECT 379.110 99.660 379.430 99.720 ;
        RECT 683.170 99.660 683.490 99.720 ;
      LAYER via ;
        RECT 379.140 99.660 379.400 99.920 ;
        RECT 683.200 99.660 683.460 99.920 ;
      LAYER met2 ;
        RECT 378.170 260.170 378.450 264.000 ;
        RECT 378.170 260.030 379.340 260.170 ;
        RECT 378.170 260.000 378.450 260.030 ;
        RECT 379.200 99.950 379.340 260.030 ;
        RECT 379.140 99.630 379.400 99.950 ;
        RECT 683.200 99.630 683.460 99.950 ;
        RECT 683.260 16.730 683.400 99.630 ;
        RECT 683.260 16.590 686.620 16.730 ;
        RECT 686.480 2.400 686.620 16.590 ;
        RECT 686.270 -4.800 686.830 2.400 ;
=======
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1041.510 93.060 1041.830 93.120 ;
        RECT 1345.570 93.060 1345.890 93.120 ;
        RECT 1041.510 92.920 1345.890 93.060 ;
        RECT 1041.510 92.860 1041.830 92.920 ;
        RECT 1345.570 92.860 1345.890 92.920 ;
      LAYER via ;
        RECT 1041.540 92.860 1041.800 93.120 ;
        RECT 1345.600 92.860 1345.860 93.120 ;
      LAYER met2 ;
        RECT 1039.650 260.170 1039.930 264.000 ;
        RECT 1039.650 260.030 1041.740 260.170 ;
        RECT 1039.650 260.000 1039.930 260.030 ;
        RECT 1041.600 93.150 1041.740 260.030 ;
        RECT 1041.540 92.830 1041.800 93.150 ;
        RECT 1345.600 92.830 1345.860 93.150 ;
        RECT 1345.660 17.410 1345.800 92.830 ;
        RECT 1345.660 17.270 1346.720 17.410 ;
        RECT 1346.580 2.400 1346.720 17.270 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
=======
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1057.610 244.020 1057.930 244.080 ;
        RECT 1062.210 244.020 1062.530 244.080 ;
        RECT 1057.610 243.880 1062.530 244.020 ;
        RECT 1057.610 243.820 1057.930 243.880 ;
        RECT 1062.210 243.820 1062.530 243.880 ;
        RECT 1062.210 107.000 1062.530 107.060 ;
        RECT 1359.370 107.000 1359.690 107.060 ;
        RECT 1062.210 106.860 1359.690 107.000 ;
        RECT 1062.210 106.800 1062.530 106.860 ;
        RECT 1359.370 106.800 1359.690 106.860 ;
      LAYER via ;
        RECT 1057.640 243.820 1057.900 244.080 ;
        RECT 1062.240 243.820 1062.500 244.080 ;
        RECT 1062.240 106.800 1062.500 107.060 ;
        RECT 1359.400 106.800 1359.660 107.060 ;
      LAYER met2 ;
        RECT 1057.590 260.000 1057.870 264.000 ;
        RECT 1057.700 244.110 1057.840 260.000 ;
        RECT 1057.640 243.790 1057.900 244.110 ;
        RECT 1062.240 243.790 1062.500 244.110 ;
        RECT 1062.300 107.090 1062.440 243.790 ;
        RECT 1062.240 106.770 1062.500 107.090 ;
        RECT 1359.400 106.770 1359.660 107.090 ;
        RECT 1359.460 17.410 1359.600 106.770 ;
        RECT 1359.460 17.270 1364.660 17.410 ;
        RECT 1364.520 2.400 1364.660 17.270 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
=======
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1075.550 113.800 1075.870 113.860 ;
        RECT 1380.070 113.800 1380.390 113.860 ;
        RECT 1075.550 113.660 1380.390 113.800 ;
        RECT 1075.550 113.600 1075.870 113.660 ;
        RECT 1380.070 113.600 1380.390 113.660 ;
      LAYER via ;
        RECT 1075.580 113.600 1075.840 113.860 ;
        RECT 1380.100 113.600 1380.360 113.860 ;
      LAYER met2 ;
        RECT 1075.530 260.000 1075.810 264.000 ;
        RECT 1075.640 113.890 1075.780 260.000 ;
        RECT 1075.580 113.570 1075.840 113.890 ;
        RECT 1380.100 113.570 1380.360 113.890 ;
        RECT 1380.160 17.410 1380.300 113.570 ;
        RECT 1380.160 17.270 1382.600 17.410 ;
        RECT 1382.460 2.400 1382.600 17.270 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
=======
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1093.030 244.020 1093.350 244.080 ;
        RECT 1096.710 244.020 1097.030 244.080 ;
        RECT 1093.030 243.880 1097.030 244.020 ;
        RECT 1093.030 243.820 1093.350 243.880 ;
        RECT 1096.710 243.820 1097.030 243.880 ;
        RECT 1096.710 31.180 1097.030 31.240 ;
        RECT 1399.850 31.180 1400.170 31.240 ;
        RECT 1096.710 31.040 1400.170 31.180 ;
        RECT 1096.710 30.980 1097.030 31.040 ;
        RECT 1399.850 30.980 1400.170 31.040 ;
      LAYER via ;
        RECT 1093.060 243.820 1093.320 244.080 ;
        RECT 1096.740 243.820 1097.000 244.080 ;
        RECT 1096.740 30.980 1097.000 31.240 ;
        RECT 1399.880 30.980 1400.140 31.240 ;
      LAYER met2 ;
        RECT 1093.010 260.000 1093.290 264.000 ;
        RECT 1093.120 244.110 1093.260 260.000 ;
        RECT 1093.060 243.790 1093.320 244.110 ;
        RECT 1096.740 243.790 1097.000 244.110 ;
        RECT 1096.800 31.270 1096.940 243.790 ;
        RECT 1096.740 30.950 1097.000 31.270 ;
        RECT 1399.880 30.950 1400.140 31.270 ;
        RECT 1399.940 30.330 1400.080 30.950 ;
        RECT 1399.940 30.190 1400.540 30.330 ;
        RECT 1400.400 2.400 1400.540 30.190 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
=======
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1110.970 244.020 1111.290 244.080 ;
        RECT 1117.410 244.020 1117.730 244.080 ;
        RECT 1110.970 243.880 1117.730 244.020 ;
        RECT 1110.970 243.820 1111.290 243.880 ;
        RECT 1117.410 243.820 1117.730 243.880 ;
        RECT 1117.410 37.980 1117.730 38.040 ;
        RECT 1418.250 37.980 1418.570 38.040 ;
        RECT 1117.410 37.840 1418.570 37.980 ;
        RECT 1117.410 37.780 1117.730 37.840 ;
        RECT 1418.250 37.780 1418.570 37.840 ;
      LAYER via ;
        RECT 1111.000 243.820 1111.260 244.080 ;
        RECT 1117.440 243.820 1117.700 244.080 ;
        RECT 1117.440 37.780 1117.700 38.040 ;
        RECT 1418.280 37.780 1418.540 38.040 ;
      LAYER met2 ;
        RECT 1110.950 260.000 1111.230 264.000 ;
        RECT 1111.060 244.110 1111.200 260.000 ;
        RECT 1111.000 243.790 1111.260 244.110 ;
        RECT 1117.440 243.790 1117.700 244.110 ;
        RECT 1117.500 38.070 1117.640 243.790 ;
        RECT 1117.440 37.750 1117.700 38.070 ;
        RECT 1418.280 37.750 1418.540 38.070 ;
        RECT 1418.340 2.400 1418.480 37.750 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
=======
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1131.210 120.600 1131.530 120.660 ;
        RECT 1435.730 120.600 1436.050 120.660 ;
        RECT 1131.210 120.460 1436.050 120.600 ;
        RECT 1131.210 120.400 1131.530 120.460 ;
        RECT 1435.730 120.400 1436.050 120.460 ;
      LAYER via ;
        RECT 1131.240 120.400 1131.500 120.660 ;
        RECT 1435.760 120.400 1436.020 120.660 ;
      LAYER met2 ;
        RECT 1128.890 260.170 1129.170 264.000 ;
        RECT 1128.890 260.030 1131.440 260.170 ;
        RECT 1128.890 260.000 1129.170 260.030 ;
        RECT 1131.300 120.690 1131.440 260.030 ;
        RECT 1131.240 120.370 1131.500 120.690 ;
        RECT 1435.760 120.370 1436.020 120.690 ;
        RECT 1435.820 2.400 1435.960 120.370 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
=======
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1146.850 244.020 1147.170 244.080 ;
        RECT 1151.910 244.020 1152.230 244.080 ;
        RECT 1146.850 243.880 1152.230 244.020 ;
        RECT 1146.850 243.820 1147.170 243.880 ;
        RECT 1151.910 243.820 1152.230 243.880 ;
        RECT 1151.910 45.120 1152.230 45.180 ;
        RECT 1453.670 45.120 1453.990 45.180 ;
        RECT 1151.910 44.980 1453.990 45.120 ;
        RECT 1151.910 44.920 1152.230 44.980 ;
        RECT 1453.670 44.920 1453.990 44.980 ;
      LAYER via ;
        RECT 1146.880 243.820 1147.140 244.080 ;
        RECT 1151.940 243.820 1152.200 244.080 ;
        RECT 1151.940 44.920 1152.200 45.180 ;
        RECT 1453.700 44.920 1453.960 45.180 ;
      LAYER met2 ;
        RECT 1146.830 260.000 1147.110 264.000 ;
        RECT 1146.940 244.110 1147.080 260.000 ;
        RECT 1146.880 243.790 1147.140 244.110 ;
        RECT 1151.940 243.790 1152.200 244.110 ;
        RECT 1152.000 45.210 1152.140 243.790 ;
        RECT 1151.940 44.890 1152.200 45.210 ;
        RECT 1453.700 44.890 1453.960 45.210 ;
        RECT 1453.760 2.400 1453.900 44.890 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
=======
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1165.710 51.580 1166.030 51.640 ;
        RECT 1469.770 51.580 1470.090 51.640 ;
        RECT 1165.710 51.440 1470.090 51.580 ;
        RECT 1165.710 51.380 1166.030 51.440 ;
        RECT 1469.770 51.380 1470.090 51.440 ;
      LAYER via ;
        RECT 1165.740 51.380 1166.000 51.640 ;
        RECT 1469.800 51.380 1470.060 51.640 ;
      LAYER met2 ;
        RECT 1164.770 260.170 1165.050 264.000 ;
        RECT 1164.770 260.030 1165.940 260.170 ;
        RECT 1164.770 260.000 1165.050 260.030 ;
        RECT 1165.800 51.670 1165.940 260.030 ;
        RECT 1165.740 51.350 1166.000 51.670 ;
        RECT 1469.800 51.350 1470.060 51.670 ;
        RECT 1469.860 16.730 1470.000 51.350 ;
        RECT 1469.860 16.590 1471.840 16.730 ;
        RECT 1471.700 2.400 1471.840 16.590 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
=======
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1186.410 128.080 1186.730 128.140 ;
        RECT 1484.030 128.080 1484.350 128.140 ;
        RECT 1186.410 127.940 1484.350 128.080 ;
        RECT 1186.410 127.880 1186.730 127.940 ;
        RECT 1484.030 127.880 1484.350 127.940 ;
      LAYER via ;
        RECT 1186.440 127.880 1186.700 128.140 ;
        RECT 1484.060 127.880 1484.320 128.140 ;
      LAYER met2 ;
        RECT 1182.710 260.170 1182.990 264.000 ;
        RECT 1182.710 260.030 1186.640 260.170 ;
        RECT 1182.710 260.000 1182.990 260.030 ;
        RECT 1186.500 128.170 1186.640 260.030 ;
        RECT 1186.440 127.850 1186.700 128.170 ;
        RECT 1484.060 127.850 1484.320 128.170 ;
        RECT 1484.120 17.410 1484.260 127.850 ;
        RECT 1484.120 17.270 1489.780 17.410 ;
        RECT 1489.640 2.400 1489.780 17.270 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
=======
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1200.670 241.640 1200.990 241.700 ;
        RECT 1207.110 241.640 1207.430 241.700 ;
        RECT 1200.670 241.500 1207.430 241.640 ;
        RECT 1200.670 241.440 1200.990 241.500 ;
        RECT 1207.110 241.440 1207.430 241.500 ;
        RECT 1207.110 58.720 1207.430 58.780 ;
        RECT 1504.270 58.720 1504.590 58.780 ;
        RECT 1207.110 58.580 1504.590 58.720 ;
        RECT 1207.110 58.520 1207.430 58.580 ;
        RECT 1504.270 58.520 1504.590 58.580 ;
      LAYER via ;
        RECT 1200.700 241.440 1200.960 241.700 ;
        RECT 1207.140 241.440 1207.400 241.700 ;
        RECT 1207.140 58.520 1207.400 58.780 ;
        RECT 1504.300 58.520 1504.560 58.780 ;
      LAYER met2 ;
        RECT 1200.650 260.000 1200.930 264.000 ;
        RECT 1200.760 241.730 1200.900 260.000 ;
        RECT 1200.700 241.410 1200.960 241.730 ;
        RECT 1207.140 241.410 1207.400 241.730 ;
        RECT 1207.200 58.810 1207.340 241.410 ;
        RECT 1207.140 58.490 1207.400 58.810 ;
        RECT 1504.300 58.490 1504.560 58.810 ;
        RECT 1504.360 17.410 1504.500 58.490 ;
        RECT 1504.360 17.270 1507.260 17.410 ;
        RECT 1507.120 2.400 1507.260 17.270 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
=======
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 399.810 107.000 400.130 107.060 ;
        RECT 704.330 107.000 704.650 107.060 ;
        RECT 399.810 106.860 704.650 107.000 ;
        RECT 399.810 106.800 400.130 106.860 ;
        RECT 704.330 106.800 704.650 106.860 ;
      LAYER via ;
        RECT 399.840 106.800 400.100 107.060 ;
        RECT 704.360 106.800 704.620 107.060 ;
      LAYER met2 ;
        RECT 396.110 260.170 396.390 264.000 ;
        RECT 396.110 260.030 400.040 260.170 ;
        RECT 396.110 260.000 396.390 260.030 ;
        RECT 399.900 107.090 400.040 260.030 ;
        RECT 399.840 106.770 400.100 107.090 ;
        RECT 704.360 106.770 704.620 107.090 ;
        RECT 704.420 2.400 704.560 106.770 ;
        RECT 704.210 -4.800 704.770 2.400 ;
=======
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1220.910 134.540 1221.230 134.600 ;
        RECT 1525.430 134.540 1525.750 134.600 ;
        RECT 1220.910 134.400 1525.750 134.540 ;
        RECT 1220.910 134.340 1221.230 134.400 ;
        RECT 1525.430 134.340 1525.750 134.400 ;
      LAYER via ;
        RECT 1220.940 134.340 1221.200 134.600 ;
        RECT 1525.460 134.340 1525.720 134.600 ;
      LAYER met2 ;
        RECT 1218.130 260.170 1218.410 264.000 ;
        RECT 1218.130 260.030 1221.140 260.170 ;
        RECT 1218.130 260.000 1218.410 260.030 ;
        RECT 1221.000 134.630 1221.140 260.030 ;
        RECT 1220.940 134.310 1221.200 134.630 ;
        RECT 1525.460 134.310 1525.720 134.630 ;
        RECT 1525.520 17.410 1525.660 134.310 ;
        RECT 1525.060 17.270 1525.660 17.410 ;
        RECT 1525.060 2.400 1525.200 17.270 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
=======
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1236.090 244.020 1236.410 244.080 ;
        RECT 1241.610 244.020 1241.930 244.080 ;
        RECT 1236.090 243.880 1241.930 244.020 ;
        RECT 1236.090 243.820 1236.410 243.880 ;
        RECT 1241.610 243.820 1241.930 243.880 ;
        RECT 1241.610 72.320 1241.930 72.380 ;
        RECT 1538.770 72.320 1539.090 72.380 ;
        RECT 1241.610 72.180 1539.090 72.320 ;
        RECT 1241.610 72.120 1241.930 72.180 ;
        RECT 1538.770 72.120 1539.090 72.180 ;
      LAYER via ;
        RECT 1236.120 243.820 1236.380 244.080 ;
        RECT 1241.640 243.820 1241.900 244.080 ;
        RECT 1241.640 72.120 1241.900 72.380 ;
        RECT 1538.800 72.120 1539.060 72.380 ;
      LAYER met2 ;
        RECT 1236.070 260.000 1236.350 264.000 ;
        RECT 1236.180 244.110 1236.320 260.000 ;
        RECT 1236.120 243.790 1236.380 244.110 ;
        RECT 1241.640 243.790 1241.900 244.110 ;
        RECT 1241.700 72.410 1241.840 243.790 ;
        RECT 1241.640 72.090 1241.900 72.410 ;
        RECT 1538.800 72.090 1539.060 72.410 ;
        RECT 1538.860 16.730 1539.000 72.090 ;
        RECT 1538.860 16.590 1543.140 16.730 ;
        RECT 1543.000 2.400 1543.140 16.590 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
=======
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1255.410 65.520 1255.730 65.580 ;
        RECT 1559.470 65.520 1559.790 65.580 ;
        RECT 1255.410 65.380 1559.790 65.520 ;
        RECT 1255.410 65.320 1255.730 65.380 ;
        RECT 1559.470 65.320 1559.790 65.380 ;
      LAYER via ;
        RECT 1255.440 65.320 1255.700 65.580 ;
        RECT 1559.500 65.320 1559.760 65.580 ;
      LAYER met2 ;
        RECT 1254.010 260.170 1254.290 264.000 ;
        RECT 1254.010 260.030 1255.640 260.170 ;
        RECT 1254.010 260.000 1254.290 260.030 ;
        RECT 1255.500 65.610 1255.640 260.030 ;
        RECT 1255.440 65.290 1255.700 65.610 ;
        RECT 1559.500 65.290 1559.760 65.610 ;
        RECT 1559.560 16.730 1559.700 65.290 ;
        RECT 1559.560 16.590 1561.080 16.730 ;
        RECT 1560.940 2.400 1561.080 16.590 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
=======
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1271.970 244.020 1272.290 244.080 ;
        RECT 1276.110 244.020 1276.430 244.080 ;
        RECT 1271.970 243.880 1276.430 244.020 ;
        RECT 1271.970 243.820 1272.290 243.880 ;
        RECT 1276.110 243.820 1276.430 243.880 ;
        RECT 1276.110 24.380 1276.430 24.440 ;
        RECT 1578.790 24.380 1579.110 24.440 ;
        RECT 1276.110 24.240 1579.110 24.380 ;
        RECT 1276.110 24.180 1276.430 24.240 ;
        RECT 1578.790 24.180 1579.110 24.240 ;
      LAYER via ;
        RECT 1272.000 243.820 1272.260 244.080 ;
        RECT 1276.140 243.820 1276.400 244.080 ;
        RECT 1276.140 24.180 1276.400 24.440 ;
        RECT 1578.820 24.180 1579.080 24.440 ;
      LAYER met2 ;
        RECT 1271.950 260.000 1272.230 264.000 ;
        RECT 1272.060 244.110 1272.200 260.000 ;
        RECT 1272.000 243.790 1272.260 244.110 ;
        RECT 1276.140 243.790 1276.400 244.110 ;
        RECT 1276.200 24.470 1276.340 243.790 ;
        RECT 1276.140 24.150 1276.400 24.470 ;
        RECT 1578.820 24.150 1579.080 24.470 ;
        RECT 1578.880 2.400 1579.020 24.150 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
=======
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1289.450 79.460 1289.770 79.520 ;
        RECT 1593.970 79.460 1594.290 79.520 ;
        RECT 1289.450 79.320 1594.290 79.460 ;
        RECT 1289.450 79.260 1289.770 79.320 ;
        RECT 1593.970 79.260 1594.290 79.320 ;
      LAYER via ;
        RECT 1289.480 79.260 1289.740 79.520 ;
        RECT 1594.000 79.260 1594.260 79.520 ;
      LAYER met2 ;
        RECT 1289.890 260.170 1290.170 264.000 ;
        RECT 1289.540 260.030 1290.170 260.170 ;
        RECT 1289.540 79.550 1289.680 260.030 ;
        RECT 1289.890 260.000 1290.170 260.030 ;
        RECT 1289.480 79.230 1289.740 79.550 ;
        RECT 1594.000 79.230 1594.260 79.550 ;
        RECT 1594.060 16.730 1594.200 79.230 ;
        RECT 1594.060 16.590 1596.500 16.730 ;
        RECT 1596.360 2.400 1596.500 16.590 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
=======
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1310.610 86.260 1310.930 86.320 ;
        RECT 1608.230 86.260 1608.550 86.320 ;
        RECT 1310.610 86.120 1608.550 86.260 ;
        RECT 1310.610 86.060 1310.930 86.120 ;
        RECT 1608.230 86.060 1608.550 86.120 ;
        RECT 1608.230 38.320 1608.550 38.380 ;
        RECT 1614.210 38.320 1614.530 38.380 ;
        RECT 1608.230 38.180 1614.530 38.320 ;
        RECT 1608.230 38.120 1608.550 38.180 ;
        RECT 1614.210 38.120 1614.530 38.180 ;
      LAYER via ;
        RECT 1310.640 86.060 1310.900 86.320 ;
        RECT 1608.260 86.060 1608.520 86.320 ;
        RECT 1608.260 38.120 1608.520 38.380 ;
        RECT 1614.240 38.120 1614.500 38.380 ;
      LAYER met2 ;
        RECT 1307.830 260.170 1308.110 264.000 ;
        RECT 1307.830 260.030 1310.840 260.170 ;
        RECT 1307.830 260.000 1308.110 260.030 ;
        RECT 1310.700 86.350 1310.840 260.030 ;
        RECT 1310.640 86.030 1310.900 86.350 ;
        RECT 1608.260 86.030 1608.520 86.350 ;
        RECT 1608.320 38.410 1608.460 86.030 ;
        RECT 1608.260 38.090 1608.520 38.410 ;
        RECT 1614.240 38.090 1614.500 38.410 ;
        RECT 1614.300 2.400 1614.440 38.090 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
=======
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1325.790 244.020 1326.110 244.080 ;
        RECT 1331.310 244.020 1331.630 244.080 ;
        RECT 1325.790 243.880 1331.630 244.020 ;
        RECT 1325.790 243.820 1326.110 243.880 ;
        RECT 1331.310 243.820 1331.630 243.880 ;
        RECT 1331.310 99.860 1331.630 99.920 ;
        RECT 1628.470 99.860 1628.790 99.920 ;
        RECT 1331.310 99.720 1628.790 99.860 ;
        RECT 1331.310 99.660 1331.630 99.720 ;
        RECT 1628.470 99.660 1628.790 99.720 ;
        RECT 1628.470 62.260 1628.790 62.520 ;
        RECT 1628.560 62.120 1628.700 62.260 ;
        RECT 1632.150 62.120 1632.470 62.180 ;
        RECT 1628.560 61.980 1632.470 62.120 ;
        RECT 1632.150 61.920 1632.470 61.980 ;
        RECT 1632.150 47.980 1632.470 48.240 ;
        RECT 1632.240 47.560 1632.380 47.980 ;
        RECT 1632.150 47.300 1632.470 47.560 ;
      LAYER via ;
        RECT 1325.820 243.820 1326.080 244.080 ;
        RECT 1331.340 243.820 1331.600 244.080 ;
        RECT 1331.340 99.660 1331.600 99.920 ;
        RECT 1628.500 99.660 1628.760 99.920 ;
        RECT 1628.500 62.260 1628.760 62.520 ;
        RECT 1632.180 61.920 1632.440 62.180 ;
        RECT 1632.180 47.980 1632.440 48.240 ;
        RECT 1632.180 47.300 1632.440 47.560 ;
      LAYER met2 ;
        RECT 1325.770 260.000 1326.050 264.000 ;
        RECT 1325.880 244.110 1326.020 260.000 ;
        RECT 1325.820 243.790 1326.080 244.110 ;
        RECT 1331.340 243.790 1331.600 244.110 ;
        RECT 1331.400 99.950 1331.540 243.790 ;
        RECT 1331.340 99.630 1331.600 99.950 ;
        RECT 1628.500 99.630 1628.760 99.950 ;
        RECT 1628.560 62.550 1628.700 99.630 ;
        RECT 1628.500 62.230 1628.760 62.550 ;
        RECT 1632.180 61.890 1632.440 62.210 ;
        RECT 1632.240 48.270 1632.380 61.890 ;
        RECT 1632.180 47.950 1632.440 48.270 ;
        RECT 1632.180 47.270 1632.440 47.590 ;
        RECT 1632.240 2.400 1632.380 47.270 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
=======
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 1650.165 48.365 1650.335 93.415 ;
      LAYER mcon ;
        RECT 1650.165 93.245 1650.335 93.415 ;
      LAYER met1 ;
        RECT 1345.110 93.400 1345.430 93.460 ;
        RECT 1650.105 93.400 1650.395 93.445 ;
        RECT 1345.110 93.260 1650.395 93.400 ;
        RECT 1345.110 93.200 1345.430 93.260 ;
        RECT 1650.105 93.215 1650.395 93.260 ;
        RECT 1650.090 48.520 1650.410 48.580 ;
        RECT 1649.895 48.380 1650.410 48.520 ;
        RECT 1650.090 48.320 1650.410 48.380 ;
      LAYER via ;
        RECT 1345.140 93.200 1345.400 93.460 ;
        RECT 1650.120 48.320 1650.380 48.580 ;
      LAYER met2 ;
        RECT 1343.250 260.170 1343.530 264.000 ;
        RECT 1343.250 260.030 1345.340 260.170 ;
        RECT 1343.250 260.000 1343.530 260.030 ;
        RECT 1345.200 93.490 1345.340 260.030 ;
        RECT 1345.140 93.170 1345.400 93.490 ;
        RECT 1650.120 48.290 1650.380 48.610 ;
        RECT 1650.180 2.400 1650.320 48.290 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
=======
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1361.210 244.020 1361.530 244.080 ;
        RECT 1365.810 244.020 1366.130 244.080 ;
        RECT 1361.210 243.880 1366.130 244.020 ;
        RECT 1361.210 243.820 1361.530 243.880 ;
        RECT 1365.810 243.820 1366.130 243.880 ;
        RECT 1365.810 107.000 1366.130 107.060 ;
        RECT 1662.970 107.000 1663.290 107.060 ;
        RECT 1365.810 106.860 1663.290 107.000 ;
        RECT 1365.810 106.800 1366.130 106.860 ;
        RECT 1662.970 106.800 1663.290 106.860 ;
      LAYER via ;
        RECT 1361.240 243.820 1361.500 244.080 ;
        RECT 1365.840 243.820 1366.100 244.080 ;
        RECT 1365.840 106.800 1366.100 107.060 ;
        RECT 1663.000 106.800 1663.260 107.060 ;
      LAYER met2 ;
        RECT 1361.190 260.000 1361.470 264.000 ;
        RECT 1361.300 244.110 1361.440 260.000 ;
        RECT 1361.240 243.790 1361.500 244.110 ;
        RECT 1365.840 243.790 1366.100 244.110 ;
        RECT 1365.900 107.090 1366.040 243.790 ;
        RECT 1365.840 106.770 1366.100 107.090 ;
        RECT 1663.000 106.770 1663.260 107.090 ;
        RECT 1663.060 16.730 1663.200 106.770 ;
        RECT 1663.060 16.590 1668.260 16.730 ;
        RECT 1668.120 2.400 1668.260 16.590 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
=======
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1379.610 237.900 1379.930 237.960 ;
        RECT 1683.670 237.900 1683.990 237.960 ;
        RECT 1379.610 237.760 1683.990 237.900 ;
        RECT 1379.610 237.700 1379.930 237.760 ;
        RECT 1683.670 237.700 1683.990 237.760 ;
      LAYER via ;
        RECT 1379.640 237.700 1379.900 237.960 ;
        RECT 1683.700 237.700 1683.960 237.960 ;
      LAYER met2 ;
        RECT 1379.130 260.170 1379.410 264.000 ;
        RECT 1379.130 260.030 1379.840 260.170 ;
        RECT 1379.130 260.000 1379.410 260.030 ;
        RECT 1379.700 237.990 1379.840 260.030 ;
        RECT 1379.640 237.670 1379.900 237.990 ;
        RECT 1683.700 237.670 1683.960 237.990 ;
        RECT 1683.760 17.410 1683.900 237.670 ;
        RECT 1683.760 17.270 1685.740 17.410 ;
        RECT 1685.600 2.400 1685.740 17.270 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
=======
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 414.070 243.340 414.390 243.400 ;
        RECT 420.050 243.340 420.370 243.400 ;
        RECT 414.070 243.200 420.370 243.340 ;
        RECT 414.070 243.140 414.390 243.200 ;
        RECT 420.050 243.140 420.370 243.200 ;
        RECT 420.050 113.800 420.370 113.860 ;
        RECT 717.670 113.800 717.990 113.860 ;
        RECT 420.050 113.660 717.990 113.800 ;
        RECT 420.050 113.600 420.370 113.660 ;
        RECT 717.670 113.600 717.990 113.660 ;
      LAYER via ;
        RECT 414.100 243.140 414.360 243.400 ;
        RECT 420.080 243.140 420.340 243.400 ;
        RECT 420.080 113.600 420.340 113.860 ;
        RECT 717.700 113.600 717.960 113.860 ;
      LAYER met2 ;
        RECT 414.050 260.000 414.330 264.000 ;
        RECT 414.160 243.430 414.300 260.000 ;
        RECT 414.100 243.110 414.360 243.430 ;
        RECT 420.080 243.110 420.340 243.430 ;
        RECT 420.140 113.890 420.280 243.110 ;
        RECT 420.080 113.570 420.340 113.890 ;
        RECT 717.700 113.570 717.960 113.890 ;
        RECT 717.760 16.730 717.900 113.570 ;
        RECT 717.760 16.590 722.500 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
=======
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1400.310 30.840 1400.630 30.900 ;
        RECT 1703.450 30.840 1703.770 30.900 ;
        RECT 1400.310 30.700 1703.770 30.840 ;
        RECT 1400.310 30.640 1400.630 30.700 ;
        RECT 1703.450 30.640 1703.770 30.700 ;
      LAYER via ;
        RECT 1400.340 30.640 1400.600 30.900 ;
        RECT 1703.480 30.640 1703.740 30.900 ;
      LAYER met2 ;
        RECT 1397.070 260.170 1397.350 264.000 ;
        RECT 1397.070 260.030 1400.540 260.170 ;
        RECT 1397.070 260.000 1397.350 260.030 ;
        RECT 1400.400 30.930 1400.540 260.030 ;
        RECT 1400.340 30.610 1400.600 30.930 ;
        RECT 1703.480 30.610 1703.740 30.930 ;
        RECT 1703.540 2.400 1703.680 30.610 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
=======
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1415.030 244.020 1415.350 244.080 ;
        RECT 1421.010 244.020 1421.330 244.080 ;
        RECT 1415.030 243.880 1421.330 244.020 ;
        RECT 1415.030 243.820 1415.350 243.880 ;
        RECT 1421.010 243.820 1421.330 243.880 ;
        RECT 1421.010 37.980 1421.330 38.040 ;
        RECT 1721.390 37.980 1721.710 38.040 ;
        RECT 1421.010 37.840 1721.710 37.980 ;
        RECT 1421.010 37.780 1421.330 37.840 ;
        RECT 1721.390 37.780 1721.710 37.840 ;
      LAYER via ;
        RECT 1415.060 243.820 1415.320 244.080 ;
        RECT 1421.040 243.820 1421.300 244.080 ;
        RECT 1421.040 37.780 1421.300 38.040 ;
        RECT 1721.420 37.780 1721.680 38.040 ;
      LAYER met2 ;
        RECT 1415.010 260.000 1415.290 264.000 ;
        RECT 1415.120 244.110 1415.260 260.000 ;
        RECT 1415.060 243.790 1415.320 244.110 ;
        RECT 1421.040 243.790 1421.300 244.110 ;
        RECT 1421.100 38.070 1421.240 243.790 ;
        RECT 1421.040 37.750 1421.300 38.070 ;
        RECT 1721.420 37.750 1721.680 38.070 ;
        RECT 1721.480 2.400 1721.620 37.750 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
=======
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1434.810 113.800 1435.130 113.860 ;
        RECT 1739.330 113.800 1739.650 113.860 ;
        RECT 1434.810 113.660 1739.650 113.800 ;
        RECT 1434.810 113.600 1435.130 113.660 ;
        RECT 1739.330 113.600 1739.650 113.660 ;
      LAYER via ;
        RECT 1434.840 113.600 1435.100 113.860 ;
        RECT 1739.360 113.600 1739.620 113.860 ;
      LAYER met2 ;
        RECT 1432.950 260.170 1433.230 264.000 ;
        RECT 1432.950 260.030 1435.040 260.170 ;
        RECT 1432.950 260.000 1433.230 260.030 ;
        RECT 1434.900 113.890 1435.040 260.030 ;
        RECT 1434.840 113.570 1435.100 113.890 ;
        RECT 1739.360 113.570 1739.620 113.890 ;
        RECT 1739.420 2.400 1739.560 113.570 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
=======
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1450.910 244.020 1451.230 244.080 ;
        RECT 1455.510 244.020 1455.830 244.080 ;
        RECT 1450.910 243.880 1455.830 244.020 ;
        RECT 1450.910 243.820 1451.230 243.880 ;
        RECT 1455.510 243.820 1455.830 243.880 ;
        RECT 1455.510 44.780 1455.830 44.840 ;
        RECT 1756.810 44.780 1757.130 44.840 ;
        RECT 1455.510 44.640 1757.130 44.780 ;
        RECT 1455.510 44.580 1455.830 44.640 ;
        RECT 1756.810 44.580 1757.130 44.640 ;
      LAYER via ;
        RECT 1450.940 243.820 1451.200 244.080 ;
        RECT 1455.540 243.820 1455.800 244.080 ;
        RECT 1455.540 44.580 1455.800 44.840 ;
        RECT 1756.840 44.580 1757.100 44.840 ;
      LAYER met2 ;
        RECT 1450.890 260.000 1451.170 264.000 ;
        RECT 1451.000 244.110 1451.140 260.000 ;
        RECT 1450.940 243.790 1451.200 244.110 ;
        RECT 1455.540 243.790 1455.800 244.110 ;
        RECT 1455.600 44.870 1455.740 243.790 ;
        RECT 1455.540 44.550 1455.800 44.870 ;
        RECT 1756.840 44.550 1757.100 44.870 ;
        RECT 1756.900 2.400 1757.040 44.550 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
=======
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1468.390 231.100 1468.710 231.160 ;
        RECT 1773.370 231.100 1773.690 231.160 ;
        RECT 1468.390 230.960 1773.690 231.100 ;
        RECT 1468.390 230.900 1468.710 230.960 ;
        RECT 1773.370 230.900 1773.690 230.960 ;
        RECT 1773.370 2.960 1773.690 3.020 ;
        RECT 1774.750 2.960 1775.070 3.020 ;
        RECT 1773.370 2.820 1775.070 2.960 ;
        RECT 1773.370 2.760 1773.690 2.820 ;
        RECT 1774.750 2.760 1775.070 2.820 ;
      LAYER via ;
        RECT 1468.420 230.900 1468.680 231.160 ;
        RECT 1773.400 230.900 1773.660 231.160 ;
        RECT 1773.400 2.760 1773.660 3.020 ;
        RECT 1774.780 2.760 1775.040 3.020 ;
      LAYER met2 ;
        RECT 1468.370 260.000 1468.650 264.000 ;
        RECT 1468.480 231.190 1468.620 260.000 ;
        RECT 1468.420 230.870 1468.680 231.190 ;
        RECT 1773.400 230.870 1773.660 231.190 ;
        RECT 1773.460 3.050 1773.600 230.870 ;
        RECT 1773.400 2.730 1773.660 3.050 ;
        RECT 1774.780 2.730 1775.040 3.050 ;
        RECT 1774.840 2.400 1774.980 2.730 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
=======
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1490.010 51.580 1490.330 51.640 ;
        RECT 1787.170 51.580 1787.490 51.640 ;
        RECT 1490.010 51.440 1787.490 51.580 ;
        RECT 1490.010 51.380 1490.330 51.440 ;
        RECT 1787.170 51.380 1787.490 51.440 ;
        RECT 1787.630 2.960 1787.950 3.020 ;
        RECT 1792.690 2.960 1793.010 3.020 ;
        RECT 1787.630 2.820 1793.010 2.960 ;
        RECT 1787.630 2.760 1787.950 2.820 ;
        RECT 1792.690 2.760 1793.010 2.820 ;
      LAYER via ;
        RECT 1490.040 51.380 1490.300 51.640 ;
        RECT 1787.200 51.380 1787.460 51.640 ;
        RECT 1787.660 2.760 1787.920 3.020 ;
        RECT 1792.720 2.760 1792.980 3.020 ;
      LAYER met2 ;
        RECT 1486.310 260.170 1486.590 264.000 ;
        RECT 1486.310 260.030 1490.240 260.170 ;
        RECT 1486.310 260.000 1486.590 260.030 ;
        RECT 1490.100 51.670 1490.240 260.030 ;
        RECT 1490.040 51.350 1490.300 51.670 ;
        RECT 1787.200 51.350 1787.460 51.670 ;
        RECT 1787.260 20.130 1787.400 51.350 ;
        RECT 1787.260 19.990 1787.860 20.130 ;
        RECT 1787.720 3.050 1787.860 19.990 ;
        RECT 1787.660 2.730 1787.920 3.050 ;
        RECT 1792.720 2.730 1792.980 3.050 ;
        RECT 1792.780 2.400 1792.920 2.730 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
=======
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1504.270 244.020 1504.590 244.080 ;
        RECT 1510.710 244.020 1511.030 244.080 ;
        RECT 1504.270 243.880 1511.030 244.020 ;
        RECT 1504.270 243.820 1504.590 243.880 ;
        RECT 1510.710 243.820 1511.030 243.880 ;
        RECT 1510.710 59.060 1511.030 59.120 ;
        RECT 1807.870 59.060 1808.190 59.120 ;
        RECT 1510.710 58.920 1808.190 59.060 ;
        RECT 1510.710 58.860 1511.030 58.920 ;
        RECT 1807.870 58.860 1808.190 58.920 ;
        RECT 1807.870 2.960 1808.190 3.020 ;
        RECT 1810.630 2.960 1810.950 3.020 ;
        RECT 1807.870 2.820 1810.950 2.960 ;
        RECT 1807.870 2.760 1808.190 2.820 ;
        RECT 1810.630 2.760 1810.950 2.820 ;
      LAYER via ;
        RECT 1504.300 243.820 1504.560 244.080 ;
        RECT 1510.740 243.820 1511.000 244.080 ;
        RECT 1510.740 58.860 1511.000 59.120 ;
        RECT 1807.900 58.860 1808.160 59.120 ;
        RECT 1807.900 2.760 1808.160 3.020 ;
        RECT 1810.660 2.760 1810.920 3.020 ;
      LAYER met2 ;
        RECT 1504.250 260.000 1504.530 264.000 ;
        RECT 1504.360 244.110 1504.500 260.000 ;
        RECT 1504.300 243.790 1504.560 244.110 ;
        RECT 1510.740 243.790 1511.000 244.110 ;
        RECT 1510.800 59.150 1510.940 243.790 ;
        RECT 1510.740 58.830 1511.000 59.150 ;
        RECT 1807.900 58.830 1808.160 59.150 ;
        RECT 1807.960 3.050 1808.100 58.830 ;
        RECT 1807.900 2.730 1808.160 3.050 ;
        RECT 1810.660 2.730 1810.920 3.050 ;
        RECT 1810.720 2.400 1810.860 2.730 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
=======
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1524.510 120.600 1524.830 120.660 ;
        RECT 1829.030 120.600 1829.350 120.660 ;
        RECT 1524.510 120.460 1829.350 120.600 ;
        RECT 1524.510 120.400 1524.830 120.460 ;
        RECT 1829.030 120.400 1829.350 120.460 ;
      LAYER via ;
        RECT 1524.540 120.400 1524.800 120.660 ;
        RECT 1829.060 120.400 1829.320 120.660 ;
      LAYER met2 ;
        RECT 1522.190 260.170 1522.470 264.000 ;
        RECT 1522.190 260.030 1524.740 260.170 ;
        RECT 1522.190 260.000 1522.470 260.030 ;
        RECT 1524.600 120.690 1524.740 260.030 ;
        RECT 1524.540 120.370 1524.800 120.690 ;
        RECT 1829.060 120.370 1829.320 120.690 ;
        RECT 1829.120 7.210 1829.260 120.370 ;
        RECT 1828.660 7.070 1829.260 7.210 ;
        RECT 1828.660 2.400 1828.800 7.070 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
=======
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1540.150 244.020 1540.470 244.080 ;
        RECT 1545.210 244.020 1545.530 244.080 ;
        RECT 1540.150 243.880 1545.530 244.020 ;
        RECT 1540.150 243.820 1540.470 243.880 ;
        RECT 1545.210 243.820 1545.530 243.880 ;
        RECT 1545.210 72.320 1545.530 72.380 ;
        RECT 1842.370 72.320 1842.690 72.380 ;
        RECT 1545.210 72.180 1842.690 72.320 ;
        RECT 1545.210 72.120 1545.530 72.180 ;
        RECT 1842.370 72.120 1842.690 72.180 ;
      LAYER via ;
        RECT 1540.180 243.820 1540.440 244.080 ;
        RECT 1545.240 243.820 1545.500 244.080 ;
        RECT 1545.240 72.120 1545.500 72.380 ;
        RECT 1842.400 72.120 1842.660 72.380 ;
      LAYER met2 ;
        RECT 1540.130 260.000 1540.410 264.000 ;
        RECT 1540.240 244.110 1540.380 260.000 ;
        RECT 1540.180 243.790 1540.440 244.110 ;
        RECT 1545.240 243.790 1545.500 244.110 ;
        RECT 1545.300 72.410 1545.440 243.790 ;
        RECT 1545.240 72.090 1545.500 72.410 ;
        RECT 1842.400 72.090 1842.660 72.410 ;
        RECT 1842.460 16.730 1842.600 72.090 ;
        RECT 1842.460 16.590 1846.280 16.730 ;
        RECT 1846.140 2.400 1846.280 16.590 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
=======
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1558.090 245.720 1558.410 245.780 ;
        RECT 1728.290 245.720 1728.610 245.780 ;
        RECT 1558.090 245.580 1728.610 245.720 ;
        RECT 1558.090 245.520 1558.410 245.580 ;
        RECT 1728.290 245.520 1728.610 245.580 ;
        RECT 1728.290 31.180 1728.610 31.240 ;
        RECT 1863.990 31.180 1864.310 31.240 ;
        RECT 1728.290 31.040 1864.310 31.180 ;
        RECT 1728.290 30.980 1728.610 31.040 ;
        RECT 1863.990 30.980 1864.310 31.040 ;
      LAYER via ;
        RECT 1558.120 245.520 1558.380 245.780 ;
        RECT 1728.320 245.520 1728.580 245.780 ;
        RECT 1728.320 30.980 1728.580 31.240 ;
        RECT 1864.020 30.980 1864.280 31.240 ;
      LAYER met2 ;
        RECT 1558.070 260.000 1558.350 264.000 ;
        RECT 1558.180 245.810 1558.320 260.000 ;
        RECT 1558.120 245.490 1558.380 245.810 ;
        RECT 1728.320 245.490 1728.580 245.810 ;
        RECT 1728.380 31.270 1728.520 245.490 ;
        RECT 1728.320 30.950 1728.580 31.270 ;
        RECT 1864.020 30.950 1864.280 31.270 ;
        RECT 1864.080 2.400 1864.220 30.950 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
=======
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 434.310 120.600 434.630 120.660 ;
        RECT 738.370 120.600 738.690 120.660 ;
        RECT 434.310 120.460 738.690 120.600 ;
        RECT 434.310 120.400 434.630 120.460 ;
        RECT 738.370 120.400 738.690 120.460 ;
      LAYER via ;
        RECT 434.340 120.400 434.600 120.660 ;
        RECT 738.400 120.400 738.660 120.660 ;
      LAYER met2 ;
        RECT 431.990 260.170 432.270 264.000 ;
        RECT 431.990 260.030 434.540 260.170 ;
        RECT 431.990 260.000 432.270 260.030 ;
        RECT 434.400 120.690 434.540 260.030 ;
        RECT 434.340 120.370 434.600 120.690 ;
        RECT 738.400 120.370 738.660 120.690 ;
        RECT 738.460 16.730 738.600 120.370 ;
        RECT 738.460 16.590 740.440 16.730 ;
        RECT 740.300 2.400 740.440 16.590 ;
        RECT 740.090 -4.800 740.650 2.400 ;
=======
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1576.030 243.680 1576.350 243.740 ;
        RECT 1579.710 243.680 1580.030 243.740 ;
        RECT 1576.030 243.540 1580.030 243.680 ;
        RECT 1576.030 243.480 1576.350 243.540 ;
        RECT 1579.710 243.480 1580.030 243.540 ;
        RECT 1579.710 65.520 1580.030 65.580 ;
        RECT 1876.870 65.520 1877.190 65.580 ;
        RECT 1579.710 65.380 1877.190 65.520 ;
        RECT 1579.710 65.320 1580.030 65.380 ;
        RECT 1876.870 65.320 1877.190 65.380 ;
        RECT 1876.870 62.120 1877.190 62.180 ;
        RECT 1881.930 62.120 1882.250 62.180 ;
        RECT 1876.870 61.980 1882.250 62.120 ;
        RECT 1876.870 61.920 1877.190 61.980 ;
        RECT 1881.930 61.920 1882.250 61.980 ;
      LAYER via ;
        RECT 1576.060 243.480 1576.320 243.740 ;
        RECT 1579.740 243.480 1580.000 243.740 ;
        RECT 1579.740 65.320 1580.000 65.580 ;
        RECT 1876.900 65.320 1877.160 65.580 ;
        RECT 1876.900 61.920 1877.160 62.180 ;
        RECT 1881.960 61.920 1882.220 62.180 ;
      LAYER met2 ;
        RECT 1576.010 260.000 1576.290 264.000 ;
        RECT 1576.120 243.770 1576.260 260.000 ;
        RECT 1576.060 243.450 1576.320 243.770 ;
        RECT 1579.740 243.450 1580.000 243.770 ;
        RECT 1579.800 65.610 1579.940 243.450 ;
        RECT 1579.740 65.290 1580.000 65.610 ;
        RECT 1876.900 65.290 1877.160 65.610 ;
        RECT 1876.960 62.210 1877.100 65.290 ;
        RECT 1876.900 61.890 1877.160 62.210 ;
        RECT 1881.960 61.890 1882.220 62.210 ;
        RECT 1882.020 2.400 1882.160 61.890 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
=======
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1593.050 79.800 1593.370 79.860 ;
        RECT 1897.570 79.800 1897.890 79.860 ;
        RECT 1593.050 79.660 1897.890 79.800 ;
        RECT 1593.050 79.600 1593.370 79.660 ;
        RECT 1897.570 79.600 1897.890 79.660 ;
      LAYER via ;
        RECT 1593.080 79.600 1593.340 79.860 ;
        RECT 1897.600 79.600 1897.860 79.860 ;
      LAYER met2 ;
        RECT 1593.490 260.170 1593.770 264.000 ;
        RECT 1593.140 260.030 1593.770 260.170 ;
        RECT 1593.140 79.890 1593.280 260.030 ;
        RECT 1593.490 260.000 1593.770 260.030 ;
        RECT 1593.080 79.570 1593.340 79.890 ;
        RECT 1897.600 79.570 1897.860 79.890 ;
        RECT 1897.660 16.730 1897.800 79.570 ;
        RECT 1897.660 16.590 1900.100 16.730 ;
        RECT 1899.960 2.400 1900.100 16.590 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
=======
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1614.210 86.260 1614.530 86.320 ;
        RECT 1911.830 86.260 1912.150 86.320 ;
        RECT 1614.210 86.120 1912.150 86.260 ;
        RECT 1614.210 86.060 1614.530 86.120 ;
        RECT 1911.830 86.060 1912.150 86.120 ;
        RECT 1911.830 17.920 1912.150 17.980 ;
        RECT 1917.810 17.920 1918.130 17.980 ;
        RECT 1911.830 17.780 1918.130 17.920 ;
        RECT 1911.830 17.720 1912.150 17.780 ;
        RECT 1917.810 17.720 1918.130 17.780 ;
      LAYER via ;
        RECT 1614.240 86.060 1614.500 86.320 ;
        RECT 1911.860 86.060 1912.120 86.320 ;
        RECT 1911.860 17.720 1912.120 17.980 ;
        RECT 1917.840 17.720 1918.100 17.980 ;
      LAYER met2 ;
        RECT 1611.430 260.170 1611.710 264.000 ;
        RECT 1611.430 260.030 1614.440 260.170 ;
        RECT 1611.430 260.000 1611.710 260.030 ;
        RECT 1614.300 86.350 1614.440 260.030 ;
        RECT 1614.240 86.030 1614.500 86.350 ;
        RECT 1911.860 86.030 1912.120 86.350 ;
        RECT 1911.920 18.010 1912.060 86.030 ;
        RECT 1911.860 17.690 1912.120 18.010 ;
        RECT 1917.840 17.690 1918.100 18.010 ;
        RECT 1917.900 2.400 1918.040 17.690 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
=======
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1629.390 244.020 1629.710 244.080 ;
        RECT 1634.910 244.020 1635.230 244.080 ;
        RECT 1629.390 243.880 1635.230 244.020 ;
        RECT 1629.390 243.820 1629.710 243.880 ;
        RECT 1634.910 243.820 1635.230 243.880 ;
        RECT 1634.910 99.860 1635.230 99.920 ;
        RECT 1932.070 99.860 1932.390 99.920 ;
        RECT 1634.910 99.720 1932.390 99.860 ;
        RECT 1634.910 99.660 1635.230 99.720 ;
        RECT 1932.070 99.660 1932.390 99.720 ;
        RECT 1932.070 2.960 1932.390 3.020 ;
        RECT 1935.290 2.960 1935.610 3.020 ;
        RECT 1932.070 2.820 1935.610 2.960 ;
        RECT 1932.070 2.760 1932.390 2.820 ;
        RECT 1935.290 2.760 1935.610 2.820 ;
      LAYER via ;
        RECT 1629.420 243.820 1629.680 244.080 ;
        RECT 1634.940 243.820 1635.200 244.080 ;
        RECT 1634.940 99.660 1635.200 99.920 ;
        RECT 1932.100 99.660 1932.360 99.920 ;
        RECT 1932.100 2.760 1932.360 3.020 ;
        RECT 1935.320 2.760 1935.580 3.020 ;
      LAYER met2 ;
        RECT 1629.370 260.000 1629.650 264.000 ;
        RECT 1629.480 244.110 1629.620 260.000 ;
        RECT 1629.420 243.790 1629.680 244.110 ;
        RECT 1634.940 243.790 1635.200 244.110 ;
        RECT 1635.000 99.950 1635.140 243.790 ;
        RECT 1634.940 99.630 1635.200 99.950 ;
        RECT 1932.100 99.630 1932.360 99.950 ;
        RECT 1932.160 3.050 1932.300 99.630 ;
        RECT 1932.100 2.730 1932.360 3.050 ;
        RECT 1935.320 2.730 1935.580 3.050 ;
        RECT 1935.380 2.400 1935.520 2.730 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
=======
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1647.330 244.020 1647.650 244.080 ;
        RECT 1652.390 244.020 1652.710 244.080 ;
        RECT 1647.330 243.880 1652.710 244.020 ;
        RECT 1647.330 243.820 1647.650 243.880 ;
        RECT 1652.390 243.820 1652.710 243.880 ;
        RECT 1652.390 93.060 1652.710 93.120 ;
        RECT 1953.230 93.060 1953.550 93.120 ;
        RECT 1652.390 92.920 1953.550 93.060 ;
        RECT 1652.390 92.860 1652.710 92.920 ;
        RECT 1953.230 92.860 1953.550 92.920 ;
      LAYER via ;
        RECT 1647.360 243.820 1647.620 244.080 ;
        RECT 1652.420 243.820 1652.680 244.080 ;
        RECT 1652.420 92.860 1652.680 93.120 ;
        RECT 1953.260 92.860 1953.520 93.120 ;
      LAYER met2 ;
        RECT 1647.310 260.000 1647.590 264.000 ;
        RECT 1647.420 244.110 1647.560 260.000 ;
        RECT 1647.360 243.790 1647.620 244.110 ;
        RECT 1652.420 243.790 1652.680 244.110 ;
        RECT 1652.480 93.150 1652.620 243.790 ;
        RECT 1652.420 92.830 1652.680 93.150 ;
        RECT 1953.260 92.830 1953.520 93.150 ;
        RECT 1953.320 2.400 1953.460 92.830 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
=======
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1665.270 244.020 1665.590 244.080 ;
        RECT 1669.410 244.020 1669.730 244.080 ;
        RECT 1665.270 243.880 1669.730 244.020 ;
        RECT 1665.270 243.820 1665.590 243.880 ;
        RECT 1669.410 243.820 1669.730 243.880 ;
        RECT 1669.410 107.000 1669.730 107.060 ;
        RECT 1966.570 107.000 1966.890 107.060 ;
        RECT 1669.410 106.860 1966.890 107.000 ;
        RECT 1669.410 106.800 1669.730 106.860 ;
        RECT 1966.570 106.800 1966.890 106.860 ;
        RECT 1966.570 62.120 1966.890 62.180 ;
        RECT 1971.170 62.120 1971.490 62.180 ;
        RECT 1966.570 61.980 1971.490 62.120 ;
        RECT 1966.570 61.920 1966.890 61.980 ;
        RECT 1971.170 61.920 1971.490 61.980 ;
      LAYER via ;
        RECT 1665.300 243.820 1665.560 244.080 ;
        RECT 1669.440 243.820 1669.700 244.080 ;
        RECT 1669.440 106.800 1669.700 107.060 ;
        RECT 1966.600 106.800 1966.860 107.060 ;
        RECT 1966.600 61.920 1966.860 62.180 ;
        RECT 1971.200 61.920 1971.460 62.180 ;
      LAYER met2 ;
        RECT 1665.250 260.000 1665.530 264.000 ;
        RECT 1665.360 244.110 1665.500 260.000 ;
        RECT 1665.300 243.790 1665.560 244.110 ;
        RECT 1669.440 243.790 1669.700 244.110 ;
        RECT 1669.500 107.090 1669.640 243.790 ;
        RECT 1669.440 106.770 1669.700 107.090 ;
        RECT 1966.600 106.770 1966.860 107.090 ;
        RECT 1966.660 62.210 1966.800 106.770 ;
        RECT 1966.600 61.890 1966.860 62.210 ;
        RECT 1971.200 61.890 1971.460 62.210 ;
        RECT 1971.260 2.400 1971.400 61.890 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
=======
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 1987.345 48.365 1987.515 96.475 ;
      LAYER mcon ;
        RECT 1987.345 96.305 1987.515 96.475 ;
      LAYER met1 ;
        RECT 1682.750 127.740 1683.070 127.800 ;
        RECT 1987.730 127.740 1988.050 127.800 ;
        RECT 1682.750 127.600 1988.050 127.740 ;
        RECT 1682.750 127.540 1683.070 127.600 ;
        RECT 1987.730 127.540 1988.050 127.600 ;
        RECT 1987.270 96.460 1987.590 96.520 ;
        RECT 1987.075 96.320 1987.590 96.460 ;
        RECT 1987.270 96.260 1987.590 96.320 ;
        RECT 1987.285 48.520 1987.575 48.565 ;
        RECT 1989.110 48.520 1989.430 48.580 ;
        RECT 1987.285 48.380 1989.430 48.520 ;
        RECT 1987.285 48.335 1987.575 48.380 ;
        RECT 1989.110 48.320 1989.430 48.380 ;
      LAYER via ;
        RECT 1682.780 127.540 1683.040 127.800 ;
        RECT 1987.760 127.540 1988.020 127.800 ;
        RECT 1987.300 96.260 1987.560 96.520 ;
        RECT 1989.140 48.320 1989.400 48.580 ;
      LAYER met2 ;
        RECT 1683.190 260.170 1683.470 264.000 ;
        RECT 1682.840 260.030 1683.470 260.170 ;
        RECT 1682.840 127.830 1682.980 260.030 ;
        RECT 1683.190 260.000 1683.470 260.030 ;
        RECT 1682.780 127.510 1683.040 127.830 ;
        RECT 1987.760 127.510 1988.020 127.830 ;
        RECT 1987.820 96.970 1987.960 127.510 ;
        RECT 1987.360 96.830 1987.960 96.970 ;
        RECT 1987.360 96.550 1987.500 96.830 ;
        RECT 1987.300 96.230 1987.560 96.550 ;
        RECT 1989.140 48.290 1989.400 48.610 ;
        RECT 1989.200 2.400 1989.340 48.290 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
=======
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1703.910 38.320 1704.230 38.380 ;
        RECT 2006.590 38.320 2006.910 38.380 ;
        RECT 1703.910 38.180 2006.910 38.320 ;
        RECT 1703.910 38.120 1704.230 38.180 ;
        RECT 2006.590 38.120 2006.910 38.180 ;
      LAYER via ;
        RECT 1703.940 38.120 1704.200 38.380 ;
        RECT 2006.620 38.120 2006.880 38.380 ;
      LAYER met2 ;
        RECT 1701.130 260.170 1701.410 264.000 ;
        RECT 1701.130 260.030 1704.140 260.170 ;
        RECT 1701.130 260.000 1701.410 260.030 ;
        RECT 1704.000 38.410 1704.140 260.030 ;
        RECT 1703.940 38.090 1704.200 38.410 ;
        RECT 2006.620 38.090 2006.880 38.410 ;
        RECT 2006.680 2.400 2006.820 38.090 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
=======
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1718.630 244.020 1718.950 244.080 ;
        RECT 1724.150 244.020 1724.470 244.080 ;
        RECT 1718.630 243.880 1724.470 244.020 ;
        RECT 1718.630 243.820 1718.950 243.880 ;
        RECT 1724.150 243.820 1724.470 243.880 ;
        RECT 1724.150 134.540 1724.470 134.600 ;
        RECT 2021.770 134.540 2022.090 134.600 ;
        RECT 1724.150 134.400 2022.090 134.540 ;
        RECT 1724.150 134.340 1724.470 134.400 ;
        RECT 2021.770 134.340 2022.090 134.400 ;
      LAYER via ;
        RECT 1718.660 243.820 1718.920 244.080 ;
        RECT 1724.180 243.820 1724.440 244.080 ;
        RECT 1724.180 134.340 1724.440 134.600 ;
        RECT 2021.800 134.340 2022.060 134.600 ;
      LAYER met2 ;
        RECT 1718.610 260.000 1718.890 264.000 ;
        RECT 1718.720 244.110 1718.860 260.000 ;
        RECT 1718.660 243.790 1718.920 244.110 ;
        RECT 1724.180 243.790 1724.440 244.110 ;
        RECT 1724.240 134.630 1724.380 243.790 ;
        RECT 1724.180 134.310 1724.440 134.630 ;
        RECT 2021.800 134.310 2022.060 134.630 ;
        RECT 2021.860 16.730 2022.000 134.310 ;
        RECT 2021.860 16.590 2024.760 16.730 ;
        RECT 2024.620 2.400 2024.760 16.590 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
=======
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1736.570 237.900 1736.890 237.960 ;
        RECT 2042.470 237.900 2042.790 237.960 ;
        RECT 1736.570 237.760 2042.790 237.900 ;
        RECT 1736.570 237.700 1736.890 237.760 ;
        RECT 2042.470 237.700 2042.790 237.760 ;
      LAYER via ;
        RECT 1736.600 237.700 1736.860 237.960 ;
        RECT 2042.500 237.700 2042.760 237.960 ;
      LAYER met2 ;
        RECT 1736.550 260.000 1736.830 264.000 ;
        RECT 1736.660 237.990 1736.800 260.000 ;
        RECT 1736.600 237.670 1736.860 237.990 ;
        RECT 2042.500 237.670 2042.760 237.990 ;
        RECT 2042.560 2.400 2042.700 237.670 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
=======
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 449.490 244.020 449.810 244.080 ;
        RECT 455.010 244.020 455.330 244.080 ;
        RECT 449.490 243.880 455.330 244.020 ;
        RECT 449.490 243.820 449.810 243.880 ;
        RECT 455.010 243.820 455.330 243.880 ;
        RECT 455.010 127.740 455.330 127.800 ;
        RECT 752.630 127.740 752.950 127.800 ;
        RECT 455.010 127.600 752.950 127.740 ;
        RECT 455.010 127.540 455.330 127.600 ;
        RECT 752.630 127.540 752.950 127.600 ;
        RECT 752.630 18.940 752.950 19.000 ;
        RECT 757.690 18.940 758.010 19.000 ;
        RECT 752.630 18.800 758.010 18.940 ;
        RECT 752.630 18.740 752.950 18.800 ;
        RECT 757.690 18.740 758.010 18.800 ;
      LAYER via ;
        RECT 449.520 243.820 449.780 244.080 ;
        RECT 455.040 243.820 455.300 244.080 ;
        RECT 455.040 127.540 455.300 127.800 ;
        RECT 752.660 127.540 752.920 127.800 ;
        RECT 752.660 18.740 752.920 19.000 ;
        RECT 757.720 18.740 757.980 19.000 ;
      LAYER met2 ;
        RECT 449.470 260.000 449.750 264.000 ;
        RECT 449.580 244.110 449.720 260.000 ;
        RECT 449.520 243.790 449.780 244.110 ;
        RECT 455.040 243.790 455.300 244.110 ;
        RECT 455.100 127.830 455.240 243.790 ;
        RECT 455.040 127.510 455.300 127.830 ;
        RECT 752.660 127.510 752.920 127.830 ;
        RECT 752.720 19.030 752.860 127.510 ;
        RECT 752.660 18.710 752.920 19.030 ;
        RECT 757.720 18.710 757.980 19.030 ;
        RECT 757.780 2.400 757.920 18.710 ;
        RECT 757.570 -4.800 758.130 2.400 ;
=======
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1754.510 244.020 1754.830 244.080 ;
        RECT 1759.110 244.020 1759.430 244.080 ;
        RECT 1754.510 243.880 1759.430 244.020 ;
        RECT 1754.510 243.820 1754.830 243.880 ;
        RECT 1759.110 243.820 1759.430 243.880 ;
        RECT 1759.110 44.780 1759.430 44.840 ;
        RECT 2060.410 44.780 2060.730 44.840 ;
        RECT 1759.110 44.640 2060.730 44.780 ;
        RECT 1759.110 44.580 1759.430 44.640 ;
        RECT 2060.410 44.580 2060.730 44.640 ;
      LAYER via ;
        RECT 1754.540 243.820 1754.800 244.080 ;
        RECT 1759.140 243.820 1759.400 244.080 ;
        RECT 1759.140 44.580 1759.400 44.840 ;
        RECT 2060.440 44.580 2060.700 44.840 ;
      LAYER met2 ;
        RECT 1754.490 260.000 1754.770 264.000 ;
        RECT 1754.600 244.110 1754.740 260.000 ;
        RECT 1754.540 243.790 1754.800 244.110 ;
        RECT 1759.140 243.790 1759.400 244.110 ;
        RECT 1759.200 44.870 1759.340 243.790 ;
        RECT 1759.140 44.550 1759.400 44.870 ;
        RECT 2060.440 44.550 2060.700 44.870 ;
        RECT 2060.500 2.400 2060.640 44.550 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
=======
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1772.450 245.040 1772.770 245.100 ;
        RECT 1838.690 245.040 1839.010 245.100 ;
        RECT 1772.450 244.900 1839.010 245.040 ;
        RECT 1772.450 244.840 1772.770 244.900 ;
        RECT 1838.690 244.840 1839.010 244.900 ;
        RECT 1838.690 51.580 1839.010 51.640 ;
        RECT 2076.970 51.580 2077.290 51.640 ;
        RECT 1838.690 51.440 2077.290 51.580 ;
        RECT 1838.690 51.380 1839.010 51.440 ;
        RECT 2076.970 51.380 2077.290 51.440 ;
      LAYER via ;
        RECT 1772.480 244.840 1772.740 245.100 ;
        RECT 1838.720 244.840 1838.980 245.100 ;
        RECT 1838.720 51.380 1838.980 51.640 ;
        RECT 2077.000 51.380 2077.260 51.640 ;
      LAYER met2 ;
        RECT 1772.430 260.000 1772.710 264.000 ;
        RECT 1772.540 245.130 1772.680 260.000 ;
        RECT 1772.480 244.810 1772.740 245.130 ;
        RECT 1838.720 244.810 1838.980 245.130 ;
        RECT 1838.780 51.670 1838.920 244.810 ;
        RECT 1838.720 51.350 1838.980 51.670 ;
        RECT 2077.000 51.350 2077.260 51.670 ;
        RECT 2077.060 4.490 2077.200 51.350 ;
        RECT 2077.060 4.350 2078.580 4.490 ;
        RECT 2078.440 2.400 2078.580 4.350 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
=======
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1793.610 25.060 1793.930 25.120 ;
        RECT 2095.830 25.060 2096.150 25.120 ;
        RECT 1793.610 24.920 2096.150 25.060 ;
        RECT 1793.610 24.860 1793.930 24.920 ;
        RECT 2095.830 24.860 2096.150 24.920 ;
      LAYER via ;
        RECT 1793.640 24.860 1793.900 25.120 ;
        RECT 2095.860 24.860 2096.120 25.120 ;
      LAYER met2 ;
        RECT 1790.370 260.170 1790.650 264.000 ;
        RECT 1790.370 260.030 1793.840 260.170 ;
        RECT 1790.370 260.000 1790.650 260.030 ;
        RECT 1793.700 25.150 1793.840 260.030 ;
        RECT 1793.640 24.830 1793.900 25.150 ;
        RECT 2095.860 24.830 2096.120 25.150 ;
        RECT 2095.920 2.400 2096.060 24.830 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
=======
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1808.330 244.020 1808.650 244.080 ;
        RECT 1814.310 244.020 1814.630 244.080 ;
        RECT 1808.330 243.880 1814.630 244.020 ;
        RECT 1808.330 243.820 1808.650 243.880 ;
        RECT 1814.310 243.820 1814.630 243.880 ;
        RECT 1814.310 26.420 1814.630 26.480 ;
        RECT 2113.770 26.420 2114.090 26.480 ;
        RECT 1814.310 26.280 2114.090 26.420 ;
        RECT 1814.310 26.220 1814.630 26.280 ;
        RECT 2113.770 26.220 2114.090 26.280 ;
      LAYER via ;
        RECT 1808.360 243.820 1808.620 244.080 ;
        RECT 1814.340 243.820 1814.600 244.080 ;
        RECT 1814.340 26.220 1814.600 26.480 ;
        RECT 2113.800 26.220 2114.060 26.480 ;
      LAYER met2 ;
        RECT 1808.310 260.000 1808.590 264.000 ;
        RECT 1808.420 244.110 1808.560 260.000 ;
        RECT 1808.360 243.790 1808.620 244.110 ;
        RECT 1814.340 243.790 1814.600 244.110 ;
        RECT 1814.400 26.510 1814.540 243.790 ;
        RECT 1814.340 26.190 1814.600 26.510 ;
        RECT 2113.800 26.190 2114.060 26.510 ;
        RECT 2113.860 2.400 2114.000 26.190 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
=======
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1826.270 231.100 1826.590 231.160 ;
        RECT 2125.270 231.100 2125.590 231.160 ;
        RECT 1826.270 230.960 2125.590 231.100 ;
        RECT 1826.270 230.900 1826.590 230.960 ;
        RECT 2125.270 230.900 2125.590 230.960 ;
        RECT 2125.270 17.580 2125.590 17.640 ;
        RECT 2131.710 17.580 2132.030 17.640 ;
        RECT 2125.270 17.440 2132.030 17.580 ;
        RECT 2125.270 17.380 2125.590 17.440 ;
        RECT 2131.710 17.380 2132.030 17.440 ;
      LAYER via ;
        RECT 1826.300 230.900 1826.560 231.160 ;
        RECT 2125.300 230.900 2125.560 231.160 ;
        RECT 2125.300 17.380 2125.560 17.640 ;
        RECT 2131.740 17.380 2132.000 17.640 ;
      LAYER met2 ;
        RECT 1826.250 260.000 1826.530 264.000 ;
        RECT 1826.360 231.190 1826.500 260.000 ;
        RECT 1826.300 230.870 1826.560 231.190 ;
        RECT 2125.300 230.870 2125.560 231.190 ;
        RECT 2125.360 17.670 2125.500 230.870 ;
        RECT 2125.300 17.350 2125.560 17.670 ;
        RECT 2131.740 17.350 2132.000 17.670 ;
        RECT 2131.800 2.400 2131.940 17.350 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
=======
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1844.210 241.640 1844.530 241.700 ;
        RECT 1848.810 241.640 1849.130 241.700 ;
        RECT 1844.210 241.500 1849.130 241.640 ;
        RECT 1844.210 241.440 1844.530 241.500 ;
        RECT 1848.810 241.440 1849.130 241.500 ;
        RECT 1848.810 26.080 1849.130 26.140 ;
        RECT 2149.650 26.080 2149.970 26.140 ;
        RECT 1848.810 25.940 2149.970 26.080 ;
        RECT 1848.810 25.880 1849.130 25.940 ;
        RECT 2149.650 25.880 2149.970 25.940 ;
      LAYER via ;
        RECT 1844.240 241.440 1844.500 241.700 ;
        RECT 1848.840 241.440 1849.100 241.700 ;
        RECT 1848.840 25.880 1849.100 26.140 ;
        RECT 2149.680 25.880 2149.940 26.140 ;
      LAYER met2 ;
        RECT 1844.190 260.000 1844.470 264.000 ;
        RECT 1844.300 241.730 1844.440 260.000 ;
        RECT 1844.240 241.410 1844.500 241.730 ;
        RECT 1848.840 241.410 1849.100 241.730 ;
        RECT 1848.900 26.170 1849.040 241.410 ;
        RECT 1848.840 25.850 1849.100 26.170 ;
        RECT 2149.680 25.850 2149.940 26.170 ;
        RECT 2149.740 2.400 2149.880 25.850 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
=======
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 1883.845 23.885 1884.015 24.735 ;
        RECT 1931.685 23.545 1931.855 24.735 ;
        RECT 1932.145 23.205 1933.235 23.375 ;
        RECT 2077.045 22.525 2077.215 23.375 ;
        RECT 2124.885 22.525 2125.055 23.715 ;
        RECT 2125.345 11.645 2125.515 23.375 ;
      LAYER mcon ;
        RECT 1883.845 24.565 1884.015 24.735 ;
        RECT 1931.685 24.565 1931.855 24.735 ;
        RECT 2124.885 23.545 2125.055 23.715 ;
        RECT 1933.065 23.205 1933.235 23.375 ;
        RECT 2077.045 23.205 2077.215 23.375 ;
        RECT 2125.345 23.205 2125.515 23.375 ;
      LAYER met1 ;
        RECT 1883.785 24.720 1884.075 24.765 ;
        RECT 1931.625 24.720 1931.915 24.765 ;
        RECT 1883.785 24.580 1931.915 24.720 ;
        RECT 1883.785 24.535 1884.075 24.580 ;
        RECT 1931.625 24.535 1931.915 24.580 ;
        RECT 1862.610 24.040 1862.930 24.100 ;
        RECT 1883.785 24.040 1884.075 24.085 ;
        RECT 1862.610 23.900 1884.075 24.040 ;
        RECT 1862.610 23.840 1862.930 23.900 ;
        RECT 1883.785 23.855 1884.075 23.900 ;
        RECT 1931.625 23.700 1931.915 23.745 ;
        RECT 2124.825 23.700 2125.115 23.745 ;
        RECT 1931.625 23.560 1932.300 23.700 ;
        RECT 1931.625 23.515 1931.915 23.560 ;
        RECT 1932.160 23.405 1932.300 23.560 ;
        RECT 2014.500 23.560 2041.780 23.700 ;
        RECT 1932.085 23.175 1932.375 23.405 ;
        RECT 1933.005 23.360 1933.295 23.405 ;
        RECT 2014.500 23.360 2014.640 23.560 ;
        RECT 1933.005 23.220 2014.640 23.360 ;
        RECT 2041.640 23.360 2041.780 23.560 ;
        RECT 2124.825 23.560 2125.500 23.700 ;
        RECT 2124.825 23.515 2125.115 23.560 ;
        RECT 2125.360 23.405 2125.500 23.560 ;
        RECT 2076.985 23.360 2077.275 23.405 ;
        RECT 2041.640 23.220 2077.275 23.360 ;
        RECT 1933.005 23.175 1933.295 23.220 ;
        RECT 2076.985 23.175 2077.275 23.220 ;
        RECT 2125.285 23.175 2125.575 23.405 ;
        RECT 2076.985 22.680 2077.275 22.725 ;
        RECT 2124.825 22.680 2125.115 22.725 ;
        RECT 2076.985 22.540 2125.115 22.680 ;
        RECT 2076.985 22.495 2077.275 22.540 ;
        RECT 2124.825 22.495 2125.115 22.540 ;
        RECT 2125.285 11.800 2125.575 11.845 ;
        RECT 2167.590 11.800 2167.910 11.860 ;
        RECT 2125.285 11.660 2167.910 11.800 ;
        RECT 2125.285 11.615 2125.575 11.660 ;
        RECT 2167.590 11.600 2167.910 11.660 ;
      LAYER via ;
        RECT 1862.640 23.840 1862.900 24.100 ;
        RECT 2167.620 11.600 2167.880 11.860 ;
      LAYER met2 ;
        RECT 1861.670 260.170 1861.950 264.000 ;
        RECT 1861.670 260.030 1862.840 260.170 ;
        RECT 1861.670 260.000 1861.950 260.030 ;
        RECT 1862.700 24.130 1862.840 260.030 ;
        RECT 1862.640 23.810 1862.900 24.130 ;
        RECT 2167.620 11.570 2167.880 11.890 ;
        RECT 2167.680 2.400 2167.820 11.570 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
=======
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1879.630 243.680 1879.950 243.740 ;
        RECT 1883.310 243.680 1883.630 243.740 ;
        RECT 1879.630 243.540 1883.630 243.680 ;
        RECT 1879.630 243.480 1879.950 243.540 ;
        RECT 1883.310 243.480 1883.630 243.540 ;
        RECT 1883.310 58.720 1883.630 58.780 ;
        RECT 2185.070 58.720 2185.390 58.780 ;
        RECT 1883.310 58.580 2185.390 58.720 ;
        RECT 1883.310 58.520 1883.630 58.580 ;
        RECT 2185.070 58.520 2185.390 58.580 ;
      LAYER via ;
        RECT 1879.660 243.480 1879.920 243.740 ;
        RECT 1883.340 243.480 1883.600 243.740 ;
        RECT 1883.340 58.520 1883.600 58.780 ;
        RECT 2185.100 58.520 2185.360 58.780 ;
      LAYER met2 ;
        RECT 1879.610 260.000 1879.890 264.000 ;
        RECT 1879.720 243.770 1879.860 260.000 ;
        RECT 1879.660 243.450 1879.920 243.770 ;
        RECT 1883.340 243.450 1883.600 243.770 ;
        RECT 1883.400 58.810 1883.540 243.450 ;
        RECT 1883.340 58.490 1883.600 58.810 ;
        RECT 2185.100 58.490 2185.360 58.810 ;
        RECT 2185.160 2.400 2185.300 58.490 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
=======
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1897.570 244.020 1897.890 244.080 ;
        RECT 1904.010 244.020 1904.330 244.080 ;
        RECT 1897.570 243.880 1904.330 244.020 ;
        RECT 1897.570 243.820 1897.890 243.880 ;
        RECT 1904.010 243.820 1904.330 243.880 ;
        RECT 1904.010 25.400 1904.330 25.460 ;
        RECT 2203.010 25.400 2203.330 25.460 ;
        RECT 1904.010 25.260 2203.330 25.400 ;
        RECT 1904.010 25.200 1904.330 25.260 ;
        RECT 2203.010 25.200 2203.330 25.260 ;
      LAYER via ;
        RECT 1897.600 243.820 1897.860 244.080 ;
        RECT 1904.040 243.820 1904.300 244.080 ;
        RECT 1904.040 25.200 1904.300 25.460 ;
        RECT 2203.040 25.200 2203.300 25.460 ;
      LAYER met2 ;
        RECT 1897.550 260.000 1897.830 264.000 ;
        RECT 1897.660 244.110 1897.800 260.000 ;
        RECT 1897.600 243.790 1897.860 244.110 ;
        RECT 1904.040 243.790 1904.300 244.110 ;
        RECT 1904.100 25.490 1904.240 243.790 ;
        RECT 1904.040 25.170 1904.300 25.490 ;
        RECT 2203.040 25.170 2203.300 25.490 ;
        RECT 2203.100 2.400 2203.240 25.170 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
=======
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1915.510 243.340 1915.830 243.400 ;
        RECT 1921.490 243.340 1921.810 243.400 ;
        RECT 1915.510 243.200 1921.810 243.340 ;
        RECT 1915.510 243.140 1915.830 243.200 ;
        RECT 1921.490 243.140 1921.810 243.200 ;
        RECT 1921.490 65.520 1921.810 65.580 ;
        RECT 2215.430 65.520 2215.750 65.580 ;
        RECT 1921.490 65.380 2215.750 65.520 ;
        RECT 1921.490 65.320 1921.810 65.380 ;
        RECT 2215.430 65.320 2215.750 65.380 ;
        RECT 2215.430 20.640 2215.750 20.700 ;
        RECT 2220.950 20.640 2221.270 20.700 ;
        RECT 2215.430 20.500 2221.270 20.640 ;
        RECT 2215.430 20.440 2215.750 20.500 ;
        RECT 2220.950 20.440 2221.270 20.500 ;
      LAYER via ;
        RECT 1915.540 243.140 1915.800 243.400 ;
        RECT 1921.520 243.140 1921.780 243.400 ;
        RECT 1921.520 65.320 1921.780 65.580 ;
        RECT 2215.460 65.320 2215.720 65.580 ;
        RECT 2215.460 20.440 2215.720 20.700 ;
        RECT 2220.980 20.440 2221.240 20.700 ;
      LAYER met2 ;
        RECT 1915.490 260.000 1915.770 264.000 ;
        RECT 1915.600 243.430 1915.740 260.000 ;
        RECT 1915.540 243.110 1915.800 243.430 ;
        RECT 1921.520 243.110 1921.780 243.430 ;
        RECT 1921.580 65.610 1921.720 243.110 ;
        RECT 1921.520 65.290 1921.780 65.610 ;
        RECT 2215.460 65.290 2215.720 65.610 ;
        RECT 2215.520 20.730 2215.660 65.290 ;
        RECT 2215.460 20.410 2215.720 20.730 ;
        RECT 2220.980 20.410 2221.240 20.730 ;
        RECT 2221.040 2.400 2221.180 20.410 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
=======
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 468.810 134.540 469.130 134.600 ;
        RECT 772.870 134.540 773.190 134.600 ;
        RECT 468.810 134.400 773.190 134.540 ;
        RECT 468.810 134.340 469.130 134.400 ;
        RECT 772.870 134.340 773.190 134.400 ;
      LAYER via ;
        RECT 468.840 134.340 469.100 134.600 ;
        RECT 772.900 134.340 773.160 134.600 ;
      LAYER met2 ;
        RECT 467.410 260.170 467.690 264.000 ;
        RECT 467.410 260.030 469.040 260.170 ;
        RECT 467.410 260.000 467.690 260.030 ;
        RECT 468.900 134.630 469.040 260.030 ;
        RECT 468.840 134.310 469.100 134.630 ;
        RECT 772.900 134.310 773.160 134.630 ;
        RECT 772.960 16.730 773.100 134.310 ;
        RECT 772.960 16.590 775.860 16.730 ;
        RECT 775.720 2.400 775.860 16.590 ;
        RECT 775.510 -4.800 776.070 2.400 ;
=======
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1933.450 244.020 1933.770 244.080 ;
        RECT 1938.510 244.020 1938.830 244.080 ;
        RECT 1933.450 243.880 1938.830 244.020 ;
        RECT 1933.450 243.820 1933.770 243.880 ;
        RECT 1938.510 243.820 1938.830 243.880 ;
        RECT 1938.510 24.720 1938.830 24.780 ;
        RECT 2238.890 24.720 2239.210 24.780 ;
        RECT 1938.510 24.580 2239.210 24.720 ;
        RECT 1938.510 24.520 1938.830 24.580 ;
        RECT 2238.890 24.520 2239.210 24.580 ;
      LAYER via ;
        RECT 1933.480 243.820 1933.740 244.080 ;
        RECT 1938.540 243.820 1938.800 244.080 ;
        RECT 1938.540 24.520 1938.800 24.780 ;
        RECT 2238.920 24.520 2239.180 24.780 ;
      LAYER met2 ;
        RECT 1933.430 260.000 1933.710 264.000 ;
        RECT 1933.540 244.110 1933.680 260.000 ;
        RECT 1933.480 243.790 1933.740 244.110 ;
        RECT 1938.540 243.790 1938.800 244.110 ;
        RECT 1938.600 24.810 1938.740 243.790 ;
        RECT 1938.540 24.490 1938.800 24.810 ;
        RECT 2238.920 24.490 2239.180 24.810 ;
        RECT 2238.980 2.400 2239.120 24.490 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
=======
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 2014.945 23.205 2015.115 24.395 ;
        RECT 2031.965 23.205 2032.135 24.395 ;
        RECT 2111.545 24.225 2111.715 25.075 ;
        RECT 2140.985 24.225 2141.155 25.075 ;
      LAYER mcon ;
        RECT 2111.545 24.905 2111.715 25.075 ;
        RECT 2014.945 24.225 2015.115 24.395 ;
        RECT 2031.965 24.225 2032.135 24.395 ;
        RECT 2140.985 24.905 2141.155 25.075 ;
      LAYER met1 ;
        RECT 2111.485 25.060 2111.775 25.105 ;
        RECT 2140.925 25.060 2141.215 25.105 ;
        RECT 2111.485 24.920 2141.215 25.060 ;
        RECT 2111.485 24.875 2111.775 24.920 ;
        RECT 2140.925 24.875 2141.215 24.920 ;
        RECT 1952.310 24.380 1952.630 24.440 ;
        RECT 2014.885 24.380 2015.175 24.425 ;
        RECT 1952.310 24.240 2015.175 24.380 ;
        RECT 1952.310 24.180 1952.630 24.240 ;
        RECT 2014.885 24.195 2015.175 24.240 ;
        RECT 2031.905 24.380 2032.195 24.425 ;
        RECT 2111.485 24.380 2111.775 24.425 ;
        RECT 2031.905 24.240 2111.775 24.380 ;
        RECT 2031.905 24.195 2032.195 24.240 ;
        RECT 2111.485 24.195 2111.775 24.240 ;
        RECT 2140.925 24.380 2141.215 24.425 ;
        RECT 2140.925 24.240 2208.300 24.380 ;
        RECT 2140.925 24.195 2141.215 24.240 ;
        RECT 2208.160 23.700 2208.300 24.240 ;
        RECT 2256.830 23.700 2257.150 23.760 ;
        RECT 2208.160 23.560 2257.150 23.700 ;
        RECT 2256.830 23.500 2257.150 23.560 ;
        RECT 2014.885 23.360 2015.175 23.405 ;
        RECT 2031.905 23.360 2032.195 23.405 ;
        RECT 2014.885 23.220 2032.195 23.360 ;
        RECT 2014.885 23.175 2015.175 23.220 ;
        RECT 2031.905 23.175 2032.195 23.220 ;
      LAYER via ;
        RECT 1952.340 24.180 1952.600 24.440 ;
        RECT 2256.860 23.500 2257.120 23.760 ;
      LAYER met2 ;
        RECT 1951.370 260.170 1951.650 264.000 ;
        RECT 1951.370 260.030 1952.540 260.170 ;
        RECT 1951.370 260.000 1951.650 260.030 ;
        RECT 1952.400 24.470 1952.540 260.030 ;
        RECT 1952.340 24.150 1952.600 24.470 ;
        RECT 2256.860 23.470 2257.120 23.790 ;
        RECT 2256.920 12.650 2257.060 23.470 ;
        RECT 2256.460 12.510 2257.060 12.650 ;
        RECT 2256.460 2.400 2256.600 12.510 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
=======
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1973.010 25.740 1973.330 25.800 ;
        RECT 2274.310 25.740 2274.630 25.800 ;
        RECT 1973.010 25.600 2274.630 25.740 ;
        RECT 1973.010 25.540 1973.330 25.600 ;
        RECT 2274.310 25.540 2274.630 25.600 ;
      LAYER via ;
        RECT 1973.040 25.540 1973.300 25.800 ;
        RECT 2274.340 25.540 2274.600 25.800 ;
      LAYER met2 ;
        RECT 1969.310 260.170 1969.590 264.000 ;
        RECT 1969.310 260.030 1973.240 260.170 ;
        RECT 1969.310 260.000 1969.590 260.030 ;
        RECT 1973.100 25.830 1973.240 260.030 ;
        RECT 1973.040 25.510 1973.300 25.830 ;
        RECT 2274.340 25.510 2274.600 25.830 ;
        RECT 2274.400 2.400 2274.540 25.510 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
=======
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1986.810 72.320 1987.130 72.380 ;
        RECT 2290.870 72.320 2291.190 72.380 ;
        RECT 1986.810 72.180 2291.190 72.320 ;
        RECT 1986.810 72.120 1987.130 72.180 ;
        RECT 2290.870 72.120 2291.190 72.180 ;
      LAYER via ;
        RECT 1986.840 72.120 1987.100 72.380 ;
        RECT 2290.900 72.120 2291.160 72.380 ;
      LAYER met2 ;
        RECT 1986.790 260.000 1987.070 264.000 ;
        RECT 1986.900 72.410 1987.040 260.000 ;
        RECT 1986.840 72.090 1987.100 72.410 ;
        RECT 2290.900 72.090 2291.160 72.410 ;
        RECT 2290.960 3.130 2291.100 72.090 ;
        RECT 2290.960 2.990 2292.480 3.130 ;
        RECT 2292.340 2.400 2292.480 2.990 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
=======
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2007.510 217.160 2007.830 217.220 ;
        RECT 2304.670 217.160 2304.990 217.220 ;
        RECT 2007.510 217.020 2304.990 217.160 ;
        RECT 2007.510 216.960 2007.830 217.020 ;
        RECT 2304.670 216.960 2304.990 217.020 ;
      LAYER via ;
        RECT 2007.540 216.960 2007.800 217.220 ;
        RECT 2304.700 216.960 2304.960 217.220 ;
      LAYER met2 ;
        RECT 2004.730 260.170 2005.010 264.000 ;
        RECT 2004.730 260.030 2007.740 260.170 ;
        RECT 2004.730 260.000 2005.010 260.030 ;
        RECT 2007.600 217.250 2007.740 260.030 ;
        RECT 2007.540 216.930 2007.800 217.250 ;
        RECT 2304.700 216.930 2304.960 217.250 ;
        RECT 2304.760 16.730 2304.900 216.930 ;
        RECT 2304.760 16.590 2310.420 16.730 ;
        RECT 2310.280 2.400 2310.420 16.590 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
=======
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2022.690 243.340 2023.010 243.400 ;
        RECT 2028.210 243.340 2028.530 243.400 ;
        RECT 2022.690 243.200 2028.530 243.340 ;
        RECT 2022.690 243.140 2023.010 243.200 ;
        RECT 2028.210 243.140 2028.530 243.200 ;
        RECT 2028.210 79.460 2028.530 79.520 ;
        RECT 2325.370 79.460 2325.690 79.520 ;
        RECT 2028.210 79.320 2325.690 79.460 ;
        RECT 2028.210 79.260 2028.530 79.320 ;
        RECT 2325.370 79.260 2325.690 79.320 ;
      LAYER via ;
        RECT 2022.720 243.140 2022.980 243.400 ;
        RECT 2028.240 243.140 2028.500 243.400 ;
        RECT 2028.240 79.260 2028.500 79.520 ;
        RECT 2325.400 79.260 2325.660 79.520 ;
      LAYER met2 ;
        RECT 2022.670 260.000 2022.950 264.000 ;
        RECT 2022.780 243.430 2022.920 260.000 ;
        RECT 2022.720 243.110 2022.980 243.430 ;
        RECT 2028.240 243.110 2028.500 243.430 ;
        RECT 2028.300 79.550 2028.440 243.110 ;
        RECT 2028.240 79.230 2028.500 79.550 ;
        RECT 2325.400 79.230 2325.660 79.550 ;
        RECT 2325.460 9.250 2325.600 79.230 ;
        RECT 2325.460 9.110 2328.360 9.250 ;
        RECT 2328.220 2.400 2328.360 9.110 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
=======
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2042.010 86.260 2042.330 86.320 ;
        RECT 2339.170 86.260 2339.490 86.320 ;
        RECT 2042.010 86.120 2339.490 86.260 ;
        RECT 2042.010 86.060 2042.330 86.120 ;
        RECT 2339.170 86.060 2339.490 86.120 ;
        RECT 2339.170 18.260 2339.490 18.320 ;
        RECT 2345.610 18.260 2345.930 18.320 ;
        RECT 2339.170 18.120 2345.930 18.260 ;
        RECT 2339.170 18.060 2339.490 18.120 ;
        RECT 2345.610 18.060 2345.930 18.120 ;
      LAYER via ;
        RECT 2042.040 86.060 2042.300 86.320 ;
        RECT 2339.200 86.060 2339.460 86.320 ;
        RECT 2339.200 18.060 2339.460 18.320 ;
        RECT 2345.640 18.060 2345.900 18.320 ;
      LAYER met2 ;
        RECT 2040.610 260.170 2040.890 264.000 ;
        RECT 2040.610 260.030 2042.240 260.170 ;
        RECT 2040.610 260.000 2040.890 260.030 ;
        RECT 2042.100 86.350 2042.240 260.030 ;
        RECT 2042.040 86.030 2042.300 86.350 ;
        RECT 2339.200 86.030 2339.460 86.350 ;
        RECT 2339.260 18.350 2339.400 86.030 ;
        RECT 2339.200 18.030 2339.460 18.350 ;
        RECT 2345.640 18.030 2345.900 18.350 ;
        RECT 2345.700 2.400 2345.840 18.030 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
=======
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2058.570 242.320 2058.890 242.380 ;
        RECT 2062.710 242.320 2063.030 242.380 ;
        RECT 2058.570 242.180 2063.030 242.320 ;
        RECT 2058.570 242.120 2058.890 242.180 ;
        RECT 2062.710 242.120 2063.030 242.180 ;
        RECT 2062.710 93.060 2063.030 93.120 ;
        RECT 2359.870 93.060 2360.190 93.120 ;
        RECT 2062.710 92.920 2360.190 93.060 ;
        RECT 2062.710 92.860 2063.030 92.920 ;
        RECT 2359.870 92.860 2360.190 92.920 ;
        RECT 2359.870 2.960 2360.190 3.020 ;
        RECT 2363.550 2.960 2363.870 3.020 ;
        RECT 2359.870 2.820 2363.870 2.960 ;
        RECT 2359.870 2.760 2360.190 2.820 ;
        RECT 2363.550 2.760 2363.870 2.820 ;
      LAYER via ;
        RECT 2058.600 242.120 2058.860 242.380 ;
        RECT 2062.740 242.120 2063.000 242.380 ;
        RECT 2062.740 92.860 2063.000 93.120 ;
        RECT 2359.900 92.860 2360.160 93.120 ;
        RECT 2359.900 2.760 2360.160 3.020 ;
        RECT 2363.580 2.760 2363.840 3.020 ;
      LAYER met2 ;
        RECT 2058.550 260.000 2058.830 264.000 ;
        RECT 2058.660 242.410 2058.800 260.000 ;
        RECT 2058.600 242.090 2058.860 242.410 ;
        RECT 2062.740 242.090 2063.000 242.410 ;
        RECT 2062.800 93.150 2062.940 242.090 ;
        RECT 2062.740 92.830 2063.000 93.150 ;
        RECT 2359.900 92.830 2360.160 93.150 ;
        RECT 2359.960 3.050 2360.100 92.830 ;
        RECT 2359.900 2.730 2360.160 3.050 ;
        RECT 2363.580 2.730 2363.840 3.050 ;
        RECT 2363.640 2.400 2363.780 2.730 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
=======
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2076.050 210.360 2076.370 210.420 ;
        RECT 2380.570 210.360 2380.890 210.420 ;
        RECT 2076.050 210.220 2380.890 210.360 ;
        RECT 2076.050 210.160 2076.370 210.220 ;
        RECT 2380.570 210.160 2380.890 210.220 ;
      LAYER via ;
        RECT 2076.080 210.160 2076.340 210.420 ;
        RECT 2380.600 210.160 2380.860 210.420 ;
      LAYER met2 ;
        RECT 2076.490 260.170 2076.770 264.000 ;
        RECT 2076.140 260.030 2076.770 260.170 ;
        RECT 2076.140 210.450 2076.280 260.030 ;
        RECT 2076.490 260.000 2076.770 260.030 ;
        RECT 2076.080 210.130 2076.340 210.450 ;
        RECT 2380.600 210.130 2380.860 210.450 ;
        RECT 2380.660 3.130 2380.800 210.130 ;
        RECT 2380.660 2.990 2381.720 3.130 ;
        RECT 2381.580 2.400 2381.720 2.990 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
=======
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2097.210 203.560 2097.530 203.620 ;
        RECT 2394.370 203.560 2394.690 203.620 ;
        RECT 2097.210 203.420 2394.690 203.560 ;
        RECT 2097.210 203.360 2097.530 203.420 ;
        RECT 2394.370 203.360 2394.690 203.420 ;
        RECT 2394.370 2.960 2394.690 3.020 ;
        RECT 2399.430 2.960 2399.750 3.020 ;
        RECT 2394.370 2.820 2399.750 2.960 ;
        RECT 2394.370 2.760 2394.690 2.820 ;
        RECT 2399.430 2.760 2399.750 2.820 ;
      LAYER via ;
        RECT 2097.240 203.360 2097.500 203.620 ;
        RECT 2394.400 203.360 2394.660 203.620 ;
        RECT 2394.400 2.760 2394.660 3.020 ;
        RECT 2399.460 2.760 2399.720 3.020 ;
      LAYER met2 ;
        RECT 2094.430 260.170 2094.710 264.000 ;
        RECT 2094.430 260.030 2097.440 260.170 ;
        RECT 2094.430 260.000 2094.710 260.030 ;
        RECT 2097.300 203.650 2097.440 260.030 ;
        RECT 2097.240 203.330 2097.500 203.650 ;
        RECT 2394.400 203.330 2394.660 203.650 ;
        RECT 2394.460 3.050 2394.600 203.330 ;
        RECT 2394.400 2.730 2394.660 3.050 ;
        RECT 2399.460 2.730 2399.720 3.050 ;
        RECT 2399.520 2.400 2399.660 2.730 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
=======
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 485.370 244.020 485.690 244.080 ;
        RECT 489.510 244.020 489.830 244.080 ;
        RECT 485.370 243.880 489.830 244.020 ;
        RECT 485.370 243.820 485.690 243.880 ;
        RECT 489.510 243.820 489.830 243.880 ;
        RECT 489.510 141.340 489.830 141.400 ;
        RECT 794.030 141.340 794.350 141.400 ;
        RECT 489.510 141.200 794.350 141.340 ;
        RECT 489.510 141.140 489.830 141.200 ;
        RECT 794.030 141.140 794.350 141.200 ;
      LAYER via ;
        RECT 485.400 243.820 485.660 244.080 ;
        RECT 489.540 243.820 489.800 244.080 ;
        RECT 489.540 141.140 489.800 141.400 ;
        RECT 794.060 141.140 794.320 141.400 ;
      LAYER met2 ;
        RECT 485.350 260.000 485.630 264.000 ;
        RECT 485.460 244.110 485.600 260.000 ;
        RECT 485.400 243.790 485.660 244.110 ;
        RECT 489.540 243.790 489.800 244.110 ;
        RECT 489.600 141.430 489.740 243.790 ;
        RECT 489.540 141.110 489.800 141.430 ;
        RECT 794.060 141.110 794.320 141.430 ;
        RECT 794.120 7.890 794.260 141.110 ;
        RECT 793.660 7.750 794.260 7.890 ;
        RECT 793.660 2.400 793.800 7.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
=======
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 330.350 244.020 330.670 244.080 ;
        RECT 334.490 244.020 334.810 244.080 ;
        RECT 330.350 243.880 334.810 244.020 ;
        RECT 330.350 243.820 330.670 243.880 ;
        RECT 334.490 243.820 334.810 243.880 ;
        RECT 334.490 79.460 334.810 79.520 ;
        RECT 634.870 79.460 635.190 79.520 ;
        RECT 334.490 79.320 635.190 79.460 ;
        RECT 334.490 79.260 334.810 79.320 ;
        RECT 634.870 79.260 635.190 79.320 ;
      LAYER via ;
        RECT 330.380 243.820 330.640 244.080 ;
        RECT 334.520 243.820 334.780 244.080 ;
        RECT 334.520 79.260 334.780 79.520 ;
        RECT 634.900 79.260 635.160 79.520 ;
      LAYER met2 ;
        RECT 330.330 260.000 330.610 264.000 ;
        RECT 330.440 244.110 330.580 260.000 ;
        RECT 330.380 243.790 330.640 244.110 ;
        RECT 334.520 243.790 334.780 244.110 ;
        RECT 334.580 79.550 334.720 243.790 ;
        RECT 334.520 79.230 334.780 79.550 ;
        RECT 634.900 79.230 635.160 79.550 ;
        RECT 634.960 17.410 635.100 79.230 ;
        RECT 634.960 17.270 639.240 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
=======
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2117.450 99.860 2117.770 99.920 ;
        RECT 2421.970 99.860 2422.290 99.920 ;
        RECT 2117.450 99.720 2422.290 99.860 ;
        RECT 2117.450 99.660 2117.770 99.720 ;
        RECT 2421.970 99.660 2422.290 99.720 ;
      LAYER via ;
        RECT 2117.480 99.660 2117.740 99.920 ;
        RECT 2422.000 99.660 2422.260 99.920 ;
      LAYER met2 ;
        RECT 2117.890 260.170 2118.170 264.000 ;
        RECT 2117.540 260.030 2118.170 260.170 ;
        RECT 2117.540 99.950 2117.680 260.030 ;
        RECT 2117.890 260.000 2118.170 260.030 ;
        RECT 2117.480 99.630 2117.740 99.950 ;
        RECT 2422.000 99.630 2422.260 99.950 ;
        RECT 2422.060 17.410 2422.200 99.630 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
=======
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2138.610 107.340 2138.930 107.400 ;
        RECT 2435.770 107.340 2436.090 107.400 ;
        RECT 2138.610 107.200 2436.090 107.340 ;
        RECT 2138.610 107.140 2138.930 107.200 ;
        RECT 2435.770 107.140 2436.090 107.200 ;
      LAYER via ;
        RECT 2138.640 107.140 2138.900 107.400 ;
        RECT 2435.800 107.140 2436.060 107.400 ;
      LAYER met2 ;
        RECT 2135.830 260.170 2136.110 264.000 ;
        RECT 2135.830 260.030 2138.840 260.170 ;
        RECT 2135.830 260.000 2136.110 260.030 ;
        RECT 2138.700 107.430 2138.840 260.030 ;
        RECT 2138.640 107.110 2138.900 107.430 ;
        RECT 2435.800 107.110 2436.060 107.430 ;
        RECT 2435.860 17.410 2436.000 107.110 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
=======
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2153.790 244.020 2154.110 244.080 ;
        RECT 2159.310 244.020 2159.630 244.080 ;
        RECT 2153.790 243.880 2159.630 244.020 ;
        RECT 2153.790 243.820 2154.110 243.880 ;
        RECT 2159.310 243.820 2159.630 243.880 ;
        RECT 2159.310 114.140 2159.630 114.200 ;
        RECT 2456.470 114.140 2456.790 114.200 ;
        RECT 2159.310 114.000 2456.790 114.140 ;
        RECT 2159.310 113.940 2159.630 114.000 ;
        RECT 2456.470 113.940 2456.790 114.000 ;
      LAYER via ;
        RECT 2153.820 243.820 2154.080 244.080 ;
        RECT 2159.340 243.820 2159.600 244.080 ;
        RECT 2159.340 113.940 2159.600 114.200 ;
        RECT 2456.500 113.940 2456.760 114.200 ;
      LAYER met2 ;
        RECT 2153.770 260.000 2154.050 264.000 ;
        RECT 2153.880 244.110 2154.020 260.000 ;
        RECT 2153.820 243.790 2154.080 244.110 ;
        RECT 2159.340 243.790 2159.600 244.110 ;
        RECT 2159.400 114.230 2159.540 243.790 ;
        RECT 2159.340 113.910 2159.600 114.230 ;
        RECT 2456.500 113.910 2456.760 114.230 ;
        RECT 2456.560 17.410 2456.700 113.910 ;
        RECT 2456.560 17.270 2459.000 17.410 ;
        RECT 2458.860 2.400 2459.000 17.270 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
=======
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2173.110 120.600 2173.430 120.660 ;
        RECT 2470.730 120.600 2471.050 120.660 ;
        RECT 2173.110 120.460 2471.050 120.600 ;
        RECT 2173.110 120.400 2173.430 120.460 ;
        RECT 2470.730 120.400 2471.050 120.460 ;
        RECT 2470.730 17.920 2471.050 17.980 ;
        RECT 2476.710 17.920 2477.030 17.980 ;
        RECT 2470.730 17.780 2477.030 17.920 ;
        RECT 2470.730 17.720 2471.050 17.780 ;
        RECT 2476.710 17.720 2477.030 17.780 ;
      LAYER via ;
        RECT 2173.140 120.400 2173.400 120.660 ;
        RECT 2470.760 120.400 2471.020 120.660 ;
        RECT 2470.760 17.720 2471.020 17.980 ;
        RECT 2476.740 17.720 2477.000 17.980 ;
      LAYER met2 ;
        RECT 2171.710 260.170 2171.990 264.000 ;
        RECT 2171.710 260.030 2173.340 260.170 ;
        RECT 2171.710 260.000 2171.990 260.030 ;
        RECT 2173.200 120.690 2173.340 260.030 ;
        RECT 2173.140 120.370 2173.400 120.690 ;
        RECT 2470.760 120.370 2471.020 120.690 ;
        RECT 2470.820 18.010 2470.960 120.370 ;
        RECT 2470.760 17.690 2471.020 18.010 ;
        RECT 2476.740 17.690 2477.000 18.010 ;
        RECT 2476.800 2.400 2476.940 17.690 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
=======
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2189.670 242.320 2189.990 242.380 ;
        RECT 2193.810 242.320 2194.130 242.380 ;
        RECT 2189.670 242.180 2194.130 242.320 ;
        RECT 2189.670 242.120 2189.990 242.180 ;
        RECT 2193.810 242.120 2194.130 242.180 ;
        RECT 2193.810 128.420 2194.130 128.480 ;
        RECT 2490.970 128.420 2491.290 128.480 ;
        RECT 2193.810 128.280 2491.290 128.420 ;
        RECT 2193.810 128.220 2194.130 128.280 ;
        RECT 2490.970 128.220 2491.290 128.280 ;
      LAYER via ;
        RECT 2189.700 242.120 2189.960 242.380 ;
        RECT 2193.840 242.120 2194.100 242.380 ;
        RECT 2193.840 128.220 2194.100 128.480 ;
        RECT 2491.000 128.220 2491.260 128.480 ;
      LAYER met2 ;
        RECT 2189.650 260.000 2189.930 264.000 ;
        RECT 2189.760 242.410 2189.900 260.000 ;
        RECT 2189.700 242.090 2189.960 242.410 ;
        RECT 2193.840 242.090 2194.100 242.410 ;
        RECT 2193.900 128.510 2194.040 242.090 ;
        RECT 2193.840 128.190 2194.100 128.510 ;
        RECT 2491.000 128.190 2491.260 128.510 ;
        RECT 2491.060 17.410 2491.200 128.190 ;
        RECT 2491.060 17.270 2494.880 17.410 ;
        RECT 2494.740 2.400 2494.880 17.270 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
=======
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2207.150 148.140 2207.470 148.200 ;
        RECT 2512.130 148.140 2512.450 148.200 ;
        RECT 2207.150 148.000 2512.450 148.140 ;
        RECT 2207.150 147.940 2207.470 148.000 ;
        RECT 2512.130 147.940 2512.450 148.000 ;
      LAYER via ;
        RECT 2207.180 147.940 2207.440 148.200 ;
        RECT 2512.160 147.940 2512.420 148.200 ;
      LAYER met2 ;
        RECT 2207.590 260.170 2207.870 264.000 ;
        RECT 2207.240 260.030 2207.870 260.170 ;
        RECT 2207.240 148.230 2207.380 260.030 ;
        RECT 2207.590 260.000 2207.870 260.030 ;
        RECT 2207.180 147.910 2207.440 148.230 ;
        RECT 2512.160 147.910 2512.420 148.230 ;
        RECT 2512.220 2.400 2512.360 147.910 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
=======
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2228.310 135.220 2228.630 135.280 ;
        RECT 2525.470 135.220 2525.790 135.280 ;
        RECT 2228.310 135.080 2525.790 135.220 ;
        RECT 2228.310 135.020 2228.630 135.080 ;
        RECT 2525.470 135.020 2525.790 135.080 ;
      LAYER via ;
        RECT 2228.340 135.020 2228.600 135.280 ;
        RECT 2525.500 135.020 2525.760 135.280 ;
      LAYER met2 ;
        RECT 2225.530 260.170 2225.810 264.000 ;
        RECT 2225.530 260.030 2228.540 260.170 ;
        RECT 2225.530 260.000 2225.810 260.030 ;
        RECT 2228.400 135.310 2228.540 260.030 ;
        RECT 2228.340 134.990 2228.600 135.310 ;
        RECT 2525.500 134.990 2525.760 135.310 ;
        RECT 2525.560 16.730 2525.700 134.990 ;
        RECT 2525.560 16.590 2530.300 16.730 ;
        RECT 2530.160 2.400 2530.300 16.590 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
=======
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2243.030 244.020 2243.350 244.080 ;
        RECT 2248.550 244.020 2248.870 244.080 ;
        RECT 2243.030 243.880 2248.870 244.020 ;
        RECT 2243.030 243.820 2243.350 243.880 ;
        RECT 2248.550 243.820 2248.870 243.880 ;
        RECT 2248.550 141.680 2248.870 141.740 ;
        RECT 2546.170 141.680 2546.490 141.740 ;
        RECT 2248.550 141.540 2546.490 141.680 ;
        RECT 2248.550 141.480 2248.870 141.540 ;
        RECT 2546.170 141.480 2546.490 141.540 ;
      LAYER via ;
        RECT 2243.060 243.820 2243.320 244.080 ;
        RECT 2248.580 243.820 2248.840 244.080 ;
        RECT 2248.580 141.480 2248.840 141.740 ;
        RECT 2546.200 141.480 2546.460 141.740 ;
      LAYER met2 ;
        RECT 2243.010 260.000 2243.290 264.000 ;
        RECT 2243.120 244.110 2243.260 260.000 ;
        RECT 2243.060 243.790 2243.320 244.110 ;
        RECT 2248.580 243.790 2248.840 244.110 ;
        RECT 2248.640 141.770 2248.780 243.790 ;
        RECT 2248.580 141.450 2248.840 141.770 ;
        RECT 2546.200 141.450 2546.460 141.770 ;
        RECT 2546.260 16.730 2546.400 141.450 ;
        RECT 2546.260 16.590 2548.240 16.730 ;
        RECT 2548.100 2.400 2548.240 16.590 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
=======
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2262.810 155.280 2263.130 155.340 ;
        RECT 2560.430 155.280 2560.750 155.340 ;
        RECT 2262.810 155.140 2560.750 155.280 ;
        RECT 2262.810 155.080 2263.130 155.140 ;
        RECT 2560.430 155.080 2560.750 155.140 ;
      LAYER via ;
        RECT 2262.840 155.080 2263.100 155.340 ;
        RECT 2560.460 155.080 2560.720 155.340 ;
      LAYER met2 ;
        RECT 2260.950 260.170 2261.230 264.000 ;
        RECT 2260.950 260.030 2263.040 260.170 ;
        RECT 2260.950 260.000 2261.230 260.030 ;
        RECT 2262.900 155.370 2263.040 260.030 ;
        RECT 2262.840 155.050 2263.100 155.370 ;
        RECT 2560.460 155.050 2560.720 155.370 ;
        RECT 2560.520 16.730 2560.660 155.050 ;
        RECT 2560.520 16.590 2566.180 16.730 ;
        RECT 2566.040 2.400 2566.180 16.590 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
=======
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2278.910 244.020 2279.230 244.080 ;
        RECT 2283.510 244.020 2283.830 244.080 ;
        RECT 2278.910 243.880 2283.830 244.020 ;
        RECT 2278.910 243.820 2279.230 243.880 ;
        RECT 2283.510 243.820 2283.830 243.880 ;
        RECT 2283.510 162.080 2283.830 162.140 ;
        RECT 2580.670 162.080 2580.990 162.140 ;
        RECT 2283.510 161.940 2580.990 162.080 ;
        RECT 2283.510 161.880 2283.830 161.940 ;
        RECT 2580.670 161.880 2580.990 161.940 ;
      LAYER via ;
        RECT 2278.940 243.820 2279.200 244.080 ;
        RECT 2283.540 243.820 2283.800 244.080 ;
        RECT 2283.540 161.880 2283.800 162.140 ;
        RECT 2580.700 161.880 2580.960 162.140 ;
      LAYER met2 ;
        RECT 2278.890 260.000 2279.170 264.000 ;
        RECT 2279.000 244.110 2279.140 260.000 ;
        RECT 2278.940 243.790 2279.200 244.110 ;
        RECT 2283.540 243.790 2283.800 244.110 ;
        RECT 2283.600 162.170 2283.740 243.790 ;
        RECT 2283.540 161.850 2283.800 162.170 ;
        RECT 2580.700 161.850 2580.960 162.170 ;
        RECT 2580.760 16.730 2580.900 161.850 ;
        RECT 2580.760 16.590 2584.120 16.730 ;
        RECT 2583.980 2.400 2584.120 16.590 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
=======
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 510.210 148.140 510.530 148.200 ;
        RECT 814.270 148.140 814.590 148.200 ;
        RECT 510.210 148.000 814.590 148.140 ;
        RECT 510.210 147.940 510.530 148.000 ;
        RECT 814.270 147.940 814.590 148.000 ;
      LAYER via ;
        RECT 510.240 147.940 510.500 148.200 ;
        RECT 814.300 147.940 814.560 148.200 ;
      LAYER met2 ;
        RECT 509.270 260.170 509.550 264.000 ;
        RECT 509.270 260.030 510.440 260.170 ;
        RECT 509.270 260.000 509.550 260.030 ;
        RECT 510.300 148.230 510.440 260.030 ;
        RECT 510.240 147.910 510.500 148.230 ;
        RECT 814.300 147.910 814.560 148.230 ;
        RECT 814.360 17.410 814.500 147.910 ;
        RECT 814.360 17.270 817.720 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
=======
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2296.850 168.880 2297.170 168.940 ;
        RECT 2601.830 168.880 2602.150 168.940 ;
        RECT 2296.850 168.740 2602.150 168.880 ;
        RECT 2296.850 168.680 2297.170 168.740 ;
        RECT 2601.830 168.680 2602.150 168.740 ;
      LAYER via ;
        RECT 2296.880 168.680 2297.140 168.940 ;
        RECT 2601.860 168.680 2602.120 168.940 ;
      LAYER met2 ;
        RECT 2296.830 260.000 2297.110 264.000 ;
        RECT 2296.940 168.970 2297.080 260.000 ;
        RECT 2296.880 168.650 2297.140 168.970 ;
        RECT 2601.860 168.650 2602.120 168.970 ;
        RECT 2601.920 17.410 2602.060 168.650 ;
        RECT 2601.460 17.270 2602.060 17.410 ;
        RECT 2601.460 2.400 2601.600 17.270 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
=======
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2318.010 25.740 2318.330 25.800 ;
        RECT 2619.310 25.740 2619.630 25.800 ;
        RECT 2318.010 25.600 2619.630 25.740 ;
        RECT 2318.010 25.540 2318.330 25.600 ;
        RECT 2619.310 25.540 2619.630 25.600 ;
      LAYER via ;
        RECT 2318.040 25.540 2318.300 25.800 ;
        RECT 2619.340 25.540 2619.600 25.800 ;
      LAYER met2 ;
        RECT 2314.770 260.170 2315.050 264.000 ;
        RECT 2314.770 260.030 2318.240 260.170 ;
        RECT 2314.770 260.000 2315.050 260.030 ;
        RECT 2318.100 25.830 2318.240 260.030 ;
        RECT 2318.040 25.510 2318.300 25.830 ;
        RECT 2619.340 25.510 2619.600 25.830 ;
        RECT 2619.400 2.400 2619.540 25.510 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
=======
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2332.730 244.020 2333.050 244.080 ;
        RECT 2338.710 244.020 2339.030 244.080 ;
        RECT 2332.730 243.880 2339.030 244.020 ;
        RECT 2332.730 243.820 2333.050 243.880 ;
        RECT 2338.710 243.820 2339.030 243.880 ;
        RECT 2338.710 176.020 2339.030 176.080 ;
        RECT 2635.870 176.020 2636.190 176.080 ;
        RECT 2338.710 175.880 2636.190 176.020 ;
        RECT 2338.710 175.820 2339.030 175.880 ;
        RECT 2635.870 175.820 2636.190 175.880 ;
      LAYER via ;
        RECT 2332.760 243.820 2333.020 244.080 ;
        RECT 2338.740 243.820 2339.000 244.080 ;
        RECT 2338.740 175.820 2339.000 176.080 ;
        RECT 2635.900 175.820 2636.160 176.080 ;
      LAYER met2 ;
        RECT 2332.710 260.000 2332.990 264.000 ;
        RECT 2332.820 244.110 2332.960 260.000 ;
        RECT 2332.760 243.790 2333.020 244.110 ;
        RECT 2338.740 243.790 2339.000 244.110 ;
        RECT 2338.800 176.110 2338.940 243.790 ;
        RECT 2338.740 175.790 2339.000 176.110 ;
        RECT 2635.900 175.790 2636.160 176.110 ;
        RECT 2635.960 16.730 2636.100 175.790 ;
        RECT 2635.960 16.590 2637.480 16.730 ;
        RECT 2637.340 2.400 2637.480 16.590 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
=======
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2352.510 182.820 2352.830 182.880 ;
        RECT 2649.670 182.820 2649.990 182.880 ;
        RECT 2352.510 182.680 2649.990 182.820 ;
        RECT 2352.510 182.620 2352.830 182.680 ;
        RECT 2649.670 182.620 2649.990 182.680 ;
      LAYER via ;
        RECT 2352.540 182.620 2352.800 182.880 ;
        RECT 2649.700 182.620 2649.960 182.880 ;
      LAYER met2 ;
        RECT 2350.650 260.170 2350.930 264.000 ;
        RECT 2350.650 260.030 2352.740 260.170 ;
        RECT 2350.650 260.000 2350.930 260.030 ;
        RECT 2352.600 182.910 2352.740 260.030 ;
        RECT 2352.540 182.590 2352.800 182.910 ;
        RECT 2649.700 182.590 2649.960 182.910 ;
        RECT 2649.760 17.410 2649.900 182.590 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
=======
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2368.150 244.020 2368.470 244.080 ;
        RECT 2373.210 244.020 2373.530 244.080 ;
        RECT 2368.150 243.880 2373.530 244.020 ;
        RECT 2368.150 243.820 2368.470 243.880 ;
        RECT 2373.210 243.820 2373.530 243.880 ;
        RECT 2373.210 93.060 2373.530 93.120 ;
        RECT 2670.370 93.060 2670.690 93.120 ;
        RECT 2373.210 92.920 2670.690 93.060 ;
        RECT 2373.210 92.860 2373.530 92.920 ;
        RECT 2670.370 92.860 2670.690 92.920 ;
      LAYER via ;
        RECT 2368.180 243.820 2368.440 244.080 ;
        RECT 2373.240 243.820 2373.500 244.080 ;
        RECT 2373.240 92.860 2373.500 93.120 ;
        RECT 2670.400 92.860 2670.660 93.120 ;
      LAYER met2 ;
        RECT 2368.130 260.000 2368.410 264.000 ;
        RECT 2368.240 244.110 2368.380 260.000 ;
        RECT 2368.180 243.790 2368.440 244.110 ;
        RECT 2373.240 243.790 2373.500 244.110 ;
        RECT 2373.300 93.150 2373.440 243.790 ;
        RECT 2373.240 92.830 2373.500 93.150 ;
        RECT 2670.400 92.830 2670.660 93.150 ;
        RECT 2670.460 17.410 2670.600 92.830 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
=======
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2386.090 248.440 2386.410 248.500 ;
        RECT 2411.390 248.440 2411.710 248.500 ;
        RECT 2386.090 248.300 2411.710 248.440 ;
        RECT 2386.090 248.240 2386.410 248.300 ;
        RECT 2411.390 248.240 2411.710 248.300 ;
        RECT 2411.390 38.320 2411.710 38.380 ;
        RECT 2690.610 38.320 2690.930 38.380 ;
        RECT 2411.390 38.180 2690.930 38.320 ;
        RECT 2411.390 38.120 2411.710 38.180 ;
        RECT 2690.610 38.120 2690.930 38.180 ;
      LAYER via ;
        RECT 2386.120 248.240 2386.380 248.500 ;
        RECT 2411.420 248.240 2411.680 248.500 ;
        RECT 2411.420 38.120 2411.680 38.380 ;
        RECT 2690.640 38.120 2690.900 38.380 ;
      LAYER met2 ;
        RECT 2386.070 260.000 2386.350 264.000 ;
        RECT 2386.180 248.530 2386.320 260.000 ;
        RECT 2386.120 248.210 2386.380 248.530 ;
        RECT 2411.420 248.210 2411.680 248.530 ;
        RECT 2411.480 38.410 2411.620 248.210 ;
        RECT 2411.420 38.090 2411.680 38.410 ;
        RECT 2690.640 38.090 2690.900 38.410 ;
        RECT 2690.700 2.400 2690.840 38.090 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
=======
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2404.030 244.020 2404.350 244.080 ;
        RECT 2407.710 244.020 2408.030 244.080 ;
        RECT 2404.030 243.880 2408.030 244.020 ;
        RECT 2404.030 243.820 2404.350 243.880 ;
        RECT 2407.710 243.820 2408.030 243.880 ;
        RECT 2407.710 100.200 2408.030 100.260 ;
        RECT 2704.870 100.200 2705.190 100.260 ;
        RECT 2407.710 100.060 2705.190 100.200 ;
        RECT 2407.710 100.000 2408.030 100.060 ;
        RECT 2704.870 100.000 2705.190 100.060 ;
      LAYER via ;
        RECT 2404.060 243.820 2404.320 244.080 ;
        RECT 2407.740 243.820 2408.000 244.080 ;
        RECT 2407.740 100.000 2408.000 100.260 ;
        RECT 2704.900 100.000 2705.160 100.260 ;
      LAYER met2 ;
        RECT 2404.010 260.000 2404.290 264.000 ;
        RECT 2404.120 244.110 2404.260 260.000 ;
        RECT 2404.060 243.790 2404.320 244.110 ;
        RECT 2407.740 243.790 2408.000 244.110 ;
        RECT 2407.800 100.290 2407.940 243.790 ;
        RECT 2407.740 99.970 2408.000 100.290 ;
        RECT 2704.900 99.970 2705.160 100.290 ;
        RECT 2704.960 17.410 2705.100 99.970 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
=======
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2421.970 241.640 2422.290 241.700 ;
        RECT 2427.950 241.640 2428.270 241.700 ;
        RECT 2421.970 241.500 2428.270 241.640 ;
        RECT 2421.970 241.440 2422.290 241.500 ;
        RECT 2427.950 241.440 2428.270 241.500 ;
        RECT 2427.950 107.000 2428.270 107.060 ;
        RECT 2725.570 107.000 2725.890 107.060 ;
        RECT 2427.950 106.860 2725.890 107.000 ;
        RECT 2427.950 106.800 2428.270 106.860 ;
        RECT 2725.570 106.800 2725.890 106.860 ;
      LAYER via ;
        RECT 2422.000 241.440 2422.260 241.700 ;
        RECT 2427.980 241.440 2428.240 241.700 ;
        RECT 2427.980 106.800 2428.240 107.060 ;
        RECT 2725.600 106.800 2725.860 107.060 ;
      LAYER met2 ;
        RECT 2421.950 260.000 2422.230 264.000 ;
        RECT 2422.060 241.730 2422.200 260.000 ;
        RECT 2422.000 241.410 2422.260 241.730 ;
        RECT 2427.980 241.410 2428.240 241.730 ;
        RECT 2428.040 107.090 2428.180 241.410 ;
        RECT 2427.980 106.770 2428.240 107.090 ;
        RECT 2725.600 106.770 2725.860 107.090 ;
        RECT 2725.660 17.410 2725.800 106.770 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
=======
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2442.210 113.800 2442.530 113.860 ;
        RECT 2739.370 113.800 2739.690 113.860 ;
        RECT 2442.210 113.660 2739.690 113.800 ;
        RECT 2442.210 113.600 2442.530 113.660 ;
        RECT 2739.370 113.600 2739.690 113.660 ;
      LAYER via ;
        RECT 2442.240 113.600 2442.500 113.860 ;
        RECT 2739.400 113.600 2739.660 113.860 ;
      LAYER met2 ;
        RECT 2439.890 260.170 2440.170 264.000 ;
        RECT 2439.890 260.030 2442.440 260.170 ;
        RECT 2439.890 260.000 2440.170 260.030 ;
        RECT 2442.300 113.890 2442.440 260.030 ;
        RECT 2442.240 113.570 2442.500 113.890 ;
        RECT 2739.400 113.570 2739.660 113.890 ;
        RECT 2739.460 17.410 2739.600 113.570 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
=======
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2457.850 244.020 2458.170 244.080 ;
        RECT 2462.910 244.020 2463.230 244.080 ;
        RECT 2457.850 243.880 2463.230 244.020 ;
        RECT 2457.850 243.820 2458.170 243.880 ;
        RECT 2462.910 243.820 2463.230 243.880 ;
        RECT 2462.910 120.940 2463.230 121.000 ;
        RECT 2760.070 120.940 2760.390 121.000 ;
        RECT 2462.910 120.800 2760.390 120.940 ;
        RECT 2462.910 120.740 2463.230 120.800 ;
        RECT 2760.070 120.740 2760.390 120.800 ;
      LAYER via ;
        RECT 2457.880 243.820 2458.140 244.080 ;
        RECT 2462.940 243.820 2463.200 244.080 ;
        RECT 2462.940 120.740 2463.200 121.000 ;
        RECT 2760.100 120.740 2760.360 121.000 ;
      LAYER met2 ;
        RECT 2457.830 260.000 2458.110 264.000 ;
        RECT 2457.940 244.110 2458.080 260.000 ;
        RECT 2457.880 243.790 2458.140 244.110 ;
        RECT 2462.940 243.790 2463.200 244.110 ;
        RECT 2463.000 121.030 2463.140 243.790 ;
        RECT 2462.940 120.710 2463.200 121.030 ;
        RECT 2760.100 120.710 2760.360 121.030 ;
        RECT 2760.160 17.410 2760.300 120.710 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
=======
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 527.230 244.020 527.550 244.080 ;
        RECT 530.910 244.020 531.230 244.080 ;
        RECT 527.230 243.880 531.230 244.020 ;
        RECT 527.230 243.820 527.550 243.880 ;
        RECT 530.910 243.820 531.230 243.880 ;
        RECT 530.910 155.280 531.230 155.340 ;
        RECT 835.430 155.280 835.750 155.340 ;
        RECT 530.910 155.140 835.750 155.280 ;
        RECT 530.910 155.080 531.230 155.140 ;
        RECT 835.430 155.080 835.750 155.140 ;
      LAYER via ;
        RECT 527.260 243.820 527.520 244.080 ;
        RECT 530.940 243.820 531.200 244.080 ;
        RECT 530.940 155.080 531.200 155.340 ;
        RECT 835.460 155.080 835.720 155.340 ;
      LAYER met2 ;
        RECT 527.210 260.000 527.490 264.000 ;
        RECT 527.320 244.110 527.460 260.000 ;
        RECT 527.260 243.790 527.520 244.110 ;
        RECT 530.940 243.790 531.200 244.110 ;
        RECT 531.000 155.370 531.140 243.790 ;
        RECT 530.940 155.050 531.200 155.370 ;
        RECT 835.460 155.050 835.720 155.370 ;
        RECT 835.520 2.400 835.660 155.050 ;
        RECT 835.310 -4.800 835.870 2.400 ;
=======
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2476.710 127.740 2477.030 127.800 ;
        RECT 2774.330 127.740 2774.650 127.800 ;
        RECT 2476.710 127.600 2774.650 127.740 ;
        RECT 2476.710 127.540 2477.030 127.600 ;
        RECT 2774.330 127.540 2774.650 127.600 ;
      LAYER via ;
        RECT 2476.740 127.540 2477.000 127.800 ;
        RECT 2774.360 127.540 2774.620 127.800 ;
      LAYER met2 ;
        RECT 2475.770 260.170 2476.050 264.000 ;
        RECT 2475.770 260.030 2476.940 260.170 ;
        RECT 2475.770 260.000 2476.050 260.030 ;
        RECT 2476.800 127.830 2476.940 260.030 ;
        RECT 2476.740 127.510 2477.000 127.830 ;
        RECT 2774.360 127.510 2774.620 127.830 ;
        RECT 2774.420 17.410 2774.560 127.510 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
=======
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2493.270 244.020 2493.590 244.080 ;
        RECT 2497.410 244.020 2497.730 244.080 ;
        RECT 2493.270 243.880 2497.730 244.020 ;
        RECT 2493.270 243.820 2493.590 243.880 ;
        RECT 2497.410 243.820 2497.730 243.880 ;
        RECT 2497.410 44.780 2497.730 44.840 ;
        RECT 2797.790 44.780 2798.110 44.840 ;
        RECT 2497.410 44.640 2798.110 44.780 ;
        RECT 2497.410 44.580 2497.730 44.640 ;
        RECT 2797.790 44.580 2798.110 44.640 ;
      LAYER via ;
        RECT 2493.300 243.820 2493.560 244.080 ;
        RECT 2497.440 243.820 2497.700 244.080 ;
        RECT 2497.440 44.580 2497.700 44.840 ;
        RECT 2797.820 44.580 2798.080 44.840 ;
      LAYER met2 ;
        RECT 2493.250 260.000 2493.530 264.000 ;
        RECT 2493.360 244.110 2493.500 260.000 ;
        RECT 2493.300 243.790 2493.560 244.110 ;
        RECT 2497.440 243.790 2497.700 244.110 ;
        RECT 2497.500 44.870 2497.640 243.790 ;
        RECT 2497.440 44.550 2497.700 44.870 ;
        RECT 2797.820 44.550 2798.080 44.870 ;
        RECT 2797.880 2.400 2798.020 44.550 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
=======
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2510.750 134.540 2511.070 134.600 ;
        RECT 2815.730 134.540 2816.050 134.600 ;
        RECT 2510.750 134.400 2816.050 134.540 ;
        RECT 2510.750 134.340 2511.070 134.400 ;
        RECT 2815.730 134.340 2816.050 134.400 ;
      LAYER via ;
        RECT 2510.780 134.340 2511.040 134.600 ;
        RECT 2815.760 134.340 2816.020 134.600 ;
      LAYER met2 ;
        RECT 2511.190 260.170 2511.470 264.000 ;
        RECT 2510.840 260.030 2511.470 260.170 ;
        RECT 2510.840 134.630 2510.980 260.030 ;
        RECT 2511.190 260.000 2511.470 260.030 ;
        RECT 2510.780 134.310 2511.040 134.630 ;
        RECT 2815.760 134.310 2816.020 134.630 ;
        RECT 2815.820 2.400 2815.960 134.310 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
=======
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2531.910 141.340 2532.230 141.400 ;
        RECT 2829.070 141.340 2829.390 141.400 ;
        RECT 2531.910 141.200 2829.390 141.340 ;
        RECT 2531.910 141.140 2532.230 141.200 ;
        RECT 2829.070 141.140 2829.390 141.200 ;
        RECT 2829.070 2.960 2829.390 3.020 ;
        RECT 2833.670 2.960 2833.990 3.020 ;
        RECT 2829.070 2.820 2833.990 2.960 ;
        RECT 2829.070 2.760 2829.390 2.820 ;
        RECT 2833.670 2.760 2833.990 2.820 ;
      LAYER via ;
        RECT 2531.940 141.140 2532.200 141.400 ;
        RECT 2829.100 141.140 2829.360 141.400 ;
        RECT 2829.100 2.760 2829.360 3.020 ;
        RECT 2833.700 2.760 2833.960 3.020 ;
      LAYER met2 ;
        RECT 2529.130 260.170 2529.410 264.000 ;
        RECT 2529.130 260.030 2532.140 260.170 ;
        RECT 2529.130 260.000 2529.410 260.030 ;
        RECT 2532.000 141.430 2532.140 260.030 ;
        RECT 2531.940 141.110 2532.200 141.430 ;
        RECT 2829.100 141.110 2829.360 141.430 ;
        RECT 2829.160 3.050 2829.300 141.110 ;
        RECT 2829.100 2.730 2829.360 3.050 ;
        RECT 2833.700 2.730 2833.960 3.050 ;
        RECT 2833.760 2.400 2833.900 2.730 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
=======
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2547.090 244.020 2547.410 244.080 ;
        RECT 2552.610 244.020 2552.930 244.080 ;
        RECT 2547.090 243.880 2552.930 244.020 ;
        RECT 2547.090 243.820 2547.410 243.880 ;
        RECT 2552.610 243.820 2552.930 243.880 ;
        RECT 2552.610 155.620 2552.930 155.680 ;
        RECT 2849.770 155.620 2850.090 155.680 ;
        RECT 2552.610 155.480 2850.090 155.620 ;
        RECT 2552.610 155.420 2552.930 155.480 ;
        RECT 2849.770 155.420 2850.090 155.480 ;
      LAYER via ;
        RECT 2547.120 243.820 2547.380 244.080 ;
        RECT 2552.640 243.820 2552.900 244.080 ;
        RECT 2552.640 155.420 2552.900 155.680 ;
        RECT 2849.800 155.420 2850.060 155.680 ;
      LAYER met2 ;
        RECT 2547.070 260.000 2547.350 264.000 ;
        RECT 2547.180 244.110 2547.320 260.000 ;
        RECT 2547.120 243.790 2547.380 244.110 ;
        RECT 2552.640 243.790 2552.900 244.110 ;
        RECT 2552.700 155.710 2552.840 243.790 ;
        RECT 2552.640 155.390 2552.900 155.710 ;
        RECT 2849.800 155.390 2850.060 155.710 ;
        RECT 2849.860 17.410 2850.000 155.390 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
=======
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2566.410 18.600 2566.730 18.660 ;
        RECT 2869.090 18.600 2869.410 18.660 ;
        RECT 2566.410 18.460 2869.410 18.600 ;
        RECT 2566.410 18.400 2566.730 18.460 ;
        RECT 2869.090 18.400 2869.410 18.460 ;
      LAYER via ;
        RECT 2566.440 18.400 2566.700 18.660 ;
        RECT 2869.120 18.400 2869.380 18.660 ;
      LAYER met2 ;
        RECT 2565.010 260.170 2565.290 264.000 ;
        RECT 2565.010 260.030 2566.640 260.170 ;
        RECT 2565.010 260.000 2565.290 260.030 ;
        RECT 2566.500 18.690 2566.640 260.030 ;
        RECT 2566.440 18.370 2566.700 18.690 ;
        RECT 2869.120 18.370 2869.380 18.690 ;
        RECT 2869.180 2.400 2869.320 18.370 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
=======
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2582.970 244.020 2583.290 244.080 ;
        RECT 2587.110 244.020 2587.430 244.080 ;
        RECT 2582.970 243.880 2587.430 244.020 ;
        RECT 2582.970 243.820 2583.290 243.880 ;
        RECT 2587.110 243.820 2587.430 243.880 ;
        RECT 2587.110 17.240 2587.430 17.300 ;
        RECT 2887.030 17.240 2887.350 17.300 ;
        RECT 2587.110 17.100 2887.350 17.240 ;
        RECT 2587.110 17.040 2587.430 17.100 ;
        RECT 2887.030 17.040 2887.350 17.100 ;
      LAYER via ;
        RECT 2583.000 243.820 2583.260 244.080 ;
        RECT 2587.140 243.820 2587.400 244.080 ;
        RECT 2587.140 17.040 2587.400 17.300 ;
        RECT 2887.060 17.040 2887.320 17.300 ;
      LAYER met2 ;
        RECT 2582.950 260.000 2583.230 264.000 ;
        RECT 2583.060 244.110 2583.200 260.000 ;
        RECT 2583.000 243.790 2583.260 244.110 ;
        RECT 2587.140 243.790 2587.400 244.110 ;
        RECT 2587.200 17.330 2587.340 243.790 ;
        RECT 2587.140 17.010 2587.400 17.330 ;
        RECT 2887.060 17.010 2887.320 17.330 ;
        RECT 2887.120 2.400 2887.260 17.010 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
=======
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2600.890 260.000 2601.170 264.000 ;
        RECT 2601.000 16.845 2601.140 260.000 ;
        RECT 2600.930 16.475 2601.210 16.845 ;
        RECT 2904.990 16.475 2905.270 16.845 ;
        RECT 2905.060 2.400 2905.200 16.475 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2600.930 16.520 2601.210 16.800 ;
        RECT 2904.990 16.520 2905.270 16.800 ;
      LAYER met3 ;
        RECT 2600.905 16.810 2601.235 16.825 ;
        RECT 2904.965 16.810 2905.295 16.825 ;
        RECT 2600.905 16.510 2905.295 16.810 ;
        RECT 2600.905 16.495 2601.235 16.510 ;
        RECT 2904.965 16.495 2905.295 16.510 ;
=======
        RECT 2904.850 -4.800 2905.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 545.170 244.020 545.490 244.080 ;
        RECT 551.610 244.020 551.930 244.080 ;
        RECT 545.170 243.880 551.930 244.020 ;
        RECT 545.170 243.820 545.490 243.880 ;
        RECT 551.610 243.820 551.930 243.880 ;
        RECT 551.610 162.080 551.930 162.140 ;
        RECT 848.770 162.080 849.090 162.140 ;
        RECT 551.610 161.940 849.090 162.080 ;
        RECT 551.610 161.880 551.930 161.940 ;
        RECT 848.770 161.880 849.090 161.940 ;
      LAYER via ;
        RECT 545.200 243.820 545.460 244.080 ;
        RECT 551.640 243.820 551.900 244.080 ;
        RECT 551.640 161.880 551.900 162.140 ;
        RECT 848.800 161.880 849.060 162.140 ;
      LAYER met2 ;
        RECT 545.150 260.000 545.430 264.000 ;
        RECT 545.260 244.110 545.400 260.000 ;
        RECT 545.200 243.790 545.460 244.110 ;
        RECT 551.640 243.790 551.900 244.110 ;
        RECT 551.700 162.170 551.840 243.790 ;
        RECT 551.640 161.850 551.900 162.170 ;
        RECT 848.800 161.850 849.060 162.170 ;
        RECT 848.860 17.410 849.000 161.850 ;
        RECT 848.860 17.270 853.140 17.410 ;
        RECT 853.000 2.400 853.140 17.270 ;
        RECT 852.790 -4.800 853.350 2.400 ;
=======
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 563.110 231.440 563.430 231.500 ;
        RECT 869.470 231.440 869.790 231.500 ;
        RECT 563.110 231.300 869.790 231.440 ;
        RECT 563.110 231.240 563.430 231.300 ;
        RECT 869.470 231.240 869.790 231.300 ;
      LAYER via ;
        RECT 563.140 231.240 563.400 231.500 ;
        RECT 869.500 231.240 869.760 231.500 ;
      LAYER met2 ;
        RECT 563.090 260.000 563.370 264.000 ;
        RECT 563.200 231.530 563.340 260.000 ;
        RECT 563.140 231.210 563.400 231.530 ;
        RECT 869.500 231.210 869.760 231.530 ;
        RECT 869.560 16.730 869.700 231.210 ;
        RECT 869.560 16.590 871.080 16.730 ;
        RECT 870.940 2.400 871.080 16.590 ;
        RECT 870.730 -4.800 871.290 2.400 ;
=======
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 580.590 244.020 580.910 244.080 ;
        RECT 586.110 244.020 586.430 244.080 ;
        RECT 580.590 243.880 586.430 244.020 ;
        RECT 580.590 243.820 580.910 243.880 ;
        RECT 586.110 243.820 586.430 243.880 ;
        RECT 586.110 168.880 586.430 168.940 ;
        RECT 883.270 168.880 883.590 168.940 ;
        RECT 586.110 168.740 883.590 168.880 ;
        RECT 586.110 168.680 586.430 168.740 ;
        RECT 883.270 168.680 883.590 168.740 ;
      LAYER via ;
        RECT 580.620 243.820 580.880 244.080 ;
        RECT 586.140 243.820 586.400 244.080 ;
        RECT 586.140 168.680 586.400 168.940 ;
        RECT 883.300 168.680 883.560 168.940 ;
      LAYER met2 ;
        RECT 580.570 260.000 580.850 264.000 ;
        RECT 580.680 244.110 580.820 260.000 ;
        RECT 580.620 243.790 580.880 244.110 ;
        RECT 586.140 243.790 586.400 244.110 ;
        RECT 586.200 168.970 586.340 243.790 ;
        RECT 586.140 168.650 586.400 168.970 ;
        RECT 883.300 168.650 883.560 168.970 ;
        RECT 883.360 16.730 883.500 168.650 ;
        RECT 883.360 16.590 889.020 16.730 ;
        RECT 888.880 2.400 889.020 16.590 ;
        RECT 888.670 -4.800 889.230 2.400 ;
=======
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 599.910 176.020 600.230 176.080 ;
        RECT 903.970 176.020 904.290 176.080 ;
        RECT 599.910 175.880 904.290 176.020 ;
        RECT 599.910 175.820 600.230 175.880 ;
        RECT 903.970 175.820 904.290 175.880 ;
      LAYER via ;
        RECT 599.940 175.820 600.200 176.080 ;
        RECT 904.000 175.820 904.260 176.080 ;
      LAYER met2 ;
        RECT 598.510 260.170 598.790 264.000 ;
        RECT 598.510 260.030 600.140 260.170 ;
        RECT 598.510 260.000 598.790 260.030 ;
        RECT 600.000 176.110 600.140 260.030 ;
        RECT 599.940 175.790 600.200 176.110 ;
        RECT 904.000 175.790 904.260 176.110 ;
        RECT 904.060 16.730 904.200 175.790 ;
        RECT 904.060 16.590 906.960 16.730 ;
        RECT 906.820 2.400 906.960 16.590 ;
        RECT 906.610 -4.800 907.170 2.400 ;
=======
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 616.470 244.020 616.790 244.080 ;
        RECT 620.610 244.020 620.930 244.080 ;
        RECT 616.470 243.880 620.930 244.020 ;
        RECT 616.470 243.820 616.790 243.880 ;
        RECT 620.610 243.820 620.930 243.880 ;
        RECT 620.610 182.820 620.930 182.880 ;
        RECT 917.770 182.820 918.090 182.880 ;
        RECT 620.610 182.680 918.090 182.820 ;
        RECT 620.610 182.620 620.930 182.680 ;
        RECT 917.770 182.620 918.090 182.680 ;
        RECT 917.770 17.920 918.090 17.980 ;
        RECT 924.210 17.920 924.530 17.980 ;
        RECT 917.770 17.780 924.530 17.920 ;
        RECT 917.770 17.720 918.090 17.780 ;
        RECT 924.210 17.720 924.530 17.780 ;
      LAYER via ;
        RECT 616.500 243.820 616.760 244.080 ;
        RECT 620.640 243.820 620.900 244.080 ;
        RECT 620.640 182.620 620.900 182.880 ;
        RECT 917.800 182.620 918.060 182.880 ;
        RECT 917.800 17.720 918.060 17.980 ;
        RECT 924.240 17.720 924.500 17.980 ;
      LAYER met2 ;
        RECT 616.450 260.000 616.730 264.000 ;
        RECT 616.560 244.110 616.700 260.000 ;
        RECT 616.500 243.790 616.760 244.110 ;
        RECT 620.640 243.790 620.900 244.110 ;
        RECT 620.700 182.910 620.840 243.790 ;
        RECT 620.640 182.590 620.900 182.910 ;
        RECT 917.800 182.590 918.060 182.910 ;
        RECT 917.860 18.010 918.000 182.590 ;
        RECT 917.800 17.690 918.060 18.010 ;
        RECT 924.240 17.690 924.500 18.010 ;
        RECT 924.300 2.400 924.440 17.690 ;
        RECT 924.090 -4.800 924.650 2.400 ;
=======
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 633.950 196.760 634.270 196.820 ;
        RECT 938.470 196.760 938.790 196.820 ;
        RECT 633.950 196.620 938.790 196.760 ;
        RECT 633.950 196.560 634.270 196.620 ;
        RECT 938.470 196.560 938.790 196.620 ;
      LAYER via ;
        RECT 633.980 196.560 634.240 196.820 ;
        RECT 938.500 196.560 938.760 196.820 ;
      LAYER met2 ;
        RECT 634.390 260.170 634.670 264.000 ;
        RECT 634.040 260.030 634.670 260.170 ;
        RECT 634.040 196.850 634.180 260.030 ;
        RECT 634.390 260.000 634.670 260.030 ;
        RECT 633.980 196.530 634.240 196.850 ;
        RECT 938.500 196.530 938.760 196.850 ;
        RECT 938.560 16.730 938.700 196.530 ;
        RECT 938.560 16.590 942.380 16.730 ;
        RECT 942.240 2.400 942.380 16.590 ;
        RECT 942.030 -4.800 942.590 2.400 ;
=======
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 655.110 224.300 655.430 224.360 ;
        RECT 959.170 224.300 959.490 224.360 ;
        RECT 655.110 224.160 959.490 224.300 ;
        RECT 655.110 224.100 655.430 224.160 ;
        RECT 959.170 224.100 959.490 224.160 ;
      LAYER via ;
        RECT 655.140 224.100 655.400 224.360 ;
        RECT 959.200 224.100 959.460 224.360 ;
      LAYER met2 ;
        RECT 652.330 260.170 652.610 264.000 ;
        RECT 652.330 260.030 655.340 260.170 ;
        RECT 652.330 260.000 652.610 260.030 ;
        RECT 655.200 224.390 655.340 260.030 ;
        RECT 655.140 224.070 655.400 224.390 ;
        RECT 959.200 224.070 959.460 224.390 ;
        RECT 959.260 16.730 959.400 224.070 ;
        RECT 959.260 16.590 960.320 16.730 ;
        RECT 960.180 2.400 960.320 16.590 ;
        RECT 959.970 -4.800 960.530 2.400 ;
=======
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 670.290 244.020 670.610 244.080 ;
        RECT 675.810 244.020 676.130 244.080 ;
        RECT 670.290 243.880 676.130 244.020 ;
        RECT 670.290 243.820 670.610 243.880 ;
        RECT 675.810 243.820 676.130 243.880 ;
        RECT 675.810 189.620 676.130 189.680 ;
        RECT 972.970 189.620 973.290 189.680 ;
        RECT 675.810 189.480 973.290 189.620 ;
        RECT 675.810 189.420 676.130 189.480 ;
        RECT 972.970 189.420 973.290 189.480 ;
      LAYER via ;
        RECT 670.320 243.820 670.580 244.080 ;
        RECT 675.840 243.820 676.100 244.080 ;
        RECT 675.840 189.420 676.100 189.680 ;
        RECT 973.000 189.420 973.260 189.680 ;
      LAYER met2 ;
        RECT 670.270 260.000 670.550 264.000 ;
        RECT 670.380 244.110 670.520 260.000 ;
        RECT 670.320 243.790 670.580 244.110 ;
        RECT 675.840 243.790 676.100 244.110 ;
        RECT 675.900 189.710 676.040 243.790 ;
        RECT 675.840 189.390 676.100 189.710 ;
        RECT 973.000 189.390 973.260 189.710 ;
        RECT 973.060 16.730 973.200 189.390 ;
        RECT 973.060 16.590 978.260 16.730 ;
        RECT 978.120 2.400 978.260 16.590 ;
        RECT 977.910 -4.800 978.470 2.400 ;
=======
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 351.510 189.620 351.830 189.680 ;
        RECT 655.570 189.620 655.890 189.680 ;
        RECT 351.510 189.480 655.890 189.620 ;
        RECT 351.510 189.420 351.830 189.480 ;
        RECT 655.570 189.420 655.890 189.480 ;
      LAYER via ;
        RECT 351.540 189.420 351.800 189.680 ;
        RECT 655.600 189.420 655.860 189.680 ;
      LAYER met2 ;
        RECT 348.270 260.170 348.550 264.000 ;
        RECT 348.270 260.030 351.740 260.170 ;
        RECT 348.270 260.000 348.550 260.030 ;
        RECT 351.600 189.710 351.740 260.030 ;
        RECT 351.540 189.390 351.800 189.710 ;
        RECT 655.600 189.390 655.860 189.710 ;
        RECT 655.660 17.410 655.800 189.390 ;
        RECT 655.660 17.270 657.180 17.410 ;
        RECT 657.040 2.400 657.180 17.270 ;
        RECT 656.830 -4.800 657.390 2.400 ;
=======
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 689.610 37.980 689.930 38.040 ;
        RECT 995.970 37.980 996.290 38.040 ;
        RECT 689.610 37.840 996.290 37.980 ;
        RECT 689.610 37.780 689.930 37.840 ;
        RECT 995.970 37.780 996.290 37.840 ;
      LAYER via ;
        RECT 689.640 37.780 689.900 38.040 ;
        RECT 996.000 37.780 996.260 38.040 ;
      LAYER met2 ;
        RECT 688.210 260.170 688.490 264.000 ;
        RECT 688.210 260.030 689.840 260.170 ;
        RECT 688.210 260.000 688.490 260.030 ;
        RECT 689.700 38.070 689.840 260.030 ;
        RECT 689.640 37.750 689.900 38.070 ;
        RECT 996.000 37.750 996.260 38.070 ;
        RECT 996.060 2.400 996.200 37.750 ;
        RECT 995.850 -4.800 996.410 2.400 ;
=======
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 705.710 244.020 706.030 244.080 ;
        RECT 710.310 244.020 710.630 244.080 ;
        RECT 705.710 243.880 710.630 244.020 ;
        RECT 705.710 243.820 706.030 243.880 ;
        RECT 710.310 243.820 710.630 243.880 ;
        RECT 710.310 203.900 710.630 203.960 ;
        RECT 1007.470 203.900 1007.790 203.960 ;
        RECT 710.310 203.760 1007.790 203.900 ;
        RECT 710.310 203.700 710.630 203.760 ;
        RECT 1007.470 203.700 1007.790 203.760 ;
        RECT 1007.470 17.920 1007.790 17.980 ;
        RECT 1013.450 17.920 1013.770 17.980 ;
        RECT 1007.470 17.780 1013.770 17.920 ;
        RECT 1007.470 17.720 1007.790 17.780 ;
        RECT 1013.450 17.720 1013.770 17.780 ;
      LAYER via ;
        RECT 705.740 243.820 706.000 244.080 ;
        RECT 710.340 243.820 710.600 244.080 ;
        RECT 710.340 203.700 710.600 203.960 ;
        RECT 1007.500 203.700 1007.760 203.960 ;
        RECT 1007.500 17.720 1007.760 17.980 ;
        RECT 1013.480 17.720 1013.740 17.980 ;
      LAYER met2 ;
        RECT 705.690 260.000 705.970 264.000 ;
        RECT 705.800 244.110 705.940 260.000 ;
        RECT 705.740 243.790 706.000 244.110 ;
        RECT 710.340 243.790 710.600 244.110 ;
        RECT 710.400 203.990 710.540 243.790 ;
        RECT 710.340 203.670 710.600 203.990 ;
        RECT 1007.500 203.670 1007.760 203.990 ;
        RECT 1007.560 18.010 1007.700 203.670 ;
        RECT 1007.500 17.690 1007.760 18.010 ;
        RECT 1013.480 17.690 1013.740 18.010 ;
        RECT 1013.540 2.400 1013.680 17.690 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
=======
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 723.650 210.360 723.970 210.420 ;
        RECT 1028.170 210.360 1028.490 210.420 ;
        RECT 723.650 210.220 1028.490 210.360 ;
        RECT 723.650 210.160 723.970 210.220 ;
        RECT 1028.170 210.160 1028.490 210.220 ;
      LAYER via ;
        RECT 723.680 210.160 723.940 210.420 ;
        RECT 1028.200 210.160 1028.460 210.420 ;
      LAYER met2 ;
        RECT 723.630 260.000 723.910 264.000 ;
        RECT 723.740 210.450 723.880 260.000 ;
        RECT 723.680 210.130 723.940 210.450 ;
        RECT 1028.200 210.130 1028.460 210.450 ;
        RECT 1028.260 16.730 1028.400 210.130 ;
        RECT 1028.260 16.590 1031.620 16.730 ;
        RECT 1031.480 2.400 1031.620 16.590 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
=======
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 744.810 217.160 745.130 217.220 ;
        RECT 1049.330 217.160 1049.650 217.220 ;
        RECT 744.810 217.020 1049.650 217.160 ;
        RECT 744.810 216.960 745.130 217.020 ;
        RECT 1049.330 216.960 1049.650 217.020 ;
      LAYER via ;
        RECT 744.840 216.960 745.100 217.220 ;
        RECT 1049.360 216.960 1049.620 217.220 ;
      LAYER met2 ;
        RECT 741.570 260.170 741.850 264.000 ;
        RECT 741.570 260.030 745.040 260.170 ;
        RECT 741.570 260.000 741.850 260.030 ;
        RECT 744.900 217.250 745.040 260.030 ;
        RECT 744.840 216.930 745.100 217.250 ;
        RECT 1049.360 216.930 1049.620 217.250 ;
        RECT 1049.420 2.400 1049.560 216.930 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
=======
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 759.530 244.020 759.850 244.080 ;
        RECT 765.050 244.020 765.370 244.080 ;
        RECT 759.530 243.880 765.370 244.020 ;
        RECT 759.530 243.820 759.850 243.880 ;
        RECT 765.050 243.820 765.370 243.880 ;
        RECT 765.050 148.480 765.370 148.540 ;
        RECT 1062.670 148.480 1062.990 148.540 ;
        RECT 765.050 148.340 1062.990 148.480 ;
        RECT 765.050 148.280 765.370 148.340 ;
        RECT 1062.670 148.280 1062.990 148.340 ;
      LAYER via ;
        RECT 759.560 243.820 759.820 244.080 ;
        RECT 765.080 243.820 765.340 244.080 ;
        RECT 765.080 148.280 765.340 148.540 ;
        RECT 1062.700 148.280 1062.960 148.540 ;
      LAYER met2 ;
        RECT 759.510 260.000 759.790 264.000 ;
        RECT 759.620 244.110 759.760 260.000 ;
        RECT 759.560 243.790 759.820 244.110 ;
        RECT 765.080 243.790 765.340 244.110 ;
        RECT 765.140 148.570 765.280 243.790 ;
        RECT 765.080 148.250 765.340 148.570 ;
        RECT 1062.700 148.250 1062.960 148.570 ;
        RECT 1062.760 16.730 1062.900 148.250 ;
        RECT 1062.760 16.590 1067.500 16.730 ;
        RECT 1067.360 2.400 1067.500 16.590 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
=======
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 779.310 155.620 779.630 155.680 ;
        RECT 1083.370 155.620 1083.690 155.680 ;
        RECT 779.310 155.480 1083.690 155.620 ;
        RECT 779.310 155.420 779.630 155.480 ;
        RECT 1083.370 155.420 1083.690 155.480 ;
      LAYER via ;
        RECT 779.340 155.420 779.600 155.680 ;
        RECT 1083.400 155.420 1083.660 155.680 ;
      LAYER met2 ;
        RECT 777.450 260.170 777.730 264.000 ;
        RECT 777.450 260.030 779.540 260.170 ;
        RECT 777.450 260.000 777.730 260.030 ;
        RECT 779.400 155.710 779.540 260.030 ;
        RECT 779.340 155.390 779.600 155.710 ;
        RECT 1083.400 155.390 1083.660 155.710 ;
        RECT 1083.460 16.730 1083.600 155.390 ;
        RECT 1083.460 16.590 1085.440 16.730 ;
        RECT 1085.300 2.400 1085.440 16.590 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
=======
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 795.410 244.020 795.730 244.080 ;
        RECT 800.010 244.020 800.330 244.080 ;
        RECT 795.410 243.880 800.330 244.020 ;
        RECT 795.410 243.820 795.730 243.880 ;
        RECT 800.010 243.820 800.330 243.880 ;
        RECT 800.010 162.420 800.330 162.480 ;
        RECT 1097.170 162.420 1097.490 162.480 ;
        RECT 800.010 162.280 1097.490 162.420 ;
        RECT 800.010 162.220 800.330 162.280 ;
        RECT 1097.170 162.220 1097.490 162.280 ;
      LAYER via ;
        RECT 795.440 243.820 795.700 244.080 ;
        RECT 800.040 243.820 800.300 244.080 ;
        RECT 800.040 162.220 800.300 162.480 ;
        RECT 1097.200 162.220 1097.460 162.480 ;
      LAYER met2 ;
        RECT 795.390 260.000 795.670 264.000 ;
        RECT 795.500 244.110 795.640 260.000 ;
        RECT 795.440 243.790 795.700 244.110 ;
        RECT 800.040 243.790 800.300 244.110 ;
        RECT 800.100 162.510 800.240 243.790 ;
        RECT 800.040 162.190 800.300 162.510 ;
        RECT 1097.200 162.190 1097.460 162.510 ;
        RECT 1097.260 16.730 1097.400 162.190 ;
        RECT 1097.260 16.590 1102.920 16.730 ;
        RECT 1102.780 2.400 1102.920 16.590 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
=======
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 813.350 231.100 813.670 231.160 ;
        RECT 1117.870 231.100 1118.190 231.160 ;
        RECT 813.350 230.960 1118.190 231.100 ;
        RECT 813.350 230.900 813.670 230.960 ;
        RECT 1117.870 230.900 1118.190 230.960 ;
      LAYER via ;
        RECT 813.380 230.900 813.640 231.160 ;
        RECT 1117.900 230.900 1118.160 231.160 ;
      LAYER met2 ;
        RECT 813.330 260.000 813.610 264.000 ;
        RECT 813.440 231.190 813.580 260.000 ;
        RECT 813.380 230.870 813.640 231.190 ;
        RECT 1117.900 230.870 1118.160 231.190 ;
        RECT 1117.960 16.730 1118.100 230.870 ;
        RECT 1117.960 16.590 1120.860 16.730 ;
        RECT 1120.720 2.400 1120.860 16.590 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
=======
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 830.830 242.660 831.150 242.720 ;
        RECT 838.190 242.660 838.510 242.720 ;
        RECT 830.830 242.520 838.510 242.660 ;
        RECT 830.830 242.460 831.150 242.520 ;
        RECT 838.190 242.460 838.510 242.520 ;
        RECT 838.190 169.220 838.510 169.280 ;
        RECT 1139.030 169.220 1139.350 169.280 ;
        RECT 838.190 169.080 1139.350 169.220 ;
        RECT 838.190 169.020 838.510 169.080 ;
        RECT 1139.030 169.020 1139.350 169.080 ;
      LAYER via ;
        RECT 830.860 242.460 831.120 242.720 ;
        RECT 838.220 242.460 838.480 242.720 ;
        RECT 838.220 169.020 838.480 169.280 ;
        RECT 1139.060 169.020 1139.320 169.280 ;
      LAYER met2 ;
        RECT 830.810 260.000 831.090 264.000 ;
        RECT 830.920 242.750 831.060 260.000 ;
        RECT 830.860 242.430 831.120 242.750 ;
        RECT 838.220 242.430 838.480 242.750 ;
        RECT 838.280 169.310 838.420 242.430 ;
        RECT 838.220 168.990 838.480 169.310 ;
        RECT 1139.060 168.990 1139.320 169.310 ;
        RECT 1139.120 17.410 1139.260 168.990 ;
        RECT 1138.660 17.270 1139.260 17.410 ;
        RECT 1138.660 2.400 1138.800 17.270 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
=======
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 848.770 244.020 849.090 244.080 ;
        RECT 854.750 244.020 855.070 244.080 ;
        RECT 848.770 243.880 855.070 244.020 ;
        RECT 848.770 243.820 849.090 243.880 ;
        RECT 854.750 243.820 855.070 243.880 ;
        RECT 854.750 176.360 855.070 176.420 ;
        RECT 1152.370 176.360 1152.690 176.420 ;
        RECT 854.750 176.220 1152.690 176.360 ;
        RECT 854.750 176.160 855.070 176.220 ;
        RECT 1152.370 176.160 1152.690 176.220 ;
      LAYER via ;
        RECT 848.800 243.820 849.060 244.080 ;
        RECT 854.780 243.820 855.040 244.080 ;
        RECT 854.780 176.160 855.040 176.420 ;
        RECT 1152.400 176.160 1152.660 176.420 ;
      LAYER met2 ;
        RECT 848.750 260.000 849.030 264.000 ;
        RECT 848.860 244.110 849.000 260.000 ;
        RECT 848.800 243.790 849.060 244.110 ;
        RECT 854.780 243.790 855.040 244.110 ;
        RECT 854.840 176.450 854.980 243.790 ;
        RECT 854.780 176.130 855.040 176.450 ;
        RECT 1152.400 176.130 1152.660 176.450 ;
        RECT 1152.460 17.410 1152.600 176.130 ;
        RECT 1152.460 17.270 1156.740 17.410 ;
        RECT 1156.600 2.400 1156.740 17.270 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
=======
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 366.230 244.020 366.550 244.080 ;
        RECT 372.210 244.020 372.530 244.080 ;
        RECT 366.230 243.880 372.530 244.020 ;
        RECT 366.230 243.820 366.550 243.880 ;
        RECT 372.210 243.820 372.530 243.880 ;
        RECT 372.210 203.560 372.530 203.620 ;
        RECT 669.370 203.560 669.690 203.620 ;
        RECT 372.210 203.420 669.690 203.560 ;
        RECT 372.210 203.360 372.530 203.420 ;
        RECT 669.370 203.360 669.690 203.420 ;
      LAYER via ;
        RECT 366.260 243.820 366.520 244.080 ;
        RECT 372.240 243.820 372.500 244.080 ;
        RECT 372.240 203.360 372.500 203.620 ;
        RECT 669.400 203.360 669.660 203.620 ;
      LAYER met2 ;
        RECT 366.210 260.000 366.490 264.000 ;
        RECT 366.320 244.110 366.460 260.000 ;
        RECT 366.260 243.790 366.520 244.110 ;
        RECT 372.240 243.790 372.500 244.110 ;
        RECT 372.300 203.650 372.440 243.790 ;
        RECT 372.240 203.330 372.500 203.650 ;
        RECT 669.400 203.330 669.660 203.650 ;
        RECT 669.460 16.730 669.600 203.330 ;
        RECT 669.460 16.590 674.660 16.730 ;
        RECT 674.520 2.400 674.660 16.590 ;
        RECT 674.310 -4.800 674.870 2.400 ;
=======
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 869.010 24.380 869.330 24.440 ;
        RECT 1173.990 24.380 1174.310 24.440 ;
        RECT 869.010 24.240 1174.310 24.380 ;
        RECT 869.010 24.180 869.330 24.240 ;
        RECT 1173.990 24.180 1174.310 24.240 ;
      LAYER via ;
        RECT 869.040 24.180 869.300 24.440 ;
        RECT 1174.020 24.180 1174.280 24.440 ;
      LAYER met2 ;
        RECT 866.690 260.170 866.970 264.000 ;
        RECT 866.690 260.030 869.240 260.170 ;
        RECT 866.690 260.000 866.970 260.030 ;
        RECT 869.100 24.470 869.240 260.030 ;
        RECT 869.040 24.150 869.300 24.470 ;
        RECT 1174.020 24.150 1174.280 24.470 ;
        RECT 1174.080 2.400 1174.220 24.150 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
=======
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 884.650 244.020 884.970 244.080 ;
        RECT 889.710 244.020 890.030 244.080 ;
        RECT 884.650 243.880 890.030 244.020 ;
        RECT 884.650 243.820 884.970 243.880 ;
        RECT 889.710 243.820 890.030 243.880 ;
        RECT 889.710 183.500 890.030 183.560 ;
        RECT 1186.870 183.500 1187.190 183.560 ;
        RECT 889.710 183.360 1187.190 183.500 ;
        RECT 889.710 183.300 890.030 183.360 ;
        RECT 1186.870 183.300 1187.190 183.360 ;
      LAYER via ;
        RECT 884.680 243.820 884.940 244.080 ;
        RECT 889.740 243.820 890.000 244.080 ;
        RECT 889.740 183.300 890.000 183.560 ;
        RECT 1186.900 183.300 1187.160 183.560 ;
      LAYER met2 ;
        RECT 884.630 260.000 884.910 264.000 ;
        RECT 884.740 244.110 884.880 260.000 ;
        RECT 884.680 243.790 884.940 244.110 ;
        RECT 889.740 243.790 890.000 244.110 ;
        RECT 889.800 183.590 889.940 243.790 ;
        RECT 889.740 183.270 890.000 183.590 ;
        RECT 1186.900 183.270 1187.160 183.590 ;
        RECT 1186.960 17.410 1187.100 183.270 ;
        RECT 1186.960 17.270 1192.160 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
=======
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 903.510 197.100 903.830 197.160 ;
        RECT 1207.570 197.100 1207.890 197.160 ;
        RECT 903.510 196.960 1207.890 197.100 ;
        RECT 903.510 196.900 903.830 196.960 ;
        RECT 1207.570 196.900 1207.890 196.960 ;
      LAYER via ;
        RECT 903.540 196.900 903.800 197.160 ;
        RECT 1207.600 196.900 1207.860 197.160 ;
      LAYER met2 ;
        RECT 902.570 260.170 902.850 264.000 ;
        RECT 902.570 260.030 903.740 260.170 ;
        RECT 902.570 260.000 902.850 260.030 ;
        RECT 903.600 197.190 903.740 260.030 ;
        RECT 903.540 196.870 903.800 197.190 ;
        RECT 1207.600 196.870 1207.860 197.190 ;
        RECT 1207.660 16.730 1207.800 196.870 ;
        RECT 1207.660 16.590 1210.100 16.730 ;
        RECT 1209.960 2.400 1210.100 16.590 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
=======
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 924.210 224.980 924.530 225.040 ;
        RECT 1221.370 224.980 1221.690 225.040 ;
        RECT 924.210 224.840 1221.690 224.980 ;
        RECT 924.210 224.780 924.530 224.840 ;
        RECT 1221.370 224.780 1221.690 224.840 ;
        RECT 1221.370 17.580 1221.690 17.640 ;
        RECT 1227.810 17.580 1228.130 17.640 ;
        RECT 1221.370 17.440 1228.130 17.580 ;
        RECT 1221.370 17.380 1221.690 17.440 ;
        RECT 1227.810 17.380 1228.130 17.440 ;
      LAYER via ;
        RECT 924.240 224.780 924.500 225.040 ;
        RECT 1221.400 224.780 1221.660 225.040 ;
        RECT 1221.400 17.380 1221.660 17.640 ;
        RECT 1227.840 17.380 1228.100 17.640 ;
      LAYER met2 ;
        RECT 920.510 260.170 920.790 264.000 ;
        RECT 920.510 260.030 924.440 260.170 ;
        RECT 920.510 260.000 920.790 260.030 ;
        RECT 924.300 225.070 924.440 260.030 ;
        RECT 924.240 224.750 924.500 225.070 ;
        RECT 1221.400 224.750 1221.660 225.070 ;
        RECT 1221.460 17.670 1221.600 224.750 ;
        RECT 1221.400 17.350 1221.660 17.670 ;
        RECT 1227.840 17.350 1228.100 17.670 ;
        RECT 1227.900 2.400 1228.040 17.350 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
=======
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 938.470 244.020 938.790 244.080 ;
        RECT 944.910 244.020 945.230 244.080 ;
        RECT 938.470 243.880 945.230 244.020 ;
        RECT 938.470 243.820 938.790 243.880 ;
        RECT 944.910 243.820 945.230 243.880 ;
        RECT 944.910 189.960 945.230 190.020 ;
        RECT 1242.070 189.960 1242.390 190.020 ;
        RECT 944.910 189.820 1242.390 189.960 ;
        RECT 944.910 189.760 945.230 189.820 ;
        RECT 1242.070 189.760 1242.390 189.820 ;
      LAYER via ;
        RECT 938.500 243.820 938.760 244.080 ;
        RECT 944.940 243.820 945.200 244.080 ;
        RECT 944.940 189.760 945.200 190.020 ;
        RECT 1242.100 189.760 1242.360 190.020 ;
      LAYER met2 ;
        RECT 938.450 260.000 938.730 264.000 ;
        RECT 938.560 244.110 938.700 260.000 ;
        RECT 938.500 243.790 938.760 244.110 ;
        RECT 944.940 243.790 945.200 244.110 ;
        RECT 945.000 190.050 945.140 243.790 ;
        RECT 944.940 189.730 945.200 190.050 ;
        RECT 1242.100 189.730 1242.360 190.050 ;
        RECT 1242.160 16.730 1242.300 189.730 ;
        RECT 1242.160 16.590 1245.980 16.730 ;
        RECT 1245.840 2.400 1245.980 16.590 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
=======
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 958.710 148.140 959.030 148.200 ;
        RECT 1263.230 148.140 1263.550 148.200 ;
        RECT 958.710 148.000 1263.550 148.140 ;
        RECT 958.710 147.940 959.030 148.000 ;
        RECT 1263.230 147.940 1263.550 148.000 ;
      LAYER via ;
        RECT 958.740 147.940 959.000 148.200 ;
        RECT 1263.260 147.940 1263.520 148.200 ;
      LAYER met2 ;
        RECT 955.930 260.170 956.210 264.000 ;
        RECT 955.930 260.030 958.940 260.170 ;
        RECT 955.930 260.000 956.210 260.030 ;
        RECT 958.800 148.230 958.940 260.030 ;
        RECT 958.740 147.910 959.000 148.230 ;
        RECT 1263.260 147.910 1263.520 148.230 ;
        RECT 1263.320 2.400 1263.460 147.910 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
=======
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 973.890 238.240 974.210 238.300 ;
        RECT 1276.570 238.240 1276.890 238.300 ;
        RECT 973.890 238.100 1276.890 238.240 ;
        RECT 973.890 238.040 974.210 238.100 ;
        RECT 1276.570 238.040 1276.890 238.100 ;
      LAYER via ;
        RECT 973.920 238.040 974.180 238.300 ;
        RECT 1276.600 238.040 1276.860 238.300 ;
      LAYER met2 ;
        RECT 973.870 260.000 974.150 264.000 ;
        RECT 973.980 238.330 974.120 260.000 ;
        RECT 973.920 238.010 974.180 238.330 ;
        RECT 1276.600 238.010 1276.860 238.330 ;
        RECT 1276.660 16.730 1276.800 238.010 ;
        RECT 1276.660 16.590 1281.400 16.730 ;
        RECT 1281.260 2.400 1281.400 16.590 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
=======
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 993.210 203.560 993.530 203.620 ;
        RECT 1297.270 203.560 1297.590 203.620 ;
        RECT 993.210 203.420 1297.590 203.560 ;
        RECT 993.210 203.360 993.530 203.420 ;
        RECT 1297.270 203.360 1297.590 203.420 ;
      LAYER via ;
        RECT 993.240 203.360 993.500 203.620 ;
        RECT 1297.300 203.360 1297.560 203.620 ;
      LAYER met2 ;
        RECT 991.810 260.170 992.090 264.000 ;
        RECT 991.810 260.030 993.440 260.170 ;
        RECT 991.810 260.000 992.090 260.030 ;
        RECT 993.300 203.650 993.440 260.030 ;
        RECT 993.240 203.330 993.500 203.650 ;
        RECT 1297.300 203.330 1297.560 203.650 ;
        RECT 1297.360 17.410 1297.500 203.330 ;
        RECT 1297.360 17.270 1299.340 17.410 ;
        RECT 1299.200 2.400 1299.340 17.270 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
=======
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1009.770 244.020 1010.090 244.080 ;
        RECT 1013.910 244.020 1014.230 244.080 ;
        RECT 1009.770 243.880 1014.230 244.020 ;
        RECT 1009.770 243.820 1010.090 243.880 ;
        RECT 1013.910 243.820 1014.230 243.880 ;
        RECT 1013.910 210.700 1014.230 210.760 ;
        RECT 1311.070 210.700 1311.390 210.760 ;
        RECT 1013.910 210.560 1311.390 210.700 ;
        RECT 1013.910 210.500 1014.230 210.560 ;
        RECT 1311.070 210.500 1311.390 210.560 ;
        RECT 1311.070 19.620 1311.390 19.680 ;
        RECT 1317.050 19.620 1317.370 19.680 ;
        RECT 1311.070 19.480 1317.370 19.620 ;
        RECT 1311.070 19.420 1311.390 19.480 ;
        RECT 1317.050 19.420 1317.370 19.480 ;
      LAYER via ;
        RECT 1009.800 243.820 1010.060 244.080 ;
        RECT 1013.940 243.820 1014.200 244.080 ;
        RECT 1013.940 210.500 1014.200 210.760 ;
        RECT 1311.100 210.500 1311.360 210.760 ;
        RECT 1311.100 19.420 1311.360 19.680 ;
        RECT 1317.080 19.420 1317.340 19.680 ;
      LAYER met2 ;
        RECT 1009.750 260.000 1010.030 264.000 ;
        RECT 1009.860 244.110 1010.000 260.000 ;
        RECT 1009.800 243.790 1010.060 244.110 ;
        RECT 1013.940 243.790 1014.200 244.110 ;
        RECT 1014.000 210.790 1014.140 243.790 ;
        RECT 1013.940 210.470 1014.200 210.790 ;
        RECT 1311.100 210.470 1311.360 210.790 ;
        RECT 1311.160 19.710 1311.300 210.470 ;
        RECT 1311.100 19.390 1311.360 19.710 ;
        RECT 1317.080 19.390 1317.340 19.710 ;
        RECT 1317.140 2.400 1317.280 19.390 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
=======
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1027.250 155.280 1027.570 155.340 ;
        RECT 1331.770 155.280 1332.090 155.340 ;
        RECT 1027.250 155.140 1332.090 155.280 ;
        RECT 1027.250 155.080 1027.570 155.140 ;
        RECT 1331.770 155.080 1332.090 155.140 ;
      LAYER via ;
        RECT 1027.280 155.080 1027.540 155.340 ;
        RECT 1331.800 155.080 1332.060 155.340 ;
      LAYER met2 ;
        RECT 1027.690 260.170 1027.970 264.000 ;
        RECT 1027.340 260.030 1027.970 260.170 ;
        RECT 1027.340 155.370 1027.480 260.030 ;
        RECT 1027.690 260.000 1027.970 260.030 ;
        RECT 1027.280 155.050 1027.540 155.370 ;
        RECT 1331.800 155.050 1332.060 155.370 ;
        RECT 1331.860 17.410 1332.000 155.050 ;
        RECT 1331.860 17.270 1335.220 17.410 ;
        RECT 1335.080 2.400 1335.220 17.270 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
=======
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 384.170 238.240 384.490 238.300 ;
        RECT 690.070 238.240 690.390 238.300 ;
        RECT 384.170 238.100 690.390 238.240 ;
        RECT 384.170 238.040 384.490 238.100 ;
        RECT 690.070 238.040 690.390 238.100 ;
      LAYER via ;
        RECT 384.200 238.040 384.460 238.300 ;
        RECT 690.100 238.040 690.360 238.300 ;
      LAYER met2 ;
        RECT 384.150 260.000 384.430 264.000 ;
        RECT 384.260 238.330 384.400 260.000 ;
        RECT 384.200 238.010 384.460 238.330 ;
        RECT 690.100 238.010 690.360 238.330 ;
        RECT 690.160 16.730 690.300 238.010 ;
        RECT 690.160 16.590 692.600 16.730 ;
        RECT 692.460 2.400 692.600 16.590 ;
        RECT 692.250 -4.800 692.810 2.400 ;
=======
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1048.410 30.840 1048.730 30.900 ;
        RECT 1352.930 30.840 1353.250 30.900 ;
        RECT 1048.410 30.700 1353.250 30.840 ;
        RECT 1048.410 30.640 1048.730 30.700 ;
        RECT 1352.930 30.640 1353.250 30.700 ;
      LAYER via ;
        RECT 1048.440 30.640 1048.700 30.900 ;
        RECT 1352.960 30.640 1353.220 30.900 ;
      LAYER met2 ;
        RECT 1045.630 260.170 1045.910 264.000 ;
        RECT 1045.630 260.030 1048.640 260.170 ;
        RECT 1045.630 260.000 1045.910 260.030 ;
        RECT 1048.500 30.930 1048.640 260.030 ;
        RECT 1048.440 30.610 1048.700 30.930 ;
        RECT 1352.960 30.610 1353.220 30.930 ;
        RECT 1353.020 16.050 1353.160 30.610 ;
        RECT 1352.560 15.910 1353.160 16.050 ;
        RECT 1352.560 2.400 1352.700 15.910 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
=======
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1063.590 244.020 1063.910 244.080 ;
        RECT 1069.110 244.020 1069.430 244.080 ;
        RECT 1063.590 243.880 1069.430 244.020 ;
        RECT 1063.590 243.820 1063.910 243.880 ;
        RECT 1069.110 243.820 1069.430 243.880 ;
        RECT 1069.110 217.160 1069.430 217.220 ;
        RECT 1366.270 217.160 1366.590 217.220 ;
        RECT 1069.110 217.020 1366.590 217.160 ;
        RECT 1069.110 216.960 1069.430 217.020 ;
        RECT 1366.270 216.960 1366.590 217.020 ;
      LAYER via ;
        RECT 1063.620 243.820 1063.880 244.080 ;
        RECT 1069.140 243.820 1069.400 244.080 ;
        RECT 1069.140 216.960 1069.400 217.220 ;
        RECT 1366.300 216.960 1366.560 217.220 ;
      LAYER met2 ;
        RECT 1063.570 260.000 1063.850 264.000 ;
        RECT 1063.680 244.110 1063.820 260.000 ;
        RECT 1063.620 243.790 1063.880 244.110 ;
        RECT 1069.140 243.790 1069.400 244.110 ;
        RECT 1069.200 217.250 1069.340 243.790 ;
        RECT 1069.140 216.930 1069.400 217.250 ;
        RECT 1366.300 216.930 1366.560 217.250 ;
        RECT 1366.360 17.410 1366.500 216.930 ;
        RECT 1366.360 17.270 1370.640 17.410 ;
        RECT 1370.500 2.400 1370.640 17.270 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
=======
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1082.910 162.080 1083.230 162.140 ;
        RECT 1386.970 162.080 1387.290 162.140 ;
        RECT 1082.910 161.940 1387.290 162.080 ;
        RECT 1082.910 161.880 1083.230 161.940 ;
        RECT 1386.970 161.880 1387.290 161.940 ;
      LAYER via ;
        RECT 1082.940 161.880 1083.200 162.140 ;
        RECT 1387.000 161.880 1387.260 162.140 ;
      LAYER met2 ;
        RECT 1081.050 260.170 1081.330 264.000 ;
        RECT 1081.050 260.030 1083.140 260.170 ;
        RECT 1081.050 260.000 1081.330 260.030 ;
        RECT 1083.000 162.170 1083.140 260.030 ;
        RECT 1082.940 161.850 1083.200 162.170 ;
        RECT 1387.000 161.850 1387.260 162.170 ;
        RECT 1387.060 16.900 1387.200 161.850 ;
        RECT 1387.060 16.760 1388.580 16.900 ;
        RECT 1388.440 2.400 1388.580 16.760 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
=======
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1099.010 231.780 1099.330 231.840 ;
        RECT 1400.770 231.780 1401.090 231.840 ;
        RECT 1099.010 231.640 1401.090 231.780 ;
        RECT 1099.010 231.580 1099.330 231.640 ;
        RECT 1400.770 231.580 1401.090 231.640 ;
      LAYER via ;
        RECT 1099.040 231.580 1099.300 231.840 ;
        RECT 1400.800 231.580 1401.060 231.840 ;
      LAYER met2 ;
        RECT 1098.990 260.000 1099.270 264.000 ;
        RECT 1099.100 231.870 1099.240 260.000 ;
        RECT 1099.040 231.550 1099.300 231.870 ;
        RECT 1400.800 231.550 1401.060 231.870 ;
        RECT 1400.860 16.900 1401.000 231.550 ;
        RECT 1400.860 16.760 1406.520 16.900 ;
        RECT 1406.380 2.400 1406.520 16.760 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
=======
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1116.950 168.880 1117.270 168.940 ;
        RECT 1421.470 168.880 1421.790 168.940 ;
        RECT 1116.950 168.740 1421.790 168.880 ;
        RECT 1116.950 168.680 1117.270 168.740 ;
        RECT 1421.470 168.680 1421.790 168.740 ;
      LAYER via ;
        RECT 1116.980 168.680 1117.240 168.940 ;
        RECT 1421.500 168.680 1421.760 168.940 ;
      LAYER met2 ;
        RECT 1116.930 260.000 1117.210 264.000 ;
        RECT 1117.040 168.970 1117.180 260.000 ;
        RECT 1116.980 168.650 1117.240 168.970 ;
        RECT 1421.500 168.650 1421.760 168.970 ;
        RECT 1421.560 16.900 1421.700 168.650 ;
        RECT 1421.560 16.760 1424.000 16.900 ;
        RECT 1423.860 2.400 1424.000 16.760 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
=======
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1138.110 176.700 1138.430 176.760 ;
        RECT 1435.270 176.700 1435.590 176.760 ;
        RECT 1138.110 176.560 1435.590 176.700 ;
        RECT 1138.110 176.500 1138.430 176.560 ;
        RECT 1435.270 176.500 1435.590 176.560 ;
        RECT 1435.270 16.900 1435.590 16.960 ;
        RECT 1441.710 16.900 1442.030 16.960 ;
        RECT 1435.270 16.760 1442.030 16.900 ;
        RECT 1435.270 16.700 1435.590 16.760 ;
        RECT 1441.710 16.700 1442.030 16.760 ;
      LAYER via ;
        RECT 1138.140 176.500 1138.400 176.760 ;
        RECT 1435.300 176.500 1435.560 176.760 ;
        RECT 1435.300 16.700 1435.560 16.960 ;
        RECT 1441.740 16.700 1442.000 16.960 ;
      LAYER met2 ;
        RECT 1134.870 260.170 1135.150 264.000 ;
        RECT 1134.870 260.030 1138.340 260.170 ;
        RECT 1134.870 260.000 1135.150 260.030 ;
        RECT 1138.200 176.790 1138.340 260.030 ;
        RECT 1138.140 176.470 1138.400 176.790 ;
        RECT 1435.300 176.470 1435.560 176.790 ;
        RECT 1435.360 16.990 1435.500 176.470 ;
        RECT 1435.300 16.670 1435.560 16.990 ;
        RECT 1441.740 16.670 1442.000 16.990 ;
        RECT 1441.800 2.400 1441.940 16.670 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
=======
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1152.830 243.340 1153.150 243.400 ;
        RECT 1158.350 243.340 1158.670 243.400 ;
        RECT 1152.830 243.200 1158.670 243.340 ;
        RECT 1152.830 243.140 1153.150 243.200 ;
        RECT 1158.350 243.140 1158.670 243.200 ;
        RECT 1158.350 183.160 1158.670 183.220 ;
        RECT 1455.970 183.160 1456.290 183.220 ;
        RECT 1158.350 183.020 1456.290 183.160 ;
        RECT 1158.350 182.960 1158.670 183.020 ;
        RECT 1455.970 182.960 1456.290 183.020 ;
      LAYER via ;
        RECT 1152.860 243.140 1153.120 243.400 ;
        RECT 1158.380 243.140 1158.640 243.400 ;
        RECT 1158.380 182.960 1158.640 183.220 ;
        RECT 1456.000 182.960 1456.260 183.220 ;
      LAYER met2 ;
        RECT 1152.810 260.000 1153.090 264.000 ;
        RECT 1152.920 243.430 1153.060 260.000 ;
        RECT 1152.860 243.110 1153.120 243.430 ;
        RECT 1158.380 243.110 1158.640 243.430 ;
        RECT 1158.440 183.250 1158.580 243.110 ;
        RECT 1158.380 182.930 1158.640 183.250 ;
        RECT 1456.000 182.930 1456.260 183.250 ;
        RECT 1456.060 16.730 1456.200 182.930 ;
        RECT 1456.060 16.590 1459.880 16.730 ;
        RECT 1459.740 2.400 1459.880 16.590 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
=======
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1172.610 196.760 1172.930 196.820 ;
        RECT 1476.670 196.760 1476.990 196.820 ;
        RECT 1172.610 196.620 1476.990 196.760 ;
        RECT 1172.610 196.560 1172.930 196.620 ;
        RECT 1476.670 196.560 1476.990 196.620 ;
      LAYER via ;
        RECT 1172.640 196.560 1172.900 196.820 ;
        RECT 1476.700 196.560 1476.960 196.820 ;
      LAYER met2 ;
        RECT 1170.750 260.170 1171.030 264.000 ;
        RECT 1170.750 260.030 1172.840 260.170 ;
        RECT 1170.750 260.000 1171.030 260.030 ;
        RECT 1172.700 196.850 1172.840 260.030 ;
        RECT 1172.640 196.530 1172.900 196.850 ;
        RECT 1476.700 196.530 1476.960 196.850 ;
        RECT 1476.760 17.240 1476.900 196.530 ;
        RECT 1476.760 17.100 1477.820 17.240 ;
        RECT 1477.680 2.400 1477.820 17.100 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
=======
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1188.710 244.020 1189.030 244.080 ;
        RECT 1193.310 244.020 1193.630 244.080 ;
        RECT 1188.710 243.880 1193.630 244.020 ;
        RECT 1188.710 243.820 1189.030 243.880 ;
        RECT 1193.310 243.820 1193.630 243.880 ;
        RECT 1193.310 224.640 1193.630 224.700 ;
        RECT 1490.470 224.640 1490.790 224.700 ;
        RECT 1193.310 224.500 1490.790 224.640 ;
        RECT 1193.310 224.440 1193.630 224.500 ;
        RECT 1490.470 224.440 1490.790 224.500 ;
      LAYER via ;
        RECT 1188.740 243.820 1189.000 244.080 ;
        RECT 1193.340 243.820 1193.600 244.080 ;
        RECT 1193.340 224.440 1193.600 224.700 ;
        RECT 1490.500 224.440 1490.760 224.700 ;
      LAYER met2 ;
        RECT 1188.690 260.000 1188.970 264.000 ;
        RECT 1188.800 244.110 1188.940 260.000 ;
        RECT 1188.740 243.790 1189.000 244.110 ;
        RECT 1193.340 243.790 1193.600 244.110 ;
        RECT 1193.400 224.730 1193.540 243.790 ;
        RECT 1193.340 224.410 1193.600 224.730 ;
        RECT 1490.500 224.410 1490.760 224.730 ;
        RECT 1490.560 17.410 1490.700 224.410 ;
        RECT 1490.560 17.270 1495.760 17.410 ;
        RECT 1495.620 2.400 1495.760 17.270 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
=======
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1206.650 189.620 1206.970 189.680 ;
        RECT 1511.170 189.620 1511.490 189.680 ;
        RECT 1206.650 189.480 1511.490 189.620 ;
        RECT 1206.650 189.420 1206.970 189.480 ;
        RECT 1511.170 189.420 1511.490 189.480 ;
      LAYER via ;
        RECT 1206.680 189.420 1206.940 189.680 ;
        RECT 1511.200 189.420 1511.460 189.680 ;
      LAYER met2 ;
        RECT 1206.630 260.000 1206.910 264.000 ;
        RECT 1206.740 189.710 1206.880 260.000 ;
        RECT 1206.680 189.390 1206.940 189.710 ;
        RECT 1511.200 189.390 1511.460 189.710 ;
        RECT 1511.260 17.410 1511.400 189.390 ;
        RECT 1511.260 17.270 1513.240 17.410 ;
        RECT 1513.100 2.400 1513.240 17.270 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
=======
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 402.110 244.020 402.430 244.080 ;
        RECT 406.710 244.020 407.030 244.080 ;
        RECT 402.110 243.880 407.030 244.020 ;
        RECT 402.110 243.820 402.430 243.880 ;
        RECT 406.710 243.820 407.030 243.880 ;
        RECT 406.710 210.360 407.030 210.420 ;
        RECT 703.870 210.360 704.190 210.420 ;
        RECT 406.710 210.220 704.190 210.360 ;
        RECT 406.710 210.160 407.030 210.220 ;
        RECT 703.870 210.160 704.190 210.220 ;
        RECT 703.870 19.280 704.190 19.340 ;
        RECT 710.310 19.280 710.630 19.340 ;
        RECT 703.870 19.140 710.630 19.280 ;
        RECT 703.870 19.080 704.190 19.140 ;
        RECT 710.310 19.080 710.630 19.140 ;
      LAYER via ;
        RECT 402.140 243.820 402.400 244.080 ;
        RECT 406.740 243.820 407.000 244.080 ;
        RECT 406.740 210.160 407.000 210.420 ;
        RECT 703.900 210.160 704.160 210.420 ;
        RECT 703.900 19.080 704.160 19.340 ;
        RECT 710.340 19.080 710.600 19.340 ;
      LAYER met2 ;
        RECT 402.090 260.000 402.370 264.000 ;
        RECT 402.200 244.110 402.340 260.000 ;
        RECT 402.140 243.790 402.400 244.110 ;
        RECT 406.740 243.790 407.000 244.110 ;
        RECT 406.800 210.450 406.940 243.790 ;
        RECT 406.740 210.130 407.000 210.450 ;
        RECT 703.900 210.130 704.160 210.450 ;
        RECT 703.960 19.370 704.100 210.130 ;
        RECT 703.900 19.050 704.160 19.370 ;
        RECT 710.340 19.050 710.600 19.370 ;
        RECT 710.400 2.400 710.540 19.050 ;
        RECT 710.190 -4.800 710.750 2.400 ;
=======
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1227.810 148.820 1228.130 148.880 ;
        RECT 1524.970 148.820 1525.290 148.880 ;
        RECT 1227.810 148.680 1525.290 148.820 ;
        RECT 1227.810 148.620 1228.130 148.680 ;
        RECT 1524.970 148.620 1525.290 148.680 ;
        RECT 1524.970 17.920 1525.290 17.980 ;
        RECT 1530.950 17.920 1531.270 17.980 ;
        RECT 1524.970 17.780 1531.270 17.920 ;
        RECT 1524.970 17.720 1525.290 17.780 ;
        RECT 1530.950 17.720 1531.270 17.780 ;
      LAYER via ;
        RECT 1227.840 148.620 1228.100 148.880 ;
        RECT 1525.000 148.620 1525.260 148.880 ;
        RECT 1525.000 17.720 1525.260 17.980 ;
        RECT 1530.980 17.720 1531.240 17.980 ;
      LAYER met2 ;
        RECT 1224.110 260.170 1224.390 264.000 ;
        RECT 1224.110 260.030 1228.040 260.170 ;
        RECT 1224.110 260.000 1224.390 260.030 ;
        RECT 1227.900 148.910 1228.040 260.030 ;
        RECT 1227.840 148.590 1228.100 148.910 ;
        RECT 1525.000 148.590 1525.260 148.910 ;
        RECT 1525.060 18.010 1525.200 148.590 ;
        RECT 1525.000 17.690 1525.260 18.010 ;
        RECT 1530.980 17.690 1531.240 18.010 ;
        RECT 1531.040 2.400 1531.180 17.690 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
=======
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1242.070 244.020 1242.390 244.080 ;
        RECT 1248.050 244.020 1248.370 244.080 ;
        RECT 1242.070 243.880 1248.370 244.020 ;
        RECT 1242.070 243.820 1242.390 243.880 ;
        RECT 1248.050 243.820 1248.370 243.880 ;
        RECT 1248.050 203.900 1248.370 203.960 ;
        RECT 1545.670 203.900 1545.990 203.960 ;
        RECT 1248.050 203.760 1545.990 203.900 ;
        RECT 1248.050 203.700 1248.370 203.760 ;
        RECT 1545.670 203.700 1545.990 203.760 ;
      LAYER via ;
        RECT 1242.100 243.820 1242.360 244.080 ;
        RECT 1248.080 243.820 1248.340 244.080 ;
        RECT 1248.080 203.700 1248.340 203.960 ;
        RECT 1545.700 203.700 1545.960 203.960 ;
      LAYER met2 ;
        RECT 1242.050 260.000 1242.330 264.000 ;
        RECT 1242.160 244.110 1242.300 260.000 ;
        RECT 1242.100 243.790 1242.360 244.110 ;
        RECT 1248.080 243.790 1248.340 244.110 ;
        RECT 1248.140 203.990 1248.280 243.790 ;
        RECT 1248.080 203.670 1248.340 203.990 ;
        RECT 1545.700 203.670 1545.960 203.990 ;
        RECT 1545.760 16.730 1545.900 203.670 ;
        RECT 1545.760 16.590 1549.120 16.730 ;
        RECT 1548.980 2.400 1549.120 16.590 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
=======
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1262.310 141.680 1262.630 141.740 ;
        RECT 1566.830 141.680 1567.150 141.740 ;
        RECT 1262.310 141.540 1567.150 141.680 ;
        RECT 1262.310 141.480 1262.630 141.540 ;
        RECT 1566.830 141.480 1567.150 141.540 ;
      LAYER via ;
        RECT 1262.340 141.480 1262.600 141.740 ;
        RECT 1566.860 141.480 1567.120 141.740 ;
      LAYER met2 ;
        RECT 1259.990 260.170 1260.270 264.000 ;
        RECT 1259.990 260.030 1262.540 260.170 ;
        RECT 1259.990 260.000 1260.270 260.030 ;
        RECT 1262.400 141.770 1262.540 260.030 ;
        RECT 1262.340 141.450 1262.600 141.770 ;
        RECT 1566.860 141.450 1567.120 141.770 ;
        RECT 1566.920 2.400 1567.060 141.450 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
=======
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1277.950 244.020 1278.270 244.080 ;
        RECT 1283.010 244.020 1283.330 244.080 ;
        RECT 1277.950 243.880 1283.330 244.020 ;
        RECT 1277.950 243.820 1278.270 243.880 ;
        RECT 1283.010 243.820 1283.330 243.880 ;
        RECT 1283.010 211.040 1283.330 211.100 ;
        RECT 1580.170 211.040 1580.490 211.100 ;
        RECT 1283.010 210.900 1580.490 211.040 ;
        RECT 1283.010 210.840 1283.330 210.900 ;
        RECT 1580.170 210.840 1580.490 210.900 ;
      LAYER via ;
        RECT 1277.980 243.820 1278.240 244.080 ;
        RECT 1283.040 243.820 1283.300 244.080 ;
        RECT 1283.040 210.840 1283.300 211.100 ;
        RECT 1580.200 210.840 1580.460 211.100 ;
      LAYER met2 ;
        RECT 1277.930 260.000 1278.210 264.000 ;
        RECT 1278.040 244.110 1278.180 260.000 ;
        RECT 1277.980 243.790 1278.240 244.110 ;
        RECT 1283.040 243.790 1283.300 244.110 ;
        RECT 1283.100 211.130 1283.240 243.790 ;
        RECT 1283.040 210.810 1283.300 211.130 ;
        RECT 1580.200 210.810 1580.460 211.130 ;
        RECT 1580.260 16.730 1580.400 210.810 ;
        RECT 1580.260 16.590 1585.000 16.730 ;
        RECT 1584.860 2.400 1585.000 16.590 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
=======
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1296.810 155.620 1297.130 155.680 ;
        RECT 1600.870 155.620 1601.190 155.680 ;
        RECT 1296.810 155.480 1601.190 155.620 ;
        RECT 1296.810 155.420 1297.130 155.480 ;
        RECT 1600.870 155.420 1601.190 155.480 ;
      LAYER via ;
        RECT 1296.840 155.420 1297.100 155.680 ;
        RECT 1600.900 155.420 1601.160 155.680 ;
      LAYER met2 ;
        RECT 1295.870 260.170 1296.150 264.000 ;
        RECT 1295.870 260.030 1297.040 260.170 ;
        RECT 1295.870 260.000 1296.150 260.030 ;
        RECT 1296.900 155.710 1297.040 260.030 ;
        RECT 1296.840 155.390 1297.100 155.710 ;
        RECT 1600.900 155.390 1601.160 155.710 ;
        RECT 1600.960 16.730 1601.100 155.390 ;
        RECT 1600.960 16.590 1602.480 16.730 ;
        RECT 1602.340 2.400 1602.480 16.590 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
=======
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1313.830 241.640 1314.150 241.700 ;
        RECT 1317.510 241.640 1317.830 241.700 ;
        RECT 1313.830 241.500 1317.830 241.640 ;
        RECT 1313.830 241.440 1314.150 241.500 ;
        RECT 1317.510 241.440 1317.830 241.500 ;
        RECT 1317.510 217.500 1317.830 217.560 ;
        RECT 1615.130 217.500 1615.450 217.560 ;
        RECT 1317.510 217.360 1615.450 217.500 ;
        RECT 1317.510 217.300 1317.830 217.360 ;
        RECT 1615.130 217.300 1615.450 217.360 ;
        RECT 1614.670 62.260 1614.990 62.520 ;
        RECT 1614.760 62.120 1614.900 62.260 ;
        RECT 1620.190 62.120 1620.510 62.180 ;
        RECT 1614.760 61.980 1620.510 62.120 ;
        RECT 1620.190 61.920 1620.510 61.980 ;
        RECT 1620.190 47.980 1620.510 48.240 ;
        RECT 1620.280 47.560 1620.420 47.980 ;
        RECT 1620.190 47.300 1620.510 47.560 ;
      LAYER via ;
        RECT 1313.860 241.440 1314.120 241.700 ;
        RECT 1317.540 241.440 1317.800 241.700 ;
        RECT 1317.540 217.300 1317.800 217.560 ;
        RECT 1615.160 217.300 1615.420 217.560 ;
        RECT 1614.700 62.260 1614.960 62.520 ;
        RECT 1620.220 61.920 1620.480 62.180 ;
        RECT 1620.220 47.980 1620.480 48.240 ;
        RECT 1620.220 47.300 1620.480 47.560 ;
      LAYER met2 ;
        RECT 1313.810 260.000 1314.090 264.000 ;
        RECT 1313.920 241.730 1314.060 260.000 ;
        RECT 1313.860 241.410 1314.120 241.730 ;
        RECT 1317.540 241.410 1317.800 241.730 ;
        RECT 1317.600 217.590 1317.740 241.410 ;
        RECT 1317.540 217.270 1317.800 217.590 ;
        RECT 1615.160 217.270 1615.420 217.590 ;
        RECT 1615.220 193.530 1615.360 217.270 ;
        RECT 1614.760 193.390 1615.360 193.530 ;
        RECT 1614.760 62.550 1614.900 193.390 ;
        RECT 1614.700 62.230 1614.960 62.550 ;
        RECT 1620.220 61.890 1620.480 62.210 ;
        RECT 1620.280 48.270 1620.420 61.890 ;
        RECT 1620.220 47.950 1620.480 48.270 ;
        RECT 1620.220 47.270 1620.480 47.590 ;
        RECT 1620.280 2.400 1620.420 47.270 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
=======
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1331.770 244.020 1332.090 244.080 ;
        RECT 1337.750 244.020 1338.070 244.080 ;
        RECT 1331.770 243.880 1338.070 244.020 ;
        RECT 1331.770 243.820 1332.090 243.880 ;
        RECT 1337.750 243.820 1338.070 243.880 ;
        RECT 1337.750 162.420 1338.070 162.480 ;
        RECT 1635.370 162.420 1635.690 162.480 ;
        RECT 1337.750 162.280 1635.690 162.420 ;
        RECT 1337.750 162.220 1338.070 162.280 ;
        RECT 1635.370 162.220 1635.690 162.280 ;
        RECT 1635.370 62.260 1635.690 62.520 ;
        RECT 1635.460 61.780 1635.600 62.260 ;
        RECT 1638.130 61.780 1638.450 61.840 ;
        RECT 1635.460 61.640 1638.450 61.780 ;
        RECT 1638.130 61.580 1638.450 61.640 ;
        RECT 1638.130 47.980 1638.450 48.240 ;
        RECT 1638.220 47.560 1638.360 47.980 ;
        RECT 1638.130 47.300 1638.450 47.560 ;
      LAYER via ;
        RECT 1331.800 243.820 1332.060 244.080 ;
        RECT 1337.780 243.820 1338.040 244.080 ;
        RECT 1337.780 162.220 1338.040 162.480 ;
        RECT 1635.400 162.220 1635.660 162.480 ;
        RECT 1635.400 62.260 1635.660 62.520 ;
        RECT 1638.160 61.580 1638.420 61.840 ;
        RECT 1638.160 47.980 1638.420 48.240 ;
        RECT 1638.160 47.300 1638.420 47.560 ;
      LAYER met2 ;
        RECT 1331.750 260.000 1332.030 264.000 ;
        RECT 1331.860 244.110 1332.000 260.000 ;
        RECT 1331.800 243.790 1332.060 244.110 ;
        RECT 1337.780 243.790 1338.040 244.110 ;
        RECT 1337.840 162.510 1337.980 243.790 ;
        RECT 1337.780 162.190 1338.040 162.510 ;
        RECT 1635.400 162.190 1635.660 162.510 ;
        RECT 1635.460 62.550 1635.600 162.190 ;
        RECT 1635.400 62.230 1635.660 62.550 ;
        RECT 1638.160 61.550 1638.420 61.870 ;
        RECT 1638.220 48.270 1638.360 61.550 ;
        RECT 1638.160 47.950 1638.420 48.270 ;
        RECT 1638.160 47.270 1638.420 47.590 ;
        RECT 1638.220 2.400 1638.360 47.270 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
=======
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1352.010 169.220 1352.330 169.280 ;
        RECT 1656.070 169.220 1656.390 169.280 ;
        RECT 1352.010 169.080 1656.390 169.220 ;
        RECT 1352.010 169.020 1352.330 169.080 ;
        RECT 1656.070 169.020 1656.390 169.080 ;
      LAYER via ;
        RECT 1352.040 169.020 1352.300 169.280 ;
        RECT 1656.100 169.020 1656.360 169.280 ;
      LAYER met2 ;
        RECT 1349.230 260.170 1349.510 264.000 ;
        RECT 1349.230 260.030 1352.240 260.170 ;
        RECT 1349.230 260.000 1349.510 260.030 ;
        RECT 1352.100 169.310 1352.240 260.030 ;
        RECT 1352.040 168.990 1352.300 169.310 ;
        RECT 1656.100 168.990 1656.360 169.310 ;
        RECT 1656.160 2.400 1656.300 168.990 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
=======
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1367.190 244.020 1367.510 244.080 ;
        RECT 1372.710 244.020 1373.030 244.080 ;
        RECT 1367.190 243.880 1373.030 244.020 ;
        RECT 1367.190 243.820 1367.510 243.880 ;
        RECT 1372.710 243.820 1373.030 243.880 ;
        RECT 1372.710 176.020 1373.030 176.080 ;
        RECT 1669.870 176.020 1670.190 176.080 ;
        RECT 1372.710 175.880 1670.190 176.020 ;
        RECT 1372.710 175.820 1373.030 175.880 ;
        RECT 1669.870 175.820 1670.190 175.880 ;
      LAYER via ;
        RECT 1367.220 243.820 1367.480 244.080 ;
        RECT 1372.740 243.820 1373.000 244.080 ;
        RECT 1372.740 175.820 1373.000 176.080 ;
        RECT 1669.900 175.820 1670.160 176.080 ;
      LAYER met2 ;
        RECT 1367.170 260.000 1367.450 264.000 ;
        RECT 1367.280 244.110 1367.420 260.000 ;
        RECT 1367.220 243.790 1367.480 244.110 ;
        RECT 1372.740 243.790 1373.000 244.110 ;
        RECT 1372.800 176.110 1372.940 243.790 ;
        RECT 1372.740 175.790 1373.000 176.110 ;
        RECT 1669.900 175.790 1670.160 176.110 ;
        RECT 1669.960 16.730 1670.100 175.790 ;
        RECT 1669.960 16.590 1673.780 16.730 ;
        RECT 1673.640 2.400 1673.780 16.590 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
=======
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1386.510 182.820 1386.830 182.880 ;
        RECT 1690.570 182.820 1690.890 182.880 ;
        RECT 1386.510 182.680 1690.890 182.820 ;
        RECT 1386.510 182.620 1386.830 182.680 ;
        RECT 1690.570 182.620 1690.890 182.680 ;
      LAYER via ;
        RECT 1386.540 182.620 1386.800 182.880 ;
        RECT 1690.600 182.620 1690.860 182.880 ;
      LAYER met2 ;
        RECT 1385.110 260.170 1385.390 264.000 ;
        RECT 1385.110 260.030 1386.740 260.170 ;
        RECT 1385.110 260.000 1385.390 260.030 ;
        RECT 1386.600 182.910 1386.740 260.030 ;
        RECT 1386.540 182.590 1386.800 182.910 ;
        RECT 1690.600 182.590 1690.860 182.910 ;
        RECT 1690.660 17.410 1690.800 182.590 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
=======
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 420.510 18.940 420.830 19.000 ;
        RECT 728.250 18.940 728.570 19.000 ;
        RECT 420.510 18.800 728.570 18.940 ;
        RECT 420.510 18.740 420.830 18.800 ;
        RECT 728.250 18.740 728.570 18.800 ;
      LAYER via ;
        RECT 420.540 18.740 420.800 19.000 ;
        RECT 728.280 18.740 728.540 19.000 ;
      LAYER met2 ;
        RECT 420.030 260.170 420.310 264.000 ;
        RECT 420.030 260.030 420.740 260.170 ;
        RECT 420.030 260.000 420.310 260.030 ;
        RECT 420.600 19.030 420.740 260.030 ;
        RECT 420.540 18.710 420.800 19.030 ;
        RECT 728.280 18.710 728.540 19.030 ;
        RECT 728.340 2.400 728.480 18.710 ;
        RECT 728.130 -4.800 728.690 2.400 ;
=======
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1403.070 244.020 1403.390 244.080 ;
        RECT 1407.210 244.020 1407.530 244.080 ;
        RECT 1403.070 243.880 1407.530 244.020 ;
        RECT 1403.070 243.820 1403.390 243.880 ;
        RECT 1407.210 243.820 1407.530 243.880 ;
        RECT 1407.210 197.100 1407.530 197.160 ;
        RECT 1704.370 197.100 1704.690 197.160 ;
        RECT 1407.210 196.960 1704.690 197.100 ;
        RECT 1407.210 196.900 1407.530 196.960 ;
        RECT 1704.370 196.900 1704.690 196.960 ;
      LAYER via ;
        RECT 1403.100 243.820 1403.360 244.080 ;
        RECT 1407.240 243.820 1407.500 244.080 ;
        RECT 1407.240 196.900 1407.500 197.160 ;
        RECT 1704.400 196.900 1704.660 197.160 ;
      LAYER met2 ;
        RECT 1403.050 260.000 1403.330 264.000 ;
        RECT 1403.160 244.110 1403.300 260.000 ;
        RECT 1403.100 243.790 1403.360 244.110 ;
        RECT 1407.240 243.790 1407.500 244.110 ;
        RECT 1407.300 197.190 1407.440 243.790 ;
        RECT 1407.240 196.870 1407.500 197.190 ;
        RECT 1704.400 196.870 1704.660 197.190 ;
        RECT 1704.460 17.410 1704.600 196.870 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
=======
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1420.550 224.300 1420.870 224.360 ;
        RECT 1725.070 224.300 1725.390 224.360 ;
        RECT 1420.550 224.160 1725.390 224.300 ;
        RECT 1420.550 224.100 1420.870 224.160 ;
        RECT 1725.070 224.100 1725.390 224.160 ;
      LAYER via ;
        RECT 1420.580 224.100 1420.840 224.360 ;
        RECT 1725.100 224.100 1725.360 224.360 ;
      LAYER met2 ;
        RECT 1420.990 260.170 1421.270 264.000 ;
        RECT 1420.640 260.030 1421.270 260.170 ;
        RECT 1420.640 224.390 1420.780 260.030 ;
        RECT 1420.990 260.000 1421.270 260.030 ;
        RECT 1420.580 224.070 1420.840 224.390 ;
        RECT 1725.100 224.070 1725.360 224.390 ;
        RECT 1725.160 17.410 1725.300 224.070 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
=======
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1441.710 189.960 1442.030 190.020 ;
        RECT 1738.870 189.960 1739.190 190.020 ;
        RECT 1441.710 189.820 1739.190 189.960 ;
        RECT 1441.710 189.760 1442.030 189.820 ;
        RECT 1738.870 189.760 1739.190 189.820 ;
        RECT 1738.870 18.940 1739.190 19.000 ;
        RECT 1745.310 18.940 1745.630 19.000 ;
        RECT 1738.870 18.800 1745.630 18.940 ;
        RECT 1738.870 18.740 1739.190 18.800 ;
        RECT 1745.310 18.740 1745.630 18.800 ;
      LAYER via ;
        RECT 1441.740 189.760 1442.000 190.020 ;
        RECT 1738.900 189.760 1739.160 190.020 ;
        RECT 1738.900 18.740 1739.160 19.000 ;
        RECT 1745.340 18.740 1745.600 19.000 ;
      LAYER met2 ;
        RECT 1438.930 260.170 1439.210 264.000 ;
        RECT 1438.930 260.030 1441.940 260.170 ;
        RECT 1438.930 260.000 1439.210 260.030 ;
        RECT 1441.800 190.050 1441.940 260.030 ;
        RECT 1441.740 189.730 1442.000 190.050 ;
        RECT 1738.900 189.730 1739.160 190.050 ;
        RECT 1738.960 19.030 1739.100 189.730 ;
        RECT 1738.900 18.710 1739.160 19.030 ;
        RECT 1745.340 18.710 1745.600 19.030 ;
        RECT 1745.400 2.400 1745.540 18.710 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
=======
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1456.890 244.020 1457.210 244.080 ;
        RECT 1462.410 244.020 1462.730 244.080 ;
        RECT 1456.890 243.880 1462.730 244.020 ;
        RECT 1456.890 243.820 1457.210 243.880 ;
        RECT 1462.410 243.820 1462.730 243.880 ;
        RECT 1462.410 148.480 1462.730 148.540 ;
        RECT 1759.570 148.480 1759.890 148.540 ;
        RECT 1462.410 148.340 1759.890 148.480 ;
        RECT 1462.410 148.280 1462.730 148.340 ;
        RECT 1759.570 148.280 1759.890 148.340 ;
      LAYER via ;
        RECT 1456.920 243.820 1457.180 244.080 ;
        RECT 1462.440 243.820 1462.700 244.080 ;
        RECT 1462.440 148.280 1462.700 148.540 ;
        RECT 1759.600 148.280 1759.860 148.540 ;
      LAYER met2 ;
        RECT 1456.870 260.000 1457.150 264.000 ;
        RECT 1456.980 244.110 1457.120 260.000 ;
        RECT 1456.920 243.790 1457.180 244.110 ;
        RECT 1462.440 243.790 1462.700 244.110 ;
        RECT 1462.500 148.570 1462.640 243.790 ;
        RECT 1462.440 148.250 1462.700 148.570 ;
        RECT 1759.600 148.250 1759.860 148.570 ;
        RECT 1759.660 17.410 1759.800 148.250 ;
        RECT 1759.660 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
=======
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1476.210 24.040 1476.530 24.100 ;
        RECT 1780.730 24.040 1781.050 24.100 ;
        RECT 1476.210 23.900 1781.050 24.040 ;
        RECT 1476.210 23.840 1476.530 23.900 ;
        RECT 1780.730 23.840 1781.050 23.900 ;
      LAYER via ;
        RECT 1476.240 23.840 1476.500 24.100 ;
        RECT 1780.760 23.840 1781.020 24.100 ;
      LAYER met2 ;
        RECT 1474.350 260.170 1474.630 264.000 ;
        RECT 1474.350 260.030 1476.440 260.170 ;
        RECT 1474.350 260.000 1474.630 260.030 ;
        RECT 1476.300 24.130 1476.440 260.030 ;
        RECT 1476.240 23.810 1476.500 24.130 ;
        RECT 1780.760 23.810 1781.020 24.130 ;
        RECT 1780.820 2.400 1780.960 23.810 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
=======
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1492.310 244.020 1492.630 244.080 ;
        RECT 1496.910 244.020 1497.230 244.080 ;
        RECT 1492.310 243.880 1497.230 244.020 ;
        RECT 1492.310 243.820 1492.630 243.880 ;
        RECT 1496.910 243.820 1497.230 243.880 ;
        RECT 1496.910 204.240 1497.230 204.300 ;
        RECT 1794.070 204.240 1794.390 204.300 ;
        RECT 1496.910 204.100 1794.390 204.240 ;
        RECT 1496.910 204.040 1497.230 204.100 ;
        RECT 1794.070 204.040 1794.390 204.100 ;
        RECT 1794.070 2.960 1794.390 3.020 ;
        RECT 1798.670 2.960 1798.990 3.020 ;
        RECT 1794.070 2.820 1798.990 2.960 ;
        RECT 1794.070 2.760 1794.390 2.820 ;
        RECT 1798.670 2.760 1798.990 2.820 ;
      LAYER via ;
        RECT 1492.340 243.820 1492.600 244.080 ;
        RECT 1496.940 243.820 1497.200 244.080 ;
        RECT 1496.940 204.040 1497.200 204.300 ;
        RECT 1794.100 204.040 1794.360 204.300 ;
        RECT 1794.100 2.760 1794.360 3.020 ;
        RECT 1798.700 2.760 1798.960 3.020 ;
      LAYER met2 ;
        RECT 1492.290 260.000 1492.570 264.000 ;
        RECT 1492.400 244.110 1492.540 260.000 ;
        RECT 1492.340 243.790 1492.600 244.110 ;
        RECT 1496.940 243.790 1497.200 244.110 ;
        RECT 1497.000 204.330 1497.140 243.790 ;
        RECT 1496.940 204.010 1497.200 204.330 ;
        RECT 1794.100 204.010 1794.360 204.330 ;
        RECT 1794.160 3.050 1794.300 204.010 ;
        RECT 1794.100 2.730 1794.360 3.050 ;
        RECT 1798.700 2.730 1798.960 3.050 ;
        RECT 1798.760 2.400 1798.900 2.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
=======
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1510.250 141.340 1510.570 141.400 ;
        RECT 1814.770 141.340 1815.090 141.400 ;
        RECT 1510.250 141.200 1815.090 141.340 ;
        RECT 1510.250 141.140 1510.570 141.200 ;
        RECT 1814.770 141.140 1815.090 141.200 ;
      LAYER via ;
        RECT 1510.280 141.140 1510.540 141.400 ;
        RECT 1814.800 141.140 1815.060 141.400 ;
      LAYER met2 ;
        RECT 1510.230 260.000 1510.510 264.000 ;
        RECT 1510.340 141.430 1510.480 260.000 ;
        RECT 1510.280 141.110 1510.540 141.430 ;
        RECT 1814.800 141.110 1815.060 141.430 ;
        RECT 1814.860 3.130 1815.000 141.110 ;
        RECT 1814.860 2.990 1816.840 3.130 ;
        RECT 1816.700 2.400 1816.840 2.990 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
=======
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1531.410 155.960 1531.730 156.020 ;
        RECT 1828.570 155.960 1828.890 156.020 ;
        RECT 1531.410 155.820 1828.890 155.960 ;
        RECT 1531.410 155.760 1531.730 155.820 ;
        RECT 1828.570 155.760 1828.890 155.820 ;
        RECT 1828.570 17.240 1828.890 17.300 ;
        RECT 1834.550 17.240 1834.870 17.300 ;
        RECT 1828.570 17.100 1834.870 17.240 ;
        RECT 1828.570 17.040 1828.890 17.100 ;
        RECT 1834.550 17.040 1834.870 17.100 ;
      LAYER via ;
        RECT 1531.440 155.760 1531.700 156.020 ;
        RECT 1828.600 155.760 1828.860 156.020 ;
        RECT 1828.600 17.040 1828.860 17.300 ;
        RECT 1834.580 17.040 1834.840 17.300 ;
      LAYER met2 ;
        RECT 1528.170 260.170 1528.450 264.000 ;
        RECT 1528.170 260.030 1531.640 260.170 ;
        RECT 1528.170 260.000 1528.450 260.030 ;
        RECT 1531.500 156.050 1531.640 260.030 ;
        RECT 1531.440 155.730 1531.700 156.050 ;
        RECT 1828.600 155.730 1828.860 156.050 ;
        RECT 1828.660 17.330 1828.800 155.730 ;
        RECT 1828.600 17.010 1828.860 17.330 ;
        RECT 1834.580 17.010 1834.840 17.330 ;
        RECT 1834.640 2.400 1834.780 17.010 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
=======
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1546.130 244.020 1546.450 244.080 ;
        RECT 1551.650 244.020 1551.970 244.080 ;
        RECT 1546.130 243.880 1551.970 244.020 ;
        RECT 1546.130 243.820 1546.450 243.880 ;
        RECT 1551.650 243.820 1551.970 243.880 ;
        RECT 1551.650 210.360 1551.970 210.420 ;
        RECT 1849.270 210.360 1849.590 210.420 ;
        RECT 1551.650 210.220 1849.590 210.360 ;
        RECT 1551.650 210.160 1551.970 210.220 ;
        RECT 1849.270 210.160 1849.590 210.220 ;
        RECT 1849.270 193.020 1849.590 193.080 ;
        RECT 1849.730 193.020 1850.050 193.080 ;
        RECT 1849.270 192.880 1850.050 193.020 ;
        RECT 1849.270 192.820 1849.590 192.880 ;
        RECT 1849.730 192.820 1850.050 192.880 ;
        RECT 1849.270 137.940 1849.590 138.000 ;
        RECT 1852.490 137.940 1852.810 138.000 ;
        RECT 1849.270 137.800 1852.810 137.940 ;
        RECT 1849.270 137.740 1849.590 137.800 ;
        RECT 1852.490 137.740 1852.810 137.800 ;
      LAYER via ;
        RECT 1546.160 243.820 1546.420 244.080 ;
        RECT 1551.680 243.820 1551.940 244.080 ;
        RECT 1551.680 210.160 1551.940 210.420 ;
        RECT 1849.300 210.160 1849.560 210.420 ;
        RECT 1849.300 192.820 1849.560 193.080 ;
        RECT 1849.760 192.820 1850.020 193.080 ;
        RECT 1849.300 137.740 1849.560 138.000 ;
        RECT 1852.520 137.740 1852.780 138.000 ;
      LAYER met2 ;
        RECT 1546.110 260.000 1546.390 264.000 ;
        RECT 1546.220 244.110 1546.360 260.000 ;
        RECT 1546.160 243.790 1546.420 244.110 ;
        RECT 1551.680 243.790 1551.940 244.110 ;
        RECT 1551.740 210.450 1551.880 243.790 ;
        RECT 1551.680 210.130 1551.940 210.450 ;
        RECT 1849.300 210.130 1849.560 210.450 ;
        RECT 1849.360 193.110 1849.500 210.130 ;
        RECT 1849.300 192.790 1849.560 193.110 ;
        RECT 1849.760 192.790 1850.020 193.110 ;
        RECT 1849.820 145.250 1849.960 192.790 ;
        RECT 1849.360 145.110 1849.960 145.250 ;
        RECT 1849.360 138.030 1849.500 145.110 ;
        RECT 1849.300 137.710 1849.560 138.030 ;
        RECT 1852.520 137.710 1852.780 138.030 ;
        RECT 1852.580 17.240 1852.720 137.710 ;
        RECT 1852.120 17.100 1852.720 17.240 ;
        RECT 1852.120 2.400 1852.260 17.100 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
=======
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1565.910 217.160 1566.230 217.220 ;
        RECT 1870.430 217.160 1870.750 217.220 ;
        RECT 1565.910 217.020 1870.750 217.160 ;
        RECT 1565.910 216.960 1566.230 217.020 ;
        RECT 1870.430 216.960 1870.750 217.020 ;
        RECT 1870.430 14.180 1870.750 14.240 ;
        RECT 1870.060 14.040 1870.750 14.180 ;
        RECT 1870.060 13.900 1870.200 14.040 ;
        RECT 1870.430 13.980 1870.750 14.040 ;
        RECT 1869.970 13.640 1870.290 13.900 ;
      LAYER via ;
        RECT 1565.940 216.960 1566.200 217.220 ;
        RECT 1870.460 216.960 1870.720 217.220 ;
        RECT 1870.460 13.980 1870.720 14.240 ;
        RECT 1870.000 13.640 1870.260 13.900 ;
      LAYER met2 ;
        RECT 1564.050 260.170 1564.330 264.000 ;
        RECT 1564.050 260.030 1566.140 260.170 ;
        RECT 1564.050 260.000 1564.330 260.030 ;
        RECT 1566.000 217.250 1566.140 260.030 ;
        RECT 1565.940 216.930 1566.200 217.250 ;
        RECT 1870.460 216.930 1870.720 217.250 ;
        RECT 1870.520 14.270 1870.660 216.930 ;
        RECT 1870.460 13.950 1870.720 14.270 ;
        RECT 1870.000 13.610 1870.260 13.930 ;
        RECT 1870.060 2.400 1870.200 13.610 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
=======
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 441.210 17.580 441.530 17.640 ;
        RECT 746.190 17.580 746.510 17.640 ;
        RECT 441.210 17.440 746.510 17.580 ;
        RECT 441.210 17.380 441.530 17.440 ;
        RECT 746.190 17.380 746.510 17.440 ;
      LAYER via ;
        RECT 441.240 17.380 441.500 17.640 ;
        RECT 746.220 17.380 746.480 17.640 ;
      LAYER met2 ;
        RECT 437.970 260.170 438.250 264.000 ;
        RECT 437.970 260.030 441.440 260.170 ;
        RECT 437.970 260.000 438.250 260.030 ;
        RECT 441.300 17.670 441.440 260.030 ;
        RECT 441.240 17.350 441.500 17.670 ;
        RECT 746.220 17.350 746.480 17.670 ;
        RECT 746.280 2.400 746.420 17.350 ;
        RECT 746.070 -4.800 746.630 2.400 ;
=======
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1582.010 244.020 1582.330 244.080 ;
        RECT 1586.610 244.020 1586.930 244.080 ;
        RECT 1582.010 243.880 1586.930 244.020 ;
        RECT 1582.010 243.820 1582.330 243.880 ;
        RECT 1586.610 243.820 1586.930 243.880 ;
        RECT 1586.610 162.760 1586.930 162.820 ;
        RECT 1883.770 162.760 1884.090 162.820 ;
        RECT 1586.610 162.620 1884.090 162.760 ;
        RECT 1586.610 162.560 1586.930 162.620 ;
        RECT 1883.770 162.560 1884.090 162.620 ;
        RECT 1883.770 62.120 1884.090 62.180 ;
        RECT 1887.910 62.120 1888.230 62.180 ;
        RECT 1883.770 61.980 1888.230 62.120 ;
        RECT 1883.770 61.920 1884.090 61.980 ;
        RECT 1887.910 61.920 1888.230 61.980 ;
      LAYER via ;
        RECT 1582.040 243.820 1582.300 244.080 ;
        RECT 1586.640 243.820 1586.900 244.080 ;
        RECT 1586.640 162.560 1586.900 162.820 ;
        RECT 1883.800 162.560 1884.060 162.820 ;
        RECT 1883.800 61.920 1884.060 62.180 ;
        RECT 1887.940 61.920 1888.200 62.180 ;
      LAYER met2 ;
        RECT 1581.990 260.000 1582.270 264.000 ;
        RECT 1582.100 244.110 1582.240 260.000 ;
        RECT 1582.040 243.790 1582.300 244.110 ;
        RECT 1586.640 243.790 1586.900 244.110 ;
        RECT 1586.700 162.850 1586.840 243.790 ;
        RECT 1586.640 162.530 1586.900 162.850 ;
        RECT 1883.800 162.530 1884.060 162.850 ;
        RECT 1883.860 62.210 1884.000 162.530 ;
        RECT 1883.800 61.890 1884.060 62.210 ;
        RECT 1887.940 61.890 1888.200 62.210 ;
        RECT 1888.000 2.400 1888.140 61.890 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
=======
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1600.410 168.880 1600.730 168.940 ;
        RECT 1904.470 168.880 1904.790 168.940 ;
        RECT 1600.410 168.740 1904.790 168.880 ;
        RECT 1600.410 168.680 1600.730 168.740 ;
        RECT 1904.470 168.680 1904.790 168.740 ;
      LAYER via ;
        RECT 1600.440 168.680 1600.700 168.940 ;
        RECT 1904.500 168.680 1904.760 168.940 ;
      LAYER met2 ;
        RECT 1599.470 260.170 1599.750 264.000 ;
        RECT 1599.470 260.030 1600.640 260.170 ;
        RECT 1599.470 260.000 1599.750 260.030 ;
        RECT 1600.500 168.970 1600.640 260.030 ;
        RECT 1600.440 168.650 1600.700 168.970 ;
        RECT 1904.500 168.650 1904.760 168.970 ;
        RECT 1904.560 16.730 1904.700 168.650 ;
        RECT 1904.560 16.590 1906.080 16.730 ;
        RECT 1905.940 2.400 1906.080 16.590 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
=======
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1617.430 244.020 1617.750 244.080 ;
        RECT 1621.110 244.020 1621.430 244.080 ;
        RECT 1617.430 243.880 1621.430 244.020 ;
        RECT 1617.430 243.820 1617.750 243.880 ;
        RECT 1621.110 243.820 1621.430 243.880 ;
        RECT 1621.110 176.700 1621.430 176.760 ;
        RECT 1918.270 176.700 1918.590 176.760 ;
        RECT 1621.110 176.560 1918.590 176.700 ;
        RECT 1621.110 176.500 1621.430 176.560 ;
        RECT 1918.270 176.500 1918.590 176.560 ;
        RECT 1918.270 2.960 1918.590 3.020 ;
        RECT 1923.330 2.960 1923.650 3.020 ;
        RECT 1918.270 2.820 1923.650 2.960 ;
        RECT 1918.270 2.760 1918.590 2.820 ;
        RECT 1923.330 2.760 1923.650 2.820 ;
      LAYER via ;
        RECT 1617.460 243.820 1617.720 244.080 ;
        RECT 1621.140 243.820 1621.400 244.080 ;
        RECT 1621.140 176.500 1621.400 176.760 ;
        RECT 1918.300 176.500 1918.560 176.760 ;
        RECT 1918.300 2.760 1918.560 3.020 ;
        RECT 1923.360 2.760 1923.620 3.020 ;
      LAYER met2 ;
        RECT 1617.410 260.000 1617.690 264.000 ;
        RECT 1617.520 244.110 1617.660 260.000 ;
        RECT 1617.460 243.790 1617.720 244.110 ;
        RECT 1621.140 243.790 1621.400 244.110 ;
        RECT 1621.200 176.790 1621.340 243.790 ;
        RECT 1621.140 176.470 1621.400 176.790 ;
        RECT 1918.300 176.470 1918.560 176.790 ;
        RECT 1918.360 3.050 1918.500 176.470 ;
        RECT 1918.300 2.730 1918.560 3.050 ;
        RECT 1923.360 2.730 1923.620 3.050 ;
        RECT 1923.420 2.400 1923.560 2.730 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
=======
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1635.370 244.020 1635.690 244.080 ;
        RECT 1641.350 244.020 1641.670 244.080 ;
        RECT 1635.370 243.880 1641.670 244.020 ;
        RECT 1635.370 243.820 1635.690 243.880 ;
        RECT 1641.350 243.820 1641.670 243.880 ;
        RECT 1641.350 183.160 1641.670 183.220 ;
        RECT 1938.970 183.160 1939.290 183.220 ;
        RECT 1641.350 183.020 1939.290 183.160 ;
        RECT 1641.350 182.960 1641.670 183.020 ;
        RECT 1938.970 182.960 1939.290 183.020 ;
        RECT 1938.970 2.960 1939.290 3.020 ;
        RECT 1941.270 2.960 1941.590 3.020 ;
        RECT 1938.970 2.820 1941.590 2.960 ;
        RECT 1938.970 2.760 1939.290 2.820 ;
        RECT 1941.270 2.760 1941.590 2.820 ;
      LAYER via ;
        RECT 1635.400 243.820 1635.660 244.080 ;
        RECT 1641.380 243.820 1641.640 244.080 ;
        RECT 1641.380 182.960 1641.640 183.220 ;
        RECT 1939.000 182.960 1939.260 183.220 ;
        RECT 1939.000 2.760 1939.260 3.020 ;
        RECT 1941.300 2.760 1941.560 3.020 ;
      LAYER met2 ;
        RECT 1635.350 260.000 1635.630 264.000 ;
        RECT 1635.460 244.110 1635.600 260.000 ;
        RECT 1635.400 243.790 1635.660 244.110 ;
        RECT 1641.380 243.790 1641.640 244.110 ;
        RECT 1641.440 183.250 1641.580 243.790 ;
        RECT 1641.380 182.930 1641.640 183.250 ;
        RECT 1939.000 182.930 1939.260 183.250 ;
        RECT 1939.060 3.050 1939.200 182.930 ;
        RECT 1939.000 2.730 1939.260 3.050 ;
        RECT 1941.300 2.730 1941.560 3.050 ;
        RECT 1941.360 2.400 1941.500 2.730 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
=======
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1655.610 197.440 1655.930 197.500 ;
        RECT 1952.770 197.440 1953.090 197.500 ;
        RECT 1655.610 197.300 1953.090 197.440 ;
        RECT 1655.610 197.240 1655.930 197.300 ;
        RECT 1952.770 197.240 1953.090 197.300 ;
        RECT 1952.770 37.980 1953.090 38.040 ;
        RECT 1959.210 37.980 1959.530 38.040 ;
        RECT 1952.770 37.840 1959.530 37.980 ;
        RECT 1952.770 37.780 1953.090 37.840 ;
        RECT 1959.210 37.780 1959.530 37.840 ;
      LAYER via ;
        RECT 1655.640 197.240 1655.900 197.500 ;
        RECT 1952.800 197.240 1953.060 197.500 ;
        RECT 1952.800 37.780 1953.060 38.040 ;
        RECT 1959.240 37.780 1959.500 38.040 ;
      LAYER met2 ;
        RECT 1653.290 260.170 1653.570 264.000 ;
        RECT 1653.290 260.030 1655.840 260.170 ;
        RECT 1653.290 260.000 1653.570 260.030 ;
        RECT 1655.700 197.530 1655.840 260.030 ;
        RECT 1655.640 197.210 1655.900 197.530 ;
        RECT 1952.800 197.210 1953.060 197.530 ;
        RECT 1952.860 38.070 1953.000 197.210 ;
        RECT 1952.800 37.750 1953.060 38.070 ;
        RECT 1959.240 37.750 1959.500 38.070 ;
        RECT 1959.300 2.400 1959.440 37.750 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
=======
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 1973.545 48.365 1973.715 96.475 ;
      LAYER mcon ;
        RECT 1973.545 96.305 1973.715 96.475 ;
      LAYER met1 ;
        RECT 1671.250 244.020 1671.570 244.080 ;
        RECT 1676.310 244.020 1676.630 244.080 ;
        RECT 1671.250 243.880 1676.630 244.020 ;
        RECT 1671.250 243.820 1671.570 243.880 ;
        RECT 1676.310 243.820 1676.630 243.880 ;
        RECT 1676.310 114.140 1676.630 114.200 ;
        RECT 1973.930 114.140 1974.250 114.200 ;
        RECT 1676.310 114.000 1974.250 114.140 ;
        RECT 1676.310 113.940 1676.630 114.000 ;
        RECT 1973.930 113.940 1974.250 114.000 ;
        RECT 1973.470 96.460 1973.790 96.520 ;
        RECT 1973.275 96.320 1973.790 96.460 ;
        RECT 1973.470 96.260 1973.790 96.320 ;
        RECT 1973.485 48.520 1973.775 48.565 ;
        RECT 1977.150 48.520 1977.470 48.580 ;
        RECT 1973.485 48.380 1977.470 48.520 ;
        RECT 1973.485 48.335 1973.775 48.380 ;
        RECT 1977.150 48.320 1977.470 48.380 ;
      LAYER via ;
        RECT 1671.280 243.820 1671.540 244.080 ;
        RECT 1676.340 243.820 1676.600 244.080 ;
        RECT 1676.340 113.940 1676.600 114.200 ;
        RECT 1973.960 113.940 1974.220 114.200 ;
        RECT 1973.500 96.260 1973.760 96.520 ;
        RECT 1977.180 48.320 1977.440 48.580 ;
      LAYER met2 ;
        RECT 1671.230 260.000 1671.510 264.000 ;
        RECT 1671.340 244.110 1671.480 260.000 ;
        RECT 1671.280 243.790 1671.540 244.110 ;
        RECT 1676.340 243.790 1676.600 244.110 ;
        RECT 1676.400 114.230 1676.540 243.790 ;
        RECT 1676.340 113.910 1676.600 114.230 ;
        RECT 1973.960 113.910 1974.220 114.230 ;
        RECT 1974.020 96.970 1974.160 113.910 ;
        RECT 1973.560 96.830 1974.160 96.970 ;
        RECT 1973.560 96.550 1973.700 96.830 ;
        RECT 1973.500 96.230 1973.760 96.550 ;
        RECT 1977.180 48.290 1977.440 48.610 ;
        RECT 1977.240 2.400 1977.380 48.290 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
=======
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1690.110 224.640 1690.430 224.700 ;
        RECT 1994.170 224.640 1994.490 224.700 ;
        RECT 1690.110 224.500 1994.490 224.640 ;
        RECT 1690.110 224.440 1690.430 224.500 ;
        RECT 1994.170 224.440 1994.490 224.500 ;
      LAYER via ;
        RECT 1690.140 224.440 1690.400 224.700 ;
        RECT 1994.200 224.440 1994.460 224.700 ;
      LAYER met2 ;
        RECT 1689.170 260.170 1689.450 264.000 ;
        RECT 1689.170 260.030 1690.340 260.170 ;
        RECT 1689.170 260.000 1689.450 260.030 ;
        RECT 1690.200 224.730 1690.340 260.030 ;
        RECT 1690.140 224.410 1690.400 224.730 ;
        RECT 1994.200 224.410 1994.460 224.730 ;
        RECT 1994.260 16.730 1994.400 224.410 ;
        RECT 1994.260 16.590 1995.320 16.730 ;
        RECT 1995.180 2.400 1995.320 16.590 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
=======
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1710.810 189.620 1711.130 189.680 ;
        RECT 2007.970 189.620 2008.290 189.680 ;
        RECT 1710.810 189.480 2008.290 189.620 ;
        RECT 1710.810 189.420 1711.130 189.480 ;
        RECT 2007.970 189.420 2008.290 189.480 ;
      LAYER via ;
        RECT 1710.840 189.420 1711.100 189.680 ;
        RECT 2008.000 189.420 2008.260 189.680 ;
      LAYER met2 ;
        RECT 1707.110 260.170 1707.390 264.000 ;
        RECT 1707.110 260.030 1711.040 260.170 ;
        RECT 1707.110 260.000 1707.390 260.030 ;
        RECT 1710.900 189.710 1711.040 260.030 ;
        RECT 1710.840 189.390 1711.100 189.710 ;
        RECT 2008.000 189.390 2008.260 189.710 ;
        RECT 2008.060 16.730 2008.200 189.390 ;
        RECT 2008.060 16.590 2012.800 16.730 ;
        RECT 2012.660 2.400 2012.800 16.590 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
=======
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1724.610 30.840 1724.930 30.900 ;
        RECT 2030.510 30.840 2030.830 30.900 ;
        RECT 1724.610 30.700 2030.830 30.840 ;
        RECT 1724.610 30.640 1724.930 30.700 ;
        RECT 2030.510 30.640 2030.830 30.700 ;
      LAYER via ;
        RECT 1724.640 30.640 1724.900 30.900 ;
        RECT 2030.540 30.640 2030.800 30.900 ;
      LAYER met2 ;
        RECT 1724.590 260.000 1724.870 264.000 ;
        RECT 1724.700 30.930 1724.840 260.000 ;
        RECT 1724.640 30.610 1724.900 30.930 ;
        RECT 2030.540 30.610 2030.800 30.930 ;
        RECT 2030.600 2.400 2030.740 30.610 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
=======
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1745.310 148.140 1745.630 148.200 ;
        RECT 2042.930 148.140 2043.250 148.200 ;
        RECT 1745.310 148.000 2043.250 148.140 ;
        RECT 1745.310 147.940 1745.630 148.000 ;
        RECT 2042.930 147.940 2043.250 148.000 ;
        RECT 2042.930 62.120 2043.250 62.180 ;
        RECT 2048.450 62.120 2048.770 62.180 ;
        RECT 2042.930 61.980 2048.770 62.120 ;
        RECT 2042.930 61.920 2043.250 61.980 ;
        RECT 2048.450 61.920 2048.770 61.980 ;
      LAYER via ;
        RECT 1745.340 147.940 1745.600 148.200 ;
        RECT 2042.960 147.940 2043.220 148.200 ;
        RECT 2042.960 61.920 2043.220 62.180 ;
        RECT 2048.480 61.920 2048.740 62.180 ;
      LAYER met2 ;
        RECT 1742.530 260.170 1742.810 264.000 ;
        RECT 1742.530 260.030 1745.540 260.170 ;
        RECT 1742.530 260.000 1742.810 260.030 ;
        RECT 1745.400 148.230 1745.540 260.030 ;
        RECT 1745.340 147.910 1745.600 148.230 ;
        RECT 2042.960 147.910 2043.220 148.230 ;
        RECT 2043.020 62.210 2043.160 147.910 ;
        RECT 2042.960 61.890 2043.220 62.210 ;
        RECT 2048.480 61.890 2048.740 62.210 ;
        RECT 2048.540 2.400 2048.680 61.890 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
=======
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 455.470 244.020 455.790 244.080 ;
        RECT 461.450 244.020 461.770 244.080 ;
        RECT 455.470 243.880 461.770 244.020 ;
        RECT 455.470 243.820 455.790 243.880 ;
        RECT 461.450 243.820 461.770 243.880 ;
        RECT 461.450 19.960 461.770 20.020 ;
        RECT 763.670 19.960 763.990 20.020 ;
        RECT 461.450 19.820 763.990 19.960 ;
        RECT 461.450 19.760 461.770 19.820 ;
        RECT 763.670 19.760 763.990 19.820 ;
      LAYER via ;
        RECT 455.500 243.820 455.760 244.080 ;
        RECT 461.480 243.820 461.740 244.080 ;
        RECT 461.480 19.760 461.740 20.020 ;
        RECT 763.700 19.760 763.960 20.020 ;
      LAYER met2 ;
        RECT 455.450 260.000 455.730 264.000 ;
        RECT 455.560 244.110 455.700 260.000 ;
        RECT 455.500 243.790 455.760 244.110 ;
        RECT 461.480 243.790 461.740 244.110 ;
        RECT 461.540 20.050 461.680 243.790 ;
        RECT 461.480 19.730 461.740 20.050 ;
        RECT 763.700 19.730 763.960 20.050 ;
        RECT 763.760 2.400 763.900 19.730 ;
        RECT 763.550 -4.800 764.110 2.400 ;
=======
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1760.490 244.020 1760.810 244.080 ;
        RECT 1766.010 244.020 1766.330 244.080 ;
        RECT 1760.490 243.880 1766.330 244.020 ;
        RECT 1760.490 243.820 1760.810 243.880 ;
        RECT 1766.010 243.820 1766.330 243.880 ;
        RECT 1766.010 141.680 1766.330 141.740 ;
        RECT 2063.170 141.680 2063.490 141.740 ;
        RECT 1766.010 141.540 2063.490 141.680 ;
        RECT 1766.010 141.480 1766.330 141.540 ;
        RECT 2063.170 141.480 2063.490 141.540 ;
        RECT 2063.170 62.120 2063.490 62.180 ;
        RECT 2066.390 62.120 2066.710 62.180 ;
        RECT 2063.170 61.980 2066.710 62.120 ;
        RECT 2063.170 61.920 2063.490 61.980 ;
        RECT 2066.390 61.920 2066.710 61.980 ;
      LAYER via ;
        RECT 1760.520 243.820 1760.780 244.080 ;
        RECT 1766.040 243.820 1766.300 244.080 ;
        RECT 1766.040 141.480 1766.300 141.740 ;
        RECT 2063.200 141.480 2063.460 141.740 ;
        RECT 2063.200 61.920 2063.460 62.180 ;
        RECT 2066.420 61.920 2066.680 62.180 ;
      LAYER met2 ;
        RECT 1760.470 260.000 1760.750 264.000 ;
        RECT 1760.580 244.110 1760.720 260.000 ;
        RECT 1760.520 243.790 1760.780 244.110 ;
        RECT 1766.040 243.790 1766.300 244.110 ;
        RECT 1766.100 141.770 1766.240 243.790 ;
        RECT 1766.040 141.450 1766.300 141.770 ;
        RECT 2063.200 141.450 2063.460 141.770 ;
        RECT 2063.260 62.210 2063.400 141.450 ;
        RECT 2063.200 61.890 2063.460 62.210 ;
        RECT 2066.420 61.890 2066.680 62.210 ;
        RECT 2066.480 2.400 2066.620 61.890 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
=======
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1779.810 203.560 1780.130 203.620 ;
        RECT 2084.330 203.560 2084.650 203.620 ;
        RECT 1779.810 203.420 2084.650 203.560 ;
        RECT 1779.810 203.360 1780.130 203.420 ;
        RECT 2084.330 203.360 2084.650 203.420 ;
      LAYER via ;
        RECT 1779.840 203.360 1780.100 203.620 ;
        RECT 2084.360 203.360 2084.620 203.620 ;
      LAYER met2 ;
        RECT 1778.410 260.170 1778.690 264.000 ;
        RECT 1778.410 260.030 1780.040 260.170 ;
        RECT 1778.410 260.000 1778.690 260.030 ;
        RECT 1779.900 203.650 1780.040 260.030 ;
        RECT 1779.840 203.330 1780.100 203.650 ;
        RECT 2084.360 203.330 2084.620 203.650 ;
        RECT 2084.420 2.400 2084.560 203.330 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
=======
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1796.370 244.020 1796.690 244.080 ;
        RECT 1800.510 244.020 1800.830 244.080 ;
        RECT 1796.370 243.880 1800.830 244.020 ;
        RECT 1796.370 243.820 1796.690 243.880 ;
        RECT 1800.510 243.820 1800.830 243.880 ;
        RECT 1800.510 120.940 1800.830 121.000 ;
        RECT 2097.670 120.940 2097.990 121.000 ;
        RECT 1800.510 120.800 2097.990 120.940 ;
        RECT 1800.510 120.740 1800.830 120.800 ;
        RECT 2097.670 120.740 2097.990 120.800 ;
      LAYER via ;
        RECT 1796.400 243.820 1796.660 244.080 ;
        RECT 1800.540 243.820 1800.800 244.080 ;
        RECT 1800.540 120.740 1800.800 121.000 ;
        RECT 2097.700 120.740 2097.960 121.000 ;
      LAYER met2 ;
        RECT 1796.350 260.000 1796.630 264.000 ;
        RECT 1796.460 244.110 1796.600 260.000 ;
        RECT 1796.400 243.790 1796.660 244.110 ;
        RECT 1800.540 243.790 1800.800 244.110 ;
        RECT 1800.600 121.030 1800.740 243.790 ;
        RECT 1800.540 120.710 1800.800 121.030 ;
        RECT 2097.700 120.710 2097.960 121.030 ;
        RECT 2097.760 16.730 2097.900 120.710 ;
        RECT 2097.760 16.590 2102.040 16.730 ;
        RECT 2101.900 2.400 2102.040 16.590 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
=======
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1813.850 155.280 1814.170 155.340 ;
        RECT 2118.370 155.280 2118.690 155.340 ;
        RECT 1813.850 155.140 2118.690 155.280 ;
        RECT 1813.850 155.080 1814.170 155.140 ;
        RECT 2118.370 155.080 2118.690 155.140 ;
      LAYER via ;
        RECT 1813.880 155.080 1814.140 155.340 ;
        RECT 2118.400 155.080 2118.660 155.340 ;
      LAYER met2 ;
        RECT 1814.290 260.170 1814.570 264.000 ;
        RECT 1813.940 260.030 1814.570 260.170 ;
        RECT 1813.940 155.370 1814.080 260.030 ;
        RECT 1814.290 260.000 1814.570 260.030 ;
        RECT 1813.880 155.050 1814.140 155.370 ;
        RECT 2118.400 155.050 2118.660 155.370 ;
        RECT 2118.460 16.730 2118.600 155.050 ;
        RECT 2118.460 16.590 2119.980 16.730 ;
        RECT 2119.840 2.400 2119.980 16.590 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
=======
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1835.010 162.080 1835.330 162.140 ;
        RECT 2132.170 162.080 2132.490 162.140 ;
        RECT 1835.010 161.940 2132.490 162.080 ;
        RECT 1835.010 161.880 1835.330 161.940 ;
        RECT 2132.170 161.880 2132.490 161.940 ;
      LAYER via ;
        RECT 1835.040 161.880 1835.300 162.140 ;
        RECT 2132.200 161.880 2132.460 162.140 ;
      LAYER met2 ;
        RECT 1832.230 260.170 1832.510 264.000 ;
        RECT 1832.230 260.030 1835.240 260.170 ;
        RECT 1832.230 260.000 1832.510 260.030 ;
        RECT 1835.100 162.170 1835.240 260.030 ;
        RECT 1835.040 161.850 1835.300 162.170 ;
        RECT 2132.200 161.850 2132.460 162.170 ;
        RECT 2132.260 16.730 2132.400 161.850 ;
        RECT 2132.260 16.590 2137.920 16.730 ;
        RECT 2137.780 2.400 2137.920 16.590 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
=======
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 2155.705 2.805 2155.875 48.195 ;
      LAYER mcon ;
        RECT 2155.705 48.025 2155.875 48.195 ;
      LAYER met1 ;
        RECT 1849.730 244.020 1850.050 244.080 ;
        RECT 1859.390 244.020 1859.710 244.080 ;
        RECT 1849.730 243.880 1859.710 244.020 ;
        RECT 1849.730 243.820 1850.050 243.880 ;
        RECT 1859.390 243.820 1859.710 243.880 ;
        RECT 1859.390 169.220 1859.710 169.280 ;
        RECT 2152.870 169.220 2153.190 169.280 ;
        RECT 1859.390 169.080 2153.190 169.220 ;
        RECT 1859.390 169.020 1859.710 169.080 ;
        RECT 2152.870 169.020 2153.190 169.080 ;
        RECT 2152.870 48.180 2153.190 48.240 ;
        RECT 2155.645 48.180 2155.935 48.225 ;
        RECT 2152.870 48.040 2155.935 48.180 ;
        RECT 2152.870 47.980 2153.190 48.040 ;
        RECT 2155.645 47.995 2155.935 48.040 ;
        RECT 2155.630 2.960 2155.950 3.020 ;
        RECT 2155.435 2.820 2155.950 2.960 ;
        RECT 2155.630 2.760 2155.950 2.820 ;
      LAYER via ;
        RECT 1849.760 243.820 1850.020 244.080 ;
        RECT 1859.420 243.820 1859.680 244.080 ;
        RECT 1859.420 169.020 1859.680 169.280 ;
        RECT 2152.900 169.020 2153.160 169.280 ;
        RECT 2152.900 47.980 2153.160 48.240 ;
        RECT 2155.660 2.760 2155.920 3.020 ;
      LAYER met2 ;
        RECT 1849.710 260.000 1849.990 264.000 ;
        RECT 1849.820 244.110 1849.960 260.000 ;
        RECT 1849.760 243.790 1850.020 244.110 ;
        RECT 1859.420 243.790 1859.680 244.110 ;
        RECT 1859.480 169.310 1859.620 243.790 ;
        RECT 1859.420 168.990 1859.680 169.310 ;
        RECT 2152.900 168.990 2153.160 169.310 ;
        RECT 2152.960 48.270 2153.100 168.990 ;
        RECT 2152.900 47.950 2153.160 48.270 ;
        RECT 2155.660 2.730 2155.920 3.050 ;
        RECT 2155.720 2.400 2155.860 2.730 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
=======
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1869.510 176.360 1869.830 176.420 ;
        RECT 2166.670 176.360 2166.990 176.420 ;
        RECT 1869.510 176.220 2166.990 176.360 ;
        RECT 1869.510 176.160 1869.830 176.220 ;
        RECT 2166.670 176.160 2166.990 176.220 ;
        RECT 2166.670 38.320 2166.990 38.380 ;
        RECT 2173.110 38.320 2173.430 38.380 ;
        RECT 2166.670 38.180 2173.430 38.320 ;
        RECT 2166.670 38.120 2166.990 38.180 ;
        RECT 2173.110 38.120 2173.430 38.180 ;
      LAYER via ;
        RECT 1869.540 176.160 1869.800 176.420 ;
        RECT 2166.700 176.160 2166.960 176.420 ;
        RECT 2166.700 38.120 2166.960 38.380 ;
        RECT 2173.140 38.120 2173.400 38.380 ;
      LAYER met2 ;
        RECT 1867.650 260.170 1867.930 264.000 ;
        RECT 1867.650 260.030 1869.740 260.170 ;
        RECT 1867.650 260.000 1867.930 260.030 ;
        RECT 1869.600 176.450 1869.740 260.030 ;
        RECT 1869.540 176.130 1869.800 176.450 ;
        RECT 2166.700 176.130 2166.960 176.450 ;
        RECT 2166.760 38.410 2166.900 176.130 ;
        RECT 2166.700 38.090 2166.960 38.410 ;
        RECT 2173.140 38.090 2173.400 38.410 ;
        RECT 2173.200 2.400 2173.340 38.090 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
=======
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1885.610 244.020 1885.930 244.080 ;
        RECT 1890.210 244.020 1890.530 244.080 ;
        RECT 1885.610 243.880 1890.530 244.020 ;
        RECT 1885.610 243.820 1885.930 243.880 ;
        RECT 1890.210 243.820 1890.530 243.880 ;
        RECT 1890.210 182.820 1890.530 182.880 ;
        RECT 2187.370 182.820 2187.690 182.880 ;
        RECT 1890.210 182.680 2187.690 182.820 ;
        RECT 1890.210 182.620 1890.530 182.680 ;
        RECT 2187.370 182.620 2187.690 182.680 ;
      LAYER via ;
        RECT 1885.640 243.820 1885.900 244.080 ;
        RECT 1890.240 243.820 1890.500 244.080 ;
        RECT 1890.240 182.620 1890.500 182.880 ;
        RECT 2187.400 182.620 2187.660 182.880 ;
      LAYER met2 ;
        RECT 1885.590 260.000 1885.870 264.000 ;
        RECT 1885.700 244.110 1885.840 260.000 ;
        RECT 1885.640 243.790 1885.900 244.110 ;
        RECT 1890.240 243.790 1890.500 244.110 ;
        RECT 1890.300 182.910 1890.440 243.790 ;
        RECT 1890.240 182.590 1890.500 182.910 ;
        RECT 2187.400 182.590 2187.660 182.910 ;
        RECT 2187.460 16.730 2187.600 182.590 ;
        RECT 2187.460 16.590 2191.280 16.730 ;
        RECT 2191.140 2.400 2191.280 16.590 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
=======
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1903.550 196.760 1903.870 196.820 ;
        RECT 2208.070 196.760 2208.390 196.820 ;
        RECT 1903.550 196.620 2208.390 196.760 ;
        RECT 1903.550 196.560 1903.870 196.620 ;
        RECT 2208.070 196.560 2208.390 196.620 ;
      LAYER via ;
        RECT 1903.580 196.560 1903.840 196.820 ;
        RECT 2208.100 196.560 2208.360 196.820 ;
      LAYER met2 ;
        RECT 1903.530 260.000 1903.810 264.000 ;
        RECT 1903.640 196.850 1903.780 260.000 ;
        RECT 1903.580 196.530 1903.840 196.850 ;
        RECT 2208.100 196.530 2208.360 196.850 ;
        RECT 2208.160 16.730 2208.300 196.530 ;
        RECT 2208.160 16.590 2209.220 16.730 ;
        RECT 2209.080 2.400 2209.220 16.590 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
=======
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1924.710 224.300 1925.030 224.360 ;
        RECT 2221.870 224.300 2222.190 224.360 ;
        RECT 1924.710 224.160 2222.190 224.300 ;
        RECT 1924.710 224.100 1925.030 224.160 ;
        RECT 2221.870 224.100 2222.190 224.160 ;
      LAYER via ;
        RECT 1924.740 224.100 1925.000 224.360 ;
        RECT 2221.900 224.100 2222.160 224.360 ;
      LAYER met2 ;
        RECT 1921.470 260.170 1921.750 264.000 ;
        RECT 1921.470 260.030 1924.940 260.170 ;
        RECT 1921.470 260.000 1921.750 260.030 ;
        RECT 1924.800 224.390 1924.940 260.030 ;
        RECT 1924.740 224.070 1925.000 224.390 ;
        RECT 2221.900 224.070 2222.160 224.390 ;
        RECT 2221.960 16.730 2222.100 224.070 ;
        RECT 2221.960 16.590 2227.160 16.730 ;
        RECT 2227.020 2.400 2227.160 16.590 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
=======
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 475.710 17.240 476.030 17.300 ;
        RECT 781.610 17.240 781.930 17.300 ;
        RECT 475.710 17.100 781.930 17.240 ;
        RECT 475.710 17.040 476.030 17.100 ;
        RECT 781.610 17.040 781.930 17.100 ;
      LAYER via ;
        RECT 475.740 17.040 476.000 17.300 ;
        RECT 781.640 17.040 781.900 17.300 ;
      LAYER met2 ;
        RECT 473.390 260.170 473.670 264.000 ;
        RECT 473.390 260.030 475.940 260.170 ;
        RECT 473.390 260.000 473.670 260.030 ;
        RECT 475.800 17.330 475.940 260.030 ;
        RECT 475.740 17.010 476.000 17.330 ;
        RECT 781.640 17.010 781.900 17.330 ;
        RECT 781.700 2.400 781.840 17.010 ;
        RECT 781.490 -4.800 782.050 2.400 ;
=======
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1939.430 243.340 1939.750 243.400 ;
        RECT 1945.410 243.340 1945.730 243.400 ;
        RECT 1939.430 243.200 1945.730 243.340 ;
        RECT 1939.430 243.140 1939.750 243.200 ;
        RECT 1945.410 243.140 1945.730 243.200 ;
        RECT 1945.410 189.960 1945.730 190.020 ;
        RECT 2242.570 189.960 2242.890 190.020 ;
        RECT 1945.410 189.820 2242.890 189.960 ;
        RECT 1945.410 189.760 1945.730 189.820 ;
        RECT 2242.570 189.760 2242.890 189.820 ;
      LAYER via ;
        RECT 1939.460 243.140 1939.720 243.400 ;
        RECT 1945.440 243.140 1945.700 243.400 ;
        RECT 1945.440 189.760 1945.700 190.020 ;
        RECT 2242.600 189.760 2242.860 190.020 ;
      LAYER met2 ;
        RECT 1939.410 260.000 1939.690 264.000 ;
        RECT 1939.520 243.430 1939.660 260.000 ;
        RECT 1939.460 243.110 1939.720 243.430 ;
        RECT 1945.440 243.110 1945.700 243.430 ;
        RECT 1945.500 190.050 1945.640 243.110 ;
        RECT 1945.440 189.730 1945.700 190.050 ;
        RECT 2242.600 189.730 2242.860 190.050 ;
        RECT 2242.660 16.730 2242.800 189.730 ;
        RECT 2242.660 16.590 2245.100 16.730 ;
        RECT 2244.960 2.400 2245.100 16.590 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
=======
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1959.210 134.880 1959.530 134.940 ;
        RECT 2256.370 134.880 2256.690 134.940 ;
        RECT 1959.210 134.740 2256.690 134.880 ;
        RECT 1959.210 134.680 1959.530 134.740 ;
        RECT 2256.370 134.680 2256.690 134.740 ;
        RECT 2256.370 18.260 2256.690 18.320 ;
        RECT 2262.350 18.260 2262.670 18.320 ;
        RECT 2256.370 18.120 2262.670 18.260 ;
        RECT 2256.370 18.060 2256.690 18.120 ;
        RECT 2262.350 18.060 2262.670 18.120 ;
      LAYER via ;
        RECT 1959.240 134.680 1959.500 134.940 ;
        RECT 2256.400 134.680 2256.660 134.940 ;
        RECT 2256.400 18.060 2256.660 18.320 ;
        RECT 2262.380 18.060 2262.640 18.320 ;
      LAYER met2 ;
        RECT 1957.350 260.170 1957.630 264.000 ;
        RECT 1957.350 260.030 1959.440 260.170 ;
        RECT 1957.350 260.000 1957.630 260.030 ;
        RECT 1959.300 134.970 1959.440 260.030 ;
        RECT 1959.240 134.650 1959.500 134.970 ;
        RECT 2256.400 134.650 2256.660 134.970 ;
        RECT 2256.460 18.350 2256.600 134.650 ;
        RECT 2256.400 18.030 2256.660 18.350 ;
        RECT 2262.380 18.030 2262.640 18.350 ;
        RECT 2262.440 2.400 2262.580 18.030 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
=======
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1974.850 244.020 1975.170 244.080 ;
        RECT 1979.910 244.020 1980.230 244.080 ;
        RECT 1974.850 243.880 1980.230 244.020 ;
        RECT 1974.850 243.820 1975.170 243.880 ;
        RECT 1979.910 243.820 1980.230 243.880 ;
        RECT 1979.910 128.080 1980.230 128.140 ;
        RECT 2277.070 128.080 2277.390 128.140 ;
        RECT 1979.910 127.940 2277.390 128.080 ;
        RECT 1979.910 127.880 1980.230 127.940 ;
        RECT 2277.070 127.880 2277.390 127.940 ;
        RECT 2277.070 2.960 2277.390 3.020 ;
        RECT 2280.290 2.960 2280.610 3.020 ;
        RECT 2277.070 2.820 2280.610 2.960 ;
        RECT 2277.070 2.760 2277.390 2.820 ;
        RECT 2280.290 2.760 2280.610 2.820 ;
      LAYER via ;
        RECT 1974.880 243.820 1975.140 244.080 ;
        RECT 1979.940 243.820 1980.200 244.080 ;
        RECT 1979.940 127.880 1980.200 128.140 ;
        RECT 2277.100 127.880 2277.360 128.140 ;
        RECT 2277.100 2.760 2277.360 3.020 ;
        RECT 2280.320 2.760 2280.580 3.020 ;
      LAYER met2 ;
        RECT 1974.830 260.000 1975.110 264.000 ;
        RECT 1974.940 244.110 1975.080 260.000 ;
        RECT 1974.880 243.790 1975.140 244.110 ;
        RECT 1979.940 243.790 1980.200 244.110 ;
        RECT 1980.000 128.170 1980.140 243.790 ;
        RECT 1979.940 127.850 1980.200 128.170 ;
        RECT 2277.100 127.850 2277.360 128.170 ;
        RECT 2277.160 3.050 2277.300 127.850 ;
        RECT 2277.100 2.730 2277.360 3.050 ;
        RECT 2280.320 2.730 2280.580 3.050 ;
        RECT 2280.380 2.400 2280.520 2.730 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
=======
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1993.710 141.340 1994.030 141.400 ;
        RECT 2298.230 141.340 2298.550 141.400 ;
        RECT 1993.710 141.200 2298.550 141.340 ;
        RECT 1993.710 141.140 1994.030 141.200 ;
        RECT 2298.230 141.140 2298.550 141.200 ;
      LAYER via ;
        RECT 1993.740 141.140 1994.000 141.400 ;
        RECT 2298.260 141.140 2298.520 141.400 ;
      LAYER met2 ;
        RECT 1992.770 260.170 1993.050 264.000 ;
        RECT 1992.770 260.030 1993.940 260.170 ;
        RECT 1992.770 260.000 1993.050 260.030 ;
        RECT 1993.800 141.430 1993.940 260.030 ;
        RECT 1993.740 141.110 1994.000 141.430 ;
        RECT 2298.260 141.110 2298.520 141.430 ;
        RECT 2298.320 2.400 2298.460 141.110 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
=======
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2014.410 148.480 2014.730 148.540 ;
        RECT 2311.570 148.480 2311.890 148.540 ;
        RECT 2014.410 148.340 2311.890 148.480 ;
        RECT 2014.410 148.280 2014.730 148.340 ;
        RECT 2311.570 148.280 2311.890 148.340 ;
      LAYER via ;
        RECT 2014.440 148.280 2014.700 148.540 ;
        RECT 2311.600 148.280 2311.860 148.540 ;
      LAYER met2 ;
        RECT 2010.710 260.170 2010.990 264.000 ;
        RECT 2010.710 260.030 2014.640 260.170 ;
        RECT 2010.710 260.000 2010.990 260.030 ;
        RECT 2014.500 148.570 2014.640 260.030 ;
        RECT 2014.440 148.250 2014.700 148.570 ;
        RECT 2311.600 148.250 2311.860 148.570 ;
        RECT 2311.660 16.730 2311.800 148.250 ;
        RECT 2311.660 16.590 2316.400 16.730 ;
        RECT 2316.260 2.400 2316.400 16.590 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
=======
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2028.670 244.020 2028.990 244.080 ;
        RECT 2034.650 244.020 2034.970 244.080 ;
        RECT 2028.670 243.880 2034.970 244.020 ;
        RECT 2028.670 243.820 2028.990 243.880 ;
        RECT 2034.650 243.820 2034.970 243.880 ;
        RECT 2034.650 176.020 2034.970 176.080 ;
        RECT 2332.270 176.020 2332.590 176.080 ;
        RECT 2034.650 175.880 2332.590 176.020 ;
        RECT 2034.650 175.820 2034.970 175.880 ;
        RECT 2332.270 175.820 2332.590 175.880 ;
      LAYER via ;
        RECT 2028.700 243.820 2028.960 244.080 ;
        RECT 2034.680 243.820 2034.940 244.080 ;
        RECT 2034.680 175.820 2034.940 176.080 ;
        RECT 2332.300 175.820 2332.560 176.080 ;
      LAYER met2 ;
        RECT 2028.650 260.000 2028.930 264.000 ;
        RECT 2028.760 244.110 2028.900 260.000 ;
        RECT 2028.700 243.790 2028.960 244.110 ;
        RECT 2034.680 243.790 2034.940 244.110 ;
        RECT 2034.740 176.110 2034.880 243.790 ;
        RECT 2034.680 175.790 2034.940 176.110 ;
        RECT 2332.300 175.790 2332.560 176.110 ;
        RECT 2332.360 16.730 2332.500 175.790 ;
        RECT 2332.360 16.590 2334.340 16.730 ;
        RECT 2334.200 2.400 2334.340 16.590 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
=======
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2048.910 183.160 2049.230 183.220 ;
        RECT 2346.070 183.160 2346.390 183.220 ;
        RECT 2048.910 183.020 2346.390 183.160 ;
        RECT 2048.910 182.960 2049.230 183.020 ;
        RECT 2346.070 182.960 2346.390 183.020 ;
      LAYER via ;
        RECT 2048.940 182.960 2049.200 183.220 ;
        RECT 2346.100 182.960 2346.360 183.220 ;
      LAYER met2 ;
        RECT 2046.590 260.170 2046.870 264.000 ;
        RECT 2046.590 260.030 2049.140 260.170 ;
        RECT 2046.590 260.000 2046.870 260.030 ;
        RECT 2049.000 183.250 2049.140 260.030 ;
        RECT 2048.940 182.930 2049.200 183.250 ;
        RECT 2346.100 182.930 2346.360 183.250 ;
        RECT 2346.160 16.730 2346.300 182.930 ;
        RECT 2346.160 16.590 2351.820 16.730 ;
        RECT 2351.680 2.400 2351.820 16.590 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
=======
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2064.550 244.020 2064.870 244.080 ;
        RECT 2069.610 244.020 2069.930 244.080 ;
        RECT 2064.550 243.880 2069.930 244.020 ;
        RECT 2064.550 243.820 2064.870 243.880 ;
        RECT 2069.610 243.820 2069.930 243.880 ;
        RECT 2069.610 162.420 2069.930 162.480 ;
        RECT 2366.770 162.420 2367.090 162.480 ;
        RECT 2069.610 162.280 2367.090 162.420 ;
        RECT 2069.610 162.220 2069.930 162.280 ;
        RECT 2366.770 162.220 2367.090 162.280 ;
        RECT 2366.770 2.960 2367.090 3.020 ;
        RECT 2369.530 2.960 2369.850 3.020 ;
        RECT 2366.770 2.820 2369.850 2.960 ;
        RECT 2366.770 2.760 2367.090 2.820 ;
        RECT 2369.530 2.760 2369.850 2.820 ;
      LAYER via ;
        RECT 2064.580 243.820 2064.840 244.080 ;
        RECT 2069.640 243.820 2069.900 244.080 ;
        RECT 2069.640 162.220 2069.900 162.480 ;
        RECT 2366.800 162.220 2367.060 162.480 ;
        RECT 2366.800 2.760 2367.060 3.020 ;
        RECT 2369.560 2.760 2369.820 3.020 ;
      LAYER met2 ;
        RECT 2064.530 260.000 2064.810 264.000 ;
        RECT 2064.640 244.110 2064.780 260.000 ;
        RECT 2064.580 243.790 2064.840 244.110 ;
        RECT 2069.640 243.790 2069.900 244.110 ;
        RECT 2069.700 162.510 2069.840 243.790 ;
        RECT 2069.640 162.190 2069.900 162.510 ;
        RECT 2366.800 162.190 2367.060 162.510 ;
        RECT 2366.860 3.050 2367.000 162.190 ;
        RECT 2366.800 2.730 2367.060 3.050 ;
        RECT 2369.560 2.730 2369.820 3.050 ;
        RECT 2369.620 2.400 2369.760 2.730 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
=======
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2083.410 51.580 2083.730 51.640 ;
        RECT 2387.930 51.580 2388.250 51.640 ;
        RECT 2083.410 51.440 2388.250 51.580 ;
        RECT 2083.410 51.380 2083.730 51.440 ;
        RECT 2387.930 51.380 2388.250 51.440 ;
      LAYER via ;
        RECT 2083.440 51.380 2083.700 51.640 ;
        RECT 2387.960 51.380 2388.220 51.640 ;
      LAYER met2 ;
        RECT 2082.470 260.170 2082.750 264.000 ;
        RECT 2082.470 260.030 2083.640 260.170 ;
        RECT 2082.470 260.000 2082.750 260.030 ;
        RECT 2083.500 51.670 2083.640 260.030 ;
        RECT 2083.440 51.350 2083.700 51.670 ;
        RECT 2387.960 51.350 2388.220 51.670 ;
        RECT 2388.020 3.130 2388.160 51.350 ;
        RECT 2387.560 2.990 2388.160 3.130 ;
        RECT 2387.560 2.400 2387.700 2.990 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
=======
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2100.430 244.020 2100.750 244.080 ;
        RECT 2104.110 244.020 2104.430 244.080 ;
        RECT 2100.430 243.880 2104.430 244.020 ;
        RECT 2100.430 243.820 2100.750 243.880 ;
        RECT 2104.110 243.820 2104.430 243.880 ;
        RECT 2104.110 197.100 2104.430 197.160 ;
        RECT 2401.270 197.100 2401.590 197.160 ;
        RECT 2104.110 196.960 2401.590 197.100 ;
        RECT 2104.110 196.900 2104.430 196.960 ;
        RECT 2401.270 196.900 2401.590 196.960 ;
      LAYER via ;
        RECT 2100.460 243.820 2100.720 244.080 ;
        RECT 2104.140 243.820 2104.400 244.080 ;
        RECT 2104.140 196.900 2104.400 197.160 ;
        RECT 2401.300 196.900 2401.560 197.160 ;
      LAYER met2 ;
        RECT 2100.410 260.000 2100.690 264.000 ;
        RECT 2100.520 244.110 2100.660 260.000 ;
        RECT 2100.460 243.790 2100.720 244.110 ;
        RECT 2104.140 243.790 2104.400 244.110 ;
        RECT 2104.200 197.190 2104.340 243.790 ;
        RECT 2104.140 196.870 2104.400 197.190 ;
        RECT 2401.300 196.870 2401.560 197.190 ;
        RECT 2401.360 17.410 2401.500 196.870 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
=======
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 491.350 244.020 491.670 244.080 ;
        RECT 496.410 244.020 496.730 244.080 ;
        RECT 491.350 243.880 496.730 244.020 ;
        RECT 491.350 243.820 491.670 243.880 ;
        RECT 496.410 243.820 496.730 243.880 ;
        RECT 496.410 15.540 496.730 15.600 ;
        RECT 799.550 15.540 799.870 15.600 ;
        RECT 496.410 15.400 799.870 15.540 ;
        RECT 496.410 15.340 496.730 15.400 ;
        RECT 799.550 15.340 799.870 15.400 ;
      LAYER via ;
        RECT 491.380 243.820 491.640 244.080 ;
        RECT 496.440 243.820 496.700 244.080 ;
        RECT 496.440 15.340 496.700 15.600 ;
        RECT 799.580 15.340 799.840 15.600 ;
      LAYER met2 ;
        RECT 491.330 260.000 491.610 264.000 ;
        RECT 491.440 244.110 491.580 260.000 ;
        RECT 491.380 243.790 491.640 244.110 ;
        RECT 496.440 243.790 496.700 244.110 ;
        RECT 496.500 15.630 496.640 243.790 ;
        RECT 496.440 15.310 496.700 15.630 ;
        RECT 799.580 15.310 799.840 15.630 ;
        RECT 799.640 2.400 799.780 15.310 ;
        RECT 799.430 -4.800 799.990 2.400 ;
=======
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 336.330 245.380 336.650 245.440 ;
        RECT 642.230 245.380 642.550 245.440 ;
        RECT 336.330 245.240 642.550 245.380 ;
        RECT 336.330 245.180 336.650 245.240 ;
        RECT 642.230 245.180 642.550 245.240 ;
      LAYER via ;
        RECT 336.360 245.180 336.620 245.440 ;
        RECT 642.260 245.180 642.520 245.440 ;
      LAYER met2 ;
        RECT 336.310 260.000 336.590 264.000 ;
        RECT 336.420 245.470 336.560 260.000 ;
        RECT 336.360 245.150 336.620 245.470 ;
        RECT 642.260 245.150 642.520 245.470 ;
        RECT 642.320 17.410 642.460 245.150 ;
        RECT 642.320 17.270 645.220 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
=======
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2124.810 189.620 2125.130 189.680 ;
        RECT 2428.870 189.620 2429.190 189.680 ;
        RECT 2124.810 189.480 2429.190 189.620 ;
        RECT 2124.810 189.420 2125.130 189.480 ;
        RECT 2428.870 189.420 2429.190 189.480 ;
      LAYER via ;
        RECT 2124.840 189.420 2125.100 189.680 ;
        RECT 2428.900 189.420 2429.160 189.680 ;
      LAYER met2 ;
        RECT 2123.870 260.170 2124.150 264.000 ;
        RECT 2123.870 260.030 2125.040 260.170 ;
        RECT 2123.870 260.000 2124.150 260.030 ;
        RECT 2124.900 189.710 2125.040 260.030 ;
        RECT 2124.840 189.390 2125.100 189.710 ;
        RECT 2428.900 189.390 2429.160 189.710 ;
        RECT 2428.960 2.400 2429.100 189.390 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
=======
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2141.830 244.020 2142.150 244.080 ;
        RECT 2145.510 244.020 2145.830 244.080 ;
        RECT 2141.830 243.880 2145.830 244.020 ;
        RECT 2141.830 243.820 2142.150 243.880 ;
        RECT 2145.510 243.820 2145.830 243.880 ;
        RECT 2145.510 17.580 2145.830 17.640 ;
        RECT 2446.810 17.580 2447.130 17.640 ;
        RECT 2145.510 17.440 2447.130 17.580 ;
        RECT 2145.510 17.380 2145.830 17.440 ;
        RECT 2446.810 17.380 2447.130 17.440 ;
      LAYER via ;
        RECT 2141.860 243.820 2142.120 244.080 ;
        RECT 2145.540 243.820 2145.800 244.080 ;
        RECT 2145.540 17.380 2145.800 17.640 ;
        RECT 2446.840 17.380 2447.100 17.640 ;
      LAYER met2 ;
        RECT 2141.810 260.000 2142.090 264.000 ;
        RECT 2141.920 244.110 2142.060 260.000 ;
        RECT 2141.860 243.790 2142.120 244.110 ;
        RECT 2145.540 243.790 2145.800 244.110 ;
        RECT 2145.600 17.670 2145.740 243.790 ;
        RECT 2145.540 17.350 2145.800 17.670 ;
        RECT 2446.840 17.350 2447.100 17.670 ;
        RECT 2446.900 2.400 2447.040 17.350 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
=======
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2159.770 244.020 2160.090 244.080 ;
        RECT 2165.750 244.020 2166.070 244.080 ;
        RECT 2159.770 243.880 2166.070 244.020 ;
        RECT 2159.770 243.820 2160.090 243.880 ;
        RECT 2165.750 243.820 2166.070 243.880 ;
        RECT 2165.750 15.540 2166.070 15.600 ;
        RECT 2464.750 15.540 2465.070 15.600 ;
        RECT 2165.750 15.400 2465.070 15.540 ;
        RECT 2165.750 15.340 2166.070 15.400 ;
        RECT 2464.750 15.340 2465.070 15.400 ;
      LAYER via ;
        RECT 2159.800 243.820 2160.060 244.080 ;
        RECT 2165.780 243.820 2166.040 244.080 ;
        RECT 2165.780 15.340 2166.040 15.600 ;
        RECT 2464.780 15.340 2465.040 15.600 ;
      LAYER met2 ;
        RECT 2159.750 260.000 2160.030 264.000 ;
        RECT 2159.860 244.110 2160.000 260.000 ;
        RECT 2159.800 243.790 2160.060 244.110 ;
        RECT 2165.780 243.790 2166.040 244.110 ;
        RECT 2165.840 15.630 2165.980 243.790 ;
        RECT 2165.780 15.310 2166.040 15.630 ;
        RECT 2464.780 15.310 2465.040 15.630 ;
        RECT 2464.840 2.400 2464.980 15.310 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
=======
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2180.010 16.900 2180.330 16.960 ;
        RECT 2482.690 16.900 2483.010 16.960 ;
        RECT 2180.010 16.760 2483.010 16.900 ;
        RECT 2180.010 16.700 2180.330 16.760 ;
        RECT 2482.690 16.700 2483.010 16.760 ;
      LAYER via ;
        RECT 2180.040 16.700 2180.300 16.960 ;
        RECT 2482.720 16.700 2482.980 16.960 ;
      LAYER met2 ;
        RECT 2177.690 260.170 2177.970 264.000 ;
        RECT 2177.690 260.030 2180.240 260.170 ;
        RECT 2177.690 260.000 2177.970 260.030 ;
        RECT 2180.100 16.990 2180.240 260.030 ;
        RECT 2180.040 16.670 2180.300 16.990 ;
        RECT 2482.720 16.670 2482.980 16.990 ;
        RECT 2482.780 2.400 2482.920 16.670 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
=======
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2195.650 244.020 2195.970 244.080 ;
        RECT 2200.710 244.020 2201.030 244.080 ;
        RECT 2195.650 243.880 2201.030 244.020 ;
        RECT 2195.650 243.820 2195.970 243.880 ;
        RECT 2200.710 243.820 2201.030 243.880 ;
        RECT 2200.710 17.240 2201.030 17.300 ;
        RECT 2500.630 17.240 2500.950 17.300 ;
        RECT 2200.710 17.100 2500.950 17.240 ;
        RECT 2200.710 17.040 2201.030 17.100 ;
        RECT 2500.630 17.040 2500.950 17.100 ;
      LAYER via ;
        RECT 2195.680 243.820 2195.940 244.080 ;
        RECT 2200.740 243.820 2201.000 244.080 ;
        RECT 2200.740 17.040 2201.000 17.300 ;
        RECT 2500.660 17.040 2500.920 17.300 ;
      LAYER met2 ;
        RECT 2195.630 260.000 2195.910 264.000 ;
        RECT 2195.740 244.110 2195.880 260.000 ;
        RECT 2195.680 243.790 2195.940 244.110 ;
        RECT 2200.740 243.790 2201.000 244.110 ;
        RECT 2200.800 17.330 2200.940 243.790 ;
        RECT 2200.740 17.010 2201.000 17.330 ;
        RECT 2500.660 17.010 2500.920 17.330 ;
        RECT 2500.720 2.400 2500.860 17.010 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
=======
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2214.510 15.880 2214.830 15.940 ;
        RECT 2518.110 15.880 2518.430 15.940 ;
        RECT 2214.510 15.740 2518.430 15.880 ;
        RECT 2214.510 15.680 2214.830 15.740 ;
        RECT 2518.110 15.680 2518.430 15.740 ;
      LAYER via ;
        RECT 2214.540 15.680 2214.800 15.940 ;
        RECT 2518.140 15.680 2518.400 15.940 ;
      LAYER met2 ;
        RECT 2213.570 260.170 2213.850 264.000 ;
        RECT 2213.570 260.030 2214.740 260.170 ;
        RECT 2213.570 260.000 2213.850 260.030 ;
        RECT 2214.600 15.970 2214.740 260.030 ;
        RECT 2214.540 15.650 2214.800 15.970 ;
        RECT 2518.140 15.650 2518.400 15.970 ;
        RECT 2518.200 2.400 2518.340 15.650 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
=======
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2231.070 244.020 2231.390 244.080 ;
        RECT 2235.210 244.020 2235.530 244.080 ;
        RECT 2231.070 243.880 2235.530 244.020 ;
        RECT 2231.070 243.820 2231.390 243.880 ;
        RECT 2235.210 243.820 2235.530 243.880 ;
        RECT 2235.210 20.640 2235.530 20.700 ;
        RECT 2536.050 20.640 2536.370 20.700 ;
        RECT 2235.210 20.500 2536.370 20.640 ;
        RECT 2235.210 20.440 2235.530 20.500 ;
        RECT 2536.050 20.440 2536.370 20.500 ;
      LAYER via ;
        RECT 2231.100 243.820 2231.360 244.080 ;
        RECT 2235.240 243.820 2235.500 244.080 ;
        RECT 2235.240 20.440 2235.500 20.700 ;
        RECT 2536.080 20.440 2536.340 20.700 ;
      LAYER met2 ;
        RECT 2231.050 260.000 2231.330 264.000 ;
        RECT 2231.160 244.110 2231.300 260.000 ;
        RECT 2231.100 243.790 2231.360 244.110 ;
        RECT 2235.240 243.790 2235.500 244.110 ;
        RECT 2235.300 20.730 2235.440 243.790 ;
        RECT 2235.240 20.410 2235.500 20.730 ;
        RECT 2536.080 20.410 2536.340 20.730 ;
        RECT 2536.140 2.400 2536.280 20.410 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
=======
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2248.990 260.000 2249.270 264.000 ;
        RECT 2249.100 17.525 2249.240 260.000 ;
        RECT 2249.030 17.155 2249.310 17.525 ;
        RECT 2554.010 17.155 2554.290 17.525 ;
        RECT 2554.080 2.400 2554.220 17.155 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
      LAYER via2 ;
        RECT 2249.030 17.200 2249.310 17.480 ;
        RECT 2554.010 17.200 2554.290 17.480 ;
      LAYER met3 ;
        RECT 2249.005 17.490 2249.335 17.505 ;
        RECT 2553.985 17.490 2554.315 17.505 ;
        RECT 2249.005 17.190 2554.315 17.490 ;
        RECT 2249.005 17.175 2249.335 17.190 ;
        RECT 2553.985 17.175 2554.315 17.190 ;
=======
        RECT 2553.870 -4.800 2554.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2269.710 16.560 2270.030 16.620 ;
        RECT 2571.930 16.560 2572.250 16.620 ;
        RECT 2269.710 16.420 2572.250 16.560 ;
        RECT 2269.710 16.360 2270.030 16.420 ;
        RECT 2571.930 16.360 2572.250 16.420 ;
      LAYER via ;
        RECT 2269.740 16.360 2270.000 16.620 ;
        RECT 2571.960 16.360 2572.220 16.620 ;
      LAYER met2 ;
        RECT 2266.930 260.170 2267.210 264.000 ;
        RECT 2266.930 260.030 2269.940 260.170 ;
        RECT 2266.930 260.000 2267.210 260.030 ;
        RECT 2269.800 16.650 2269.940 260.030 ;
        RECT 2269.740 16.330 2270.000 16.650 ;
        RECT 2571.960 16.330 2572.220 16.650 ;
        RECT 2572.020 2.400 2572.160 16.330 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
=======
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2284.890 244.020 2285.210 244.080 ;
        RECT 2290.410 244.020 2290.730 244.080 ;
        RECT 2284.890 243.880 2290.730 244.020 ;
        RECT 2284.890 243.820 2285.210 243.880 ;
        RECT 2290.410 243.820 2290.730 243.880 ;
        RECT 2290.410 16.220 2290.730 16.280 ;
        RECT 2589.410 16.220 2589.730 16.280 ;
        RECT 2290.410 16.080 2589.730 16.220 ;
        RECT 2290.410 16.020 2290.730 16.080 ;
        RECT 2589.410 16.020 2589.730 16.080 ;
      LAYER via ;
        RECT 2284.920 243.820 2285.180 244.080 ;
        RECT 2290.440 243.820 2290.700 244.080 ;
        RECT 2290.440 16.020 2290.700 16.280 ;
        RECT 2589.440 16.020 2589.700 16.280 ;
      LAYER met2 ;
        RECT 2284.870 260.000 2285.150 264.000 ;
        RECT 2284.980 244.110 2285.120 260.000 ;
        RECT 2284.920 243.790 2285.180 244.110 ;
        RECT 2290.440 243.790 2290.700 244.110 ;
        RECT 2290.500 16.310 2290.640 243.790 ;
        RECT 2290.440 15.990 2290.700 16.310 ;
        RECT 2589.440 15.990 2589.700 16.310 ;
        RECT 2589.500 2.400 2589.640 15.990 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
=======
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 515.270 246.400 515.590 246.460 ;
        RECT 821.630 246.400 821.950 246.460 ;
        RECT 515.270 246.260 821.950 246.400 ;
        RECT 515.270 246.200 515.590 246.260 ;
        RECT 821.630 246.200 821.950 246.260 ;
      LAYER via ;
        RECT 515.300 246.200 515.560 246.460 ;
        RECT 821.660 246.200 821.920 246.460 ;
      LAYER met2 ;
        RECT 515.250 260.000 515.530 264.000 ;
        RECT 515.360 246.490 515.500 260.000 ;
        RECT 515.300 246.170 515.560 246.490 ;
        RECT 821.660 246.170 821.920 246.490 ;
        RECT 821.720 17.410 821.860 246.170 ;
        RECT 821.720 17.270 823.700 17.410 ;
        RECT 823.560 2.400 823.700 17.270 ;
        RECT 823.350 -4.800 823.910 2.400 ;
=======
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2304.210 19.960 2304.530 20.020 ;
        RECT 2607.350 19.960 2607.670 20.020 ;
        RECT 2304.210 19.820 2607.670 19.960 ;
        RECT 2304.210 19.760 2304.530 19.820 ;
        RECT 2607.350 19.760 2607.670 19.820 ;
      LAYER via ;
        RECT 2304.240 19.760 2304.500 20.020 ;
        RECT 2607.380 19.760 2607.640 20.020 ;
      LAYER met2 ;
        RECT 2302.810 260.170 2303.090 264.000 ;
        RECT 2302.810 260.030 2304.440 260.170 ;
        RECT 2302.810 260.000 2303.090 260.030 ;
        RECT 2304.300 20.050 2304.440 260.030 ;
        RECT 2304.240 19.730 2304.500 20.050 ;
        RECT 2607.380 19.730 2607.640 20.050 ;
        RECT 2607.440 2.400 2607.580 19.730 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
=======
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2320.770 244.020 2321.090 244.080 ;
        RECT 2324.910 244.020 2325.230 244.080 ;
        RECT 2320.770 243.880 2325.230 244.020 ;
        RECT 2320.770 243.820 2321.090 243.880 ;
        RECT 2324.910 243.820 2325.230 243.880 ;
        RECT 2324.910 19.620 2325.230 19.680 ;
        RECT 2625.290 19.620 2625.610 19.680 ;
        RECT 2324.910 19.480 2625.610 19.620 ;
        RECT 2324.910 19.420 2325.230 19.480 ;
        RECT 2625.290 19.420 2625.610 19.480 ;
      LAYER via ;
        RECT 2320.800 243.820 2321.060 244.080 ;
        RECT 2324.940 243.820 2325.200 244.080 ;
        RECT 2324.940 19.420 2325.200 19.680 ;
        RECT 2625.320 19.420 2625.580 19.680 ;
      LAYER met2 ;
        RECT 2320.750 260.000 2321.030 264.000 ;
        RECT 2320.860 244.110 2321.000 260.000 ;
        RECT 2320.800 243.790 2321.060 244.110 ;
        RECT 2324.940 243.790 2325.200 244.110 ;
        RECT 2325.000 19.710 2325.140 243.790 ;
        RECT 2324.940 19.390 2325.200 19.710 ;
        RECT 2625.320 19.390 2625.580 19.710 ;
        RECT 2625.380 2.400 2625.520 19.390 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
=======
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2338.710 245.040 2339.030 245.100 ;
        RECT 2642.770 245.040 2643.090 245.100 ;
        RECT 2338.710 244.900 2643.090 245.040 ;
        RECT 2338.710 244.840 2339.030 244.900 ;
        RECT 2642.770 244.840 2643.090 244.900 ;
      LAYER via ;
        RECT 2338.740 244.840 2339.000 245.100 ;
        RECT 2642.800 244.840 2643.060 245.100 ;
      LAYER met2 ;
        RECT 2338.690 260.000 2338.970 264.000 ;
        RECT 2338.800 245.130 2338.940 260.000 ;
        RECT 2338.740 244.810 2339.000 245.130 ;
        RECT 2642.800 244.810 2643.060 245.130 ;
        RECT 2642.860 17.410 2643.000 244.810 ;
        RECT 2642.860 17.270 2643.460 17.410 ;
        RECT 2643.320 2.400 2643.460 17.270 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
=======
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 2642.845 15.725 2643.015 18.955 ;
      LAYER mcon ;
        RECT 2642.845 18.785 2643.015 18.955 ;
      LAYER met1 ;
        RECT 2359.410 18.940 2359.730 19.000 ;
        RECT 2642.785 18.940 2643.075 18.985 ;
        RECT 2359.410 18.800 2643.075 18.940 ;
        RECT 2359.410 18.740 2359.730 18.800 ;
        RECT 2642.785 18.755 2643.075 18.800 ;
        RECT 2642.785 15.880 2643.075 15.925 ;
        RECT 2661.170 15.880 2661.490 15.940 ;
        RECT 2642.785 15.740 2661.490 15.880 ;
        RECT 2642.785 15.695 2643.075 15.740 ;
        RECT 2661.170 15.680 2661.490 15.740 ;
      LAYER via ;
        RECT 2359.440 18.740 2359.700 19.000 ;
        RECT 2661.200 15.680 2661.460 15.940 ;
      LAYER met2 ;
        RECT 2356.630 260.170 2356.910 264.000 ;
        RECT 2356.630 260.030 2359.640 260.170 ;
        RECT 2356.630 260.000 2356.910 260.030 ;
        RECT 2359.500 19.030 2359.640 260.030 ;
        RECT 2359.440 18.710 2359.700 19.030 ;
        RECT 2661.200 15.650 2661.460 15.970 ;
        RECT 2661.260 2.400 2661.400 15.650 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
=======
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2374.130 246.060 2374.450 246.120 ;
        RECT 2677.270 246.060 2677.590 246.120 ;
        RECT 2374.130 245.920 2677.590 246.060 ;
        RECT 2374.130 245.860 2374.450 245.920 ;
        RECT 2677.270 245.860 2677.590 245.920 ;
      LAYER via ;
        RECT 2374.160 245.860 2374.420 246.120 ;
        RECT 2677.300 245.860 2677.560 246.120 ;
      LAYER met2 ;
        RECT 2374.110 260.000 2374.390 264.000 ;
        RECT 2374.220 246.150 2374.360 260.000 ;
        RECT 2374.160 245.830 2374.420 246.150 ;
        RECT 2677.300 245.830 2677.560 246.150 ;
        RECT 2677.360 17.410 2677.500 245.830 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
=======
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2393.910 18.260 2394.230 18.320 ;
        RECT 2696.590 18.260 2696.910 18.320 ;
        RECT 2393.910 18.120 2696.910 18.260 ;
        RECT 2393.910 18.060 2394.230 18.120 ;
        RECT 2696.590 18.060 2696.910 18.120 ;
      LAYER via ;
        RECT 2393.940 18.060 2394.200 18.320 ;
        RECT 2696.620 18.060 2696.880 18.320 ;
      LAYER met2 ;
        RECT 2392.050 260.170 2392.330 264.000 ;
        RECT 2392.050 260.030 2394.140 260.170 ;
        RECT 2392.050 260.000 2392.330 260.030 ;
        RECT 2394.000 18.350 2394.140 260.030 ;
        RECT 2393.940 18.030 2394.200 18.350 ;
        RECT 2696.620 18.030 2696.880 18.350 ;
        RECT 2696.680 2.400 2696.820 18.030 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
=======
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2410.010 245.720 2410.330 245.780 ;
        RECT 2711.770 245.720 2712.090 245.780 ;
        RECT 2410.010 245.580 2712.090 245.720 ;
        RECT 2410.010 245.520 2410.330 245.580 ;
        RECT 2711.770 245.520 2712.090 245.580 ;
      LAYER via ;
        RECT 2410.040 245.520 2410.300 245.780 ;
        RECT 2711.800 245.520 2712.060 245.780 ;
      LAYER met2 ;
        RECT 2409.990 260.000 2410.270 264.000 ;
        RECT 2410.100 245.810 2410.240 260.000 ;
        RECT 2410.040 245.490 2410.300 245.810 ;
        RECT 2711.800 245.490 2712.060 245.810 ;
        RECT 2711.860 17.410 2712.000 245.490 ;
        RECT 2711.860 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
=======
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2427.930 260.170 2428.210 264.000 ;
        RECT 2427.930 260.030 2428.640 260.170 ;
        RECT 2427.930 260.000 2428.210 260.030 ;
        RECT 2428.500 18.205 2428.640 260.030 ;
        RECT 2428.430 17.835 2428.710 18.205 ;
        RECT 2732.490 17.835 2732.770 18.205 ;
        RECT 2732.560 2.400 2732.700 17.835 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 2428.430 17.880 2428.710 18.160 ;
        RECT 2732.490 17.880 2732.770 18.160 ;
      LAYER met3 ;
        RECT 2428.405 18.170 2428.735 18.185 ;
        RECT 2732.465 18.170 2732.795 18.185 ;
        RECT 2428.405 17.870 2732.795 18.170 ;
        RECT 2428.405 17.855 2428.735 17.870 ;
        RECT 2732.465 17.855 2732.795 17.870 ;
=======
        RECT 2732.350 -4.800 2732.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2445.890 245.380 2446.210 245.440 ;
        RECT 2746.270 245.380 2746.590 245.440 ;
        RECT 2445.890 245.240 2746.590 245.380 ;
        RECT 2445.890 245.180 2446.210 245.240 ;
        RECT 2746.270 245.180 2746.590 245.240 ;
      LAYER via ;
        RECT 2445.920 245.180 2446.180 245.440 ;
        RECT 2746.300 245.180 2746.560 245.440 ;
      LAYER met2 ;
        RECT 2445.870 260.000 2446.150 264.000 ;
        RECT 2445.980 245.470 2446.120 260.000 ;
        RECT 2445.920 245.150 2446.180 245.470 ;
        RECT 2746.300 245.150 2746.560 245.470 ;
        RECT 2746.360 17.410 2746.500 245.150 ;
        RECT 2746.360 17.270 2750.640 17.410 ;
        RECT 2750.500 2.400 2750.640 17.270 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
=======
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2463.830 244.020 2464.150 244.080 ;
        RECT 2469.810 244.020 2470.130 244.080 ;
        RECT 2463.830 243.880 2470.130 244.020 ;
        RECT 2463.830 243.820 2464.150 243.880 ;
        RECT 2469.810 243.820 2470.130 243.880 ;
        RECT 2469.810 17.580 2470.130 17.640 ;
        RECT 2767.890 17.580 2768.210 17.640 ;
        RECT 2469.810 17.440 2768.210 17.580 ;
        RECT 2469.810 17.380 2470.130 17.440 ;
        RECT 2767.890 17.380 2768.210 17.440 ;
      LAYER via ;
        RECT 2463.860 243.820 2464.120 244.080 ;
        RECT 2469.840 243.820 2470.100 244.080 ;
        RECT 2469.840 17.380 2470.100 17.640 ;
        RECT 2767.920 17.380 2768.180 17.640 ;
      LAYER met2 ;
        RECT 2463.810 260.000 2464.090 264.000 ;
        RECT 2463.920 244.110 2464.060 260.000 ;
        RECT 2463.860 243.790 2464.120 244.110 ;
        RECT 2469.840 243.790 2470.100 244.110 ;
        RECT 2469.900 17.670 2470.040 243.790 ;
        RECT 2469.840 17.350 2470.100 17.670 ;
        RECT 2767.920 17.350 2768.180 17.670 ;
        RECT 2767.980 2.400 2768.120 17.350 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
=======
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 533.210 244.020 533.530 244.080 ;
        RECT 537.810 244.020 538.130 244.080 ;
        RECT 533.210 243.880 538.130 244.020 ;
        RECT 533.210 243.820 533.530 243.880 ;
        RECT 537.810 243.820 538.130 243.880 ;
        RECT 537.810 16.220 538.130 16.280 ;
        RECT 840.950 16.220 841.270 16.280 ;
        RECT 537.810 16.080 841.270 16.220 ;
        RECT 537.810 16.020 538.130 16.080 ;
        RECT 840.950 16.020 841.270 16.080 ;
      LAYER via ;
        RECT 533.240 243.820 533.500 244.080 ;
        RECT 537.840 243.820 538.100 244.080 ;
        RECT 537.840 16.020 538.100 16.280 ;
        RECT 840.980 16.020 841.240 16.280 ;
      LAYER met2 ;
        RECT 533.190 260.000 533.470 264.000 ;
        RECT 533.300 244.110 533.440 260.000 ;
        RECT 533.240 243.790 533.500 244.110 ;
        RECT 537.840 243.790 538.100 244.110 ;
        RECT 537.900 16.310 538.040 243.790 ;
        RECT 537.840 15.990 538.100 16.310 ;
        RECT 840.980 15.990 841.240 16.310 ;
        RECT 841.040 2.400 841.180 15.990 ;
        RECT 840.830 -4.800 841.390 2.400 ;
=======
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2483.610 17.920 2483.930 17.980 ;
        RECT 2785.830 17.920 2786.150 17.980 ;
        RECT 2483.610 17.780 2786.150 17.920 ;
        RECT 2483.610 17.720 2483.930 17.780 ;
        RECT 2785.830 17.720 2786.150 17.780 ;
      LAYER via ;
        RECT 2483.640 17.720 2483.900 17.980 ;
        RECT 2785.860 17.720 2786.120 17.980 ;
      LAYER met2 ;
        RECT 2481.750 260.170 2482.030 264.000 ;
        RECT 2481.750 260.030 2483.840 260.170 ;
        RECT 2481.750 260.000 2482.030 260.030 ;
        RECT 2483.700 18.010 2483.840 260.030 ;
        RECT 2483.640 17.690 2483.900 18.010 ;
        RECT 2785.860 17.690 2786.120 18.010 ;
        RECT 2785.920 2.400 2786.060 17.690 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
=======
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2499.250 244.020 2499.570 244.080 ;
        RECT 2504.310 244.020 2504.630 244.080 ;
        RECT 2499.250 243.880 2504.630 244.020 ;
        RECT 2499.250 243.820 2499.570 243.880 ;
        RECT 2504.310 243.820 2504.630 243.880 ;
        RECT 2504.310 19.280 2504.630 19.340 ;
        RECT 2803.770 19.280 2804.090 19.340 ;
        RECT 2504.310 19.140 2804.090 19.280 ;
        RECT 2504.310 19.080 2504.630 19.140 ;
        RECT 2803.770 19.080 2804.090 19.140 ;
      LAYER via ;
        RECT 2499.280 243.820 2499.540 244.080 ;
        RECT 2504.340 243.820 2504.600 244.080 ;
        RECT 2504.340 19.080 2504.600 19.340 ;
        RECT 2803.800 19.080 2804.060 19.340 ;
      LAYER met2 ;
        RECT 2499.230 260.000 2499.510 264.000 ;
        RECT 2499.340 244.110 2499.480 260.000 ;
        RECT 2499.280 243.790 2499.540 244.110 ;
        RECT 2504.340 243.790 2504.600 244.110 ;
        RECT 2504.400 19.370 2504.540 243.790 ;
        RECT 2504.340 19.050 2504.600 19.370 ;
        RECT 2803.800 19.050 2804.060 19.370 ;
        RECT 2803.860 2.400 2804.000 19.050 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
=======
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2518.110 20.300 2518.430 20.360 ;
        RECT 2821.710 20.300 2822.030 20.360 ;
        RECT 2518.110 20.160 2822.030 20.300 ;
        RECT 2518.110 20.100 2518.430 20.160 ;
        RECT 2821.710 20.100 2822.030 20.160 ;
      LAYER via ;
        RECT 2518.140 20.100 2518.400 20.360 ;
        RECT 2821.740 20.100 2822.000 20.360 ;
      LAYER met2 ;
        RECT 2517.170 260.170 2517.450 264.000 ;
        RECT 2517.170 260.030 2518.340 260.170 ;
        RECT 2517.170 260.000 2517.450 260.030 ;
        RECT 2518.200 20.390 2518.340 260.030 ;
        RECT 2518.140 20.070 2518.400 20.390 ;
        RECT 2821.740 20.070 2822.000 20.390 ;
        RECT 2821.800 2.400 2821.940 20.070 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
=======
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2538.810 20.640 2539.130 20.700 ;
        RECT 2839.190 20.640 2839.510 20.700 ;
        RECT 2538.810 20.500 2839.510 20.640 ;
        RECT 2538.810 20.440 2539.130 20.500 ;
        RECT 2839.190 20.440 2839.510 20.500 ;
      LAYER via ;
        RECT 2538.840 20.440 2539.100 20.700 ;
        RECT 2839.220 20.440 2839.480 20.700 ;
      LAYER met2 ;
        RECT 2535.110 260.170 2535.390 264.000 ;
        RECT 2535.110 260.030 2539.040 260.170 ;
        RECT 2535.110 260.000 2535.390 260.030 ;
        RECT 2538.900 20.730 2539.040 260.030 ;
        RECT 2538.840 20.410 2539.100 20.730 ;
        RECT 2839.220 20.410 2839.480 20.730 ;
        RECT 2839.280 2.400 2839.420 20.410 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
=======
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2553.070 242.660 2553.390 242.720 ;
        RECT 2559.510 242.660 2559.830 242.720 ;
        RECT 2553.070 242.520 2559.830 242.660 ;
        RECT 2553.070 242.460 2553.390 242.520 ;
        RECT 2559.510 242.460 2559.830 242.520 ;
        RECT 2559.510 16.900 2559.830 16.960 ;
        RECT 2857.130 16.900 2857.450 16.960 ;
        RECT 2559.510 16.760 2857.450 16.900 ;
        RECT 2559.510 16.700 2559.830 16.760 ;
        RECT 2857.130 16.700 2857.450 16.760 ;
      LAYER via ;
        RECT 2553.100 242.460 2553.360 242.720 ;
        RECT 2559.540 242.460 2559.800 242.720 ;
        RECT 2559.540 16.700 2559.800 16.960 ;
        RECT 2857.160 16.700 2857.420 16.960 ;
      LAYER met2 ;
        RECT 2553.050 260.000 2553.330 264.000 ;
        RECT 2553.160 242.750 2553.300 260.000 ;
        RECT 2553.100 242.430 2553.360 242.750 ;
        RECT 2559.540 242.430 2559.800 242.750 ;
        RECT 2559.600 16.990 2559.740 242.430 ;
        RECT 2559.540 16.670 2559.800 16.990 ;
        RECT 2857.160 16.670 2857.420 16.990 ;
        RECT 2857.220 2.400 2857.360 16.670 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
=======
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2573.310 16.560 2573.630 16.620 ;
        RECT 2875.070 16.560 2875.390 16.620 ;
        RECT 2573.310 16.420 2875.390 16.560 ;
        RECT 2573.310 16.360 2573.630 16.420 ;
        RECT 2875.070 16.360 2875.390 16.420 ;
      LAYER via ;
        RECT 2573.340 16.360 2573.600 16.620 ;
        RECT 2875.100 16.360 2875.360 16.620 ;
      LAYER met2 ;
        RECT 2570.990 260.170 2571.270 264.000 ;
        RECT 2570.990 260.030 2573.540 260.170 ;
        RECT 2570.990 260.000 2571.270 260.030 ;
        RECT 2573.400 16.650 2573.540 260.030 ;
        RECT 2573.340 16.330 2573.600 16.650 ;
        RECT 2875.100 16.330 2875.360 16.650 ;
        RECT 2875.160 2.400 2875.300 16.330 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
=======
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2588.950 244.020 2589.270 244.080 ;
        RECT 2594.010 244.020 2594.330 244.080 ;
        RECT 2588.950 243.880 2594.330 244.020 ;
        RECT 2588.950 243.820 2589.270 243.880 ;
        RECT 2594.010 243.820 2594.330 243.880 ;
        RECT 2594.010 16.220 2594.330 16.280 ;
        RECT 2893.010 16.220 2893.330 16.280 ;
        RECT 2594.010 16.080 2893.330 16.220 ;
        RECT 2594.010 16.020 2594.330 16.080 ;
        RECT 2893.010 16.020 2893.330 16.080 ;
      LAYER via ;
        RECT 2588.980 243.820 2589.240 244.080 ;
        RECT 2594.040 243.820 2594.300 244.080 ;
        RECT 2594.040 16.020 2594.300 16.280 ;
        RECT 2893.040 16.020 2893.300 16.280 ;
      LAYER met2 ;
        RECT 2588.930 260.000 2589.210 264.000 ;
        RECT 2589.040 244.110 2589.180 260.000 ;
        RECT 2588.980 243.790 2589.240 244.110 ;
        RECT 2594.040 243.790 2594.300 244.110 ;
        RECT 2594.100 16.310 2594.240 243.790 ;
        RECT 2594.040 15.990 2594.300 16.310 ;
        RECT 2893.040 15.990 2893.300 16.310 ;
        RECT 2893.100 2.400 2893.240 15.990 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
=======
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2607.810 19.960 2608.130 20.020 ;
        RECT 2910.950 19.960 2911.270 20.020 ;
        RECT 2607.810 19.820 2911.270 19.960 ;
        RECT 2607.810 19.760 2608.130 19.820 ;
        RECT 2910.950 19.760 2911.270 19.820 ;
      LAYER via ;
        RECT 2607.840 19.760 2608.100 20.020 ;
        RECT 2910.980 19.760 2911.240 20.020 ;
      LAYER met2 ;
        RECT 2606.870 260.170 2607.150 264.000 ;
        RECT 2606.870 260.030 2608.040 260.170 ;
        RECT 2606.870 260.000 2607.150 260.030 ;
        RECT 2607.900 20.050 2608.040 260.030 ;
        RECT 2607.840 19.730 2608.100 20.050 ;
        RECT 2910.980 19.730 2911.240 20.050 ;
        RECT 2911.040 2.400 2911.180 19.730 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
=======
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 551.150 247.080 551.470 247.140 ;
        RECT 856.130 247.080 856.450 247.140 ;
        RECT 551.150 246.940 856.450 247.080 ;
        RECT 551.150 246.880 551.470 246.940 ;
        RECT 856.130 246.880 856.450 246.940 ;
      LAYER via ;
        RECT 551.180 246.880 551.440 247.140 ;
        RECT 856.160 246.880 856.420 247.140 ;
      LAYER met2 ;
        RECT 551.130 260.000 551.410 264.000 ;
        RECT 551.240 247.170 551.380 260.000 ;
        RECT 551.180 246.850 551.440 247.170 ;
        RECT 856.160 246.850 856.420 247.170 ;
        RECT 856.220 16.730 856.360 246.850 ;
        RECT 856.220 16.590 859.120 16.730 ;
        RECT 858.980 2.400 859.120 16.590 ;
        RECT 858.770 -4.800 859.330 2.400 ;
=======
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 568.630 244.020 568.950 244.080 ;
        RECT 572.310 244.020 572.630 244.080 ;
        RECT 568.630 243.880 572.630 244.020 ;
        RECT 568.630 243.820 568.950 243.880 ;
        RECT 572.310 243.820 572.630 243.880 ;
        RECT 572.310 18.600 572.630 18.660 ;
        RECT 876.370 18.600 876.690 18.660 ;
        RECT 572.310 18.460 876.690 18.600 ;
        RECT 572.310 18.400 572.630 18.460 ;
        RECT 876.370 18.400 876.690 18.460 ;
      LAYER via ;
        RECT 568.660 243.820 568.920 244.080 ;
        RECT 572.340 243.820 572.600 244.080 ;
        RECT 572.340 18.400 572.600 18.660 ;
        RECT 876.400 18.400 876.660 18.660 ;
      LAYER met2 ;
        RECT 568.610 260.000 568.890 264.000 ;
        RECT 568.720 244.110 568.860 260.000 ;
        RECT 568.660 243.790 568.920 244.110 ;
        RECT 572.340 243.790 572.600 244.110 ;
        RECT 572.400 18.690 572.540 243.790 ;
        RECT 572.340 18.370 572.600 18.690 ;
        RECT 876.400 18.370 876.660 18.690 ;
        RECT 876.460 16.050 876.600 18.370 ;
        RECT 876.460 15.910 877.060 16.050 ;
        RECT 876.920 2.400 877.060 15.910 ;
        RECT 876.710 -4.800 877.270 2.400 ;
=======
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 586.570 244.020 586.890 244.080 ;
        RECT 593.010 244.020 593.330 244.080 ;
        RECT 586.570 243.880 593.330 244.020 ;
        RECT 586.570 243.820 586.890 243.880 ;
        RECT 593.010 243.820 593.330 243.880 ;
        RECT 593.010 16.560 593.330 16.620 ;
        RECT 593.010 16.420 865.100 16.560 ;
        RECT 593.010 16.360 593.330 16.420 ;
        RECT 864.960 16.220 865.100 16.420 ;
        RECT 894.770 16.220 895.090 16.280 ;
        RECT 864.960 16.080 895.090 16.220 ;
        RECT 894.770 16.020 895.090 16.080 ;
      LAYER via ;
        RECT 586.600 243.820 586.860 244.080 ;
        RECT 593.040 243.820 593.300 244.080 ;
        RECT 593.040 16.360 593.300 16.620 ;
        RECT 894.800 16.020 895.060 16.280 ;
      LAYER met2 ;
        RECT 586.550 260.000 586.830 264.000 ;
        RECT 586.660 244.110 586.800 260.000 ;
        RECT 586.600 243.790 586.860 244.110 ;
        RECT 593.040 243.790 593.300 244.110 ;
        RECT 593.100 16.650 593.240 243.790 ;
        RECT 593.040 16.330 593.300 16.650 ;
        RECT 894.800 15.990 895.060 16.310 ;
        RECT 894.860 2.400 895.000 15.990 ;
        RECT 894.650 -4.800 895.210 2.400 ;
=======
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 606.810 18.260 607.130 18.320 ;
        RECT 912.710 18.260 913.030 18.320 ;
        RECT 606.810 18.120 913.030 18.260 ;
        RECT 606.810 18.060 607.130 18.120 ;
        RECT 912.710 18.060 913.030 18.120 ;
      LAYER via ;
        RECT 606.840 18.060 607.100 18.320 ;
        RECT 912.740 18.060 913.000 18.320 ;
      LAYER met2 ;
        RECT 604.490 260.170 604.770 264.000 ;
        RECT 604.490 260.030 607.040 260.170 ;
        RECT 604.490 260.000 604.770 260.030 ;
        RECT 606.900 18.350 607.040 260.030 ;
        RECT 606.840 18.030 607.100 18.350 ;
        RECT 912.740 18.030 913.000 18.350 ;
        RECT 912.800 2.400 912.940 18.030 ;
        RECT 912.590 -4.800 913.150 2.400 ;
=======
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 622.450 244.020 622.770 244.080 ;
        RECT 627.510 244.020 627.830 244.080 ;
        RECT 622.450 243.880 627.830 244.020 ;
        RECT 622.450 243.820 622.770 243.880 ;
        RECT 627.510 243.820 627.830 243.880 ;
        RECT 627.510 16.900 627.830 16.960 ;
        RECT 930.190 16.900 930.510 16.960 ;
        RECT 627.510 16.760 930.510 16.900 ;
        RECT 627.510 16.700 627.830 16.760 ;
        RECT 930.190 16.700 930.510 16.760 ;
      LAYER via ;
        RECT 622.480 243.820 622.740 244.080 ;
        RECT 627.540 243.820 627.800 244.080 ;
        RECT 627.540 16.700 627.800 16.960 ;
        RECT 930.220 16.700 930.480 16.960 ;
      LAYER met2 ;
        RECT 622.430 260.000 622.710 264.000 ;
        RECT 622.540 244.110 622.680 260.000 ;
        RECT 622.480 243.790 622.740 244.110 ;
        RECT 627.540 243.790 627.800 244.110 ;
        RECT 627.600 16.990 627.740 243.790 ;
        RECT 627.540 16.670 627.800 16.990 ;
        RECT 930.220 16.670 930.480 16.990 ;
        RECT 930.280 2.400 930.420 16.670 ;
        RECT 930.070 -4.800 930.630 2.400 ;
=======
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 948.130 18.260 948.450 18.320 ;
        RECT 917.400 18.120 948.450 18.260 ;
        RECT 641.310 17.920 641.630 17.980 ;
        RECT 917.400 17.920 917.540 18.120 ;
        RECT 948.130 18.060 948.450 18.120 ;
        RECT 641.310 17.780 917.540 17.920 ;
        RECT 641.310 17.720 641.630 17.780 ;
      LAYER via ;
        RECT 641.340 17.720 641.600 17.980 ;
        RECT 948.160 18.060 948.420 18.320 ;
      LAYER met2 ;
        RECT 640.370 260.170 640.650 264.000 ;
        RECT 640.370 260.030 641.540 260.170 ;
        RECT 640.370 260.000 640.650 260.030 ;
        RECT 641.400 18.010 641.540 260.030 ;
        RECT 948.160 18.030 948.420 18.350 ;
        RECT 641.340 17.690 641.600 18.010 ;
        RECT 948.220 2.400 948.360 18.030 ;
        RECT 948.010 -4.800 948.570 2.400 ;
=======
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 658.330 245.380 658.650 245.440 ;
        RECT 966.990 245.380 967.310 245.440 ;
        RECT 658.330 245.240 967.310 245.380 ;
        RECT 658.330 245.180 658.650 245.240 ;
        RECT 966.990 245.180 967.310 245.240 ;
      LAYER via ;
        RECT 658.360 245.180 658.620 245.440 ;
        RECT 967.020 245.180 967.280 245.440 ;
      LAYER met2 ;
        RECT 658.310 260.000 658.590 264.000 ;
        RECT 658.420 245.470 658.560 260.000 ;
        RECT 658.360 245.150 658.620 245.470 ;
        RECT 967.020 245.150 967.280 245.470 ;
        RECT 967.080 16.730 967.220 245.150 ;
        RECT 966.160 16.590 967.220 16.730 ;
        RECT 966.160 2.400 966.300 16.590 ;
        RECT 965.950 -4.800 966.510 2.400 ;
=======
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 676.270 242.660 676.590 242.720 ;
        RECT 682.250 242.660 682.570 242.720 ;
        RECT 676.270 242.520 682.570 242.660 ;
        RECT 676.270 242.460 676.590 242.520 ;
        RECT 682.250 242.460 682.570 242.520 ;
        RECT 682.250 19.620 682.570 19.680 ;
        RECT 984.010 19.620 984.330 19.680 ;
        RECT 682.250 19.480 984.330 19.620 ;
        RECT 682.250 19.420 682.570 19.480 ;
        RECT 984.010 19.420 984.330 19.480 ;
      LAYER via ;
        RECT 676.300 242.460 676.560 242.720 ;
        RECT 682.280 242.460 682.540 242.720 ;
        RECT 682.280 19.420 682.540 19.680 ;
        RECT 984.040 19.420 984.300 19.680 ;
      LAYER met2 ;
        RECT 676.250 260.000 676.530 264.000 ;
        RECT 676.360 242.750 676.500 260.000 ;
        RECT 676.300 242.430 676.560 242.750 ;
        RECT 682.280 242.430 682.540 242.750 ;
        RECT 682.340 19.710 682.480 242.430 ;
        RECT 682.280 19.390 682.540 19.710 ;
        RECT 984.040 19.390 984.300 19.710 ;
        RECT 984.100 2.400 984.240 19.390 ;
        RECT 983.890 -4.800 984.450 2.400 ;
=======
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 354.270 244.020 354.590 244.080 ;
        RECT 358.410 244.020 358.730 244.080 ;
        RECT 354.270 243.880 358.730 244.020 ;
        RECT 354.270 243.820 354.590 243.880 ;
        RECT 358.410 243.820 358.730 243.880 ;
        RECT 358.410 19.620 358.730 19.680 ;
        RECT 662.470 19.620 662.790 19.680 ;
        RECT 358.410 19.480 662.790 19.620 ;
        RECT 358.410 19.420 358.730 19.480 ;
        RECT 662.470 19.420 662.790 19.480 ;
      LAYER via ;
        RECT 354.300 243.820 354.560 244.080 ;
        RECT 358.440 243.820 358.700 244.080 ;
        RECT 358.440 19.420 358.700 19.680 ;
        RECT 662.500 19.420 662.760 19.680 ;
      LAYER met2 ;
        RECT 354.250 260.000 354.530 264.000 ;
        RECT 354.360 244.110 354.500 260.000 ;
        RECT 354.300 243.790 354.560 244.110 ;
        RECT 358.440 243.790 358.700 244.110 ;
        RECT 358.500 19.710 358.640 243.790 ;
        RECT 358.440 19.390 358.700 19.710 ;
        RECT 662.500 19.390 662.760 19.710 ;
        RECT 662.560 18.770 662.700 19.390 ;
        RECT 662.560 18.630 663.160 18.770 ;
        RECT 663.020 2.400 663.160 18.630 ;
        RECT 662.810 -4.800 663.370 2.400 ;
=======
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 694.210 245.720 694.530 245.780 ;
        RECT 1001.030 245.720 1001.350 245.780 ;
        RECT 694.210 245.580 1001.350 245.720 ;
        RECT 694.210 245.520 694.530 245.580 ;
        RECT 1001.030 245.520 1001.350 245.580 ;
      LAYER via ;
        RECT 694.240 245.520 694.500 245.780 ;
        RECT 1001.060 245.520 1001.320 245.780 ;
      LAYER met2 ;
        RECT 694.190 260.000 694.470 264.000 ;
        RECT 694.300 245.810 694.440 260.000 ;
        RECT 694.240 245.490 694.500 245.810 ;
        RECT 1001.060 245.490 1001.320 245.810 ;
        RECT 1001.120 16.730 1001.260 245.490 ;
        RECT 1001.120 16.590 1002.180 16.730 ;
        RECT 1002.040 2.400 1002.180 16.590 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
=======
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 711.690 244.020 712.010 244.080 ;
        RECT 717.210 244.020 717.530 244.080 ;
        RECT 711.690 243.880 717.530 244.020 ;
        RECT 711.690 243.820 712.010 243.880 ;
        RECT 717.210 243.820 717.530 243.880 ;
        RECT 717.210 20.640 717.530 20.700 ;
        RECT 1019.430 20.640 1019.750 20.700 ;
        RECT 717.210 20.500 1019.750 20.640 ;
        RECT 717.210 20.440 717.530 20.500 ;
        RECT 1019.430 20.440 1019.750 20.500 ;
      LAYER via ;
        RECT 711.720 243.820 711.980 244.080 ;
        RECT 717.240 243.820 717.500 244.080 ;
        RECT 717.240 20.440 717.500 20.700 ;
        RECT 1019.460 20.440 1019.720 20.700 ;
      LAYER met2 ;
        RECT 711.670 260.000 711.950 264.000 ;
        RECT 711.780 244.110 711.920 260.000 ;
        RECT 711.720 243.790 711.980 244.110 ;
        RECT 717.240 243.790 717.500 244.110 ;
        RECT 717.300 20.730 717.440 243.790 ;
        RECT 717.240 20.410 717.500 20.730 ;
        RECT 1019.460 20.410 1019.720 20.730 ;
        RECT 1019.520 2.400 1019.660 20.410 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
=======
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 729.630 246.060 729.950 246.120 ;
        RECT 1035.530 246.060 1035.850 246.120 ;
        RECT 729.630 245.920 1035.850 246.060 ;
        RECT 729.630 245.860 729.950 245.920 ;
        RECT 1035.530 245.860 1035.850 245.920 ;
      LAYER via ;
        RECT 729.660 245.860 729.920 246.120 ;
        RECT 1035.560 245.860 1035.820 246.120 ;
      LAYER met2 ;
        RECT 729.610 260.000 729.890 264.000 ;
        RECT 729.720 246.150 729.860 260.000 ;
        RECT 729.660 245.830 729.920 246.150 ;
        RECT 1035.560 245.830 1035.820 246.150 ;
        RECT 1035.620 16.730 1035.760 245.830 ;
        RECT 1035.620 16.590 1037.600 16.730 ;
        RECT 1037.460 2.400 1037.600 16.590 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
=======
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 747.570 244.020 747.890 244.080 ;
        RECT 751.710 244.020 752.030 244.080 ;
        RECT 747.570 243.880 752.030 244.020 ;
        RECT 747.570 243.820 747.890 243.880 ;
        RECT 751.710 243.820 752.030 243.880 ;
        RECT 751.710 20.300 752.030 20.360 ;
        RECT 1055.310 20.300 1055.630 20.360 ;
        RECT 751.710 20.160 1055.630 20.300 ;
        RECT 751.710 20.100 752.030 20.160 ;
        RECT 1055.310 20.100 1055.630 20.160 ;
      LAYER via ;
        RECT 747.600 243.820 747.860 244.080 ;
        RECT 751.740 243.820 752.000 244.080 ;
        RECT 751.740 20.100 752.000 20.360 ;
        RECT 1055.340 20.100 1055.600 20.360 ;
      LAYER met2 ;
        RECT 747.550 260.000 747.830 264.000 ;
        RECT 747.660 244.110 747.800 260.000 ;
        RECT 747.600 243.790 747.860 244.110 ;
        RECT 751.740 243.790 752.000 244.110 ;
        RECT 751.800 20.390 751.940 243.790 ;
        RECT 751.740 20.070 752.000 20.390 ;
        RECT 1055.340 20.070 1055.600 20.390 ;
        RECT 1055.400 2.400 1055.540 20.070 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
=======
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 765.510 18.940 765.830 19.000 ;
        RECT 1073.250 18.940 1073.570 19.000 ;
        RECT 765.510 18.800 1073.570 18.940 ;
        RECT 765.510 18.740 765.830 18.800 ;
        RECT 1073.250 18.740 1073.570 18.800 ;
      LAYER via ;
        RECT 765.540 18.740 765.800 19.000 ;
        RECT 1073.280 18.740 1073.540 19.000 ;
      LAYER met2 ;
        RECT 765.490 260.000 765.770 264.000 ;
        RECT 765.600 19.030 765.740 260.000 ;
        RECT 765.540 18.710 765.800 19.030 ;
        RECT 1073.280 18.710 1073.540 19.030 ;
        RECT 1073.340 2.400 1073.480 18.710 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
=======
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 786.210 19.280 786.530 19.340 ;
        RECT 1090.270 19.280 1090.590 19.340 ;
        RECT 786.210 19.140 1090.590 19.280 ;
        RECT 786.210 19.080 786.530 19.140 ;
        RECT 1090.270 19.080 1090.590 19.140 ;
      LAYER via ;
        RECT 786.240 19.080 786.500 19.340 ;
        RECT 1090.300 19.080 1090.560 19.340 ;
      LAYER met2 ;
        RECT 783.430 260.170 783.710 264.000 ;
        RECT 783.430 260.030 786.440 260.170 ;
        RECT 783.430 260.000 783.710 260.030 ;
        RECT 786.300 19.370 786.440 260.030 ;
        RECT 786.240 19.050 786.500 19.370 ;
        RECT 1090.300 19.050 1090.560 19.370 ;
        RECT 1090.360 17.410 1090.500 19.050 ;
        RECT 1090.360 17.270 1090.960 17.410 ;
        RECT 1090.820 2.400 1090.960 17.270 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
=======
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 801.390 244.020 801.710 244.080 ;
        RECT 806.910 244.020 807.230 244.080 ;
        RECT 801.390 243.880 807.230 244.020 ;
        RECT 801.390 243.820 801.710 243.880 ;
        RECT 806.910 243.820 807.230 243.880 ;
        RECT 806.910 19.960 807.230 20.020 ;
        RECT 1108.670 19.960 1108.990 20.020 ;
        RECT 806.910 19.820 1108.990 19.960 ;
        RECT 806.910 19.760 807.230 19.820 ;
        RECT 1108.670 19.760 1108.990 19.820 ;
      LAYER via ;
        RECT 801.420 243.820 801.680 244.080 ;
        RECT 806.940 243.820 807.200 244.080 ;
        RECT 806.940 19.760 807.200 20.020 ;
        RECT 1108.700 19.760 1108.960 20.020 ;
      LAYER met2 ;
        RECT 801.370 260.000 801.650 264.000 ;
        RECT 801.480 244.110 801.620 260.000 ;
        RECT 801.420 243.790 801.680 244.110 ;
        RECT 806.940 243.790 807.200 244.110 ;
        RECT 807.000 20.050 807.140 243.790 ;
        RECT 806.940 19.730 807.200 20.050 ;
        RECT 1108.700 19.730 1108.960 20.050 ;
        RECT 1108.760 2.400 1108.900 19.730 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
=======
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 820.710 17.240 821.030 17.300 ;
        RECT 1126.610 17.240 1126.930 17.300 ;
        RECT 820.710 17.100 1126.930 17.240 ;
        RECT 820.710 17.040 821.030 17.100 ;
        RECT 1126.610 17.040 1126.930 17.100 ;
      LAYER via ;
        RECT 820.740 17.040 821.000 17.300 ;
        RECT 1126.640 17.040 1126.900 17.300 ;
      LAYER met2 ;
        RECT 819.310 260.170 819.590 264.000 ;
        RECT 819.310 260.030 820.940 260.170 ;
        RECT 819.310 260.000 819.590 260.030 ;
        RECT 820.800 17.330 820.940 260.030 ;
        RECT 820.740 17.010 821.000 17.330 ;
        RECT 1126.640 17.010 1126.900 17.330 ;
        RECT 1126.700 2.400 1126.840 17.010 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
=======
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 836.810 247.420 837.130 247.480 ;
        RECT 1139.490 247.420 1139.810 247.480 ;
        RECT 836.810 247.280 1139.810 247.420 ;
        RECT 836.810 247.220 837.130 247.280 ;
        RECT 1139.490 247.220 1139.810 247.280 ;
      LAYER via ;
        RECT 836.840 247.220 837.100 247.480 ;
        RECT 1139.520 247.220 1139.780 247.480 ;
      LAYER met2 ;
        RECT 836.790 260.000 837.070 264.000 ;
        RECT 836.900 247.510 837.040 260.000 ;
        RECT 836.840 247.190 837.100 247.510 ;
        RECT 1139.520 247.190 1139.780 247.510 ;
        RECT 1139.580 16.730 1139.720 247.190 ;
        RECT 1139.580 16.590 1144.780 16.730 ;
        RECT 1144.640 2.400 1144.780 16.590 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
=======
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 855.210 17.580 855.530 17.640 ;
        RECT 1162.490 17.580 1162.810 17.640 ;
        RECT 855.210 17.440 1162.810 17.580 ;
        RECT 855.210 17.380 855.530 17.440 ;
        RECT 1162.490 17.380 1162.810 17.440 ;
      LAYER via ;
        RECT 855.240 17.380 855.500 17.640 ;
        RECT 1162.520 17.380 1162.780 17.640 ;
      LAYER met2 ;
        RECT 854.730 260.170 855.010 264.000 ;
        RECT 854.730 260.030 855.440 260.170 ;
        RECT 854.730 260.000 855.010 260.030 ;
        RECT 855.300 17.670 855.440 260.030 ;
        RECT 855.240 17.350 855.500 17.670 ;
        RECT 1162.520 17.350 1162.780 17.670 ;
        RECT 1162.580 2.400 1162.720 17.350 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
=======
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 372.210 245.720 372.530 245.780 ;
        RECT 677.190 245.720 677.510 245.780 ;
        RECT 372.210 245.580 677.510 245.720 ;
        RECT 372.210 245.520 372.530 245.580 ;
        RECT 677.190 245.520 677.510 245.580 ;
      LAYER via ;
        RECT 372.240 245.520 372.500 245.780 ;
        RECT 677.220 245.520 677.480 245.780 ;
      LAYER met2 ;
        RECT 372.190 260.000 372.470 264.000 ;
        RECT 372.300 245.810 372.440 260.000 ;
        RECT 372.240 245.490 372.500 245.810 ;
        RECT 677.220 245.490 677.480 245.810 ;
        RECT 677.280 16.730 677.420 245.490 ;
        RECT 677.280 16.590 680.640 16.730 ;
        RECT 680.500 2.400 680.640 16.590 ;
        RECT 680.290 -4.800 680.850 2.400 ;
=======
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 872.690 246.400 873.010 246.460 ;
        RECT 1180.890 246.400 1181.210 246.460 ;
        RECT 872.690 246.260 1181.210 246.400 ;
        RECT 872.690 246.200 873.010 246.260 ;
        RECT 1180.890 246.200 1181.210 246.260 ;
      LAYER via ;
        RECT 872.720 246.200 872.980 246.460 ;
        RECT 1180.920 246.200 1181.180 246.460 ;
      LAYER met2 ;
        RECT 872.670 260.000 872.950 264.000 ;
        RECT 872.780 246.490 872.920 260.000 ;
        RECT 872.720 246.170 872.980 246.490 ;
        RECT 1180.920 246.170 1181.180 246.490 ;
        RECT 1180.980 17.410 1181.120 246.170 ;
        RECT 1180.060 17.270 1181.120 17.410 ;
        RECT 1180.060 2.400 1180.200 17.270 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
=======
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 890.630 244.020 890.950 244.080 ;
        RECT 896.610 244.020 896.930 244.080 ;
        RECT 890.630 243.880 896.930 244.020 ;
        RECT 890.630 243.820 890.950 243.880 ;
        RECT 896.610 243.820 896.930 243.880 ;
        RECT 896.610 15.540 896.930 15.600 ;
        RECT 1197.910 15.540 1198.230 15.600 ;
        RECT 896.610 15.400 1198.230 15.540 ;
        RECT 896.610 15.340 896.930 15.400 ;
        RECT 1197.910 15.340 1198.230 15.400 ;
      LAYER via ;
        RECT 890.660 243.820 890.920 244.080 ;
        RECT 896.640 243.820 896.900 244.080 ;
        RECT 896.640 15.340 896.900 15.600 ;
        RECT 1197.940 15.340 1198.200 15.600 ;
      LAYER met2 ;
        RECT 890.610 260.000 890.890 264.000 ;
        RECT 890.720 244.110 890.860 260.000 ;
        RECT 890.660 243.790 890.920 244.110 ;
        RECT 896.640 243.790 896.900 244.110 ;
        RECT 896.700 15.630 896.840 243.790 ;
        RECT 896.640 15.310 896.900 15.630 ;
        RECT 1197.940 15.310 1198.200 15.630 ;
        RECT 1198.000 2.400 1198.140 15.310 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
=======
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 908.570 245.040 908.890 245.100 ;
        RECT 1214.930 245.040 1215.250 245.100 ;
        RECT 908.570 244.900 1215.250 245.040 ;
        RECT 908.570 244.840 908.890 244.900 ;
        RECT 1214.930 244.840 1215.250 244.900 ;
      LAYER via ;
        RECT 908.600 244.840 908.860 245.100 ;
        RECT 1214.960 244.840 1215.220 245.100 ;
      LAYER met2 ;
        RECT 908.550 260.000 908.830 264.000 ;
        RECT 908.660 245.130 908.800 260.000 ;
        RECT 908.600 244.810 908.860 245.130 ;
        RECT 1214.960 244.810 1215.220 245.130 ;
        RECT 1215.020 16.730 1215.160 244.810 ;
        RECT 1215.020 16.590 1216.080 16.730 ;
        RECT 1215.940 2.400 1216.080 16.590 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
=======
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 926.510 244.020 926.830 244.080 ;
        RECT 931.110 244.020 931.430 244.080 ;
        RECT 926.510 243.880 931.430 244.020 ;
        RECT 926.510 243.820 926.830 243.880 ;
        RECT 931.110 243.820 931.430 243.880 ;
        RECT 931.110 15.200 931.430 15.260 ;
        RECT 1233.790 15.200 1234.110 15.260 ;
        RECT 931.110 15.060 1234.110 15.200 ;
        RECT 931.110 15.000 931.430 15.060 ;
        RECT 1233.790 15.000 1234.110 15.060 ;
      LAYER via ;
        RECT 926.540 243.820 926.800 244.080 ;
        RECT 931.140 243.820 931.400 244.080 ;
        RECT 931.140 15.000 931.400 15.260 ;
        RECT 1233.820 15.000 1234.080 15.260 ;
      LAYER met2 ;
        RECT 926.490 260.000 926.770 264.000 ;
        RECT 926.600 244.110 926.740 260.000 ;
        RECT 926.540 243.790 926.800 244.110 ;
        RECT 931.140 243.790 931.400 244.110 ;
        RECT 931.200 15.290 931.340 243.790 ;
        RECT 931.140 14.970 931.400 15.290 ;
        RECT 1233.820 14.970 1234.080 15.290 ;
        RECT 1233.880 2.400 1234.020 14.970 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
=======
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 944.450 246.740 944.770 246.800 ;
        RECT 1249.430 246.740 1249.750 246.800 ;
        RECT 944.450 246.600 1249.750 246.740 ;
        RECT 944.450 246.540 944.770 246.600 ;
        RECT 1249.430 246.540 1249.750 246.600 ;
      LAYER via ;
        RECT 944.480 246.540 944.740 246.800 ;
        RECT 1249.460 246.540 1249.720 246.800 ;
      LAYER met2 ;
        RECT 944.430 260.000 944.710 264.000 ;
        RECT 944.540 246.830 944.680 260.000 ;
        RECT 944.480 246.510 944.740 246.830 ;
        RECT 1249.460 246.510 1249.720 246.830 ;
        RECT 1249.520 16.730 1249.660 246.510 ;
        RECT 1249.520 16.590 1251.960 16.730 ;
        RECT 1251.820 2.400 1251.960 16.590 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
=======
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 965.610 15.880 965.930 15.940 ;
        RECT 1269.210 15.880 1269.530 15.940 ;
        RECT 965.610 15.740 1269.530 15.880 ;
        RECT 965.610 15.680 965.930 15.740 ;
        RECT 1269.210 15.680 1269.530 15.740 ;
      LAYER via ;
        RECT 965.640 15.680 965.900 15.940 ;
        RECT 1269.240 15.680 1269.500 15.940 ;
      LAYER met2 ;
        RECT 961.910 260.170 962.190 264.000 ;
        RECT 961.910 260.030 965.840 260.170 ;
        RECT 961.910 260.000 962.190 260.030 ;
        RECT 965.700 15.970 965.840 260.030 ;
        RECT 965.640 15.650 965.900 15.970 ;
        RECT 1269.240 15.650 1269.500 15.970 ;
        RECT 1269.300 2.400 1269.440 15.650 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
=======
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 979.870 243.340 980.190 243.400 ;
        RECT 986.310 243.340 986.630 243.400 ;
        RECT 979.870 243.200 986.630 243.340 ;
        RECT 979.870 243.140 980.190 243.200 ;
        RECT 986.310 243.140 986.630 243.200 ;
        RECT 986.310 16.220 986.630 16.280 ;
        RECT 1287.150 16.220 1287.470 16.280 ;
        RECT 986.310 16.080 1287.470 16.220 ;
        RECT 986.310 16.020 986.630 16.080 ;
        RECT 1287.150 16.020 1287.470 16.080 ;
      LAYER via ;
        RECT 979.900 243.140 980.160 243.400 ;
        RECT 986.340 243.140 986.600 243.400 ;
        RECT 986.340 16.020 986.600 16.280 ;
        RECT 1287.180 16.020 1287.440 16.280 ;
      LAYER met2 ;
        RECT 979.850 260.000 980.130 264.000 ;
        RECT 979.960 243.430 980.100 260.000 ;
        RECT 979.900 243.110 980.160 243.430 ;
        RECT 986.340 243.110 986.600 243.430 ;
        RECT 986.400 16.310 986.540 243.110 ;
        RECT 986.340 15.990 986.600 16.310 ;
        RECT 1287.180 15.990 1287.440 16.310 ;
        RECT 1287.240 2.400 1287.380 15.990 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
=======
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1000.110 19.620 1000.430 19.680 ;
        RECT 1305.090 19.620 1305.410 19.680 ;
        RECT 1000.110 19.480 1305.410 19.620 ;
        RECT 1000.110 19.420 1000.430 19.480 ;
        RECT 1305.090 19.420 1305.410 19.480 ;
      LAYER via ;
        RECT 1000.140 19.420 1000.400 19.680 ;
        RECT 1305.120 19.420 1305.380 19.680 ;
      LAYER met2 ;
        RECT 997.790 260.170 998.070 264.000 ;
        RECT 997.790 260.030 1000.340 260.170 ;
        RECT 997.790 260.000 998.070 260.030 ;
        RECT 1000.200 19.710 1000.340 260.030 ;
        RECT 1000.140 19.390 1000.400 19.710 ;
        RECT 1305.120 19.390 1305.380 19.710 ;
        RECT 1305.180 2.400 1305.320 19.390 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
=======
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1015.750 244.020 1016.070 244.080 ;
        RECT 1020.810 244.020 1021.130 244.080 ;
        RECT 1015.750 243.880 1021.130 244.020 ;
        RECT 1015.750 243.820 1016.070 243.880 ;
        RECT 1020.810 243.820 1021.130 243.880 ;
        RECT 1020.810 16.560 1021.130 16.620 ;
        RECT 1323.030 16.560 1323.350 16.620 ;
        RECT 1020.810 16.420 1323.350 16.560 ;
        RECT 1020.810 16.360 1021.130 16.420 ;
        RECT 1323.030 16.360 1323.350 16.420 ;
      LAYER via ;
        RECT 1015.780 243.820 1016.040 244.080 ;
        RECT 1020.840 243.820 1021.100 244.080 ;
        RECT 1020.840 16.360 1021.100 16.620 ;
        RECT 1323.060 16.360 1323.320 16.620 ;
      LAYER met2 ;
        RECT 1015.730 260.000 1016.010 264.000 ;
        RECT 1015.840 244.110 1015.980 260.000 ;
        RECT 1015.780 243.790 1016.040 244.110 ;
        RECT 1020.840 243.790 1021.100 244.110 ;
        RECT 1020.900 16.650 1021.040 243.790 ;
        RECT 1020.840 16.330 1021.100 16.650 ;
        RECT 1323.060 16.330 1323.320 16.650 ;
        RECT 1323.120 2.400 1323.260 16.330 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
=======
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1034.610 18.600 1034.930 18.660 ;
        RECT 1340.510 18.600 1340.830 18.660 ;
        RECT 1034.610 18.460 1340.830 18.600 ;
        RECT 1034.610 18.400 1034.930 18.460 ;
        RECT 1340.510 18.400 1340.830 18.460 ;
      LAYER via ;
        RECT 1034.640 18.400 1034.900 18.660 ;
        RECT 1340.540 18.400 1340.800 18.660 ;
      LAYER met2 ;
        RECT 1033.670 260.170 1033.950 264.000 ;
        RECT 1033.670 260.030 1034.840 260.170 ;
        RECT 1033.670 260.000 1033.950 260.030 ;
        RECT 1034.700 18.690 1034.840 260.030 ;
        RECT 1034.640 18.370 1034.900 18.690 ;
        RECT 1340.540 18.370 1340.800 18.690 ;
        RECT 1340.600 2.400 1340.740 18.370 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
=======
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 663.020 19.480 669.600 19.620 ;
        RECT 392.910 19.280 393.230 19.340 ;
        RECT 663.020 19.280 663.160 19.480 ;
        RECT 392.910 19.140 663.160 19.280 ;
        RECT 669.460 19.280 669.600 19.480 ;
        RECT 698.350 19.280 698.670 19.340 ;
        RECT 669.460 19.140 698.670 19.280 ;
        RECT 392.910 19.080 393.230 19.140 ;
        RECT 698.350 19.080 698.670 19.140 ;
      LAYER via ;
        RECT 392.940 19.080 393.200 19.340 ;
        RECT 698.380 19.080 698.640 19.340 ;
      LAYER met2 ;
        RECT 390.130 260.170 390.410 264.000 ;
        RECT 390.130 260.030 393.140 260.170 ;
        RECT 390.130 260.000 390.410 260.030 ;
        RECT 393.000 19.370 393.140 260.030 ;
        RECT 392.940 19.050 393.200 19.370 ;
        RECT 698.380 19.050 698.640 19.370 ;
        RECT 698.440 2.400 698.580 19.050 ;
        RECT 698.230 -4.800 698.790 2.400 ;
=======
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1051.630 246.060 1051.950 246.120 ;
        RECT 1352.470 246.060 1352.790 246.120 ;
        RECT 1051.630 245.920 1352.790 246.060 ;
        RECT 1051.630 245.860 1051.950 245.920 ;
        RECT 1352.470 245.860 1352.790 245.920 ;
        RECT 1352.470 16.900 1352.790 16.960 ;
        RECT 1358.450 16.900 1358.770 16.960 ;
        RECT 1352.470 16.760 1358.770 16.900 ;
        RECT 1352.470 16.700 1352.790 16.760 ;
        RECT 1358.450 16.700 1358.770 16.760 ;
      LAYER via ;
        RECT 1051.660 245.860 1051.920 246.120 ;
        RECT 1352.500 245.860 1352.760 246.120 ;
        RECT 1352.500 16.700 1352.760 16.960 ;
        RECT 1358.480 16.700 1358.740 16.960 ;
      LAYER met2 ;
        RECT 1051.610 260.000 1051.890 264.000 ;
        RECT 1051.720 246.150 1051.860 260.000 ;
        RECT 1051.660 245.830 1051.920 246.150 ;
        RECT 1352.500 245.830 1352.760 246.150 ;
        RECT 1352.560 16.990 1352.700 245.830 ;
        RECT 1352.500 16.670 1352.760 16.990 ;
        RECT 1358.480 16.670 1358.740 16.990 ;
        RECT 1358.540 2.400 1358.680 16.670 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
=======
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1069.570 244.020 1069.890 244.080 ;
        RECT 1076.010 244.020 1076.330 244.080 ;
        RECT 1069.570 243.880 1076.330 244.020 ;
        RECT 1069.570 243.820 1069.890 243.880 ;
        RECT 1076.010 243.820 1076.330 243.880 ;
        RECT 1076.010 16.900 1076.330 16.960 ;
        RECT 1076.010 16.760 1338.900 16.900 ;
        RECT 1076.010 16.700 1076.330 16.760 ;
        RECT 1338.760 16.220 1338.900 16.760 ;
        RECT 1376.390 16.220 1376.710 16.280 ;
        RECT 1338.760 16.080 1376.710 16.220 ;
        RECT 1376.390 16.020 1376.710 16.080 ;
      LAYER via ;
        RECT 1069.600 243.820 1069.860 244.080 ;
        RECT 1076.040 243.820 1076.300 244.080 ;
        RECT 1076.040 16.700 1076.300 16.960 ;
        RECT 1376.420 16.020 1376.680 16.280 ;
      LAYER met2 ;
        RECT 1069.550 260.000 1069.830 264.000 ;
        RECT 1069.660 244.110 1069.800 260.000 ;
        RECT 1069.600 243.790 1069.860 244.110 ;
        RECT 1076.040 243.790 1076.300 244.110 ;
        RECT 1076.100 16.990 1076.240 243.790 ;
        RECT 1076.040 16.670 1076.300 16.990 ;
        RECT 1376.420 15.990 1376.680 16.310 ;
        RECT 1376.480 2.400 1376.620 15.990 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
=======
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1087.050 245.380 1087.370 245.440 ;
        RECT 1394.790 245.380 1395.110 245.440 ;
        RECT 1087.050 245.240 1395.110 245.380 ;
        RECT 1087.050 245.180 1087.370 245.240 ;
        RECT 1394.790 245.180 1395.110 245.240 ;
      LAYER via ;
        RECT 1087.080 245.180 1087.340 245.440 ;
        RECT 1394.820 245.180 1395.080 245.440 ;
      LAYER met2 ;
        RECT 1087.030 260.000 1087.310 264.000 ;
        RECT 1087.140 245.470 1087.280 260.000 ;
        RECT 1087.080 245.150 1087.340 245.470 ;
        RECT 1394.820 245.150 1395.080 245.470 ;
        RECT 1394.880 17.410 1395.020 245.150 ;
        RECT 1394.420 17.270 1395.020 17.410 ;
        RECT 1394.420 2.400 1394.560 17.270 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
=======
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1104.990 244.020 1105.310 244.080 ;
        RECT 1110.510 244.020 1110.830 244.080 ;
        RECT 1104.990 243.880 1110.830 244.020 ;
        RECT 1104.990 243.820 1105.310 243.880 ;
        RECT 1110.510 243.820 1110.830 243.880 ;
        RECT 1110.510 18.940 1110.830 19.000 ;
        RECT 1412.270 18.940 1412.590 19.000 ;
        RECT 1110.510 18.800 1412.590 18.940 ;
        RECT 1110.510 18.740 1110.830 18.800 ;
        RECT 1412.270 18.740 1412.590 18.800 ;
      LAYER via ;
        RECT 1105.020 243.820 1105.280 244.080 ;
        RECT 1110.540 243.820 1110.800 244.080 ;
        RECT 1110.540 18.740 1110.800 19.000 ;
        RECT 1412.300 18.740 1412.560 19.000 ;
      LAYER met2 ;
        RECT 1104.970 260.000 1105.250 264.000 ;
        RECT 1105.080 244.110 1105.220 260.000 ;
        RECT 1105.020 243.790 1105.280 244.110 ;
        RECT 1110.540 243.790 1110.800 244.110 ;
        RECT 1110.600 19.030 1110.740 243.790 ;
        RECT 1110.540 18.710 1110.800 19.030 ;
        RECT 1412.300 18.710 1412.560 19.030 ;
        RECT 1412.360 2.400 1412.500 18.710 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
=======
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1122.930 245.720 1123.250 245.780 ;
        RECT 1428.830 245.720 1429.150 245.780 ;
        RECT 1122.930 245.580 1429.150 245.720 ;
        RECT 1122.930 245.520 1123.250 245.580 ;
        RECT 1428.830 245.520 1429.150 245.580 ;
      LAYER via ;
        RECT 1122.960 245.520 1123.220 245.780 ;
        RECT 1428.860 245.520 1429.120 245.780 ;
      LAYER met2 ;
        RECT 1122.910 260.000 1123.190 264.000 ;
        RECT 1123.020 245.810 1123.160 260.000 ;
        RECT 1122.960 245.490 1123.220 245.810 ;
        RECT 1428.860 245.490 1429.120 245.810 ;
        RECT 1428.920 16.900 1429.060 245.490 ;
        RECT 1428.920 16.760 1429.980 16.900 ;
        RECT 1429.840 2.400 1429.980 16.760 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
=======
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1140.870 244.020 1141.190 244.080 ;
        RECT 1145.010 244.020 1145.330 244.080 ;
        RECT 1140.870 243.880 1145.330 244.020 ;
        RECT 1140.870 243.820 1141.190 243.880 ;
        RECT 1145.010 243.820 1145.330 243.880 ;
        RECT 1145.010 19.280 1145.330 19.340 ;
        RECT 1447.690 19.280 1448.010 19.340 ;
        RECT 1145.010 19.140 1448.010 19.280 ;
        RECT 1145.010 19.080 1145.330 19.140 ;
        RECT 1447.690 19.080 1448.010 19.140 ;
      LAYER via ;
        RECT 1140.900 243.820 1141.160 244.080 ;
        RECT 1145.040 243.820 1145.300 244.080 ;
        RECT 1145.040 19.080 1145.300 19.340 ;
        RECT 1447.720 19.080 1447.980 19.340 ;
      LAYER met2 ;
        RECT 1140.850 260.000 1141.130 264.000 ;
        RECT 1140.960 244.110 1141.100 260.000 ;
        RECT 1140.900 243.790 1141.160 244.110 ;
        RECT 1145.040 243.790 1145.300 244.110 ;
        RECT 1145.100 19.370 1145.240 243.790 ;
        RECT 1145.040 19.050 1145.300 19.370 ;
        RECT 1447.720 19.050 1447.980 19.370 ;
        RECT 1447.780 2.400 1447.920 19.050 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
=======
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1158.810 18.260 1159.130 18.320 ;
        RECT 1465.630 18.260 1465.950 18.320 ;
        RECT 1158.810 18.120 1465.950 18.260 ;
        RECT 1158.810 18.060 1159.130 18.120 ;
        RECT 1465.630 18.060 1465.950 18.120 ;
      LAYER via ;
        RECT 1158.840 18.060 1159.100 18.320 ;
        RECT 1465.660 18.060 1465.920 18.320 ;
      LAYER met2 ;
        RECT 1158.790 260.000 1159.070 264.000 ;
        RECT 1158.900 18.350 1159.040 260.000 ;
        RECT 1158.840 18.030 1159.100 18.350 ;
        RECT 1465.660 18.030 1465.920 18.350 ;
        RECT 1465.720 2.400 1465.860 18.030 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
=======
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1179.510 17.240 1179.830 17.300 ;
        RECT 1483.570 17.240 1483.890 17.300 ;
        RECT 1179.510 17.100 1483.890 17.240 ;
        RECT 1179.510 17.040 1179.830 17.100 ;
        RECT 1483.570 17.040 1483.890 17.100 ;
      LAYER via ;
        RECT 1179.540 17.040 1179.800 17.300 ;
        RECT 1483.600 17.040 1483.860 17.300 ;
      LAYER met2 ;
        RECT 1176.730 260.170 1177.010 264.000 ;
        RECT 1176.730 260.030 1179.740 260.170 ;
        RECT 1176.730 260.000 1177.010 260.030 ;
        RECT 1179.600 17.330 1179.740 260.030 ;
        RECT 1179.540 17.010 1179.800 17.330 ;
        RECT 1483.600 17.010 1483.860 17.330 ;
        RECT 1483.660 2.400 1483.800 17.010 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
=======
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1194.690 243.680 1195.010 243.740 ;
        RECT 1200.210 243.680 1200.530 243.740 ;
        RECT 1194.690 243.540 1200.530 243.680 ;
        RECT 1194.690 243.480 1195.010 243.540 ;
        RECT 1200.210 243.480 1200.530 243.540 ;
        RECT 1200.210 20.640 1200.530 20.700 ;
        RECT 1501.510 20.640 1501.830 20.700 ;
        RECT 1200.210 20.500 1501.830 20.640 ;
        RECT 1200.210 20.440 1200.530 20.500 ;
        RECT 1501.510 20.440 1501.830 20.500 ;
      LAYER via ;
        RECT 1194.720 243.480 1194.980 243.740 ;
        RECT 1200.240 243.480 1200.500 243.740 ;
        RECT 1200.240 20.440 1200.500 20.700 ;
        RECT 1501.540 20.440 1501.800 20.700 ;
      LAYER met2 ;
        RECT 1194.670 260.000 1194.950 264.000 ;
        RECT 1194.780 243.770 1194.920 260.000 ;
        RECT 1194.720 243.450 1194.980 243.770 ;
        RECT 1200.240 243.450 1200.500 243.770 ;
        RECT 1200.300 20.730 1200.440 243.450 ;
        RECT 1200.240 20.410 1200.500 20.730 ;
        RECT 1501.540 20.410 1501.800 20.730 ;
        RECT 1501.600 2.400 1501.740 20.410 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
=======
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1214.010 17.920 1214.330 17.980 ;
        RECT 1518.990 17.920 1519.310 17.980 ;
        RECT 1214.010 17.780 1519.310 17.920 ;
        RECT 1214.010 17.720 1214.330 17.780 ;
        RECT 1518.990 17.720 1519.310 17.780 ;
      LAYER via ;
        RECT 1214.040 17.720 1214.300 17.980 ;
        RECT 1519.020 17.720 1519.280 17.980 ;
      LAYER met2 ;
        RECT 1212.150 260.170 1212.430 264.000 ;
        RECT 1212.150 260.030 1214.240 260.170 ;
        RECT 1212.150 260.000 1212.430 260.030 ;
        RECT 1214.100 18.010 1214.240 260.030 ;
        RECT 1214.040 17.690 1214.300 18.010 ;
        RECT 1519.020 17.690 1519.280 18.010 ;
        RECT 1519.080 2.400 1519.220 17.690 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
=======
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 408.090 246.060 408.410 246.120 ;
        RECT 711.230 246.060 711.550 246.120 ;
        RECT 408.090 245.920 711.550 246.060 ;
        RECT 408.090 245.860 408.410 245.920 ;
        RECT 711.230 245.860 711.550 245.920 ;
      LAYER via ;
        RECT 408.120 245.860 408.380 246.120 ;
        RECT 711.260 245.860 711.520 246.120 ;
      LAYER met2 ;
        RECT 408.070 260.000 408.350 264.000 ;
        RECT 408.180 246.150 408.320 260.000 ;
        RECT 408.120 245.830 408.380 246.150 ;
        RECT 711.260 245.830 711.520 246.150 ;
        RECT 711.320 16.730 711.460 245.830 ;
        RECT 711.320 16.590 716.520 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
=======
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1230.110 244.020 1230.430 244.080 ;
        RECT 1234.710 244.020 1235.030 244.080 ;
        RECT 1230.110 243.880 1235.030 244.020 ;
        RECT 1230.110 243.820 1230.430 243.880 ;
        RECT 1234.710 243.820 1235.030 243.880 ;
        RECT 1234.710 19.960 1235.030 20.020 ;
        RECT 1536.930 19.960 1537.250 20.020 ;
        RECT 1234.710 19.820 1537.250 19.960 ;
        RECT 1234.710 19.760 1235.030 19.820 ;
        RECT 1536.930 19.760 1537.250 19.820 ;
      LAYER via ;
        RECT 1230.140 243.820 1230.400 244.080 ;
        RECT 1234.740 243.820 1235.000 244.080 ;
        RECT 1234.740 19.760 1235.000 20.020 ;
        RECT 1536.960 19.760 1537.220 20.020 ;
      LAYER met2 ;
        RECT 1230.090 260.000 1230.370 264.000 ;
        RECT 1230.200 244.110 1230.340 260.000 ;
        RECT 1230.140 243.790 1230.400 244.110 ;
        RECT 1234.740 243.790 1235.000 244.110 ;
        RECT 1234.800 20.050 1234.940 243.790 ;
        RECT 1234.740 19.730 1235.000 20.050 ;
        RECT 1536.960 19.730 1537.220 20.050 ;
        RECT 1537.020 2.400 1537.160 19.730 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
=======
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1248.510 17.580 1248.830 17.640 ;
        RECT 1554.870 17.580 1555.190 17.640 ;
        RECT 1248.510 17.440 1555.190 17.580 ;
        RECT 1248.510 17.380 1248.830 17.440 ;
        RECT 1554.870 17.380 1555.190 17.440 ;
      LAYER via ;
        RECT 1248.540 17.380 1248.800 17.640 ;
        RECT 1554.900 17.380 1555.160 17.640 ;
      LAYER met2 ;
        RECT 1248.030 260.170 1248.310 264.000 ;
        RECT 1248.030 260.030 1248.740 260.170 ;
        RECT 1248.030 260.000 1248.310 260.030 ;
        RECT 1248.600 17.670 1248.740 260.030 ;
        RECT 1248.540 17.350 1248.800 17.670 ;
        RECT 1554.900 17.350 1555.160 17.670 ;
        RECT 1554.960 2.400 1555.100 17.350 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
=======
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1265.990 246.400 1266.310 246.460 ;
        RECT 1567.290 246.400 1567.610 246.460 ;
        RECT 1265.990 246.260 1567.610 246.400 ;
        RECT 1265.990 246.200 1266.310 246.260 ;
        RECT 1567.290 246.200 1567.610 246.260 ;
      LAYER via ;
        RECT 1266.020 246.200 1266.280 246.460 ;
        RECT 1567.320 246.200 1567.580 246.460 ;
      LAYER met2 ;
        RECT 1265.970 260.000 1266.250 264.000 ;
        RECT 1266.080 246.490 1266.220 260.000 ;
        RECT 1266.020 246.170 1266.280 246.490 ;
        RECT 1567.320 246.170 1567.580 246.490 ;
        RECT 1567.380 16.730 1567.520 246.170 ;
        RECT 1567.380 16.590 1573.040 16.730 ;
        RECT 1572.900 2.400 1573.040 16.590 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
=======
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1283.930 244.020 1284.250 244.080 ;
        RECT 1289.910 244.020 1290.230 244.080 ;
        RECT 1283.930 243.880 1290.230 244.020 ;
        RECT 1283.930 243.820 1284.250 243.880 ;
        RECT 1289.910 243.820 1290.230 243.880 ;
        RECT 1289.910 20.300 1290.230 20.360 ;
        RECT 1590.290 20.300 1590.610 20.360 ;
        RECT 1289.910 20.160 1590.610 20.300 ;
        RECT 1289.910 20.100 1290.230 20.160 ;
        RECT 1590.290 20.100 1590.610 20.160 ;
      LAYER via ;
        RECT 1283.960 243.820 1284.220 244.080 ;
        RECT 1289.940 243.820 1290.200 244.080 ;
        RECT 1289.940 20.100 1290.200 20.360 ;
        RECT 1590.320 20.100 1590.580 20.360 ;
      LAYER met2 ;
        RECT 1283.910 260.000 1284.190 264.000 ;
        RECT 1284.020 244.110 1284.160 260.000 ;
        RECT 1283.960 243.790 1284.220 244.110 ;
        RECT 1289.940 243.790 1290.200 244.110 ;
        RECT 1290.000 20.390 1290.140 243.790 ;
        RECT 1289.940 20.070 1290.200 20.390 ;
        RECT 1590.320 20.070 1590.580 20.390 ;
        RECT 1590.380 2.400 1590.520 20.070 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
=======
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1301.870 245.040 1302.190 245.100 ;
        RECT 1608.690 245.040 1609.010 245.100 ;
        RECT 1301.870 244.900 1609.010 245.040 ;
        RECT 1301.870 244.840 1302.190 244.900 ;
        RECT 1608.690 244.840 1609.010 244.900 ;
      LAYER via ;
        RECT 1301.900 244.840 1302.160 245.100 ;
        RECT 1608.720 244.840 1608.980 245.100 ;
      LAYER met2 ;
        RECT 1301.850 260.000 1302.130 264.000 ;
        RECT 1301.960 245.130 1302.100 260.000 ;
        RECT 1301.900 244.810 1302.160 245.130 ;
        RECT 1608.720 244.810 1608.980 245.130 ;
        RECT 1608.780 37.810 1608.920 244.810 ;
        RECT 1608.320 37.670 1608.920 37.810 ;
        RECT 1608.320 2.400 1608.460 37.670 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
=======
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1319.810 244.020 1320.130 244.080 ;
        RECT 1324.410 244.020 1324.730 244.080 ;
        RECT 1319.810 243.880 1324.730 244.020 ;
        RECT 1319.810 243.820 1320.130 243.880 ;
        RECT 1324.410 243.820 1324.730 243.880 ;
        RECT 1626.170 38.660 1626.490 38.720 ;
        RECT 1607.860 38.520 1626.490 38.660 ;
        RECT 1324.410 38.320 1324.730 38.380 ;
        RECT 1607.860 38.320 1608.000 38.520 ;
        RECT 1626.170 38.460 1626.490 38.520 ;
        RECT 1324.410 38.180 1608.000 38.320 ;
        RECT 1324.410 38.120 1324.730 38.180 ;
      LAYER via ;
        RECT 1319.840 243.820 1320.100 244.080 ;
        RECT 1324.440 243.820 1324.700 244.080 ;
        RECT 1324.440 38.120 1324.700 38.380 ;
        RECT 1626.200 38.460 1626.460 38.720 ;
      LAYER met2 ;
        RECT 1319.790 260.000 1320.070 264.000 ;
        RECT 1319.900 244.110 1320.040 260.000 ;
        RECT 1319.840 243.790 1320.100 244.110 ;
        RECT 1324.440 243.790 1324.700 244.110 ;
        RECT 1324.500 38.410 1324.640 243.790 ;
        RECT 1626.200 38.430 1626.460 38.750 ;
        RECT 1324.440 38.090 1324.700 38.410 ;
        RECT 1626.260 2.400 1626.400 38.430 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
=======
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 1642.345 48.365 1642.515 96.475 ;
      LAYER mcon ;
        RECT 1642.345 96.305 1642.515 96.475 ;
      LAYER met1 ;
        RECT 1338.210 127.740 1338.530 127.800 ;
        RECT 1642.730 127.740 1643.050 127.800 ;
        RECT 1338.210 127.600 1643.050 127.740 ;
        RECT 1338.210 127.540 1338.530 127.600 ;
        RECT 1642.730 127.540 1643.050 127.600 ;
        RECT 1642.270 96.460 1642.590 96.520 ;
        RECT 1642.270 96.320 1642.785 96.460 ;
        RECT 1642.270 96.260 1642.590 96.320 ;
        RECT 1642.285 48.520 1642.575 48.565 ;
        RECT 1644.110 48.520 1644.430 48.580 ;
        RECT 1642.285 48.380 1644.430 48.520 ;
        RECT 1642.285 48.335 1642.575 48.380 ;
        RECT 1644.110 48.320 1644.430 48.380 ;
        RECT 1644.110 2.960 1644.430 3.020 ;
        RECT 1644.570 2.960 1644.890 3.020 ;
        RECT 1644.110 2.820 1644.890 2.960 ;
        RECT 1644.110 2.760 1644.430 2.820 ;
        RECT 1644.570 2.760 1644.890 2.820 ;
      LAYER via ;
        RECT 1338.240 127.540 1338.500 127.800 ;
        RECT 1642.760 127.540 1643.020 127.800 ;
        RECT 1642.300 96.260 1642.560 96.520 ;
        RECT 1644.140 48.320 1644.400 48.580 ;
        RECT 1644.140 2.760 1644.400 3.020 ;
        RECT 1644.600 2.760 1644.860 3.020 ;
      LAYER met2 ;
        RECT 1337.270 260.170 1337.550 264.000 ;
        RECT 1337.270 260.030 1338.440 260.170 ;
        RECT 1337.270 260.000 1337.550 260.030 ;
        RECT 1338.300 127.830 1338.440 260.030 ;
        RECT 1338.240 127.510 1338.500 127.830 ;
        RECT 1642.760 127.510 1643.020 127.830 ;
        RECT 1642.820 96.970 1642.960 127.510 ;
        RECT 1642.360 96.830 1642.960 96.970 ;
        RECT 1642.360 96.550 1642.500 96.830 ;
        RECT 1642.300 96.230 1642.560 96.550 ;
        RECT 1644.140 48.290 1644.400 48.610 ;
        RECT 1644.200 48.010 1644.340 48.290 ;
        RECT 1644.200 47.870 1644.800 48.010 ;
        RECT 1644.660 3.050 1644.800 47.870 ;
        RECT 1644.140 2.730 1644.400 3.050 ;
        RECT 1644.600 2.730 1644.860 3.050 ;
        RECT 1644.200 2.400 1644.340 2.730 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
=======
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1355.230 243.680 1355.550 243.740 ;
        RECT 1362.590 243.680 1362.910 243.740 ;
        RECT 1355.230 243.540 1362.910 243.680 ;
        RECT 1355.230 243.480 1355.550 243.540 ;
        RECT 1362.590 243.480 1362.910 243.540 ;
        RECT 1362.590 134.880 1362.910 134.940 ;
        RECT 1656.530 134.880 1656.850 134.940 ;
        RECT 1362.590 134.740 1656.850 134.880 ;
        RECT 1362.590 134.680 1362.910 134.740 ;
        RECT 1656.530 134.680 1656.850 134.740 ;
      LAYER via ;
        RECT 1355.260 243.480 1355.520 243.740 ;
        RECT 1362.620 243.480 1362.880 243.740 ;
        RECT 1362.620 134.680 1362.880 134.940 ;
        RECT 1656.560 134.680 1656.820 134.940 ;
      LAYER met2 ;
        RECT 1355.210 260.000 1355.490 264.000 ;
        RECT 1355.320 243.770 1355.460 260.000 ;
        RECT 1355.260 243.450 1355.520 243.770 ;
        RECT 1362.620 243.450 1362.880 243.770 ;
        RECT 1362.680 134.970 1362.820 243.450 ;
        RECT 1362.620 134.650 1362.880 134.970 ;
        RECT 1656.560 134.650 1656.820 134.970 ;
        RECT 1656.620 16.730 1656.760 134.650 ;
        RECT 1656.620 16.590 1662.280 16.730 ;
        RECT 1662.140 2.400 1662.280 16.590 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
=======
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1373.170 244.020 1373.490 244.080 ;
        RECT 1379.150 244.020 1379.470 244.080 ;
        RECT 1373.170 243.880 1379.470 244.020 ;
        RECT 1373.170 243.820 1373.490 243.880 ;
        RECT 1379.150 243.820 1379.470 243.880 ;
        RECT 1379.150 120.940 1379.470 121.000 ;
        RECT 1676.770 120.940 1677.090 121.000 ;
        RECT 1379.150 120.800 1677.090 120.940 ;
        RECT 1379.150 120.740 1379.470 120.800 ;
        RECT 1676.770 120.740 1677.090 120.800 ;
      LAYER via ;
        RECT 1373.200 243.820 1373.460 244.080 ;
        RECT 1379.180 243.820 1379.440 244.080 ;
        RECT 1379.180 120.740 1379.440 121.000 ;
        RECT 1676.800 120.740 1677.060 121.000 ;
      LAYER met2 ;
        RECT 1373.150 260.000 1373.430 264.000 ;
        RECT 1373.260 244.110 1373.400 260.000 ;
        RECT 1373.200 243.790 1373.460 244.110 ;
        RECT 1379.180 243.790 1379.440 244.110 ;
        RECT 1379.240 121.030 1379.380 243.790 ;
        RECT 1379.180 120.710 1379.440 121.030 ;
        RECT 1676.800 120.710 1677.060 121.030 ;
        RECT 1676.860 17.410 1677.000 120.710 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
=======
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1391.110 231.440 1391.430 231.500 ;
        RECT 1697.470 231.440 1697.790 231.500 ;
        RECT 1391.110 231.300 1697.790 231.440 ;
        RECT 1391.110 231.240 1391.430 231.300 ;
        RECT 1697.470 231.240 1697.790 231.300 ;
      LAYER via ;
        RECT 1391.140 231.240 1391.400 231.500 ;
        RECT 1697.500 231.240 1697.760 231.500 ;
      LAYER met2 ;
        RECT 1391.090 260.000 1391.370 264.000 ;
        RECT 1391.200 231.530 1391.340 260.000 ;
        RECT 1391.140 231.210 1391.400 231.530 ;
        RECT 1697.500 231.210 1697.760 231.530 ;
        RECT 1697.560 2.400 1697.700 231.210 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
=======
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 426.010 260.170 426.290 264.000 ;
        RECT 426.010 260.030 427.640 260.170 ;
        RECT 426.010 260.000 426.290 260.030 ;
        RECT 427.500 17.525 427.640 260.030 ;
        RECT 427.430 17.155 427.710 17.525 ;
        RECT 734.250 17.155 734.530 17.525 ;
        RECT 734.320 2.400 734.460 17.155 ;
        RECT 734.110 -4.800 734.670 2.400 ;
      LAYER via2 ;
        RECT 427.430 17.200 427.710 17.480 ;
        RECT 734.250 17.200 734.530 17.480 ;
      LAYER met3 ;
        RECT 427.405 17.490 427.735 17.505 ;
        RECT 734.225 17.490 734.555 17.505 ;
        RECT 427.405 17.190 734.555 17.490 ;
        RECT 427.405 17.175 427.735 17.190 ;
        RECT 734.225 17.175 734.555 17.190 ;
=======
        RECT 734.110 -4.800 734.670 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1409.050 244.020 1409.370 244.080 ;
        RECT 1414.110 244.020 1414.430 244.080 ;
        RECT 1409.050 243.880 1414.430 244.020 ;
        RECT 1409.050 243.820 1409.370 243.880 ;
        RECT 1414.110 243.820 1414.430 243.880 ;
        RECT 1414.110 31.180 1414.430 31.240 ;
        RECT 1715.410 31.180 1715.730 31.240 ;
        RECT 1414.110 31.040 1715.730 31.180 ;
        RECT 1414.110 30.980 1414.430 31.040 ;
        RECT 1715.410 30.980 1715.730 31.040 ;
      LAYER via ;
        RECT 1409.080 243.820 1409.340 244.080 ;
        RECT 1414.140 243.820 1414.400 244.080 ;
        RECT 1414.140 30.980 1414.400 31.240 ;
        RECT 1715.440 30.980 1715.700 31.240 ;
      LAYER met2 ;
        RECT 1409.030 260.000 1409.310 264.000 ;
        RECT 1409.140 244.110 1409.280 260.000 ;
        RECT 1409.080 243.790 1409.340 244.110 ;
        RECT 1414.140 243.790 1414.400 244.110 ;
        RECT 1414.200 31.270 1414.340 243.790 ;
        RECT 1414.140 30.950 1414.400 31.270 ;
        RECT 1715.440 30.950 1715.700 31.270 ;
        RECT 1715.500 2.400 1715.640 30.950 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
=======
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1427.910 51.920 1428.230 51.980 ;
        RECT 1731.970 51.920 1732.290 51.980 ;
        RECT 1427.910 51.780 1732.290 51.920 ;
        RECT 1427.910 51.720 1428.230 51.780 ;
        RECT 1731.970 51.720 1732.290 51.780 ;
      LAYER via ;
        RECT 1427.940 51.720 1428.200 51.980 ;
        RECT 1732.000 51.720 1732.260 51.980 ;
      LAYER met2 ;
        RECT 1426.970 260.170 1427.250 264.000 ;
        RECT 1426.970 260.030 1428.140 260.170 ;
        RECT 1426.970 260.000 1427.250 260.030 ;
        RECT 1428.000 52.010 1428.140 260.030 ;
        RECT 1427.940 51.690 1428.200 52.010 ;
        RECT 1732.000 51.690 1732.260 52.010 ;
        RECT 1732.060 17.410 1732.200 51.690 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
=======
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1751.290 19.280 1751.610 19.340 ;
        RECT 1738.040 19.140 1751.610 19.280 ;
        RECT 1448.610 18.940 1448.930 19.000 ;
        RECT 1738.040 18.940 1738.180 19.140 ;
        RECT 1751.290 19.080 1751.610 19.140 ;
        RECT 1448.610 18.800 1738.180 18.940 ;
        RECT 1448.610 18.740 1448.930 18.800 ;
      LAYER via ;
        RECT 1448.640 18.740 1448.900 19.000 ;
        RECT 1751.320 19.080 1751.580 19.340 ;
      LAYER met2 ;
        RECT 1444.910 260.170 1445.190 264.000 ;
        RECT 1444.910 260.030 1448.840 260.170 ;
        RECT 1444.910 260.000 1445.190 260.030 ;
        RECT 1448.700 19.030 1448.840 260.030 ;
        RECT 1751.320 19.050 1751.580 19.370 ;
        RECT 1448.640 18.710 1448.900 19.030 ;
        RECT 1751.380 2.400 1751.520 19.050 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
=======
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 1737.565 19.125 1737.735 20.655 ;
      LAYER mcon ;
        RECT 1737.565 20.485 1737.735 20.655 ;
      LAYER met1 ;
        RECT 1462.870 244.020 1463.190 244.080 ;
        RECT 1469.310 244.020 1469.630 244.080 ;
        RECT 1462.870 243.880 1469.630 244.020 ;
        RECT 1462.870 243.820 1463.190 243.880 ;
        RECT 1469.310 243.820 1469.630 243.880 ;
        RECT 1737.505 20.640 1737.795 20.685 ;
        RECT 1768.770 20.640 1769.090 20.700 ;
        RECT 1737.505 20.500 1769.090 20.640 ;
        RECT 1737.505 20.455 1737.795 20.500 ;
        RECT 1768.770 20.440 1769.090 20.500 ;
        RECT 1469.310 19.280 1469.630 19.340 ;
        RECT 1737.505 19.280 1737.795 19.325 ;
        RECT 1469.310 19.140 1737.795 19.280 ;
        RECT 1469.310 19.080 1469.630 19.140 ;
        RECT 1737.505 19.095 1737.795 19.140 ;
      LAYER via ;
        RECT 1462.900 243.820 1463.160 244.080 ;
        RECT 1469.340 243.820 1469.600 244.080 ;
        RECT 1768.800 20.440 1769.060 20.700 ;
        RECT 1469.340 19.080 1469.600 19.340 ;
      LAYER met2 ;
        RECT 1462.850 260.000 1463.130 264.000 ;
        RECT 1462.960 244.110 1463.100 260.000 ;
        RECT 1462.900 243.790 1463.160 244.110 ;
        RECT 1469.340 243.790 1469.600 244.110 ;
        RECT 1469.400 19.370 1469.540 243.790 ;
        RECT 1768.800 20.410 1769.060 20.730 ;
        RECT 1469.340 19.050 1469.600 19.370 ;
        RECT 1768.860 2.400 1769.000 20.410 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
=======
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1483.110 18.600 1483.430 18.660 ;
        RECT 1786.710 18.600 1787.030 18.660 ;
        RECT 1483.110 18.460 1787.030 18.600 ;
        RECT 1483.110 18.400 1483.430 18.460 ;
        RECT 1786.710 18.400 1787.030 18.460 ;
      LAYER via ;
        RECT 1483.140 18.400 1483.400 18.660 ;
        RECT 1786.740 18.400 1787.000 18.660 ;
      LAYER met2 ;
        RECT 1480.330 260.170 1480.610 264.000 ;
        RECT 1480.330 260.030 1483.340 260.170 ;
        RECT 1480.330 260.000 1480.610 260.030 ;
        RECT 1483.200 18.690 1483.340 260.030 ;
        RECT 1483.140 18.370 1483.400 18.690 ;
        RECT 1786.740 18.370 1787.000 18.690 ;
        RECT 1786.800 2.400 1786.940 18.370 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
=======
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1498.290 244.020 1498.610 244.080 ;
        RECT 1503.810 244.020 1504.130 244.080 ;
        RECT 1498.290 243.880 1504.130 244.020 ;
        RECT 1498.290 243.820 1498.610 243.880 ;
        RECT 1503.810 243.820 1504.130 243.880 ;
        RECT 1503.810 17.240 1504.130 17.300 ;
        RECT 1804.650 17.240 1804.970 17.300 ;
        RECT 1503.810 17.100 1804.970 17.240 ;
        RECT 1503.810 17.040 1504.130 17.100 ;
        RECT 1804.650 17.040 1804.970 17.100 ;
      LAYER via ;
        RECT 1498.320 243.820 1498.580 244.080 ;
        RECT 1503.840 243.820 1504.100 244.080 ;
        RECT 1503.840 17.040 1504.100 17.300 ;
        RECT 1804.680 17.040 1804.940 17.300 ;
      LAYER met2 ;
        RECT 1498.270 260.000 1498.550 264.000 ;
        RECT 1498.380 244.110 1498.520 260.000 ;
        RECT 1498.320 243.790 1498.580 244.110 ;
        RECT 1503.840 243.790 1504.100 244.110 ;
        RECT 1503.900 17.330 1504.040 243.790 ;
        RECT 1503.840 17.010 1504.100 17.330 ;
        RECT 1804.680 17.010 1804.940 17.330 ;
        RECT 1804.740 2.400 1804.880 17.010 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
=======
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1517.610 58.720 1517.930 58.780 ;
        RECT 1821.670 58.720 1821.990 58.780 ;
        RECT 1517.610 58.580 1821.990 58.720 ;
        RECT 1517.610 58.520 1517.930 58.580 ;
        RECT 1821.670 58.520 1821.990 58.580 ;
      LAYER via ;
        RECT 1517.640 58.520 1517.900 58.780 ;
        RECT 1821.700 58.520 1821.960 58.780 ;
      LAYER met2 ;
        RECT 1516.210 260.170 1516.490 264.000 ;
        RECT 1516.210 260.030 1517.840 260.170 ;
        RECT 1516.210 260.000 1516.490 260.030 ;
        RECT 1517.700 58.810 1517.840 260.030 ;
        RECT 1517.640 58.490 1517.900 58.810 ;
        RECT 1821.700 58.490 1821.960 58.810 ;
        RECT 1821.760 16.730 1821.900 58.490 ;
        RECT 1821.760 16.590 1822.820 16.730 ;
        RECT 1822.680 2.400 1822.820 16.590 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
=======
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1534.170 244.020 1534.490 244.080 ;
        RECT 1538.310 244.020 1538.630 244.080 ;
        RECT 1534.170 243.880 1538.630 244.020 ;
        RECT 1534.170 243.820 1534.490 243.880 ;
        RECT 1538.310 243.820 1538.630 243.880 ;
        RECT 1538.310 19.620 1538.630 19.680 ;
        RECT 1840.070 19.620 1840.390 19.680 ;
        RECT 1538.310 19.480 1840.390 19.620 ;
        RECT 1538.310 19.420 1538.630 19.480 ;
        RECT 1840.070 19.420 1840.390 19.480 ;
      LAYER via ;
        RECT 1534.200 243.820 1534.460 244.080 ;
        RECT 1538.340 243.820 1538.600 244.080 ;
        RECT 1538.340 19.420 1538.600 19.680 ;
        RECT 1840.100 19.420 1840.360 19.680 ;
      LAYER met2 ;
        RECT 1534.150 260.000 1534.430 264.000 ;
        RECT 1534.260 244.110 1534.400 260.000 ;
        RECT 1534.200 243.790 1534.460 244.110 ;
        RECT 1538.340 243.790 1538.600 244.110 ;
        RECT 1538.400 19.710 1538.540 243.790 ;
        RECT 1538.340 19.390 1538.600 19.710 ;
        RECT 1840.100 19.390 1840.360 19.710 ;
        RECT 1840.160 2.400 1840.300 19.390 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
=======
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 1631.305 17.765 1632.395 17.935 ;
      LAYER mcon ;
        RECT 1632.225 17.765 1632.395 17.935 ;
      LAYER met1 ;
        RECT 1552.110 17.920 1552.430 17.980 ;
        RECT 1631.245 17.920 1631.535 17.965 ;
        RECT 1552.110 17.780 1631.535 17.920 ;
        RECT 1552.110 17.720 1552.430 17.780 ;
        RECT 1631.245 17.735 1631.535 17.780 ;
        RECT 1632.165 17.920 1632.455 17.965 ;
        RECT 1858.010 17.920 1858.330 17.980 ;
        RECT 1632.165 17.780 1858.330 17.920 ;
        RECT 1632.165 17.735 1632.455 17.780 ;
        RECT 1858.010 17.720 1858.330 17.780 ;
      LAYER via ;
        RECT 1552.140 17.720 1552.400 17.980 ;
        RECT 1858.040 17.720 1858.300 17.980 ;
      LAYER met2 ;
        RECT 1552.090 260.000 1552.370 264.000 ;
        RECT 1552.200 18.010 1552.340 260.000 ;
        RECT 1552.140 17.690 1552.400 18.010 ;
        RECT 1858.040 17.690 1858.300 18.010 ;
        RECT 1858.100 2.400 1858.240 17.690 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
=======
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1572.810 19.960 1573.130 20.020 ;
        RECT 1875.950 19.960 1876.270 20.020 ;
        RECT 1572.810 19.820 1876.270 19.960 ;
        RECT 1572.810 19.760 1573.130 19.820 ;
        RECT 1875.950 19.760 1876.270 19.820 ;
      LAYER via ;
        RECT 1572.840 19.760 1573.100 20.020 ;
        RECT 1875.980 19.760 1876.240 20.020 ;
      LAYER met2 ;
        RECT 1570.030 260.170 1570.310 264.000 ;
        RECT 1570.030 260.030 1573.040 260.170 ;
        RECT 1570.030 260.000 1570.310 260.030 ;
        RECT 1572.900 20.050 1573.040 260.030 ;
        RECT 1572.840 19.730 1573.100 20.050 ;
        RECT 1875.980 19.730 1876.240 20.050 ;
        RECT 1876.040 2.400 1876.180 19.730 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
=======
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 443.510 246.740 443.830 246.800 ;
        RECT 753.090 246.740 753.410 246.800 ;
        RECT 443.510 246.600 753.410 246.740 ;
        RECT 443.510 246.540 443.830 246.600 ;
        RECT 753.090 246.540 753.410 246.600 ;
      LAYER via ;
        RECT 443.540 246.540 443.800 246.800 ;
        RECT 753.120 246.540 753.380 246.800 ;
      LAYER met2 ;
        RECT 443.490 260.000 443.770 264.000 ;
        RECT 443.600 246.830 443.740 260.000 ;
        RECT 443.540 246.510 443.800 246.830 ;
        RECT 753.120 246.510 753.380 246.830 ;
        RECT 753.180 17.410 753.320 246.510 ;
        RECT 752.260 17.270 753.320 17.410 ;
        RECT 752.260 2.400 752.400 17.270 ;
        RECT 752.050 -4.800 752.610 2.400 ;
=======
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1587.990 241.640 1588.310 241.700 ;
        RECT 1593.510 241.640 1593.830 241.700 ;
        RECT 1587.990 241.500 1593.830 241.640 ;
        RECT 1587.990 241.440 1588.310 241.500 ;
        RECT 1593.510 241.440 1593.830 241.500 ;
        RECT 1593.510 16.560 1593.830 16.620 ;
        RECT 1893.890 16.560 1894.210 16.620 ;
        RECT 1593.510 16.420 1894.210 16.560 ;
        RECT 1593.510 16.360 1593.830 16.420 ;
        RECT 1893.890 16.360 1894.210 16.420 ;
      LAYER via ;
        RECT 1588.020 241.440 1588.280 241.700 ;
        RECT 1593.540 241.440 1593.800 241.700 ;
        RECT 1593.540 16.360 1593.800 16.620 ;
        RECT 1893.920 16.360 1894.180 16.620 ;
      LAYER met2 ;
        RECT 1587.970 260.000 1588.250 264.000 ;
        RECT 1588.080 241.730 1588.220 260.000 ;
        RECT 1588.020 241.410 1588.280 241.730 ;
        RECT 1593.540 241.410 1593.800 241.730 ;
        RECT 1593.600 16.650 1593.740 241.410 ;
        RECT 1593.540 16.330 1593.800 16.650 ;
        RECT 1893.920 16.330 1894.180 16.650 ;
        RECT 1893.980 2.400 1894.120 16.330 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
=======
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1911.370 18.260 1911.690 18.320 ;
        RECT 1631.780 18.120 1911.690 18.260 ;
        RECT 1607.310 17.580 1607.630 17.640 ;
        RECT 1631.780 17.580 1631.920 18.120 ;
        RECT 1911.370 18.060 1911.690 18.120 ;
        RECT 1607.310 17.440 1631.920 17.580 ;
        RECT 1607.310 17.380 1607.630 17.440 ;
      LAYER via ;
        RECT 1607.340 17.380 1607.600 17.640 ;
        RECT 1911.400 18.060 1911.660 18.320 ;
      LAYER met2 ;
        RECT 1605.450 260.170 1605.730 264.000 ;
        RECT 1605.450 260.030 1607.540 260.170 ;
        RECT 1605.450 260.000 1605.730 260.030 ;
        RECT 1607.400 17.670 1607.540 260.030 ;
        RECT 1911.400 18.030 1911.660 18.350 ;
        RECT 1607.340 17.350 1607.600 17.670 ;
        RECT 1911.460 17.410 1911.600 18.030 ;
        RECT 1911.460 17.270 1912.060 17.410 ;
        RECT 1911.920 2.400 1912.060 17.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
=======
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1623.410 244.020 1623.730 244.080 ;
        RECT 1628.010 244.020 1628.330 244.080 ;
        RECT 1623.410 243.880 1628.330 244.020 ;
        RECT 1623.410 243.820 1623.730 243.880 ;
        RECT 1628.010 243.820 1628.330 243.880 ;
        RECT 1628.010 16.220 1628.330 16.280 ;
        RECT 1929.310 16.220 1929.630 16.280 ;
        RECT 1628.010 16.080 1929.630 16.220 ;
        RECT 1628.010 16.020 1628.330 16.080 ;
        RECT 1929.310 16.020 1929.630 16.080 ;
      LAYER via ;
        RECT 1623.440 243.820 1623.700 244.080 ;
        RECT 1628.040 243.820 1628.300 244.080 ;
        RECT 1628.040 16.020 1628.300 16.280 ;
        RECT 1929.340 16.020 1929.600 16.280 ;
      LAYER met2 ;
        RECT 1623.390 260.000 1623.670 264.000 ;
        RECT 1623.500 244.110 1623.640 260.000 ;
        RECT 1623.440 243.790 1623.700 244.110 ;
        RECT 1628.040 243.790 1628.300 244.110 ;
        RECT 1628.100 16.310 1628.240 243.790 ;
        RECT 1628.040 15.990 1628.300 16.310 ;
        RECT 1929.340 15.990 1929.600 16.310 ;
        RECT 1929.400 2.400 1929.540 15.990 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
=======
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1641.810 17.580 1642.130 17.640 ;
        RECT 1947.250 17.580 1947.570 17.640 ;
        RECT 1641.810 17.440 1947.570 17.580 ;
        RECT 1641.810 17.380 1642.130 17.440 ;
        RECT 1947.250 17.380 1947.570 17.440 ;
      LAYER via ;
        RECT 1641.840 17.380 1642.100 17.640 ;
        RECT 1947.280 17.380 1947.540 17.640 ;
      LAYER met2 ;
        RECT 1641.330 260.170 1641.610 264.000 ;
        RECT 1641.330 260.030 1642.040 260.170 ;
        RECT 1641.330 260.000 1641.610 260.030 ;
        RECT 1641.900 17.670 1642.040 260.030 ;
        RECT 1641.840 17.350 1642.100 17.670 ;
        RECT 1947.280 17.350 1947.540 17.670 ;
        RECT 1947.340 2.400 1947.480 17.350 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
=======
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1662.510 15.880 1662.830 15.940 ;
        RECT 1965.190 15.880 1965.510 15.940 ;
        RECT 1662.510 15.740 1965.510 15.880 ;
        RECT 1662.510 15.680 1662.830 15.740 ;
        RECT 1965.190 15.680 1965.510 15.740 ;
      LAYER via ;
        RECT 1662.540 15.680 1662.800 15.940 ;
        RECT 1965.220 15.680 1965.480 15.940 ;
      LAYER met2 ;
        RECT 1659.270 260.170 1659.550 264.000 ;
        RECT 1659.270 260.030 1662.740 260.170 ;
        RECT 1659.270 260.000 1659.550 260.030 ;
        RECT 1662.600 15.970 1662.740 260.030 ;
        RECT 1662.540 15.650 1662.800 15.970 ;
        RECT 1965.220 15.650 1965.480 15.970 ;
        RECT 1965.280 2.400 1965.420 15.650 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
=======
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1677.230 244.020 1677.550 244.080 ;
        RECT 1683.210 244.020 1683.530 244.080 ;
        RECT 1677.230 243.880 1683.530 244.020 ;
        RECT 1677.230 243.820 1677.550 243.880 ;
        RECT 1683.210 243.820 1683.530 243.880 ;
        RECT 1683.210 16.900 1683.530 16.960 ;
        RECT 1983.130 16.900 1983.450 16.960 ;
        RECT 1683.210 16.760 1983.450 16.900 ;
        RECT 1683.210 16.700 1683.530 16.760 ;
        RECT 1983.130 16.700 1983.450 16.760 ;
      LAYER via ;
        RECT 1677.260 243.820 1677.520 244.080 ;
        RECT 1683.240 243.820 1683.500 244.080 ;
        RECT 1683.240 16.700 1683.500 16.960 ;
        RECT 1983.160 16.700 1983.420 16.960 ;
      LAYER met2 ;
        RECT 1677.210 260.000 1677.490 264.000 ;
        RECT 1677.320 244.110 1677.460 260.000 ;
        RECT 1677.260 243.790 1677.520 244.110 ;
        RECT 1683.240 243.790 1683.500 244.110 ;
        RECT 1683.300 16.990 1683.440 243.790 ;
        RECT 1683.240 16.670 1683.500 16.990 ;
        RECT 1983.160 16.670 1983.420 16.990 ;
        RECT 1983.220 2.400 1983.360 16.670 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
=======
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1695.150 260.170 1695.430 264.000 ;
        RECT 1695.150 260.030 1697.240 260.170 ;
        RECT 1695.150 260.000 1695.430 260.030 ;
        RECT 1697.100 16.845 1697.240 260.030 ;
        RECT 1697.030 16.475 1697.310 16.845 ;
        RECT 2001.090 16.475 2001.370 16.845 ;
        RECT 2001.160 2.400 2001.300 16.475 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
      LAYER via2 ;
        RECT 1697.030 16.520 1697.310 16.800 ;
        RECT 2001.090 16.520 2001.370 16.800 ;
      LAYER met3 ;
        RECT 1697.005 16.810 1697.335 16.825 ;
        RECT 2001.065 16.810 2001.395 16.825 ;
        RECT 1697.005 16.510 2001.395 16.810 ;
        RECT 1697.005 16.495 1697.335 16.510 ;
        RECT 2001.065 16.495 2001.395 16.510 ;
=======
        RECT 2000.950 -4.800 2001.510 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1713.110 244.020 1713.430 244.080 ;
        RECT 1717.710 244.020 1718.030 244.080 ;
        RECT 1713.110 243.880 1718.030 244.020 ;
        RECT 1713.110 243.820 1713.430 243.880 ;
        RECT 1717.710 243.820 1718.030 243.880 ;
        RECT 1717.710 15.540 1718.030 15.600 ;
        RECT 2018.550 15.540 2018.870 15.600 ;
        RECT 1717.710 15.400 2018.870 15.540 ;
        RECT 1717.710 15.340 1718.030 15.400 ;
        RECT 2018.550 15.340 2018.870 15.400 ;
      LAYER via ;
        RECT 1713.140 243.820 1713.400 244.080 ;
        RECT 1717.740 243.820 1718.000 244.080 ;
        RECT 1717.740 15.340 1718.000 15.600 ;
        RECT 2018.580 15.340 2018.840 15.600 ;
      LAYER met2 ;
        RECT 1713.090 260.000 1713.370 264.000 ;
        RECT 1713.200 244.110 1713.340 260.000 ;
        RECT 1713.140 243.790 1713.400 244.110 ;
        RECT 1717.740 243.790 1718.000 244.110 ;
        RECT 1717.800 15.630 1717.940 243.790 ;
        RECT 1717.740 15.310 1718.000 15.630 ;
        RECT 2018.580 15.310 2018.840 15.630 ;
        RECT 2018.640 2.400 2018.780 15.310 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
=======
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1730.590 245.380 1730.910 245.440 ;
        RECT 2036.030 245.380 2036.350 245.440 ;
        RECT 1730.590 245.240 2036.350 245.380 ;
        RECT 1730.590 245.180 1730.910 245.240 ;
        RECT 2036.030 245.180 2036.350 245.240 ;
      LAYER via ;
        RECT 1730.620 245.180 1730.880 245.440 ;
        RECT 2036.060 245.180 2036.320 245.440 ;
      LAYER met2 ;
        RECT 1730.570 260.000 1730.850 264.000 ;
        RECT 1730.680 245.470 1730.820 260.000 ;
        RECT 1730.620 245.150 1730.880 245.470 ;
        RECT 2036.060 245.150 2036.320 245.470 ;
        RECT 2036.120 17.410 2036.260 245.150 ;
        RECT 2036.120 17.270 2036.720 17.410 ;
        RECT 2036.580 2.400 2036.720 17.270 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
=======
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1752.210 20.300 1752.530 20.360 ;
        RECT 2054.430 20.300 2054.750 20.360 ;
        RECT 1752.210 20.160 2054.750 20.300 ;
        RECT 1752.210 20.100 1752.530 20.160 ;
        RECT 2054.430 20.100 2054.750 20.160 ;
      LAYER via ;
        RECT 1752.240 20.100 1752.500 20.360 ;
        RECT 2054.460 20.100 2054.720 20.360 ;
      LAYER met2 ;
        RECT 1748.510 260.170 1748.790 264.000 ;
        RECT 1748.510 260.030 1752.440 260.170 ;
        RECT 1748.510 260.000 1748.790 260.030 ;
        RECT 1752.300 20.390 1752.440 260.030 ;
        RECT 1752.240 20.070 1752.500 20.390 ;
        RECT 2054.460 20.070 2054.720 20.390 ;
        RECT 2054.520 2.400 2054.660 20.070 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
=======
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 461.430 260.170 461.710 264.000 ;
        RECT 461.430 260.030 462.140 260.170 ;
        RECT 461.430 260.000 461.710 260.030 ;
        RECT 462.000 16.845 462.140 260.030 ;
        RECT 461.930 16.475 462.210 16.845 ;
        RECT 769.670 16.475 769.950 16.845 ;
        RECT 769.740 2.400 769.880 16.475 ;
        RECT 769.530 -4.800 770.090 2.400 ;
      LAYER via2 ;
        RECT 461.930 16.520 462.210 16.800 ;
        RECT 769.670 16.520 769.950 16.800 ;
      LAYER met3 ;
        RECT 461.905 16.810 462.235 16.825 ;
        RECT 769.645 16.810 769.975 16.825 ;
        RECT 461.905 16.510 769.975 16.810 ;
        RECT 461.905 16.495 462.235 16.510 ;
        RECT 769.645 16.495 769.975 16.510 ;
=======
        RECT 769.530 -4.800 770.090 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1766.470 244.020 1766.790 244.080 ;
        RECT 1772.910 244.020 1773.230 244.080 ;
        RECT 1766.470 243.880 1773.230 244.020 ;
        RECT 1766.470 243.820 1766.790 243.880 ;
        RECT 1772.910 243.820 1773.230 243.880 ;
        RECT 1772.910 19.280 1773.230 19.340 ;
        RECT 2072.370 19.280 2072.690 19.340 ;
        RECT 1772.910 19.140 2072.690 19.280 ;
        RECT 1772.910 19.080 1773.230 19.140 ;
        RECT 2072.370 19.080 2072.690 19.140 ;
      LAYER via ;
        RECT 1766.500 243.820 1766.760 244.080 ;
        RECT 1772.940 243.820 1773.200 244.080 ;
        RECT 1772.940 19.080 1773.200 19.340 ;
        RECT 2072.400 19.080 2072.660 19.340 ;
      LAYER met2 ;
        RECT 1766.450 260.000 1766.730 264.000 ;
        RECT 1766.560 244.110 1766.700 260.000 ;
        RECT 1766.500 243.790 1766.760 244.110 ;
        RECT 1772.940 243.790 1773.200 244.110 ;
        RECT 1773.000 19.370 1773.140 243.790 ;
        RECT 1772.940 19.050 1773.200 19.370 ;
        RECT 2072.400 19.050 2072.660 19.370 ;
        RECT 2072.460 2.400 2072.600 19.050 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
=======
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1787.170 18.600 1787.490 18.660 ;
        RECT 2089.850 18.600 2090.170 18.660 ;
        RECT 1787.170 18.460 2090.170 18.600 ;
        RECT 1787.170 18.400 1787.490 18.460 ;
        RECT 2089.850 18.400 2090.170 18.460 ;
      LAYER via ;
        RECT 1787.200 18.400 1787.460 18.660 ;
        RECT 2089.880 18.400 2090.140 18.660 ;
      LAYER met2 ;
        RECT 1784.390 260.170 1784.670 264.000 ;
        RECT 1784.390 260.030 1786.940 260.170 ;
        RECT 1784.390 260.000 1784.670 260.030 ;
        RECT 1786.800 19.280 1786.940 260.030 ;
        RECT 1786.800 19.140 1787.400 19.280 ;
        RECT 1787.260 18.690 1787.400 19.140 ;
        RECT 1787.200 18.370 1787.460 18.690 ;
        RECT 2089.880 18.370 2090.140 18.690 ;
        RECT 2089.940 2.400 2090.080 18.370 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
=======
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1802.350 244.020 1802.670 244.080 ;
        RECT 1807.410 244.020 1807.730 244.080 ;
        RECT 1802.350 243.880 1807.730 244.020 ;
        RECT 1802.350 243.820 1802.670 243.880 ;
        RECT 1807.410 243.820 1807.730 243.880 ;
        RECT 1807.410 20.640 1807.730 20.700 ;
        RECT 2107.790 20.640 2108.110 20.700 ;
        RECT 1807.410 20.500 2108.110 20.640 ;
        RECT 1807.410 20.440 1807.730 20.500 ;
        RECT 2107.790 20.440 2108.110 20.500 ;
      LAYER via ;
        RECT 1802.380 243.820 1802.640 244.080 ;
        RECT 1807.440 243.820 1807.700 244.080 ;
        RECT 1807.440 20.440 1807.700 20.700 ;
        RECT 2107.820 20.440 2108.080 20.700 ;
      LAYER met2 ;
        RECT 1802.330 260.000 1802.610 264.000 ;
        RECT 1802.440 244.110 1802.580 260.000 ;
        RECT 1802.380 243.790 1802.640 244.110 ;
        RECT 1807.440 243.790 1807.700 244.110 ;
        RECT 1807.500 20.730 1807.640 243.790 ;
        RECT 1807.440 20.410 1807.700 20.730 ;
        RECT 2107.820 20.410 2108.080 20.730 ;
        RECT 2107.880 2.400 2108.020 20.410 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
=======
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1820.270 260.170 1820.550 264.000 ;
        RECT 1820.270 260.030 1821.440 260.170 ;
        RECT 1820.270 260.000 1820.550 260.030 ;
        RECT 1821.300 17.525 1821.440 260.030 ;
        RECT 1821.230 17.155 1821.510 17.525 ;
        RECT 2125.750 17.155 2126.030 17.525 ;
        RECT 2125.820 2.400 2125.960 17.155 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
      LAYER via2 ;
        RECT 1821.230 17.200 1821.510 17.480 ;
        RECT 2125.750 17.200 2126.030 17.480 ;
      LAYER met3 ;
        RECT 1821.205 17.490 1821.535 17.505 ;
        RECT 2125.725 17.490 2126.055 17.505 ;
        RECT 1821.205 17.190 2126.055 17.490 ;
        RECT 1821.205 17.175 1821.535 17.190 ;
        RECT 2125.725 17.175 2126.055 17.190 ;
=======
        RECT 2125.610 -4.800 2126.170 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 2139.605 241.485 2139.775 246.075 ;
        RECT 2139.605 144.925 2139.775 193.035 ;
        RECT 2139.605 48.365 2139.775 96.475 ;
      LAYER mcon ;
        RECT 2139.605 245.905 2139.775 246.075 ;
        RECT 2139.605 192.865 2139.775 193.035 ;
        RECT 2139.605 96.305 2139.775 96.475 ;
      LAYER met1 ;
        RECT 1838.230 246.060 1838.550 246.120 ;
        RECT 2139.545 246.060 2139.835 246.105 ;
        RECT 1838.230 245.920 2139.835 246.060 ;
        RECT 1838.230 245.860 1838.550 245.920 ;
        RECT 2139.545 245.875 2139.835 245.920 ;
        RECT 2139.530 241.640 2139.850 241.700 ;
        RECT 2139.335 241.500 2139.850 241.640 ;
        RECT 2139.530 241.440 2139.850 241.500 ;
        RECT 2139.530 193.020 2139.850 193.080 ;
        RECT 2139.335 192.880 2139.850 193.020 ;
        RECT 2139.530 192.820 2139.850 192.880 ;
        RECT 2139.530 145.080 2139.850 145.140 ;
        RECT 2139.335 144.940 2139.850 145.080 ;
        RECT 2139.530 144.880 2139.850 144.940 ;
        RECT 2139.530 96.460 2139.850 96.520 ;
        RECT 2139.335 96.320 2139.850 96.460 ;
        RECT 2139.530 96.260 2139.850 96.320 ;
        RECT 2139.530 48.520 2139.850 48.580 ;
        RECT 2139.335 48.380 2139.850 48.520 ;
        RECT 2139.530 48.320 2139.850 48.380 ;
        RECT 2139.530 14.180 2139.850 14.240 ;
        RECT 2139.530 14.040 2143.900 14.180 ;
        RECT 2139.530 13.980 2139.850 14.040 ;
        RECT 2143.760 13.900 2143.900 14.040 ;
        RECT 2143.670 13.640 2143.990 13.900 ;
      LAYER via ;
        RECT 1838.260 245.860 1838.520 246.120 ;
        RECT 2139.560 241.440 2139.820 241.700 ;
        RECT 2139.560 192.820 2139.820 193.080 ;
        RECT 2139.560 144.880 2139.820 145.140 ;
        RECT 2139.560 96.260 2139.820 96.520 ;
        RECT 2139.560 48.320 2139.820 48.580 ;
        RECT 2139.560 13.980 2139.820 14.240 ;
        RECT 2143.700 13.640 2143.960 13.900 ;
      LAYER met2 ;
        RECT 1838.210 260.000 1838.490 264.000 ;
        RECT 1838.320 246.150 1838.460 260.000 ;
        RECT 1838.260 245.830 1838.520 246.150 ;
        RECT 2139.560 241.410 2139.820 241.730 ;
        RECT 2139.620 193.110 2139.760 241.410 ;
        RECT 2139.560 192.790 2139.820 193.110 ;
        RECT 2139.560 144.850 2139.820 145.170 ;
        RECT 2139.620 96.550 2139.760 144.850 ;
        RECT 2139.560 96.230 2139.820 96.550 ;
        RECT 2139.560 48.290 2139.820 48.610 ;
        RECT 2139.620 14.270 2139.760 48.290 ;
        RECT 2139.560 13.950 2139.820 14.270 ;
        RECT 2143.700 13.610 2143.960 13.930 ;
        RECT 2143.760 2.400 2143.900 13.610 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
=======
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1855.710 17.240 1856.030 17.300 ;
        RECT 2161.610 17.240 2161.930 17.300 ;
        RECT 1855.710 17.100 2161.930 17.240 ;
        RECT 1855.710 17.040 1856.030 17.100 ;
        RECT 2161.610 17.040 2161.930 17.100 ;
      LAYER via ;
        RECT 1855.740 17.040 1856.000 17.300 ;
        RECT 2161.640 17.040 2161.900 17.300 ;
      LAYER met2 ;
        RECT 1855.690 260.000 1855.970 264.000 ;
        RECT 1855.800 17.330 1855.940 260.000 ;
        RECT 1855.740 17.010 1856.000 17.330 ;
        RECT 2161.640 17.010 2161.900 17.330 ;
        RECT 2161.700 2.400 2161.840 17.010 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
=======
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 2174.105 241.485 2174.275 246.415 ;
        RECT 2174.105 144.925 2174.275 193.035 ;
        RECT 2174.105 48.705 2174.275 96.475 ;
        RECT 2179.165 2.805 2179.335 48.195 ;
      LAYER mcon ;
        RECT 2174.105 246.245 2174.275 246.415 ;
        RECT 2174.105 192.865 2174.275 193.035 ;
        RECT 2174.105 96.305 2174.275 96.475 ;
        RECT 2179.165 48.025 2179.335 48.195 ;
      LAYER met1 ;
        RECT 1873.650 246.400 1873.970 246.460 ;
        RECT 2174.045 246.400 2174.335 246.445 ;
        RECT 1873.650 246.260 2174.335 246.400 ;
        RECT 1873.650 246.200 1873.970 246.260 ;
        RECT 2174.045 246.215 2174.335 246.260 ;
        RECT 2174.030 241.640 2174.350 241.700 ;
        RECT 2173.835 241.500 2174.350 241.640 ;
        RECT 2174.030 241.440 2174.350 241.500 ;
        RECT 2174.030 193.020 2174.350 193.080 ;
        RECT 2173.835 192.880 2174.350 193.020 ;
        RECT 2174.030 192.820 2174.350 192.880 ;
        RECT 2174.030 145.080 2174.350 145.140 ;
        RECT 2173.835 144.940 2174.350 145.080 ;
        RECT 2174.030 144.880 2174.350 144.940 ;
        RECT 2174.030 96.460 2174.350 96.520 ;
        RECT 2173.835 96.320 2174.350 96.460 ;
        RECT 2174.030 96.260 2174.350 96.320 ;
        RECT 2174.030 48.860 2174.350 48.920 ;
        RECT 2173.835 48.720 2174.350 48.860 ;
        RECT 2174.030 48.660 2174.350 48.720 ;
        RECT 2174.030 48.180 2174.350 48.240 ;
        RECT 2179.105 48.180 2179.395 48.225 ;
        RECT 2174.030 48.040 2179.395 48.180 ;
        RECT 2174.030 47.980 2174.350 48.040 ;
        RECT 2179.105 47.995 2179.395 48.040 ;
        RECT 2179.090 2.960 2179.410 3.020 ;
        RECT 2178.895 2.820 2179.410 2.960 ;
        RECT 2179.090 2.760 2179.410 2.820 ;
      LAYER via ;
        RECT 1873.680 246.200 1873.940 246.460 ;
        RECT 2174.060 241.440 2174.320 241.700 ;
        RECT 2174.060 192.820 2174.320 193.080 ;
        RECT 2174.060 144.880 2174.320 145.140 ;
        RECT 2174.060 96.260 2174.320 96.520 ;
        RECT 2174.060 48.660 2174.320 48.920 ;
        RECT 2174.060 47.980 2174.320 48.240 ;
        RECT 2179.120 2.760 2179.380 3.020 ;
      LAYER met2 ;
        RECT 1873.630 260.000 1873.910 264.000 ;
        RECT 1873.740 246.490 1873.880 260.000 ;
        RECT 1873.680 246.170 1873.940 246.490 ;
        RECT 2174.060 241.410 2174.320 241.730 ;
        RECT 2174.120 193.110 2174.260 241.410 ;
        RECT 2174.060 192.790 2174.320 193.110 ;
        RECT 2174.060 144.850 2174.320 145.170 ;
        RECT 2174.120 96.550 2174.260 144.850 ;
        RECT 2174.060 96.230 2174.320 96.550 ;
        RECT 2174.060 48.630 2174.320 48.950 ;
        RECT 2174.120 48.270 2174.260 48.630 ;
        RECT 2174.060 47.950 2174.320 48.270 ;
        RECT 2179.120 2.730 2179.380 3.050 ;
        RECT 2179.180 2.400 2179.320 2.730 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
=======
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1891.590 244.020 1891.910 244.080 ;
        RECT 1897.110 244.020 1897.430 244.080 ;
        RECT 1891.590 243.880 1897.430 244.020 ;
        RECT 1891.590 243.820 1891.910 243.880 ;
        RECT 1897.110 243.820 1897.430 243.880 ;
        RECT 1897.110 18.940 1897.430 19.000 ;
        RECT 2197.030 18.940 2197.350 19.000 ;
        RECT 1897.110 18.800 2197.350 18.940 ;
        RECT 1897.110 18.740 1897.430 18.800 ;
        RECT 2197.030 18.740 2197.350 18.800 ;
      LAYER via ;
        RECT 1891.620 243.820 1891.880 244.080 ;
        RECT 1897.140 243.820 1897.400 244.080 ;
        RECT 1897.140 18.740 1897.400 19.000 ;
        RECT 2197.060 18.740 2197.320 19.000 ;
      LAYER met2 ;
        RECT 1891.570 260.000 1891.850 264.000 ;
        RECT 1891.680 244.110 1891.820 260.000 ;
        RECT 1891.620 243.790 1891.880 244.110 ;
        RECT 1897.140 243.790 1897.400 244.110 ;
        RECT 1897.200 19.030 1897.340 243.790 ;
        RECT 1897.140 18.710 1897.400 19.030 ;
        RECT 2197.060 18.710 2197.320 19.030 ;
        RECT 2197.120 2.400 2197.260 18.710 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
=======
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1909.530 245.040 1909.850 245.100 ;
        RECT 2215.890 245.040 2216.210 245.100 ;
        RECT 1909.530 244.900 2216.210 245.040 ;
        RECT 1909.530 244.840 1909.850 244.900 ;
        RECT 2215.890 244.840 2216.210 244.900 ;
      LAYER via ;
        RECT 1909.560 244.840 1909.820 245.100 ;
        RECT 2215.920 244.840 2216.180 245.100 ;
      LAYER met2 ;
        RECT 1909.510 260.000 1909.790 264.000 ;
        RECT 1909.620 245.130 1909.760 260.000 ;
        RECT 1909.560 244.810 1909.820 245.130 ;
        RECT 2215.920 244.810 2216.180 245.130 ;
        RECT 2215.980 17.410 2216.120 244.810 ;
        RECT 2215.060 17.270 2216.120 17.410 ;
        RECT 2215.060 2.400 2215.200 17.270 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
=======
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1927.470 241.980 1927.790 242.040 ;
        RECT 1931.610 241.980 1931.930 242.040 ;
        RECT 1927.470 241.840 1931.930 241.980 ;
        RECT 1927.470 241.780 1927.790 241.840 ;
        RECT 1931.610 241.780 1931.930 241.840 ;
        RECT 2232.910 18.940 2233.230 19.000 ;
        RECT 2215.520 18.800 2233.230 18.940 ;
        RECT 1931.610 18.260 1931.930 18.320 ;
        RECT 2215.520 18.260 2215.660 18.800 ;
        RECT 2232.910 18.740 2233.230 18.800 ;
        RECT 1931.610 18.120 2215.660 18.260 ;
        RECT 1931.610 18.060 1931.930 18.120 ;
      LAYER via ;
        RECT 1927.500 241.780 1927.760 242.040 ;
        RECT 1931.640 241.780 1931.900 242.040 ;
        RECT 1931.640 18.060 1931.900 18.320 ;
        RECT 2232.940 18.740 2233.200 19.000 ;
      LAYER met2 ;
        RECT 1927.450 260.000 1927.730 264.000 ;
        RECT 1927.560 242.070 1927.700 260.000 ;
        RECT 1927.500 241.750 1927.760 242.070 ;
        RECT 1931.640 241.750 1931.900 242.070 ;
        RECT 1931.700 18.350 1931.840 241.750 ;
        RECT 2232.940 18.710 2233.200 19.030 ;
        RECT 1931.640 18.030 1931.900 18.350 ;
        RECT 2233.000 2.400 2233.140 18.710 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
=======
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 479.390 245.040 479.710 245.100 ;
        RECT 787.130 245.040 787.450 245.100 ;
        RECT 479.390 244.900 787.450 245.040 ;
        RECT 479.390 244.840 479.710 244.900 ;
        RECT 787.130 244.840 787.450 244.900 ;
      LAYER via ;
        RECT 479.420 244.840 479.680 245.100 ;
        RECT 787.160 244.840 787.420 245.100 ;
      LAYER met2 ;
        RECT 479.370 260.000 479.650 264.000 ;
        RECT 479.480 245.130 479.620 260.000 ;
        RECT 479.420 244.810 479.680 245.130 ;
        RECT 787.160 244.810 787.420 245.130 ;
        RECT 787.220 7.890 787.360 244.810 ;
        RECT 787.220 7.750 787.820 7.890 ;
        RECT 787.680 2.400 787.820 7.750 ;
        RECT 787.470 -4.800 788.030 2.400 ;
=======
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1945.410 245.720 1945.730 245.780 ;
        RECT 2249.930 245.720 2250.250 245.780 ;
        RECT 1945.410 245.580 2250.250 245.720 ;
        RECT 1945.410 245.520 1945.730 245.580 ;
        RECT 2249.930 245.520 2250.250 245.580 ;
      LAYER via ;
        RECT 1945.440 245.520 1945.700 245.780 ;
        RECT 2249.960 245.520 2250.220 245.780 ;
      LAYER met2 ;
        RECT 1945.390 260.000 1945.670 264.000 ;
        RECT 1945.500 245.810 1945.640 260.000 ;
        RECT 1945.440 245.490 1945.700 245.810 ;
        RECT 2249.960 245.490 2250.220 245.810 ;
        RECT 2250.020 16.730 2250.160 245.490 ;
        RECT 2250.020 16.590 2251.080 16.730 ;
        RECT 2250.940 2.400 2251.080 16.590 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
=======
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1966.110 19.620 1966.430 19.680 ;
        RECT 2268.330 19.620 2268.650 19.680 ;
        RECT 1966.110 19.480 2268.650 19.620 ;
        RECT 1966.110 19.420 1966.430 19.480 ;
        RECT 2268.330 19.420 2268.650 19.480 ;
      LAYER via ;
        RECT 1966.140 19.420 1966.400 19.680 ;
        RECT 2268.360 19.420 2268.620 19.680 ;
      LAYER met2 ;
        RECT 1963.330 260.170 1963.610 264.000 ;
        RECT 1963.330 260.030 1966.340 260.170 ;
        RECT 1963.330 260.000 1963.610 260.030 ;
        RECT 1966.200 19.710 1966.340 260.030 ;
        RECT 1966.140 19.390 1966.400 19.710 ;
        RECT 2268.360 19.390 2268.620 19.710 ;
        RECT 2268.420 2.400 2268.560 19.390 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
=======
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 1980.830 247.080 1981.150 247.140 ;
        RECT 2284.430 247.080 2284.750 247.140 ;
        RECT 1980.830 246.940 2284.750 247.080 ;
        RECT 1980.830 246.880 1981.150 246.940 ;
        RECT 2284.430 246.880 2284.750 246.940 ;
        RECT 2284.430 2.960 2284.750 3.020 ;
        RECT 2286.270 2.960 2286.590 3.020 ;
        RECT 2284.430 2.820 2286.590 2.960 ;
        RECT 2284.430 2.760 2284.750 2.820 ;
        RECT 2286.270 2.760 2286.590 2.820 ;
      LAYER via ;
        RECT 1980.860 246.880 1981.120 247.140 ;
        RECT 2284.460 246.880 2284.720 247.140 ;
        RECT 2284.460 2.760 2284.720 3.020 ;
        RECT 2286.300 2.760 2286.560 3.020 ;
      LAYER met2 ;
        RECT 1980.810 260.000 1981.090 264.000 ;
        RECT 1980.920 247.170 1981.060 260.000 ;
        RECT 1980.860 246.850 1981.120 247.170 ;
        RECT 2284.460 246.850 2284.720 247.170 ;
        RECT 2284.520 3.050 2284.660 246.850 ;
        RECT 2284.460 2.730 2284.720 3.050 ;
        RECT 2286.300 2.730 2286.560 3.050 ;
        RECT 2286.360 2.400 2286.500 2.730 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
=======
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2000.610 19.960 2000.930 20.020 ;
        RECT 2303.750 19.960 2304.070 20.020 ;
        RECT 2000.610 19.820 2304.070 19.960 ;
        RECT 2000.610 19.760 2000.930 19.820 ;
        RECT 2303.750 19.760 2304.070 19.820 ;
      LAYER via ;
        RECT 2000.640 19.760 2000.900 20.020 ;
        RECT 2303.780 19.760 2304.040 20.020 ;
      LAYER met2 ;
        RECT 1998.750 260.170 1999.030 264.000 ;
        RECT 1998.750 260.030 2000.840 260.170 ;
        RECT 1998.750 260.000 1999.030 260.030 ;
        RECT 2000.700 20.050 2000.840 260.030 ;
        RECT 2000.640 19.730 2000.900 20.050 ;
        RECT 2303.780 19.730 2304.040 20.050 ;
        RECT 2303.840 19.450 2303.980 19.730 ;
        RECT 2303.840 19.310 2304.440 19.450 ;
        RECT 2304.300 2.400 2304.440 19.310 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
=======
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2016.710 246.740 2017.030 246.800 ;
        RECT 2318.930 246.740 2319.250 246.800 ;
        RECT 2016.710 246.600 2319.250 246.740 ;
        RECT 2016.710 246.540 2017.030 246.600 ;
        RECT 2318.930 246.540 2319.250 246.600 ;
      LAYER via ;
        RECT 2016.740 246.540 2017.000 246.800 ;
        RECT 2318.960 246.540 2319.220 246.800 ;
      LAYER met2 ;
        RECT 2016.690 260.000 2016.970 264.000 ;
        RECT 2016.800 246.830 2016.940 260.000 ;
        RECT 2016.740 246.510 2017.000 246.830 ;
        RECT 2318.960 246.510 2319.220 246.830 ;
        RECT 2319.020 16.730 2319.160 246.510 ;
        RECT 2319.020 16.590 2322.380 16.730 ;
        RECT 2322.240 2.400 2322.380 16.590 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
=======
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 2034.630 260.170 2034.910 264.000 ;
        RECT 2034.630 260.030 2035.340 260.170 ;
        RECT 2034.630 260.000 2034.910 260.030 ;
        RECT 2035.200 16.845 2035.340 260.030 ;
        RECT 2035.130 16.475 2035.410 16.845 ;
        RECT 2339.650 16.475 2339.930 16.845 ;
        RECT 2339.720 2.400 2339.860 16.475 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
      LAYER via2 ;
        RECT 2035.130 16.520 2035.410 16.800 ;
        RECT 2339.650 16.520 2339.930 16.800 ;
      LAYER met3 ;
        RECT 2035.105 16.810 2035.435 16.825 ;
        RECT 2339.625 16.810 2339.955 16.825 ;
        RECT 2035.105 16.510 2339.955 16.810 ;
        RECT 2035.105 16.495 2035.435 16.510 ;
        RECT 2339.625 16.495 2339.955 16.510 ;
=======
        RECT 2339.510 -4.800 2340.070 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2055.810 20.300 2056.130 20.360 ;
        RECT 2357.570 20.300 2357.890 20.360 ;
        RECT 2055.810 20.160 2357.890 20.300 ;
        RECT 2055.810 20.100 2056.130 20.160 ;
        RECT 2357.570 20.100 2357.890 20.160 ;
      LAYER via ;
        RECT 2055.840 20.100 2056.100 20.360 ;
        RECT 2357.600 20.100 2357.860 20.360 ;
      LAYER met2 ;
        RECT 2052.570 260.170 2052.850 264.000 ;
        RECT 2052.570 260.030 2056.040 260.170 ;
        RECT 2052.570 260.000 2052.850 260.030 ;
        RECT 2055.900 20.390 2056.040 260.030 ;
        RECT 2055.840 20.070 2056.100 20.390 ;
        RECT 2357.600 20.070 2357.860 20.390 ;
        RECT 2357.660 2.400 2357.800 20.070 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
=======
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2070.530 244.020 2070.850 244.080 ;
        RECT 2076.510 244.020 2076.830 244.080 ;
        RECT 2070.530 243.880 2076.830 244.020 ;
        RECT 2070.530 243.820 2070.850 243.880 ;
        RECT 2076.510 243.820 2076.830 243.880 ;
        RECT 2076.510 19.280 2076.830 19.340 ;
        RECT 2375.510 19.280 2375.830 19.340 ;
        RECT 2076.510 19.140 2375.830 19.280 ;
        RECT 2076.510 19.080 2076.830 19.140 ;
        RECT 2375.510 19.080 2375.830 19.140 ;
      LAYER via ;
        RECT 2070.560 243.820 2070.820 244.080 ;
        RECT 2076.540 243.820 2076.800 244.080 ;
        RECT 2076.540 19.080 2076.800 19.340 ;
        RECT 2375.540 19.080 2375.800 19.340 ;
      LAYER met2 ;
        RECT 2070.510 260.000 2070.790 264.000 ;
        RECT 2070.620 244.110 2070.760 260.000 ;
        RECT 2070.560 243.790 2070.820 244.110 ;
        RECT 2076.540 243.790 2076.800 244.110 ;
        RECT 2076.600 19.370 2076.740 243.790 ;
        RECT 2076.540 19.050 2076.800 19.370 ;
        RECT 2375.540 19.050 2375.800 19.370 ;
        RECT 2375.600 2.400 2375.740 19.050 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
=======
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER li1 ;
        RECT 2214.585 18.445 2216.135 18.615 ;
      LAYER mcon ;
        RECT 2215.965 18.445 2216.135 18.615 ;
      LAYER met1 ;
        RECT 2090.310 18.600 2090.630 18.660 ;
        RECT 2214.525 18.600 2214.815 18.645 ;
        RECT 2090.310 18.460 2214.815 18.600 ;
        RECT 2090.310 18.400 2090.630 18.460 ;
        RECT 2214.525 18.415 2214.815 18.460 ;
        RECT 2215.905 18.600 2216.195 18.645 ;
        RECT 2393.450 18.600 2393.770 18.660 ;
        RECT 2215.905 18.460 2393.770 18.600 ;
        RECT 2215.905 18.415 2216.195 18.460 ;
        RECT 2393.450 18.400 2393.770 18.460 ;
      LAYER via ;
        RECT 2090.340 18.400 2090.600 18.660 ;
        RECT 2393.480 18.400 2393.740 18.660 ;
      LAYER met2 ;
        RECT 2088.450 260.170 2088.730 264.000 ;
        RECT 2088.450 260.030 2090.540 260.170 ;
        RECT 2088.450 260.000 2088.730 260.030 ;
        RECT 2090.400 18.690 2090.540 260.030 ;
        RECT 2090.340 18.370 2090.600 18.690 ;
        RECT 2393.480 18.370 2393.740 18.690 ;
        RECT 2393.540 2.400 2393.680 18.370 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
=======
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2105.950 244.020 2106.270 244.080 ;
        RECT 2111.010 244.020 2111.330 244.080 ;
        RECT 2105.950 243.880 2111.330 244.020 ;
        RECT 2105.950 243.820 2106.270 243.880 ;
        RECT 2111.010 243.820 2111.330 243.880 ;
        RECT 2111.010 17.920 2111.330 17.980 ;
        RECT 2411.390 17.920 2411.710 17.980 ;
        RECT 2111.010 17.780 2411.710 17.920 ;
        RECT 2111.010 17.720 2111.330 17.780 ;
        RECT 2411.390 17.720 2411.710 17.780 ;
      LAYER via ;
        RECT 2105.980 243.820 2106.240 244.080 ;
        RECT 2111.040 243.820 2111.300 244.080 ;
        RECT 2111.040 17.720 2111.300 17.980 ;
        RECT 2411.420 17.720 2411.680 17.980 ;
      LAYER met2 ;
        RECT 2105.930 260.000 2106.210 264.000 ;
        RECT 2106.040 244.110 2106.180 260.000 ;
        RECT 2105.980 243.790 2106.240 244.110 ;
        RECT 2111.040 243.790 2111.300 244.110 ;
        RECT 2111.100 18.010 2111.240 243.790 ;
        RECT 2111.040 17.690 2111.300 18.010 ;
        RECT 2411.420 17.690 2411.680 18.010 ;
        RECT 2411.480 2.400 2411.620 17.690 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
=======
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 497.330 244.020 497.650 244.080 ;
        RECT 503.310 244.020 503.630 244.080 ;
        RECT 497.330 243.880 503.630 244.020 ;
        RECT 497.330 243.820 497.650 243.880 ;
        RECT 503.310 243.820 503.630 243.880 ;
        RECT 503.310 15.880 503.630 15.940 ;
        RECT 805.530 15.880 805.850 15.940 ;
        RECT 503.310 15.740 805.850 15.880 ;
        RECT 503.310 15.680 503.630 15.740 ;
        RECT 805.530 15.680 805.850 15.740 ;
      LAYER via ;
        RECT 497.360 243.820 497.620 244.080 ;
        RECT 503.340 243.820 503.600 244.080 ;
        RECT 503.340 15.680 503.600 15.940 ;
        RECT 805.560 15.680 805.820 15.940 ;
      LAYER met2 ;
        RECT 497.310 260.000 497.590 264.000 ;
        RECT 497.420 244.110 497.560 260.000 ;
        RECT 497.360 243.790 497.620 244.110 ;
        RECT 503.340 243.790 503.600 244.110 ;
        RECT 503.400 15.970 503.540 243.790 ;
        RECT 503.340 15.650 503.600 15.970 ;
        RECT 805.560 15.650 805.820 15.970 ;
        RECT 805.620 2.400 805.760 15.650 ;
        RECT 805.410 -4.800 805.970 2.400 ;
=======
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 0.300 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 310.570 17.240 310.890 17.300 ;
        RECT 2.830 17.100 310.890 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 310.570 17.040 310.890 17.100 ;
      LAYER via ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 310.600 17.040 310.860 17.300 ;
      LAYER met2 ;
        RECT 312.850 260.170 313.130 264.000 ;
        RECT 310.660 260.030 313.130 260.170 ;
        RECT 310.660 17.330 310.800 260.030 ;
        RECT 312.850 260.000 313.130 260.030 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 310.600 17.010 310.860 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
=======
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met1 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 317.470 17.580 317.790 17.640 ;
        RECT 8.350 17.440 317.790 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 317.470 17.380 317.790 17.440 ;
      LAYER via ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 317.500 17.380 317.760 17.640 ;
      LAYER met2 ;
        RECT 318.370 260.170 318.650 264.000 ;
        RECT 317.560 260.030 318.650 260.170 ;
        RECT 317.560 17.670 317.700 260.030 ;
        RECT 318.370 260.000 318.650 260.030 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 317.500 17.350 317.760 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
=======
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 0.300 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 0.300 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 0.300 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 0.300 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 0.300 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 0.300 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 0.300 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 0.300 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 0.300 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 0.300 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 0.300 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 0.300 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 0.300 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 0.300 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 0.300 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 0.300 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 0.300 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 0.300 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 0.300 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 0.300 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 0.300 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 0.300 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 0.300 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 0.300 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 0.300 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 0.300 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 0.300 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 0.300 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 0.300 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 0.300 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 0.300 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 0.300 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 0.300 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 0.300 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 0.300 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 0.300 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 0.300 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 0.300 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 0.300 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 0.300 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 0.300 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 0.300 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 0.300 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 0.300 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 0.300 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 0.300 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 0.300 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 0.300 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 0.300 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 0.300 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 0.300 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 0.300 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 0.300 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 0.300 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 0.300 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 0.300 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 0.300 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 0.300 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 0.300 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 0.300 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 0.300 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 0.300 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 0.300 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 0.300 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 0.300 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 0.300 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 0.300 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 0.300 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 0.300 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 0.300 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 0.300 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 0.300 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 0.300 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 0.300 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 0.300 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 0.300 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 0.300 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 0.300 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 0.300 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 0.300 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 0.300 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 0.300 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 0.300 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 0.300 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 0.300 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 0.300 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 0.300 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 0.300 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 0.300 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 0.300 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 0.300 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 0.300 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 0.300 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 0.300 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 0.300 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 0.300 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 0.300 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 0.300 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 0.300 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 0.300 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 0.300 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 0.300 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 0.300 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 0.300 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.580 -14.220 -16.580 3533.900 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
<<<<<<< HEAD
        RECT 4.020 -9.420 7.020 3529.100 ;
        RECT 22.020 -19.020 25.020 3538.700 ;
        RECT 184.020 -9.420 187.020 3529.100 ;
        RECT 202.020 -19.020 205.020 3538.700 ;
        RECT 364.020 3260.000 367.020 3529.100 ;
        RECT 382.020 3260.000 385.020 3538.700 ;
        RECT 544.020 3260.000 547.020 3529.100 ;
        RECT 562.020 3260.000 565.020 3538.700 ;
        RECT 724.020 3260.000 727.020 3529.100 ;
        RECT 742.020 3260.000 745.020 3538.700 ;
        RECT 904.020 3260.000 907.020 3529.100 ;
        RECT 922.020 3260.000 925.020 3538.700 ;
        RECT 1084.020 3260.000 1087.020 3529.100 ;
        RECT 1102.020 3260.000 1105.020 3538.700 ;
        RECT 1264.020 3260.000 1267.020 3529.100 ;
        RECT 1282.020 3260.000 1285.020 3538.700 ;
        RECT 1444.020 3260.000 1447.020 3529.100 ;
        RECT 1462.020 3260.000 1465.020 3538.700 ;
        RECT 1624.020 3260.000 1627.020 3529.100 ;
        RECT 1642.020 3260.000 1645.020 3538.700 ;
        RECT 1804.020 3260.000 1807.020 3529.100 ;
        RECT 1822.020 3260.000 1825.020 3538.700 ;
        RECT 1984.020 3260.000 1987.020 3529.100 ;
        RECT 2002.020 3260.000 2005.020 3538.700 ;
        RECT 2164.020 3260.000 2167.020 3529.100 ;
        RECT 2182.020 3260.000 2185.020 3538.700 ;
        RECT 2344.020 3260.000 2347.020 3529.100 ;
        RECT 2362.020 3260.000 2365.020 3538.700 ;
        RECT 2524.020 3260.000 2527.020 3529.100 ;
        RECT 2542.020 3260.000 2545.020 3538.700 ;
        RECT 331.040 270.640 332.640 3246.800 ;
        RECT 364.020 -9.420 367.020 260.000 ;
        RECT 382.020 -19.020 385.020 260.000 ;
        RECT 544.020 -9.420 547.020 260.000 ;
        RECT 562.020 -19.020 565.020 260.000 ;
        RECT 724.020 -9.420 727.020 260.000 ;
        RECT 742.020 -19.020 745.020 260.000 ;
        RECT 904.020 -9.420 907.020 260.000 ;
        RECT 922.020 -19.020 925.020 260.000 ;
        RECT 1084.020 -9.420 1087.020 260.000 ;
        RECT 1102.020 -19.020 1105.020 260.000 ;
        RECT 1264.020 -9.420 1267.020 260.000 ;
        RECT 1282.020 -19.020 1285.020 260.000 ;
        RECT 1444.020 -9.420 1447.020 260.000 ;
        RECT 1462.020 -19.020 1465.020 260.000 ;
        RECT 1624.020 -9.420 1627.020 260.000 ;
        RECT 1642.020 -19.020 1645.020 260.000 ;
        RECT 1804.020 -9.420 1807.020 260.000 ;
        RECT 1822.020 -19.020 1825.020 260.000 ;
        RECT 1984.020 -9.420 1987.020 260.000 ;
        RECT 2002.020 -19.020 2005.020 260.000 ;
        RECT 2164.020 -9.420 2167.020 260.000 ;
        RECT 2182.020 -19.020 2185.020 260.000 ;
        RECT 2344.020 -9.420 2347.020 260.000 ;
        RECT 2362.020 -19.020 2365.020 260.000 ;
        RECT 2524.020 -9.420 2527.020 260.000 ;
        RECT 2542.020 -19.020 2545.020 260.000 ;
        RECT 2704.020 -9.420 2707.020 3529.100 ;
        RECT 2722.020 -19.020 2725.020 3538.700 ;
        RECT 2884.020 -9.420 2887.020 3529.100 ;
        RECT 2902.020 -19.020 2905.020 3538.700 ;
=======
        RECT 4.020 3519.700 7.020 3529.000 ;
        RECT 184.020 3519.700 187.020 3529.000 ;
        RECT 364.020 3519.700 367.020 3529.000 ;
        RECT 544.020 3519.700 547.020 3529.000 ;
        RECT 724.020 3519.700 727.020 3529.000 ;
        RECT 904.020 3519.700 907.020 3529.000 ;
        RECT 1084.020 3519.700 1087.020 3529.000 ;
        RECT 1264.020 3519.700 1267.020 3529.000 ;
        RECT 1444.020 3519.700 1447.020 3529.000 ;
        RECT 1624.020 3519.700 1627.020 3529.000 ;
        RECT 1804.020 3519.700 1807.020 3529.000 ;
        RECT 1984.020 3519.700 1987.020 3529.000 ;
        RECT 2164.020 3519.700 2167.020 3529.000 ;
        RECT 2344.020 3519.700 2347.020 3529.000 ;
        RECT 2524.020 3519.700 2527.020 3529.000 ;
        RECT 2704.020 3519.700 2707.020 3529.000 ;
        RECT 2884.020 3519.700 2887.020 3529.000 ;
        RECT 4.020 -9.320 7.020 0.300 ;
        RECT 184.020 -9.320 187.020 0.300 ;
        RECT 364.020 -9.320 367.020 0.300 ;
        RECT 544.020 -9.320 547.020 0.300 ;
        RECT 724.020 -9.320 727.020 0.300 ;
        RECT 904.020 -9.320 907.020 0.300 ;
        RECT 1084.020 -9.320 1087.020 0.300 ;
        RECT 1264.020 -9.320 1267.020 0.300 ;
        RECT 1444.020 -9.320 1447.020 0.300 ;
        RECT 1624.020 -9.320 1627.020 0.300 ;
        RECT 1804.020 -9.320 1807.020 0.300 ;
        RECT 1984.020 -9.320 1987.020 0.300 ;
        RECT 2164.020 -9.320 2167.020 0.300 ;
        RECT 2344.020 -9.320 2347.020 0.300 ;
        RECT 2524.020 -9.320 2527.020 0.300 ;
        RECT 2704.020 -9.320 2707.020 0.300 ;
        RECT 2884.020 -9.320 2887.020 0.300 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.200 -14.220 2939.200 3533.900 ;
      LAYER via4 ;
        RECT -18.670 3532.610 -17.490 3533.790 ;
        RECT -18.670 3531.010 -17.490 3532.190 ;
        RECT 22.930 3532.610 24.110 3533.790 ;
        RECT 22.930 3531.010 24.110 3532.190 ;
        RECT -18.670 3449.090 -17.490 3450.270 ;
        RECT -18.670 3447.490 -17.490 3448.670 ;
        RECT -18.670 3269.090 -17.490 3270.270 ;
        RECT -18.670 3267.490 -17.490 3268.670 ;
        RECT -18.670 3089.090 -17.490 3090.270 ;
        RECT -18.670 3087.490 -17.490 3088.670 ;
        RECT -18.670 2909.090 -17.490 2910.270 ;
        RECT -18.670 2907.490 -17.490 2908.670 ;
        RECT -18.670 2729.090 -17.490 2730.270 ;
        RECT -18.670 2727.490 -17.490 2728.670 ;
        RECT -18.670 2549.090 -17.490 2550.270 ;
        RECT -18.670 2547.490 -17.490 2548.670 ;
        RECT -18.670 2369.090 -17.490 2370.270 ;
        RECT -18.670 2367.490 -17.490 2368.670 ;
        RECT -18.670 2189.090 -17.490 2190.270 ;
        RECT -18.670 2187.490 -17.490 2188.670 ;
        RECT -18.670 2009.090 -17.490 2010.270 ;
        RECT -18.670 2007.490 -17.490 2008.670 ;
        RECT -18.670 1829.090 -17.490 1830.270 ;
        RECT -18.670 1827.490 -17.490 1828.670 ;
        RECT -18.670 1649.090 -17.490 1650.270 ;
        RECT -18.670 1647.490 -17.490 1648.670 ;
        RECT -18.670 1469.090 -17.490 1470.270 ;
        RECT -18.670 1467.490 -17.490 1468.670 ;
        RECT -18.670 1289.090 -17.490 1290.270 ;
        RECT -18.670 1287.490 -17.490 1288.670 ;
        RECT -18.670 1109.090 -17.490 1110.270 ;
        RECT -18.670 1107.490 -17.490 1108.670 ;
        RECT -18.670 929.090 -17.490 930.270 ;
        RECT -18.670 927.490 -17.490 928.670 ;
        RECT -18.670 749.090 -17.490 750.270 ;
        RECT -18.670 747.490 -17.490 748.670 ;
        RECT -18.670 569.090 -17.490 570.270 ;
        RECT -18.670 567.490 -17.490 568.670 ;
        RECT -18.670 389.090 -17.490 390.270 ;
        RECT -18.670 387.490 -17.490 388.670 ;
        RECT -18.670 209.090 -17.490 210.270 ;
        RECT -18.670 207.490 -17.490 208.670 ;
        RECT -18.670 29.090 -17.490 30.270 ;
        RECT -18.670 27.490 -17.490 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
<<<<<<< HEAD
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 202.930 3532.610 204.110 3533.790 ;
        RECT 202.930 3531.010 204.110 3532.190 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.670 -12.510 -17.490 -11.330 ;
        RECT -18.670 -14.110 -17.490 -12.930 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 382.930 3532.610 384.110 3533.790 ;
        RECT 382.930 3531.010 384.110 3532.190 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 562.930 3532.610 564.110 3533.790 ;
        RECT 562.930 3531.010 564.110 3532.190 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 742.930 3532.610 744.110 3533.790 ;
        RECT 742.930 3531.010 744.110 3532.190 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 922.930 3532.610 924.110 3533.790 ;
        RECT 922.930 3531.010 924.110 3532.190 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 1102.930 3532.610 1104.110 3533.790 ;
        RECT 1102.930 3531.010 1104.110 3532.190 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1282.930 3532.610 1284.110 3533.790 ;
        RECT 1282.930 3531.010 1284.110 3532.190 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1462.930 3532.610 1464.110 3533.790 ;
        RECT 1462.930 3531.010 1464.110 3532.190 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1642.930 3532.610 1644.110 3533.790 ;
        RECT 1642.930 3531.010 1644.110 3532.190 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1822.930 3532.610 1824.110 3533.790 ;
        RECT 1822.930 3531.010 1824.110 3532.190 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 2002.930 3532.610 2004.110 3533.790 ;
        RECT 2002.930 3531.010 2004.110 3532.190 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 2182.930 3532.610 2184.110 3533.790 ;
        RECT 2182.930 3531.010 2184.110 3532.190 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2362.930 3532.610 2364.110 3533.790 ;
        RECT 2362.930 3531.010 2364.110 3532.190 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2542.930 3532.610 2544.110 3533.790 ;
        RECT 2542.930 3531.010 2544.110 3532.190 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2722.930 3532.610 2724.110 3533.790 ;
        RECT 2722.930 3531.010 2724.110 3532.190 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 331.250 3089.090 332.430 3090.270 ;
        RECT 331.250 3087.490 332.430 3088.670 ;
        RECT 331.250 3071.090 332.430 3072.270 ;
        RECT 331.250 3069.490 332.430 3070.670 ;
        RECT 331.250 2909.090 332.430 2910.270 ;
        RECT 331.250 2907.490 332.430 2908.670 ;
        RECT 331.250 2891.090 332.430 2892.270 ;
        RECT 331.250 2889.490 332.430 2890.670 ;
        RECT 331.250 2729.090 332.430 2730.270 ;
        RECT 331.250 2727.490 332.430 2728.670 ;
        RECT 331.250 2711.090 332.430 2712.270 ;
        RECT 331.250 2709.490 332.430 2710.670 ;
        RECT 331.250 2549.090 332.430 2550.270 ;
        RECT 331.250 2547.490 332.430 2548.670 ;
        RECT 331.250 2531.090 332.430 2532.270 ;
        RECT 331.250 2529.490 332.430 2530.670 ;
        RECT 331.250 2369.090 332.430 2370.270 ;
        RECT 331.250 2367.490 332.430 2368.670 ;
        RECT 331.250 2351.090 332.430 2352.270 ;
        RECT 331.250 2349.490 332.430 2350.670 ;
        RECT 331.250 2189.090 332.430 2190.270 ;
        RECT 331.250 2187.490 332.430 2188.670 ;
        RECT 331.250 2171.090 332.430 2172.270 ;
        RECT 331.250 2169.490 332.430 2170.670 ;
        RECT 331.250 2009.090 332.430 2010.270 ;
        RECT 331.250 2007.490 332.430 2008.670 ;
        RECT 331.250 1991.090 332.430 1992.270 ;
        RECT 331.250 1989.490 332.430 1990.670 ;
        RECT 331.250 1829.090 332.430 1830.270 ;
        RECT 331.250 1827.490 332.430 1828.670 ;
        RECT 331.250 1811.090 332.430 1812.270 ;
        RECT 331.250 1809.490 332.430 1810.670 ;
        RECT 331.250 1649.090 332.430 1650.270 ;
        RECT 331.250 1647.490 332.430 1648.670 ;
        RECT 331.250 1631.090 332.430 1632.270 ;
        RECT 331.250 1629.490 332.430 1630.670 ;
        RECT 331.250 1469.090 332.430 1470.270 ;
        RECT 331.250 1467.490 332.430 1468.670 ;
        RECT 331.250 1451.090 332.430 1452.270 ;
        RECT 331.250 1449.490 332.430 1450.670 ;
        RECT 331.250 1289.090 332.430 1290.270 ;
        RECT 331.250 1287.490 332.430 1288.670 ;
        RECT 331.250 1271.090 332.430 1272.270 ;
        RECT 331.250 1269.490 332.430 1270.670 ;
        RECT 331.250 1109.090 332.430 1110.270 ;
        RECT 331.250 1107.490 332.430 1108.670 ;
        RECT 331.250 1091.090 332.430 1092.270 ;
        RECT 331.250 1089.490 332.430 1090.670 ;
        RECT 331.250 929.090 332.430 930.270 ;
        RECT 331.250 927.490 332.430 928.670 ;
        RECT 331.250 911.090 332.430 912.270 ;
        RECT 331.250 909.490 332.430 910.670 ;
        RECT 331.250 749.090 332.430 750.270 ;
        RECT 331.250 747.490 332.430 748.670 ;
        RECT 331.250 731.090 332.430 732.270 ;
        RECT 331.250 729.490 332.430 730.670 ;
        RECT 331.250 569.090 332.430 570.270 ;
        RECT 331.250 567.490 332.430 568.670 ;
        RECT 331.250 551.090 332.430 552.270 ;
        RECT 331.250 549.490 332.430 550.670 ;
        RECT 331.250 389.090 332.430 390.270 ;
        RECT 331.250 387.490 332.430 388.670 ;
        RECT 331.250 371.090 332.430 372.270 ;
        RECT 331.250 369.490 332.430 370.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 22.930 -12.510 24.110 -11.330 ;
        RECT 22.930 -14.110 24.110 -12.930 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 202.930 -12.510 204.110 -11.330 ;
        RECT 202.930 -14.110 204.110 -12.930 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 382.930 -12.510 384.110 -11.330 ;
        RECT 382.930 -14.110 384.110 -12.930 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 562.930 -12.510 564.110 -11.330 ;
        RECT 562.930 -14.110 564.110 -12.930 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 742.930 -12.510 744.110 -11.330 ;
        RECT 742.930 -14.110 744.110 -12.930 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 922.930 -12.510 924.110 -11.330 ;
        RECT 922.930 -14.110 924.110 -12.930 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1102.930 -12.510 1104.110 -11.330 ;
        RECT 1102.930 -14.110 1104.110 -12.930 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1282.930 -12.510 1284.110 -11.330 ;
        RECT 1282.930 -14.110 1284.110 -12.930 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1462.930 -12.510 1464.110 -11.330 ;
        RECT 1462.930 -14.110 1464.110 -12.930 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1642.930 -12.510 1644.110 -11.330 ;
        RECT 1642.930 -14.110 1644.110 -12.930 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 1822.930 -12.510 1824.110 -11.330 ;
        RECT 1822.930 -14.110 1824.110 -12.930 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2002.930 -12.510 2004.110 -11.330 ;
        RECT 2002.930 -14.110 2004.110 -12.930 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2182.930 -12.510 2184.110 -11.330 ;
        RECT 2182.930 -14.110 2184.110 -12.930 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2362.930 -12.510 2364.110 -11.330 ;
        RECT 2362.930 -14.110 2364.110 -12.930 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2902.930 3532.610 2904.110 3533.790 ;
        RECT 2902.930 3531.010 2904.110 3532.190 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2542.930 -12.510 2544.110 -11.330 ;
        RECT 2542.930 -14.110 2544.110 -12.930 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2937.110 3532.610 2938.290 3533.790 ;
        RECT 2937.110 3531.010 2938.290 3532.190 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2722.930 -12.510 2724.110 -11.330 ;
        RECT 2722.930 -14.110 2724.110 -12.930 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
=======
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT -9.070 3430.850 -7.890 3432.030 ;
        RECT -9.070 3429.250 -7.890 3430.430 ;
        RECT -9.070 3250.850 -7.890 3252.030 ;
        RECT -9.070 3249.250 -7.890 3250.430 ;
        RECT -9.070 3070.850 -7.890 3072.030 ;
        RECT -9.070 3069.250 -7.890 3070.430 ;
        RECT -9.070 2890.850 -7.890 2892.030 ;
        RECT -9.070 2889.250 -7.890 2890.430 ;
        RECT -9.070 2710.850 -7.890 2712.030 ;
        RECT -9.070 2709.250 -7.890 2710.430 ;
        RECT -9.070 2530.850 -7.890 2532.030 ;
        RECT -9.070 2529.250 -7.890 2530.430 ;
        RECT -9.070 2350.850 -7.890 2352.030 ;
        RECT -9.070 2349.250 -7.890 2350.430 ;
        RECT -9.070 2170.850 -7.890 2172.030 ;
        RECT -9.070 2169.250 -7.890 2170.430 ;
        RECT -9.070 1990.850 -7.890 1992.030 ;
        RECT -9.070 1989.250 -7.890 1990.430 ;
        RECT -9.070 1810.850 -7.890 1812.030 ;
        RECT -9.070 1809.250 -7.890 1810.430 ;
        RECT -9.070 1630.850 -7.890 1632.030 ;
        RECT -9.070 1629.250 -7.890 1630.430 ;
        RECT -9.070 1450.850 -7.890 1452.030 ;
        RECT -9.070 1449.250 -7.890 1450.430 ;
        RECT -9.070 1270.850 -7.890 1272.030 ;
        RECT -9.070 1269.250 -7.890 1270.430 ;
        RECT -9.070 1090.850 -7.890 1092.030 ;
        RECT -9.070 1089.250 -7.890 1090.430 ;
        RECT -9.070 910.850 -7.890 912.030 ;
        RECT -9.070 909.250 -7.890 910.430 ;
        RECT -9.070 730.850 -7.890 732.030 ;
        RECT -9.070 729.250 -7.890 730.430 ;
        RECT -9.070 550.850 -7.890 552.030 ;
        RECT -9.070 549.250 -7.890 550.430 ;
        RECT -9.070 370.850 -7.890 372.030 ;
        RECT -9.070 369.250 -7.890 370.430 ;
        RECT -9.070 190.850 -7.890 192.030 ;
        RECT -9.070 189.250 -7.890 190.430 ;
        RECT -9.070 10.850 -7.890 12.030 ;
        RECT -9.070 9.250 -7.890 10.430 ;
        RECT 2927.510 3430.850 2928.690 3432.030 ;
        RECT 2927.510 3429.250 2928.690 3430.430 ;
        RECT 2927.510 3250.850 2928.690 3252.030 ;
        RECT 2927.510 3249.250 2928.690 3250.430 ;
        RECT 2927.510 3070.850 2928.690 3072.030 ;
        RECT 2927.510 3069.250 2928.690 3070.430 ;
        RECT 2927.510 2890.850 2928.690 2892.030 ;
        RECT 2927.510 2889.250 2928.690 2890.430 ;
        RECT 2927.510 2710.850 2928.690 2712.030 ;
        RECT 2927.510 2709.250 2928.690 2710.430 ;
        RECT 2927.510 2530.850 2928.690 2532.030 ;
        RECT 2927.510 2529.250 2928.690 2530.430 ;
        RECT 2927.510 2350.850 2928.690 2352.030 ;
        RECT 2927.510 2349.250 2928.690 2350.430 ;
        RECT 2927.510 2170.850 2928.690 2172.030 ;
        RECT 2927.510 2169.250 2928.690 2170.430 ;
        RECT 2927.510 1990.850 2928.690 1992.030 ;
        RECT 2927.510 1989.250 2928.690 1990.430 ;
        RECT 2927.510 1810.850 2928.690 1812.030 ;
        RECT 2927.510 1809.250 2928.690 1810.430 ;
        RECT 2927.510 1630.850 2928.690 1632.030 ;
        RECT 2927.510 1629.250 2928.690 1630.430 ;
        RECT 2927.510 1450.850 2928.690 1452.030 ;
        RECT 2927.510 1449.250 2928.690 1450.430 ;
        RECT 2927.510 1270.850 2928.690 1272.030 ;
        RECT 2927.510 1269.250 2928.690 1270.430 ;
        RECT 2927.510 1090.850 2928.690 1092.030 ;
        RECT 2927.510 1089.250 2928.690 1090.430 ;
        RECT 2927.510 910.850 2928.690 912.030 ;
        RECT 2927.510 909.250 2928.690 910.430 ;
        RECT 2927.510 730.850 2928.690 732.030 ;
        RECT 2927.510 729.250 2928.690 730.430 ;
        RECT 2927.510 550.850 2928.690 552.030 ;
        RECT 2927.510 549.250 2928.690 550.430 ;
        RECT 2927.510 370.850 2928.690 372.030 ;
        RECT 2927.510 369.250 2928.690 370.430 ;
        RECT 2927.510 190.850 2928.690 192.030 ;
        RECT 2927.510 189.250 2928.690 190.430 ;
        RECT 2927.510 10.850 2928.690 12.030 ;
        RECT 2927.510 9.250 2928.690 10.430 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2937.110 3449.090 2938.290 3450.270 ;
        RECT 2937.110 3447.490 2938.290 3448.670 ;
        RECT 2937.110 3269.090 2938.290 3270.270 ;
        RECT 2937.110 3267.490 2938.290 3268.670 ;
        RECT 2937.110 3089.090 2938.290 3090.270 ;
        RECT 2937.110 3087.490 2938.290 3088.670 ;
        RECT 2937.110 2909.090 2938.290 2910.270 ;
        RECT 2937.110 2907.490 2938.290 2908.670 ;
        RECT 2937.110 2729.090 2938.290 2730.270 ;
        RECT 2937.110 2727.490 2938.290 2728.670 ;
        RECT 2937.110 2549.090 2938.290 2550.270 ;
        RECT 2937.110 2547.490 2938.290 2548.670 ;
        RECT 2937.110 2369.090 2938.290 2370.270 ;
        RECT 2937.110 2367.490 2938.290 2368.670 ;
        RECT 2937.110 2189.090 2938.290 2190.270 ;
        RECT 2937.110 2187.490 2938.290 2188.670 ;
        RECT 2937.110 2009.090 2938.290 2010.270 ;
        RECT 2937.110 2007.490 2938.290 2008.670 ;
        RECT 2937.110 1829.090 2938.290 1830.270 ;
        RECT 2937.110 1827.490 2938.290 1828.670 ;
        RECT 2937.110 1649.090 2938.290 1650.270 ;
        RECT 2937.110 1647.490 2938.290 1648.670 ;
        RECT 2937.110 1469.090 2938.290 1470.270 ;
        RECT 2937.110 1467.490 2938.290 1468.670 ;
        RECT 2937.110 1289.090 2938.290 1290.270 ;
        RECT 2937.110 1287.490 2938.290 1288.670 ;
        RECT 2937.110 1109.090 2938.290 1110.270 ;
        RECT 2937.110 1107.490 2938.290 1108.670 ;
        RECT 2937.110 929.090 2938.290 930.270 ;
        RECT 2937.110 927.490 2938.290 928.670 ;
        RECT 2937.110 749.090 2938.290 750.270 ;
        RECT 2937.110 747.490 2938.290 748.670 ;
        RECT 2937.110 569.090 2938.290 570.270 ;
        RECT 2937.110 567.490 2938.290 568.670 ;
        RECT 2937.110 389.090 2938.290 390.270 ;
        RECT 2937.110 387.490 2938.290 388.670 ;
        RECT 2937.110 209.090 2938.290 210.270 ;
        RECT 2937.110 207.490 2938.290 208.670 ;
        RECT 2937.110 29.090 2938.290 30.270 ;
        RECT 2937.110 27.490 2938.290 28.670 ;
        RECT 2902.930 -12.510 2904.110 -11.330 ;
        RECT 2902.930 -14.110 2904.110 -12.930 ;
        RECT 2937.110 -12.510 2938.290 -11.330 ;
        RECT 2937.110 -14.110 2938.290 -12.930 ;
      LAYER met5 ;
        RECT -19.580 3533.900 -16.580 3533.910 ;
        RECT 22.020 3533.900 25.020 3533.910 ;
        RECT 202.020 3533.900 205.020 3533.910 ;
        RECT 382.020 3533.900 385.020 3533.910 ;
        RECT 562.020 3533.900 565.020 3533.910 ;
        RECT 742.020 3533.900 745.020 3533.910 ;
        RECT 922.020 3533.900 925.020 3533.910 ;
        RECT 1102.020 3533.900 1105.020 3533.910 ;
        RECT 1282.020 3533.900 1285.020 3533.910 ;
        RECT 1462.020 3533.900 1465.020 3533.910 ;
        RECT 1642.020 3533.900 1645.020 3533.910 ;
        RECT 1822.020 3533.900 1825.020 3533.910 ;
        RECT 2002.020 3533.900 2005.020 3533.910 ;
        RECT 2182.020 3533.900 2185.020 3533.910 ;
        RECT 2362.020 3533.900 2365.020 3533.910 ;
        RECT 2542.020 3533.900 2545.020 3533.910 ;
        RECT 2722.020 3533.900 2725.020 3533.910 ;
        RECT 2902.020 3533.900 2905.020 3533.910 ;
        RECT 2936.200 3533.900 2939.200 3533.910 ;
        RECT -19.580 3530.900 2939.200 3533.900 ;
        RECT -19.580 3530.890 -16.580 3530.900 ;
        RECT 22.020 3530.890 25.020 3530.900 ;
        RECT 202.020 3530.890 205.020 3530.900 ;
        RECT 382.020 3530.890 385.020 3530.900 ;
        RECT 562.020 3530.890 565.020 3530.900 ;
        RECT 742.020 3530.890 745.020 3530.900 ;
        RECT 922.020 3530.890 925.020 3530.900 ;
        RECT 1102.020 3530.890 1105.020 3530.900 ;
        RECT 1282.020 3530.890 1285.020 3530.900 ;
        RECT 1462.020 3530.890 1465.020 3530.900 ;
        RECT 1642.020 3530.890 1645.020 3530.900 ;
        RECT 1822.020 3530.890 1825.020 3530.900 ;
        RECT 2002.020 3530.890 2005.020 3530.900 ;
        RECT 2182.020 3530.890 2185.020 3530.900 ;
        RECT 2362.020 3530.890 2365.020 3530.900 ;
        RECT 2542.020 3530.890 2545.020 3530.900 ;
        RECT 2722.020 3530.890 2725.020 3530.900 ;
        RECT 2902.020 3530.890 2905.020 3530.900 ;
        RECT 2936.200 3530.890 2939.200 3530.900 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
<<<<<<< HEAD
        RECT -19.580 3450.380 -16.580 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.200 3450.380 2939.200 3450.390 ;
        RECT -24.380 3447.380 2944.000 3450.380 ;
        RECT -19.580 3447.370 -16.580 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.200 3447.370 2939.200 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.780 3429.380 2934.400 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -19.580 3270.380 -16.580 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.200 3270.380 2939.200 3270.390 ;
        RECT -24.380 3267.380 2944.000 3270.380 ;
        RECT -19.580 3267.370 -16.580 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.200 3267.370 2939.200 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.780 3249.380 2934.400 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -19.580 3090.380 -16.580 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 331.040 3090.380 332.640 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.200 3090.380 2939.200 3090.390 ;
        RECT -24.380 3087.380 2944.000 3090.380 ;
        RECT -19.580 3087.370 -16.580 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 331.040 3087.370 332.640 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.200 3087.370 2939.200 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 331.040 3072.380 332.640 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.780 3069.380 2934.400 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 331.040 3069.370 332.640 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -19.580 2910.380 -16.580 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 331.040 2910.380 332.640 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.200 2910.380 2939.200 2910.390 ;
        RECT -24.380 2907.380 2944.000 2910.380 ;
        RECT -19.580 2907.370 -16.580 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 331.040 2907.370 332.640 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.200 2907.370 2939.200 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 331.040 2892.380 332.640 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.780 2889.380 2934.400 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 331.040 2889.370 332.640 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -19.580 2730.380 -16.580 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 331.040 2730.380 332.640 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.200 2730.380 2939.200 2730.390 ;
        RECT -24.380 2727.380 2944.000 2730.380 ;
        RECT -19.580 2727.370 -16.580 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 331.040 2727.370 332.640 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.200 2727.370 2939.200 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 331.040 2712.380 332.640 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.780 2709.380 2934.400 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 331.040 2709.370 332.640 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -19.580 2550.380 -16.580 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 331.040 2550.380 332.640 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.200 2550.380 2939.200 2550.390 ;
        RECT -24.380 2547.380 2944.000 2550.380 ;
        RECT -19.580 2547.370 -16.580 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 331.040 2547.370 332.640 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.200 2547.370 2939.200 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 331.040 2532.380 332.640 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.780 2529.380 2934.400 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 331.040 2529.370 332.640 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -19.580 2370.380 -16.580 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 331.040 2370.380 332.640 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.200 2370.380 2939.200 2370.390 ;
        RECT -24.380 2367.380 2944.000 2370.380 ;
        RECT -19.580 2367.370 -16.580 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 331.040 2367.370 332.640 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.200 2367.370 2939.200 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 331.040 2352.380 332.640 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.780 2349.380 2934.400 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 331.040 2349.370 332.640 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -19.580 2190.380 -16.580 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 331.040 2190.380 332.640 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.200 2190.380 2939.200 2190.390 ;
        RECT -24.380 2187.380 2944.000 2190.380 ;
        RECT -19.580 2187.370 -16.580 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 331.040 2187.370 332.640 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.200 2187.370 2939.200 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 331.040 2172.380 332.640 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.780 2169.380 2934.400 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 331.040 2169.370 332.640 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -19.580 2010.380 -16.580 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 331.040 2010.380 332.640 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.200 2010.380 2939.200 2010.390 ;
        RECT -24.380 2007.380 2944.000 2010.380 ;
        RECT -19.580 2007.370 -16.580 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 331.040 2007.370 332.640 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.200 2007.370 2939.200 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 331.040 1992.380 332.640 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.780 1989.380 2934.400 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 331.040 1989.370 332.640 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -19.580 1830.380 -16.580 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 331.040 1830.380 332.640 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.200 1830.380 2939.200 1830.390 ;
        RECT -24.380 1827.380 2944.000 1830.380 ;
        RECT -19.580 1827.370 -16.580 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 331.040 1827.370 332.640 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.200 1827.370 2939.200 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 331.040 1812.380 332.640 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.780 1809.380 2934.400 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 331.040 1809.370 332.640 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -19.580 1650.380 -16.580 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 331.040 1650.380 332.640 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.200 1650.380 2939.200 1650.390 ;
        RECT -24.380 1647.380 2944.000 1650.380 ;
        RECT -19.580 1647.370 -16.580 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 331.040 1647.370 332.640 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.200 1647.370 2939.200 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 331.040 1632.380 332.640 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.780 1629.380 2934.400 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 331.040 1629.370 332.640 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -19.580 1470.380 -16.580 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 331.040 1470.380 332.640 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.200 1470.380 2939.200 1470.390 ;
        RECT -24.380 1467.380 2944.000 1470.380 ;
        RECT -19.580 1467.370 -16.580 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 331.040 1467.370 332.640 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.200 1467.370 2939.200 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 331.040 1452.380 332.640 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.780 1449.380 2934.400 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 331.040 1449.370 332.640 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -19.580 1290.380 -16.580 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 331.040 1290.380 332.640 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.200 1290.380 2939.200 1290.390 ;
        RECT -24.380 1287.380 2944.000 1290.380 ;
        RECT -19.580 1287.370 -16.580 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 331.040 1287.370 332.640 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.200 1287.370 2939.200 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 331.040 1272.380 332.640 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.780 1269.380 2934.400 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 331.040 1269.370 332.640 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -19.580 1110.380 -16.580 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 331.040 1110.380 332.640 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.200 1110.380 2939.200 1110.390 ;
        RECT -24.380 1107.380 2944.000 1110.380 ;
        RECT -19.580 1107.370 -16.580 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 331.040 1107.370 332.640 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.200 1107.370 2939.200 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 331.040 1092.380 332.640 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.780 1089.380 2934.400 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 331.040 1089.370 332.640 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -19.580 930.380 -16.580 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 331.040 930.380 332.640 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.200 930.380 2939.200 930.390 ;
        RECT -24.380 927.380 2944.000 930.380 ;
        RECT -19.580 927.370 -16.580 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 331.040 927.370 332.640 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.200 927.370 2939.200 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 331.040 912.380 332.640 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.780 909.380 2934.400 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 331.040 909.370 332.640 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -19.580 750.380 -16.580 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 331.040 750.380 332.640 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.200 750.380 2939.200 750.390 ;
        RECT -24.380 747.380 2944.000 750.380 ;
        RECT -19.580 747.370 -16.580 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 331.040 747.370 332.640 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.200 747.370 2939.200 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 331.040 732.380 332.640 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.780 729.380 2934.400 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 331.040 729.370 332.640 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -19.580 570.380 -16.580 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 331.040 570.380 332.640 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.200 570.380 2939.200 570.390 ;
        RECT -24.380 567.380 2944.000 570.380 ;
        RECT -19.580 567.370 -16.580 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 331.040 567.370 332.640 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.200 567.370 2939.200 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 331.040 552.380 332.640 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.780 549.380 2934.400 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 331.040 549.370 332.640 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -19.580 390.380 -16.580 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 331.040 390.380 332.640 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.200 390.380 2939.200 390.390 ;
        RECT -24.380 387.380 2944.000 390.380 ;
        RECT -19.580 387.370 -16.580 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 331.040 387.370 332.640 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.200 387.370 2939.200 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 331.040 372.380 332.640 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.780 369.380 2934.400 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 331.040 369.370 332.640 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -19.580 210.380 -16.580 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.200 210.380 2939.200 210.390 ;
        RECT -24.380 207.380 2944.000 210.380 ;
        RECT -19.580 207.370 -16.580 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.200 207.370 2939.200 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.780 189.380 2934.400 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -19.580 30.380 -16.580 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.200 30.380 2939.200 30.390 ;
        RECT -24.380 27.380 2944.000 30.380 ;
        RECT -19.580 27.370 -16.580 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.200 27.370 2939.200 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.780 9.380 2934.400 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
=======
        RECT -9.980 3432.140 -6.980 3432.150 ;
        RECT 2926.600 3432.140 2929.600 3432.150 ;
        RECT -14.680 3429.140 0.300 3432.140 ;
        RECT 2919.700 3429.140 2934.300 3432.140 ;
        RECT -9.980 3429.130 -6.980 3429.140 ;
        RECT 2926.600 3429.130 2929.600 3429.140 ;
        RECT -9.980 3252.140 -6.980 3252.150 ;
        RECT 2926.600 3252.140 2929.600 3252.150 ;
        RECT -14.680 3249.140 0.300 3252.140 ;
        RECT 2919.700 3249.140 2934.300 3252.140 ;
        RECT -9.980 3249.130 -6.980 3249.140 ;
        RECT 2926.600 3249.130 2929.600 3249.140 ;
        RECT -9.980 3072.140 -6.980 3072.150 ;
        RECT 2926.600 3072.140 2929.600 3072.150 ;
        RECT -14.680 3069.140 0.300 3072.140 ;
        RECT 2919.700 3069.140 2934.300 3072.140 ;
        RECT -9.980 3069.130 -6.980 3069.140 ;
        RECT 2926.600 3069.130 2929.600 3069.140 ;
        RECT -9.980 2892.140 -6.980 2892.150 ;
        RECT 2926.600 2892.140 2929.600 2892.150 ;
        RECT -14.680 2889.140 0.300 2892.140 ;
        RECT 2919.700 2889.140 2934.300 2892.140 ;
        RECT -9.980 2889.130 -6.980 2889.140 ;
        RECT 2926.600 2889.130 2929.600 2889.140 ;
        RECT -9.980 2712.140 -6.980 2712.150 ;
        RECT 2926.600 2712.140 2929.600 2712.150 ;
        RECT -14.680 2709.140 0.300 2712.140 ;
        RECT 2919.700 2709.140 2934.300 2712.140 ;
        RECT -9.980 2709.130 -6.980 2709.140 ;
        RECT 2926.600 2709.130 2929.600 2709.140 ;
        RECT -9.980 2532.140 -6.980 2532.150 ;
        RECT 2926.600 2532.140 2929.600 2532.150 ;
        RECT -14.680 2529.140 0.300 2532.140 ;
        RECT 2919.700 2529.140 2934.300 2532.140 ;
        RECT -9.980 2529.130 -6.980 2529.140 ;
        RECT 2926.600 2529.130 2929.600 2529.140 ;
        RECT -9.980 2352.140 -6.980 2352.150 ;
        RECT 2926.600 2352.140 2929.600 2352.150 ;
        RECT -14.680 2349.140 0.300 2352.140 ;
        RECT 2919.700 2349.140 2934.300 2352.140 ;
        RECT -9.980 2349.130 -6.980 2349.140 ;
        RECT 2926.600 2349.130 2929.600 2349.140 ;
        RECT -9.980 2172.140 -6.980 2172.150 ;
        RECT 2926.600 2172.140 2929.600 2172.150 ;
        RECT -14.680 2169.140 0.300 2172.140 ;
        RECT 2919.700 2169.140 2934.300 2172.140 ;
        RECT -9.980 2169.130 -6.980 2169.140 ;
        RECT 2926.600 2169.130 2929.600 2169.140 ;
        RECT -9.980 1992.140 -6.980 1992.150 ;
        RECT 2926.600 1992.140 2929.600 1992.150 ;
        RECT -14.680 1989.140 0.300 1992.140 ;
        RECT 2919.700 1989.140 2934.300 1992.140 ;
        RECT -9.980 1989.130 -6.980 1989.140 ;
        RECT 2926.600 1989.130 2929.600 1989.140 ;
        RECT -9.980 1812.140 -6.980 1812.150 ;
        RECT 2926.600 1812.140 2929.600 1812.150 ;
        RECT -14.680 1809.140 0.300 1812.140 ;
        RECT 2919.700 1809.140 2934.300 1812.140 ;
        RECT -9.980 1809.130 -6.980 1809.140 ;
        RECT 2926.600 1809.130 2929.600 1809.140 ;
        RECT -9.980 1632.140 -6.980 1632.150 ;
        RECT 2926.600 1632.140 2929.600 1632.150 ;
        RECT -14.680 1629.140 0.300 1632.140 ;
        RECT 2919.700 1629.140 2934.300 1632.140 ;
        RECT -9.980 1629.130 -6.980 1629.140 ;
        RECT 2926.600 1629.130 2929.600 1629.140 ;
        RECT -9.980 1452.140 -6.980 1452.150 ;
        RECT 2926.600 1452.140 2929.600 1452.150 ;
        RECT -14.680 1449.140 0.300 1452.140 ;
        RECT 2919.700 1449.140 2934.300 1452.140 ;
        RECT -9.980 1449.130 -6.980 1449.140 ;
        RECT 2926.600 1449.130 2929.600 1449.140 ;
        RECT -9.980 1272.140 -6.980 1272.150 ;
        RECT 2926.600 1272.140 2929.600 1272.150 ;
        RECT -14.680 1269.140 0.300 1272.140 ;
        RECT 2919.700 1269.140 2934.300 1272.140 ;
        RECT -9.980 1269.130 -6.980 1269.140 ;
        RECT 2926.600 1269.130 2929.600 1269.140 ;
        RECT -9.980 1092.140 -6.980 1092.150 ;
        RECT 2926.600 1092.140 2929.600 1092.150 ;
        RECT -14.680 1089.140 0.300 1092.140 ;
        RECT 2919.700 1089.140 2934.300 1092.140 ;
        RECT -9.980 1089.130 -6.980 1089.140 ;
        RECT 2926.600 1089.130 2929.600 1089.140 ;
        RECT -9.980 912.140 -6.980 912.150 ;
        RECT 2926.600 912.140 2929.600 912.150 ;
        RECT -14.680 909.140 0.300 912.140 ;
        RECT 2919.700 909.140 2934.300 912.140 ;
        RECT -9.980 909.130 -6.980 909.140 ;
        RECT 2926.600 909.130 2929.600 909.140 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 2926.600 732.140 2929.600 732.150 ;
        RECT -14.680 729.140 0.300 732.140 ;
        RECT 2919.700 729.140 2934.300 732.140 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 2926.600 729.130 2929.600 729.140 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 2926.600 552.140 2929.600 552.150 ;
        RECT -14.680 549.140 0.300 552.140 ;
        RECT 2919.700 549.140 2934.300 552.140 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 2926.600 549.130 2929.600 549.140 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 2926.600 372.140 2929.600 372.150 ;
        RECT -14.680 369.140 0.300 372.140 ;
        RECT 2919.700 369.140 2934.300 372.140 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 2926.600 369.130 2929.600 369.140 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 2926.600 192.140 2929.600 192.150 ;
        RECT -14.680 189.140 0.300 192.140 ;
        RECT 2919.700 189.140 2934.300 192.140 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 2926.600 189.130 2929.600 189.140 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 2926.600 12.140 2929.600 12.150 ;
        RECT -14.680 9.140 0.300 12.140 ;
        RECT 2919.700 9.140 2934.300 12.140 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 2926.600 9.130 2929.600 9.140 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.580 -11.220 -16.580 -11.210 ;
        RECT 22.020 -11.220 25.020 -11.210 ;
        RECT 202.020 -11.220 205.020 -11.210 ;
        RECT 382.020 -11.220 385.020 -11.210 ;
        RECT 562.020 -11.220 565.020 -11.210 ;
        RECT 742.020 -11.220 745.020 -11.210 ;
        RECT 922.020 -11.220 925.020 -11.210 ;
        RECT 1102.020 -11.220 1105.020 -11.210 ;
        RECT 1282.020 -11.220 1285.020 -11.210 ;
        RECT 1462.020 -11.220 1465.020 -11.210 ;
        RECT 1642.020 -11.220 1645.020 -11.210 ;
        RECT 1822.020 -11.220 1825.020 -11.210 ;
        RECT 2002.020 -11.220 2005.020 -11.210 ;
        RECT 2182.020 -11.220 2185.020 -11.210 ;
        RECT 2362.020 -11.220 2365.020 -11.210 ;
        RECT 2542.020 -11.220 2545.020 -11.210 ;
        RECT 2722.020 -11.220 2725.020 -11.210 ;
        RECT 2902.020 -11.220 2905.020 -11.210 ;
        RECT 2936.200 -11.220 2939.200 -11.210 ;
        RECT -19.580 -14.220 2939.200 -11.220 ;
        RECT -19.580 -14.230 -16.580 -14.220 ;
        RECT 22.020 -14.230 25.020 -14.220 ;
        RECT 202.020 -14.230 205.020 -14.220 ;
        RECT 382.020 -14.230 385.020 -14.220 ;
        RECT 562.020 -14.230 565.020 -14.220 ;
        RECT 742.020 -14.230 745.020 -14.220 ;
        RECT 922.020 -14.230 925.020 -14.220 ;
        RECT 1102.020 -14.230 1105.020 -14.220 ;
        RECT 1282.020 -14.230 1285.020 -14.220 ;
        RECT 1462.020 -14.230 1465.020 -14.220 ;
        RECT 1642.020 -14.230 1645.020 -14.220 ;
        RECT 1822.020 -14.230 1825.020 -14.220 ;
        RECT 2002.020 -14.230 2005.020 -14.220 ;
        RECT 2182.020 -14.230 2185.020 -14.220 ;
        RECT 2362.020 -14.230 2365.020 -14.220 ;
        RECT 2542.020 -14.230 2545.020 -14.220 ;
        RECT 2722.020 -14.230 2725.020 -14.220 ;
        RECT 2902.020 -14.230 2905.020 -14.220 ;
        RECT 2936.200 -14.230 2939.200 -14.220 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
<<<<<<< HEAD
        RECT -24.380 -19.020 -21.380 3538.700 ;
        RECT -14.780 -9.420 -11.780 3529.100 ;
        RECT 94.020 -9.420 97.020 3529.100 ;
        RECT 112.020 -19.020 115.020 3538.700 ;
        RECT 274.020 -9.420 277.020 3529.100 ;
        RECT 292.020 -19.020 295.020 3538.700 ;
        RECT 454.020 3260.000 457.020 3529.100 ;
        RECT 472.020 3260.000 475.020 3538.700 ;
        RECT 634.020 3260.000 637.020 3529.100 ;
        RECT 652.020 3260.000 655.020 3538.700 ;
        RECT 814.020 3260.000 817.020 3529.100 ;
        RECT 832.020 3260.000 835.020 3538.700 ;
        RECT 994.020 3260.000 997.020 3529.100 ;
        RECT 1012.020 3260.000 1015.020 3538.700 ;
        RECT 1174.020 3260.000 1177.020 3529.100 ;
        RECT 1192.020 3260.000 1195.020 3538.700 ;
        RECT 1354.020 3260.000 1357.020 3529.100 ;
        RECT 1372.020 3260.000 1375.020 3538.700 ;
        RECT 1534.020 3260.000 1537.020 3529.100 ;
        RECT 1552.020 3260.000 1555.020 3538.700 ;
        RECT 1714.020 3260.000 1717.020 3529.100 ;
        RECT 1732.020 3260.000 1735.020 3538.700 ;
        RECT 1894.020 3260.000 1897.020 3529.100 ;
        RECT 1912.020 3260.000 1915.020 3538.700 ;
        RECT 2074.020 3260.000 2077.020 3529.100 ;
        RECT 2092.020 3260.000 2095.020 3538.700 ;
        RECT 2254.020 3260.000 2257.020 3529.100 ;
        RECT 2272.020 3260.000 2275.020 3538.700 ;
        RECT 2434.020 3260.000 2437.020 3529.100 ;
        RECT 2452.020 3260.000 2455.020 3538.700 ;
        RECT 407.840 270.640 409.440 3246.800 ;
        RECT 454.020 -9.420 457.020 260.000 ;
        RECT 472.020 -19.020 475.020 260.000 ;
        RECT 634.020 -9.420 637.020 260.000 ;
        RECT 652.020 -19.020 655.020 260.000 ;
        RECT 814.020 -9.420 817.020 260.000 ;
        RECT 832.020 -19.020 835.020 260.000 ;
        RECT 994.020 -9.420 997.020 260.000 ;
        RECT 1012.020 -19.020 1015.020 260.000 ;
        RECT 1174.020 -9.420 1177.020 260.000 ;
        RECT 1192.020 -19.020 1195.020 260.000 ;
        RECT 1354.020 -9.420 1357.020 260.000 ;
        RECT 1372.020 -19.020 1375.020 260.000 ;
        RECT 1534.020 -9.420 1537.020 260.000 ;
        RECT 1552.020 -19.020 1555.020 260.000 ;
        RECT 1714.020 -9.420 1717.020 260.000 ;
        RECT 1732.020 -19.020 1735.020 260.000 ;
        RECT 1894.020 -9.420 1897.020 260.000 ;
        RECT 1912.020 -19.020 1915.020 260.000 ;
        RECT 2074.020 -9.420 2077.020 260.000 ;
        RECT 2092.020 -19.020 2095.020 260.000 ;
        RECT 2254.020 -9.420 2257.020 260.000 ;
        RECT 2272.020 -19.020 2275.020 260.000 ;
        RECT 2434.020 -9.420 2437.020 260.000 ;
        RECT 2452.020 -19.020 2455.020 260.000 ;
        RECT 2614.020 -9.420 2617.020 3529.100 ;
        RECT 2632.020 -19.020 2635.020 3538.700 ;
        RECT 2794.020 -9.420 2797.020 3529.100 ;
        RECT 2812.020 -19.020 2815.020 3538.700 ;
        RECT 2931.400 -9.420 2934.400 3529.100 ;
        RECT 2941.000 -19.020 2944.000 3538.700 ;
      LAYER via4 ;
        RECT -23.470 3537.410 -22.290 3538.590 ;
        RECT -23.470 3535.810 -22.290 3536.990 ;
        RECT 112.930 3537.410 114.110 3538.590 ;
        RECT 112.930 3535.810 114.110 3536.990 ;
        RECT -23.470 3359.090 -22.290 3360.270 ;
        RECT -23.470 3357.490 -22.290 3358.670 ;
        RECT -23.470 3179.090 -22.290 3180.270 ;
        RECT -23.470 3177.490 -22.290 3178.670 ;
        RECT -23.470 2999.090 -22.290 3000.270 ;
        RECT -23.470 2997.490 -22.290 2998.670 ;
        RECT -23.470 2819.090 -22.290 2820.270 ;
        RECT -23.470 2817.490 -22.290 2818.670 ;
        RECT -23.470 2639.090 -22.290 2640.270 ;
        RECT -23.470 2637.490 -22.290 2638.670 ;
        RECT -23.470 2459.090 -22.290 2460.270 ;
        RECT -23.470 2457.490 -22.290 2458.670 ;
        RECT -23.470 2279.090 -22.290 2280.270 ;
        RECT -23.470 2277.490 -22.290 2278.670 ;
        RECT -23.470 2099.090 -22.290 2100.270 ;
        RECT -23.470 2097.490 -22.290 2098.670 ;
        RECT -23.470 1919.090 -22.290 1920.270 ;
        RECT -23.470 1917.490 -22.290 1918.670 ;
        RECT -23.470 1739.090 -22.290 1740.270 ;
        RECT -23.470 1737.490 -22.290 1738.670 ;
        RECT -23.470 1559.090 -22.290 1560.270 ;
        RECT -23.470 1557.490 -22.290 1558.670 ;
        RECT -23.470 1379.090 -22.290 1380.270 ;
        RECT -23.470 1377.490 -22.290 1378.670 ;
        RECT -23.470 1199.090 -22.290 1200.270 ;
        RECT -23.470 1197.490 -22.290 1198.670 ;
        RECT -23.470 1019.090 -22.290 1020.270 ;
        RECT -23.470 1017.490 -22.290 1018.670 ;
        RECT -23.470 839.090 -22.290 840.270 ;
        RECT -23.470 837.490 -22.290 838.670 ;
        RECT -23.470 659.090 -22.290 660.270 ;
        RECT -23.470 657.490 -22.290 658.670 ;
        RECT -23.470 479.090 -22.290 480.270 ;
        RECT -23.470 477.490 -22.290 478.670 ;
        RECT -23.470 299.090 -22.290 300.270 ;
        RECT -23.470 297.490 -22.290 298.670 ;
        RECT -23.470 119.090 -22.290 120.270 ;
        RECT -23.470 117.490 -22.290 118.670 ;
        RECT -13.870 3527.810 -12.690 3528.990 ;
        RECT -13.870 3526.210 -12.690 3527.390 ;
        RECT -13.870 3341.090 -12.690 3342.270 ;
        RECT -13.870 3339.490 -12.690 3340.670 ;
        RECT -13.870 3161.090 -12.690 3162.270 ;
        RECT -13.870 3159.490 -12.690 3160.670 ;
        RECT -13.870 2981.090 -12.690 2982.270 ;
        RECT -13.870 2979.490 -12.690 2980.670 ;
        RECT -13.870 2801.090 -12.690 2802.270 ;
        RECT -13.870 2799.490 -12.690 2800.670 ;
        RECT -13.870 2621.090 -12.690 2622.270 ;
        RECT -13.870 2619.490 -12.690 2620.670 ;
        RECT -13.870 2441.090 -12.690 2442.270 ;
        RECT -13.870 2439.490 -12.690 2440.670 ;
        RECT -13.870 2261.090 -12.690 2262.270 ;
        RECT -13.870 2259.490 -12.690 2260.670 ;
        RECT -13.870 2081.090 -12.690 2082.270 ;
        RECT -13.870 2079.490 -12.690 2080.670 ;
        RECT -13.870 1901.090 -12.690 1902.270 ;
        RECT -13.870 1899.490 -12.690 1900.670 ;
        RECT -13.870 1721.090 -12.690 1722.270 ;
        RECT -13.870 1719.490 -12.690 1720.670 ;
        RECT -13.870 1541.090 -12.690 1542.270 ;
        RECT -13.870 1539.490 -12.690 1540.670 ;
        RECT -13.870 1361.090 -12.690 1362.270 ;
        RECT -13.870 1359.490 -12.690 1360.670 ;
        RECT -13.870 1181.090 -12.690 1182.270 ;
        RECT -13.870 1179.490 -12.690 1180.670 ;
        RECT -13.870 1001.090 -12.690 1002.270 ;
        RECT -13.870 999.490 -12.690 1000.670 ;
        RECT -13.870 821.090 -12.690 822.270 ;
        RECT -13.870 819.490 -12.690 820.670 ;
        RECT -13.870 641.090 -12.690 642.270 ;
        RECT -13.870 639.490 -12.690 640.670 ;
        RECT -13.870 461.090 -12.690 462.270 ;
        RECT -13.870 459.490 -12.690 460.670 ;
        RECT -13.870 281.090 -12.690 282.270 ;
        RECT -13.870 279.490 -12.690 280.670 ;
        RECT -13.870 101.090 -12.690 102.270 ;
        RECT -13.870 99.490 -12.690 100.670 ;
        RECT -13.870 -7.710 -12.690 -6.530 ;
        RECT -13.870 -9.310 -12.690 -8.130 ;
        RECT 94.930 3527.810 96.110 3528.990 ;
        RECT 94.930 3526.210 96.110 3527.390 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.710 96.110 -6.530 ;
        RECT 94.930 -9.310 96.110 -8.130 ;
        RECT 292.930 3537.410 294.110 3538.590 ;
        RECT 292.930 3535.810 294.110 3536.990 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.470 -17.310 -22.290 -16.130 ;
        RECT -23.470 -18.910 -22.290 -17.730 ;
        RECT 274.930 3527.810 276.110 3528.990 ;
        RECT 274.930 3526.210 276.110 3527.390 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.710 276.110 -6.530 ;
        RECT 274.930 -9.310 276.110 -8.130 ;
        RECT 472.930 3537.410 474.110 3538.590 ;
        RECT 472.930 3535.810 474.110 3536.990 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 454.930 3527.810 456.110 3528.990 ;
        RECT 454.930 3526.210 456.110 3527.390 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 652.930 3537.410 654.110 3538.590 ;
        RECT 652.930 3535.810 654.110 3536.990 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 634.930 3527.810 636.110 3528.990 ;
        RECT 634.930 3526.210 636.110 3527.390 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 832.930 3537.410 834.110 3538.590 ;
        RECT 832.930 3535.810 834.110 3536.990 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 814.930 3527.810 816.110 3528.990 ;
        RECT 814.930 3526.210 816.110 3527.390 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 1012.930 3537.410 1014.110 3538.590 ;
        RECT 1012.930 3535.810 1014.110 3536.990 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 994.930 3527.810 996.110 3528.990 ;
        RECT 994.930 3526.210 996.110 3527.390 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1192.930 3537.410 1194.110 3538.590 ;
        RECT 1192.930 3535.810 1194.110 3536.990 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1174.930 3527.810 1176.110 3528.990 ;
        RECT 1174.930 3526.210 1176.110 3527.390 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1372.930 3537.410 1374.110 3538.590 ;
        RECT 1372.930 3535.810 1374.110 3536.990 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1354.930 3527.810 1356.110 3528.990 ;
        RECT 1354.930 3526.210 1356.110 3527.390 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1552.930 3537.410 1554.110 3538.590 ;
        RECT 1552.930 3535.810 1554.110 3536.990 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1534.930 3527.810 1536.110 3528.990 ;
        RECT 1534.930 3526.210 1536.110 3527.390 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1732.930 3537.410 1734.110 3538.590 ;
        RECT 1732.930 3535.810 1734.110 3536.990 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1714.930 3527.810 1716.110 3528.990 ;
        RECT 1714.930 3526.210 1716.110 3527.390 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1912.930 3537.410 1914.110 3538.590 ;
        RECT 1912.930 3535.810 1914.110 3536.990 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1894.930 3527.810 1896.110 3528.990 ;
        RECT 1894.930 3526.210 1896.110 3527.390 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 2092.930 3537.410 2094.110 3538.590 ;
        RECT 2092.930 3535.810 2094.110 3536.990 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 2074.930 3527.810 2076.110 3528.990 ;
        RECT 2074.930 3526.210 2076.110 3527.390 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2272.930 3537.410 2274.110 3538.590 ;
        RECT 2272.930 3535.810 2274.110 3536.990 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2254.930 3527.810 2256.110 3528.990 ;
        RECT 2254.930 3526.210 2256.110 3527.390 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2452.930 3537.410 2454.110 3538.590 ;
        RECT 2452.930 3535.810 2454.110 3536.990 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2434.930 3527.810 2436.110 3528.990 ;
        RECT 2434.930 3526.210 2436.110 3527.390 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2632.930 3537.410 2634.110 3538.590 ;
        RECT 2632.930 3535.810 2634.110 3536.990 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2614.930 3527.810 2616.110 3528.990 ;
        RECT 2614.930 3526.210 2616.110 3527.390 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 408.050 3179.090 409.230 3180.270 ;
        RECT 408.050 3177.490 409.230 3178.670 ;
        RECT 408.050 3161.090 409.230 3162.270 ;
        RECT 408.050 3159.490 409.230 3160.670 ;
        RECT 408.050 2999.090 409.230 3000.270 ;
        RECT 408.050 2997.490 409.230 2998.670 ;
        RECT 408.050 2981.090 409.230 2982.270 ;
        RECT 408.050 2979.490 409.230 2980.670 ;
        RECT 408.050 2819.090 409.230 2820.270 ;
        RECT 408.050 2817.490 409.230 2818.670 ;
        RECT 408.050 2801.090 409.230 2802.270 ;
        RECT 408.050 2799.490 409.230 2800.670 ;
        RECT 408.050 2639.090 409.230 2640.270 ;
        RECT 408.050 2637.490 409.230 2638.670 ;
        RECT 408.050 2621.090 409.230 2622.270 ;
        RECT 408.050 2619.490 409.230 2620.670 ;
        RECT 408.050 2459.090 409.230 2460.270 ;
        RECT 408.050 2457.490 409.230 2458.670 ;
        RECT 408.050 2441.090 409.230 2442.270 ;
        RECT 408.050 2439.490 409.230 2440.670 ;
        RECT 408.050 2279.090 409.230 2280.270 ;
        RECT 408.050 2277.490 409.230 2278.670 ;
        RECT 408.050 2261.090 409.230 2262.270 ;
        RECT 408.050 2259.490 409.230 2260.670 ;
        RECT 408.050 2099.090 409.230 2100.270 ;
        RECT 408.050 2097.490 409.230 2098.670 ;
        RECT 408.050 2081.090 409.230 2082.270 ;
        RECT 408.050 2079.490 409.230 2080.670 ;
        RECT 408.050 1919.090 409.230 1920.270 ;
        RECT 408.050 1917.490 409.230 1918.670 ;
        RECT 408.050 1901.090 409.230 1902.270 ;
        RECT 408.050 1899.490 409.230 1900.670 ;
        RECT 408.050 1739.090 409.230 1740.270 ;
        RECT 408.050 1737.490 409.230 1738.670 ;
        RECT 408.050 1721.090 409.230 1722.270 ;
        RECT 408.050 1719.490 409.230 1720.670 ;
        RECT 408.050 1559.090 409.230 1560.270 ;
        RECT 408.050 1557.490 409.230 1558.670 ;
        RECT 408.050 1541.090 409.230 1542.270 ;
        RECT 408.050 1539.490 409.230 1540.670 ;
        RECT 408.050 1379.090 409.230 1380.270 ;
        RECT 408.050 1377.490 409.230 1378.670 ;
        RECT 408.050 1361.090 409.230 1362.270 ;
        RECT 408.050 1359.490 409.230 1360.670 ;
        RECT 408.050 1199.090 409.230 1200.270 ;
        RECT 408.050 1197.490 409.230 1198.670 ;
        RECT 408.050 1181.090 409.230 1182.270 ;
        RECT 408.050 1179.490 409.230 1180.670 ;
        RECT 408.050 1019.090 409.230 1020.270 ;
        RECT 408.050 1017.490 409.230 1018.670 ;
        RECT 408.050 1001.090 409.230 1002.270 ;
        RECT 408.050 999.490 409.230 1000.670 ;
        RECT 408.050 839.090 409.230 840.270 ;
        RECT 408.050 837.490 409.230 838.670 ;
        RECT 408.050 821.090 409.230 822.270 ;
        RECT 408.050 819.490 409.230 820.670 ;
        RECT 408.050 659.090 409.230 660.270 ;
        RECT 408.050 657.490 409.230 658.670 ;
        RECT 408.050 641.090 409.230 642.270 ;
        RECT 408.050 639.490 409.230 640.670 ;
        RECT 408.050 479.090 409.230 480.270 ;
        RECT 408.050 477.490 409.230 478.670 ;
        RECT 408.050 461.090 409.230 462.270 ;
        RECT 408.050 459.490 409.230 460.670 ;
        RECT 408.050 299.090 409.230 300.270 ;
        RECT 408.050 297.490 409.230 298.670 ;
        RECT 408.050 281.090 409.230 282.270 ;
        RECT 408.050 279.490 409.230 280.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 112.930 -17.310 114.110 -16.130 ;
        RECT 112.930 -18.910 114.110 -17.730 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.710 456.110 -6.530 ;
        RECT 454.930 -9.310 456.110 -8.130 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 292.930 -17.310 294.110 -16.130 ;
        RECT 292.930 -18.910 294.110 -17.730 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.710 636.110 -6.530 ;
        RECT 634.930 -9.310 636.110 -8.130 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 472.930 -17.310 474.110 -16.130 ;
        RECT 472.930 -18.910 474.110 -17.730 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.710 816.110 -6.530 ;
        RECT 814.930 -9.310 816.110 -8.130 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 652.930 -17.310 654.110 -16.130 ;
        RECT 652.930 -18.910 654.110 -17.730 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.710 996.110 -6.530 ;
        RECT 994.930 -9.310 996.110 -8.130 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 832.930 -17.310 834.110 -16.130 ;
        RECT 832.930 -18.910 834.110 -17.730 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.710 1176.110 -6.530 ;
        RECT 1174.930 -9.310 1176.110 -8.130 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1012.930 -17.310 1014.110 -16.130 ;
        RECT 1012.930 -18.910 1014.110 -17.730 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.710 1356.110 -6.530 ;
        RECT 1354.930 -9.310 1356.110 -8.130 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1192.930 -17.310 1194.110 -16.130 ;
        RECT 1192.930 -18.910 1194.110 -17.730 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.710 1536.110 -6.530 ;
        RECT 1534.930 -9.310 1536.110 -8.130 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1372.930 -17.310 1374.110 -16.130 ;
        RECT 1372.930 -18.910 1374.110 -17.730 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.710 1716.110 -6.530 ;
        RECT 1714.930 -9.310 1716.110 -8.130 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1552.930 -17.310 1554.110 -16.130 ;
        RECT 1552.930 -18.910 1554.110 -17.730 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.710 1896.110 -6.530 ;
        RECT 1894.930 -9.310 1896.110 -8.130 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1732.930 -17.310 1734.110 -16.130 ;
        RECT 1732.930 -18.910 1734.110 -17.730 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.710 2076.110 -6.530 ;
        RECT 2074.930 -9.310 2076.110 -8.130 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 1912.930 -17.310 1914.110 -16.130 ;
        RECT 1912.930 -18.910 1914.110 -17.730 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.710 2256.110 -6.530 ;
        RECT 2254.930 -9.310 2256.110 -8.130 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2092.930 -17.310 2094.110 -16.130 ;
        RECT 2092.930 -18.910 2094.110 -17.730 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.710 2436.110 -6.530 ;
        RECT 2434.930 -9.310 2436.110 -8.130 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2272.930 -17.310 2274.110 -16.130 ;
        RECT 2272.930 -18.910 2274.110 -17.730 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.710 2616.110 -6.530 ;
        RECT 2614.930 -9.310 2616.110 -8.130 ;
        RECT 2812.930 3537.410 2814.110 3538.590 ;
        RECT 2812.930 3535.810 2814.110 3536.990 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2452.930 -17.310 2454.110 -16.130 ;
        RECT 2452.930 -18.910 2454.110 -17.730 ;
        RECT 2794.930 3527.810 2796.110 3528.990 ;
        RECT 2794.930 3526.210 2796.110 3527.390 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.710 2796.110 -6.530 ;
        RECT 2794.930 -9.310 2796.110 -8.130 ;
        RECT 2941.910 3537.410 2943.090 3538.590 ;
        RECT 2941.910 3535.810 2943.090 3536.990 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2632.930 -17.310 2634.110 -16.130 ;
        RECT 2632.930 -18.910 2634.110 -17.730 ;
        RECT 2932.310 3527.810 2933.490 3528.990 ;
        RECT 2932.310 3526.210 2933.490 3527.390 ;
        RECT 2932.310 3341.090 2933.490 3342.270 ;
        RECT 2932.310 3339.490 2933.490 3340.670 ;
        RECT 2932.310 3161.090 2933.490 3162.270 ;
        RECT 2932.310 3159.490 2933.490 3160.670 ;
        RECT 2932.310 2981.090 2933.490 2982.270 ;
        RECT 2932.310 2979.490 2933.490 2980.670 ;
        RECT 2932.310 2801.090 2933.490 2802.270 ;
        RECT 2932.310 2799.490 2933.490 2800.670 ;
        RECT 2932.310 2621.090 2933.490 2622.270 ;
        RECT 2932.310 2619.490 2933.490 2620.670 ;
        RECT 2932.310 2441.090 2933.490 2442.270 ;
        RECT 2932.310 2439.490 2933.490 2440.670 ;
        RECT 2932.310 2261.090 2933.490 2262.270 ;
        RECT 2932.310 2259.490 2933.490 2260.670 ;
        RECT 2932.310 2081.090 2933.490 2082.270 ;
        RECT 2932.310 2079.490 2933.490 2080.670 ;
        RECT 2932.310 1901.090 2933.490 1902.270 ;
        RECT 2932.310 1899.490 2933.490 1900.670 ;
        RECT 2932.310 1721.090 2933.490 1722.270 ;
        RECT 2932.310 1719.490 2933.490 1720.670 ;
        RECT 2932.310 1541.090 2933.490 1542.270 ;
        RECT 2932.310 1539.490 2933.490 1540.670 ;
        RECT 2932.310 1361.090 2933.490 1362.270 ;
        RECT 2932.310 1359.490 2933.490 1360.670 ;
        RECT 2932.310 1181.090 2933.490 1182.270 ;
        RECT 2932.310 1179.490 2933.490 1180.670 ;
        RECT 2932.310 1001.090 2933.490 1002.270 ;
        RECT 2932.310 999.490 2933.490 1000.670 ;
        RECT 2932.310 821.090 2933.490 822.270 ;
        RECT 2932.310 819.490 2933.490 820.670 ;
        RECT 2932.310 641.090 2933.490 642.270 ;
        RECT 2932.310 639.490 2933.490 640.670 ;
        RECT 2932.310 461.090 2933.490 462.270 ;
        RECT 2932.310 459.490 2933.490 460.670 ;
        RECT 2932.310 281.090 2933.490 282.270 ;
        RECT 2932.310 279.490 2933.490 280.670 ;
        RECT 2932.310 101.090 2933.490 102.270 ;
        RECT 2932.310 99.490 2933.490 100.670 ;
        RECT 2932.310 -7.710 2933.490 -6.530 ;
        RECT 2932.310 -9.310 2933.490 -8.130 ;
        RECT 2941.910 3359.090 2943.090 3360.270 ;
        RECT 2941.910 3357.490 2943.090 3358.670 ;
        RECT 2941.910 3179.090 2943.090 3180.270 ;
        RECT 2941.910 3177.490 2943.090 3178.670 ;
        RECT 2941.910 2999.090 2943.090 3000.270 ;
        RECT 2941.910 2997.490 2943.090 2998.670 ;
        RECT 2941.910 2819.090 2943.090 2820.270 ;
        RECT 2941.910 2817.490 2943.090 2818.670 ;
        RECT 2941.910 2639.090 2943.090 2640.270 ;
        RECT 2941.910 2637.490 2943.090 2638.670 ;
        RECT 2941.910 2459.090 2943.090 2460.270 ;
        RECT 2941.910 2457.490 2943.090 2458.670 ;
        RECT 2941.910 2279.090 2943.090 2280.270 ;
        RECT 2941.910 2277.490 2943.090 2278.670 ;
        RECT 2941.910 2099.090 2943.090 2100.270 ;
        RECT 2941.910 2097.490 2943.090 2098.670 ;
        RECT 2941.910 1919.090 2943.090 1920.270 ;
        RECT 2941.910 1917.490 2943.090 1918.670 ;
        RECT 2941.910 1739.090 2943.090 1740.270 ;
        RECT 2941.910 1737.490 2943.090 1738.670 ;
        RECT 2941.910 1559.090 2943.090 1560.270 ;
        RECT 2941.910 1557.490 2943.090 1558.670 ;
        RECT 2941.910 1379.090 2943.090 1380.270 ;
        RECT 2941.910 1377.490 2943.090 1378.670 ;
        RECT 2941.910 1199.090 2943.090 1200.270 ;
        RECT 2941.910 1197.490 2943.090 1198.670 ;
        RECT 2941.910 1019.090 2943.090 1020.270 ;
        RECT 2941.910 1017.490 2943.090 1018.670 ;
        RECT 2941.910 839.090 2943.090 840.270 ;
        RECT 2941.910 837.490 2943.090 838.670 ;
        RECT 2941.910 659.090 2943.090 660.270 ;
        RECT 2941.910 657.490 2943.090 658.670 ;
        RECT 2941.910 479.090 2943.090 480.270 ;
        RECT 2941.910 477.490 2943.090 478.670 ;
        RECT 2941.910 299.090 2943.090 300.270 ;
        RECT 2941.910 297.490 2943.090 298.670 ;
        RECT 2941.910 119.090 2943.090 120.270 ;
        RECT 2941.910 117.490 2943.090 118.670 ;
        RECT 2812.930 -17.310 2814.110 -16.130 ;
        RECT 2812.930 -18.910 2814.110 -17.730 ;
        RECT 2941.910 -17.310 2943.090 -16.130 ;
        RECT 2941.910 -18.910 2943.090 -17.730 ;
      LAYER met5 ;
        RECT -24.380 3538.700 -21.380 3538.710 ;
        RECT 112.020 3538.700 115.020 3538.710 ;
        RECT 292.020 3538.700 295.020 3538.710 ;
        RECT 472.020 3538.700 475.020 3538.710 ;
        RECT 652.020 3538.700 655.020 3538.710 ;
        RECT 832.020 3538.700 835.020 3538.710 ;
        RECT 1012.020 3538.700 1015.020 3538.710 ;
        RECT 1192.020 3538.700 1195.020 3538.710 ;
        RECT 1372.020 3538.700 1375.020 3538.710 ;
        RECT 1552.020 3538.700 1555.020 3538.710 ;
        RECT 1732.020 3538.700 1735.020 3538.710 ;
        RECT 1912.020 3538.700 1915.020 3538.710 ;
        RECT 2092.020 3538.700 2095.020 3538.710 ;
        RECT 2272.020 3538.700 2275.020 3538.710 ;
        RECT 2452.020 3538.700 2455.020 3538.710 ;
        RECT 2632.020 3538.700 2635.020 3538.710 ;
        RECT 2812.020 3538.700 2815.020 3538.710 ;
        RECT 2941.000 3538.700 2944.000 3538.710 ;
        RECT -24.380 3535.700 2944.000 3538.700 ;
        RECT -24.380 3535.690 -21.380 3535.700 ;
        RECT 112.020 3535.690 115.020 3535.700 ;
        RECT 292.020 3535.690 295.020 3535.700 ;
        RECT 472.020 3535.690 475.020 3535.700 ;
        RECT 652.020 3535.690 655.020 3535.700 ;
        RECT 832.020 3535.690 835.020 3535.700 ;
        RECT 1012.020 3535.690 1015.020 3535.700 ;
        RECT 1192.020 3535.690 1195.020 3535.700 ;
        RECT 1372.020 3535.690 1375.020 3535.700 ;
        RECT 1552.020 3535.690 1555.020 3535.700 ;
        RECT 1732.020 3535.690 1735.020 3535.700 ;
        RECT 1912.020 3535.690 1915.020 3535.700 ;
        RECT 2092.020 3535.690 2095.020 3535.700 ;
        RECT 2272.020 3535.690 2275.020 3535.700 ;
        RECT 2452.020 3535.690 2455.020 3535.700 ;
        RECT 2632.020 3535.690 2635.020 3535.700 ;
        RECT 2812.020 3535.690 2815.020 3535.700 ;
        RECT 2941.000 3535.690 2944.000 3535.700 ;
        RECT -14.780 3529.100 -11.780 3529.110 ;
        RECT 94.020 3529.100 97.020 3529.110 ;
        RECT 274.020 3529.100 277.020 3529.110 ;
        RECT 454.020 3529.100 457.020 3529.110 ;
        RECT 634.020 3529.100 637.020 3529.110 ;
        RECT 814.020 3529.100 817.020 3529.110 ;
        RECT 994.020 3529.100 997.020 3529.110 ;
        RECT 1174.020 3529.100 1177.020 3529.110 ;
        RECT 1354.020 3529.100 1357.020 3529.110 ;
        RECT 1534.020 3529.100 1537.020 3529.110 ;
        RECT 1714.020 3529.100 1717.020 3529.110 ;
        RECT 1894.020 3529.100 1897.020 3529.110 ;
        RECT 2074.020 3529.100 2077.020 3529.110 ;
        RECT 2254.020 3529.100 2257.020 3529.110 ;
        RECT 2434.020 3529.100 2437.020 3529.110 ;
        RECT 2614.020 3529.100 2617.020 3529.110 ;
        RECT 2794.020 3529.100 2797.020 3529.110 ;
        RECT 2931.400 3529.100 2934.400 3529.110 ;
        RECT -14.780 3526.100 2934.400 3529.100 ;
        RECT -14.780 3526.090 -11.780 3526.100 ;
        RECT 94.020 3526.090 97.020 3526.100 ;
        RECT 274.020 3526.090 277.020 3526.100 ;
        RECT 454.020 3526.090 457.020 3526.100 ;
        RECT 634.020 3526.090 637.020 3526.100 ;
        RECT 814.020 3526.090 817.020 3526.100 ;
        RECT 994.020 3526.090 997.020 3526.100 ;
        RECT 1174.020 3526.090 1177.020 3526.100 ;
        RECT 1354.020 3526.090 1357.020 3526.100 ;
        RECT 1534.020 3526.090 1537.020 3526.100 ;
        RECT 1714.020 3526.090 1717.020 3526.100 ;
        RECT 1894.020 3526.090 1897.020 3526.100 ;
        RECT 2074.020 3526.090 2077.020 3526.100 ;
        RECT 2254.020 3526.090 2257.020 3526.100 ;
        RECT 2434.020 3526.090 2437.020 3526.100 ;
        RECT 2614.020 3526.090 2617.020 3526.100 ;
        RECT 2794.020 3526.090 2797.020 3526.100 ;
        RECT 2931.400 3526.090 2934.400 3526.100 ;
        RECT -24.380 3360.380 -21.380 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2941.000 3360.380 2944.000 3360.390 ;
        RECT -24.380 3357.380 2944.000 3360.380 ;
        RECT -24.380 3357.370 -21.380 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2941.000 3357.370 2944.000 3357.380 ;
        RECT -14.780 3342.380 -11.780 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.400 3342.380 2934.400 3342.390 ;
        RECT -14.780 3339.380 2934.400 3342.380 ;
        RECT -14.780 3339.370 -11.780 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.400 3339.370 2934.400 3339.380 ;
        RECT -24.380 3180.380 -21.380 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 407.840 3180.380 409.440 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2941.000 3180.380 2944.000 3180.390 ;
        RECT -24.380 3177.380 2944.000 3180.380 ;
        RECT -24.380 3177.370 -21.380 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 407.840 3177.370 409.440 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2941.000 3177.370 2944.000 3177.380 ;
        RECT -14.780 3162.380 -11.780 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 407.840 3162.380 409.440 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.400 3162.380 2934.400 3162.390 ;
        RECT -14.780 3159.380 2934.400 3162.380 ;
        RECT -14.780 3159.370 -11.780 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 407.840 3159.370 409.440 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.400 3159.370 2934.400 3159.380 ;
        RECT -24.380 3000.380 -21.380 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 407.840 3000.380 409.440 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2941.000 3000.380 2944.000 3000.390 ;
        RECT -24.380 2997.380 2944.000 3000.380 ;
        RECT -24.380 2997.370 -21.380 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 407.840 2997.370 409.440 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2941.000 2997.370 2944.000 2997.380 ;
        RECT -14.780 2982.380 -11.780 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 407.840 2982.380 409.440 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.400 2982.380 2934.400 2982.390 ;
        RECT -14.780 2979.380 2934.400 2982.380 ;
        RECT -14.780 2979.370 -11.780 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 407.840 2979.370 409.440 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.400 2979.370 2934.400 2979.380 ;
        RECT -24.380 2820.380 -21.380 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 407.840 2820.380 409.440 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2941.000 2820.380 2944.000 2820.390 ;
        RECT -24.380 2817.380 2944.000 2820.380 ;
        RECT -24.380 2817.370 -21.380 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 407.840 2817.370 409.440 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2941.000 2817.370 2944.000 2817.380 ;
        RECT -14.780 2802.380 -11.780 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 407.840 2802.380 409.440 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.400 2802.380 2934.400 2802.390 ;
        RECT -14.780 2799.380 2934.400 2802.380 ;
        RECT -14.780 2799.370 -11.780 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 407.840 2799.370 409.440 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.400 2799.370 2934.400 2799.380 ;
        RECT -24.380 2640.380 -21.380 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 407.840 2640.380 409.440 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2941.000 2640.380 2944.000 2640.390 ;
        RECT -24.380 2637.380 2944.000 2640.380 ;
        RECT -24.380 2637.370 -21.380 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 407.840 2637.370 409.440 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2941.000 2637.370 2944.000 2637.380 ;
        RECT -14.780 2622.380 -11.780 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 407.840 2622.380 409.440 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.400 2622.380 2934.400 2622.390 ;
        RECT -14.780 2619.380 2934.400 2622.380 ;
        RECT -14.780 2619.370 -11.780 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 407.840 2619.370 409.440 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.400 2619.370 2934.400 2619.380 ;
        RECT -24.380 2460.380 -21.380 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 407.840 2460.380 409.440 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2941.000 2460.380 2944.000 2460.390 ;
        RECT -24.380 2457.380 2944.000 2460.380 ;
        RECT -24.380 2457.370 -21.380 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 407.840 2457.370 409.440 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2941.000 2457.370 2944.000 2457.380 ;
        RECT -14.780 2442.380 -11.780 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 407.840 2442.380 409.440 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.400 2442.380 2934.400 2442.390 ;
        RECT -14.780 2439.380 2934.400 2442.380 ;
        RECT -14.780 2439.370 -11.780 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 407.840 2439.370 409.440 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.400 2439.370 2934.400 2439.380 ;
        RECT -24.380 2280.380 -21.380 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 407.840 2280.380 409.440 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2941.000 2280.380 2944.000 2280.390 ;
        RECT -24.380 2277.380 2944.000 2280.380 ;
        RECT -24.380 2277.370 -21.380 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 407.840 2277.370 409.440 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2941.000 2277.370 2944.000 2277.380 ;
        RECT -14.780 2262.380 -11.780 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 407.840 2262.380 409.440 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.400 2262.380 2934.400 2262.390 ;
        RECT -14.780 2259.380 2934.400 2262.380 ;
        RECT -14.780 2259.370 -11.780 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 407.840 2259.370 409.440 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.400 2259.370 2934.400 2259.380 ;
        RECT -24.380 2100.380 -21.380 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 407.840 2100.380 409.440 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2941.000 2100.380 2944.000 2100.390 ;
        RECT -24.380 2097.380 2944.000 2100.380 ;
        RECT -24.380 2097.370 -21.380 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 407.840 2097.370 409.440 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2941.000 2097.370 2944.000 2097.380 ;
        RECT -14.780 2082.380 -11.780 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 407.840 2082.380 409.440 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.400 2082.380 2934.400 2082.390 ;
        RECT -14.780 2079.380 2934.400 2082.380 ;
        RECT -14.780 2079.370 -11.780 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 407.840 2079.370 409.440 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.400 2079.370 2934.400 2079.380 ;
        RECT -24.380 1920.380 -21.380 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 407.840 1920.380 409.440 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2941.000 1920.380 2944.000 1920.390 ;
        RECT -24.380 1917.380 2944.000 1920.380 ;
        RECT -24.380 1917.370 -21.380 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 407.840 1917.370 409.440 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2941.000 1917.370 2944.000 1917.380 ;
        RECT -14.780 1902.380 -11.780 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 407.840 1902.380 409.440 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.400 1902.380 2934.400 1902.390 ;
        RECT -14.780 1899.380 2934.400 1902.380 ;
        RECT -14.780 1899.370 -11.780 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 407.840 1899.370 409.440 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.400 1899.370 2934.400 1899.380 ;
        RECT -24.380 1740.380 -21.380 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 407.840 1740.380 409.440 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2941.000 1740.380 2944.000 1740.390 ;
        RECT -24.380 1737.380 2944.000 1740.380 ;
        RECT -24.380 1737.370 -21.380 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 407.840 1737.370 409.440 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2941.000 1737.370 2944.000 1737.380 ;
        RECT -14.780 1722.380 -11.780 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 407.840 1722.380 409.440 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.400 1722.380 2934.400 1722.390 ;
        RECT -14.780 1719.380 2934.400 1722.380 ;
        RECT -14.780 1719.370 -11.780 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 407.840 1719.370 409.440 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.400 1719.370 2934.400 1719.380 ;
        RECT -24.380 1560.380 -21.380 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 407.840 1560.380 409.440 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2941.000 1560.380 2944.000 1560.390 ;
        RECT -24.380 1557.380 2944.000 1560.380 ;
        RECT -24.380 1557.370 -21.380 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 407.840 1557.370 409.440 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2941.000 1557.370 2944.000 1557.380 ;
        RECT -14.780 1542.380 -11.780 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 407.840 1542.380 409.440 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.400 1542.380 2934.400 1542.390 ;
        RECT -14.780 1539.380 2934.400 1542.380 ;
        RECT -14.780 1539.370 -11.780 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 407.840 1539.370 409.440 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.400 1539.370 2934.400 1539.380 ;
        RECT -24.380 1380.380 -21.380 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 407.840 1380.380 409.440 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2941.000 1380.380 2944.000 1380.390 ;
        RECT -24.380 1377.380 2944.000 1380.380 ;
        RECT -24.380 1377.370 -21.380 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 407.840 1377.370 409.440 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2941.000 1377.370 2944.000 1377.380 ;
        RECT -14.780 1362.380 -11.780 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 407.840 1362.380 409.440 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.400 1362.380 2934.400 1362.390 ;
        RECT -14.780 1359.380 2934.400 1362.380 ;
        RECT -14.780 1359.370 -11.780 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 407.840 1359.370 409.440 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.400 1359.370 2934.400 1359.380 ;
        RECT -24.380 1200.380 -21.380 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 407.840 1200.380 409.440 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2941.000 1200.380 2944.000 1200.390 ;
        RECT -24.380 1197.380 2944.000 1200.380 ;
        RECT -24.380 1197.370 -21.380 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 407.840 1197.370 409.440 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2941.000 1197.370 2944.000 1197.380 ;
        RECT -14.780 1182.380 -11.780 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 407.840 1182.380 409.440 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.400 1182.380 2934.400 1182.390 ;
        RECT -14.780 1179.380 2934.400 1182.380 ;
        RECT -14.780 1179.370 -11.780 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 407.840 1179.370 409.440 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.400 1179.370 2934.400 1179.380 ;
        RECT -24.380 1020.380 -21.380 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 407.840 1020.380 409.440 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2941.000 1020.380 2944.000 1020.390 ;
        RECT -24.380 1017.380 2944.000 1020.380 ;
        RECT -24.380 1017.370 -21.380 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 407.840 1017.370 409.440 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2941.000 1017.370 2944.000 1017.380 ;
        RECT -14.780 1002.380 -11.780 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 407.840 1002.380 409.440 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.400 1002.380 2934.400 1002.390 ;
        RECT -14.780 999.380 2934.400 1002.380 ;
        RECT -14.780 999.370 -11.780 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 407.840 999.370 409.440 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.400 999.370 2934.400 999.380 ;
        RECT -24.380 840.380 -21.380 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 407.840 840.380 409.440 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2941.000 840.380 2944.000 840.390 ;
        RECT -24.380 837.380 2944.000 840.380 ;
        RECT -24.380 837.370 -21.380 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 407.840 837.370 409.440 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2941.000 837.370 2944.000 837.380 ;
        RECT -14.780 822.380 -11.780 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 407.840 822.380 409.440 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.400 822.380 2934.400 822.390 ;
        RECT -14.780 819.380 2934.400 822.380 ;
        RECT -14.780 819.370 -11.780 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 407.840 819.370 409.440 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.400 819.370 2934.400 819.380 ;
        RECT -24.380 660.380 -21.380 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 407.840 660.380 409.440 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2941.000 660.380 2944.000 660.390 ;
        RECT -24.380 657.380 2944.000 660.380 ;
        RECT -24.380 657.370 -21.380 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 407.840 657.370 409.440 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2941.000 657.370 2944.000 657.380 ;
        RECT -14.780 642.380 -11.780 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 407.840 642.380 409.440 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.400 642.380 2934.400 642.390 ;
        RECT -14.780 639.380 2934.400 642.380 ;
        RECT -14.780 639.370 -11.780 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 407.840 639.370 409.440 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.400 639.370 2934.400 639.380 ;
        RECT -24.380 480.380 -21.380 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 407.840 480.380 409.440 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2941.000 480.380 2944.000 480.390 ;
        RECT -24.380 477.380 2944.000 480.380 ;
        RECT -24.380 477.370 -21.380 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 407.840 477.370 409.440 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2941.000 477.370 2944.000 477.380 ;
        RECT -14.780 462.380 -11.780 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 407.840 462.380 409.440 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.400 462.380 2934.400 462.390 ;
        RECT -14.780 459.380 2934.400 462.380 ;
        RECT -14.780 459.370 -11.780 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 407.840 459.370 409.440 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.400 459.370 2934.400 459.380 ;
        RECT -24.380 300.380 -21.380 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 407.840 300.380 409.440 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2941.000 300.380 2944.000 300.390 ;
        RECT -24.380 297.380 2944.000 300.380 ;
        RECT -24.380 297.370 -21.380 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 407.840 297.370 409.440 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2941.000 297.370 2944.000 297.380 ;
        RECT -14.780 282.380 -11.780 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 407.840 282.380 409.440 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.400 282.380 2934.400 282.390 ;
        RECT -14.780 279.380 2934.400 282.380 ;
        RECT -14.780 279.370 -11.780 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 407.840 279.370 409.440 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.400 279.370 2934.400 279.380 ;
        RECT -24.380 120.380 -21.380 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2941.000 120.380 2944.000 120.390 ;
        RECT -24.380 117.380 2944.000 120.380 ;
        RECT -24.380 117.370 -21.380 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2941.000 117.370 2944.000 117.380 ;
        RECT -14.780 102.380 -11.780 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.400 102.380 2934.400 102.390 ;
        RECT -14.780 99.380 2934.400 102.380 ;
        RECT -14.780 99.370 -11.780 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.400 99.370 2934.400 99.380 ;
        RECT -14.780 -6.420 -11.780 -6.410 ;
        RECT 94.020 -6.420 97.020 -6.410 ;
        RECT 274.020 -6.420 277.020 -6.410 ;
        RECT 454.020 -6.420 457.020 -6.410 ;
        RECT 634.020 -6.420 637.020 -6.410 ;
        RECT 814.020 -6.420 817.020 -6.410 ;
        RECT 994.020 -6.420 997.020 -6.410 ;
        RECT 1174.020 -6.420 1177.020 -6.410 ;
        RECT 1354.020 -6.420 1357.020 -6.410 ;
        RECT 1534.020 -6.420 1537.020 -6.410 ;
        RECT 1714.020 -6.420 1717.020 -6.410 ;
        RECT 1894.020 -6.420 1897.020 -6.410 ;
        RECT 2074.020 -6.420 2077.020 -6.410 ;
        RECT 2254.020 -6.420 2257.020 -6.410 ;
        RECT 2434.020 -6.420 2437.020 -6.410 ;
        RECT 2614.020 -6.420 2617.020 -6.410 ;
        RECT 2794.020 -6.420 2797.020 -6.410 ;
        RECT 2931.400 -6.420 2934.400 -6.410 ;
        RECT -14.780 -9.420 2934.400 -6.420 ;
        RECT -14.780 -9.430 -11.780 -9.420 ;
        RECT 94.020 -9.430 97.020 -9.420 ;
        RECT 274.020 -9.430 277.020 -9.420 ;
        RECT 454.020 -9.430 457.020 -9.420 ;
        RECT 634.020 -9.430 637.020 -9.420 ;
        RECT 814.020 -9.430 817.020 -9.420 ;
        RECT 994.020 -9.430 997.020 -9.420 ;
        RECT 1174.020 -9.430 1177.020 -9.420 ;
        RECT 1354.020 -9.430 1357.020 -9.420 ;
        RECT 1534.020 -9.430 1537.020 -9.420 ;
        RECT 1714.020 -9.430 1717.020 -9.420 ;
        RECT 1894.020 -9.430 1897.020 -9.420 ;
        RECT 2074.020 -9.430 2077.020 -9.420 ;
        RECT 2254.020 -9.430 2257.020 -9.420 ;
        RECT 2434.020 -9.430 2437.020 -9.420 ;
        RECT 2614.020 -9.430 2617.020 -9.420 ;
        RECT 2794.020 -9.430 2797.020 -9.420 ;
        RECT 2931.400 -9.430 2934.400 -9.420 ;
        RECT -24.380 -16.020 -21.380 -16.010 ;
        RECT 112.020 -16.020 115.020 -16.010 ;
        RECT 292.020 -16.020 295.020 -16.010 ;
        RECT 472.020 -16.020 475.020 -16.010 ;
        RECT 652.020 -16.020 655.020 -16.010 ;
        RECT 832.020 -16.020 835.020 -16.010 ;
        RECT 1012.020 -16.020 1015.020 -16.010 ;
        RECT 1192.020 -16.020 1195.020 -16.010 ;
        RECT 1372.020 -16.020 1375.020 -16.010 ;
        RECT 1552.020 -16.020 1555.020 -16.010 ;
        RECT 1732.020 -16.020 1735.020 -16.010 ;
        RECT 1912.020 -16.020 1915.020 -16.010 ;
        RECT 2092.020 -16.020 2095.020 -16.010 ;
        RECT 2272.020 -16.020 2275.020 -16.010 ;
        RECT 2452.020 -16.020 2455.020 -16.010 ;
        RECT 2632.020 -16.020 2635.020 -16.010 ;
        RECT 2812.020 -16.020 2815.020 -16.010 ;
        RECT 2941.000 -16.020 2944.000 -16.010 ;
        RECT -24.380 -19.020 2944.000 -16.020 ;
        RECT -24.380 -19.030 -21.380 -19.020 ;
        RECT 112.020 -19.030 115.020 -19.020 ;
        RECT 292.020 -19.030 295.020 -19.020 ;
        RECT 472.020 -19.030 475.020 -19.020 ;
        RECT 652.020 -19.030 655.020 -19.020 ;
        RECT 832.020 -19.030 835.020 -19.020 ;
        RECT 1012.020 -19.030 1015.020 -19.020 ;
        RECT 1192.020 -19.030 1195.020 -19.020 ;
        RECT 1372.020 -19.030 1375.020 -19.020 ;
        RECT 1552.020 -19.030 1555.020 -19.020 ;
        RECT 1732.020 -19.030 1735.020 -19.020 ;
        RECT 1912.020 -19.030 1915.020 -19.020 ;
        RECT 2092.020 -19.030 2095.020 -19.020 ;
        RECT 2272.020 -19.030 2275.020 -19.020 ;
        RECT 2452.020 -19.030 2455.020 -19.020 ;
        RECT 2632.020 -19.030 2635.020 -19.020 ;
        RECT 2812.020 -19.030 2815.020 -19.020 ;
        RECT 2941.000 -19.030 2944.000 -19.020 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 315.520 270.795 2604.480 3246.645 ;
      LAYER met1 ;
        RECT 315.520 268.540 2604.480 3246.800 ;
      LAYER met2 ;
        RECT 312.850 3255.720 352.130 3256.000 ;
        RECT 352.970 3255.720 437.230 3256.000 ;
        RECT 438.070 3255.720 522.330 3256.000 ;
        RECT 523.170 3255.720 607.430 3256.000 ;
        RECT 608.270 3255.720 692.530 3256.000 ;
        RECT 693.370 3255.720 777.630 3256.000 ;
        RECT 778.470 3255.720 863.190 3256.000 ;
        RECT 864.030 3255.720 948.290 3256.000 ;
        RECT 949.130 3255.720 1033.390 3256.000 ;
        RECT 1034.230 3255.720 1118.490 3256.000 ;
        RECT 1119.330 3255.720 1203.590 3256.000 ;
        RECT 1204.430 3255.720 1289.150 3256.000 ;
        RECT 1289.990 3255.720 1374.250 3256.000 ;
        RECT 1375.090 3255.720 1459.350 3256.000 ;
        RECT 1460.190 3255.720 1544.450 3256.000 ;
        RECT 1545.290 3255.720 1629.550 3256.000 ;
        RECT 1630.390 3255.720 1714.650 3256.000 ;
        RECT 1715.490 3255.720 1800.210 3256.000 ;
        RECT 1801.050 3255.720 1885.310 3256.000 ;
        RECT 1886.150 3255.720 1970.410 3256.000 ;
        RECT 1971.250 3255.720 2055.510 3256.000 ;
        RECT 2056.350 3255.720 2140.610 3256.000 ;
        RECT 2141.450 3255.720 2226.170 3256.000 ;
        RECT 2227.010 3255.720 2311.270 3256.000 ;
        RECT 2312.110 3255.720 2396.370 3256.000 ;
        RECT 2397.210 3255.720 2481.470 3256.000 ;
        RECT 2482.310 3255.720 2566.570 3256.000 ;
        RECT 2567.410 3255.720 2602.540 3256.000 ;
        RECT 312.850 264.280 2602.540 3255.720 ;
        RECT 313.410 264.000 318.090 264.280 ;
        RECT 318.930 264.000 324.070 264.280 ;
        RECT 324.910 264.000 330.050 264.280 ;
        RECT 330.890 264.000 336.030 264.280 ;
        RECT 336.870 264.000 342.010 264.280 ;
        RECT 342.850 264.000 347.990 264.280 ;
        RECT 348.830 264.000 353.970 264.280 ;
        RECT 354.810 264.000 359.950 264.280 ;
        RECT 360.790 264.000 365.930 264.280 ;
        RECT 366.770 264.000 371.910 264.280 ;
        RECT 372.750 264.000 377.890 264.280 ;
        RECT 378.730 264.000 383.870 264.280 ;
        RECT 384.710 264.000 389.850 264.280 ;
        RECT 390.690 264.000 395.830 264.280 ;
        RECT 396.670 264.000 401.810 264.280 ;
        RECT 402.650 264.000 407.790 264.280 ;
        RECT 408.630 264.000 413.770 264.280 ;
        RECT 414.610 264.000 419.750 264.280 ;
        RECT 420.590 264.000 425.730 264.280 ;
        RECT 426.570 264.000 431.710 264.280 ;
        RECT 432.550 264.000 437.690 264.280 ;
        RECT 438.530 264.000 443.210 264.280 ;
        RECT 444.050 264.000 449.190 264.280 ;
        RECT 450.030 264.000 455.170 264.280 ;
        RECT 456.010 264.000 461.150 264.280 ;
        RECT 461.990 264.000 467.130 264.280 ;
        RECT 467.970 264.000 473.110 264.280 ;
        RECT 473.950 264.000 479.090 264.280 ;
        RECT 479.930 264.000 485.070 264.280 ;
        RECT 485.910 264.000 491.050 264.280 ;
        RECT 491.890 264.000 497.030 264.280 ;
        RECT 497.870 264.000 503.010 264.280 ;
        RECT 503.850 264.000 508.990 264.280 ;
        RECT 509.830 264.000 514.970 264.280 ;
        RECT 515.810 264.000 520.950 264.280 ;
        RECT 521.790 264.000 526.930 264.280 ;
        RECT 527.770 264.000 532.910 264.280 ;
        RECT 533.750 264.000 538.890 264.280 ;
        RECT 539.730 264.000 544.870 264.280 ;
        RECT 545.710 264.000 550.850 264.280 ;
        RECT 551.690 264.000 556.830 264.280 ;
        RECT 557.670 264.000 562.810 264.280 ;
        RECT 563.650 264.000 568.330 264.280 ;
        RECT 569.170 264.000 574.310 264.280 ;
        RECT 575.150 264.000 580.290 264.280 ;
        RECT 581.130 264.000 586.270 264.280 ;
        RECT 587.110 264.000 592.250 264.280 ;
        RECT 593.090 264.000 598.230 264.280 ;
        RECT 599.070 264.000 604.210 264.280 ;
        RECT 605.050 264.000 610.190 264.280 ;
        RECT 611.030 264.000 616.170 264.280 ;
        RECT 617.010 264.000 622.150 264.280 ;
        RECT 622.990 264.000 628.130 264.280 ;
        RECT 628.970 264.000 634.110 264.280 ;
        RECT 634.950 264.000 640.090 264.280 ;
        RECT 640.930 264.000 646.070 264.280 ;
        RECT 646.910 264.000 652.050 264.280 ;
        RECT 652.890 264.000 658.030 264.280 ;
        RECT 658.870 264.000 664.010 264.280 ;
        RECT 664.850 264.000 669.990 264.280 ;
        RECT 670.830 264.000 675.970 264.280 ;
        RECT 676.810 264.000 681.950 264.280 ;
        RECT 682.790 264.000 687.930 264.280 ;
        RECT 688.770 264.000 693.910 264.280 ;
        RECT 694.750 264.000 699.430 264.280 ;
        RECT 700.270 264.000 705.410 264.280 ;
        RECT 706.250 264.000 711.390 264.280 ;
        RECT 712.230 264.000 717.370 264.280 ;
        RECT 718.210 264.000 723.350 264.280 ;
        RECT 724.190 264.000 729.330 264.280 ;
        RECT 730.170 264.000 735.310 264.280 ;
        RECT 736.150 264.000 741.290 264.280 ;
        RECT 742.130 264.000 747.270 264.280 ;
        RECT 748.110 264.000 753.250 264.280 ;
        RECT 754.090 264.000 759.230 264.280 ;
        RECT 760.070 264.000 765.210 264.280 ;
        RECT 766.050 264.000 771.190 264.280 ;
        RECT 772.030 264.000 777.170 264.280 ;
        RECT 778.010 264.000 783.150 264.280 ;
        RECT 783.990 264.000 789.130 264.280 ;
        RECT 789.970 264.000 795.110 264.280 ;
        RECT 795.950 264.000 801.090 264.280 ;
        RECT 801.930 264.000 807.070 264.280 ;
        RECT 807.910 264.000 813.050 264.280 ;
        RECT 813.890 264.000 819.030 264.280 ;
        RECT 819.870 264.000 824.550 264.280 ;
        RECT 825.390 264.000 830.530 264.280 ;
        RECT 831.370 264.000 836.510 264.280 ;
        RECT 837.350 264.000 842.490 264.280 ;
        RECT 843.330 264.000 848.470 264.280 ;
        RECT 849.310 264.000 854.450 264.280 ;
        RECT 855.290 264.000 860.430 264.280 ;
        RECT 861.270 264.000 866.410 264.280 ;
        RECT 867.250 264.000 872.390 264.280 ;
        RECT 873.230 264.000 878.370 264.280 ;
        RECT 879.210 264.000 884.350 264.280 ;
        RECT 885.190 264.000 890.330 264.280 ;
        RECT 891.170 264.000 896.310 264.280 ;
        RECT 897.150 264.000 902.290 264.280 ;
        RECT 903.130 264.000 908.270 264.280 ;
        RECT 909.110 264.000 914.250 264.280 ;
        RECT 915.090 264.000 920.230 264.280 ;
        RECT 921.070 264.000 926.210 264.280 ;
        RECT 927.050 264.000 932.190 264.280 ;
        RECT 933.030 264.000 938.170 264.280 ;
        RECT 939.010 264.000 944.150 264.280 ;
        RECT 944.990 264.000 950.130 264.280 ;
        RECT 950.970 264.000 955.650 264.280 ;
        RECT 956.490 264.000 961.630 264.280 ;
        RECT 962.470 264.000 967.610 264.280 ;
        RECT 968.450 264.000 973.590 264.280 ;
        RECT 974.430 264.000 979.570 264.280 ;
        RECT 980.410 264.000 985.550 264.280 ;
        RECT 986.390 264.000 991.530 264.280 ;
        RECT 992.370 264.000 997.510 264.280 ;
        RECT 998.350 264.000 1003.490 264.280 ;
        RECT 1004.330 264.000 1009.470 264.280 ;
        RECT 1010.310 264.000 1015.450 264.280 ;
        RECT 1016.290 264.000 1021.430 264.280 ;
        RECT 1022.270 264.000 1027.410 264.280 ;
        RECT 1028.250 264.000 1033.390 264.280 ;
        RECT 1034.230 264.000 1039.370 264.280 ;
        RECT 1040.210 264.000 1045.350 264.280 ;
        RECT 1046.190 264.000 1051.330 264.280 ;
        RECT 1052.170 264.000 1057.310 264.280 ;
        RECT 1058.150 264.000 1063.290 264.280 ;
        RECT 1064.130 264.000 1069.270 264.280 ;
        RECT 1070.110 264.000 1075.250 264.280 ;
        RECT 1076.090 264.000 1080.770 264.280 ;
        RECT 1081.610 264.000 1086.750 264.280 ;
        RECT 1087.590 264.000 1092.730 264.280 ;
        RECT 1093.570 264.000 1098.710 264.280 ;
        RECT 1099.550 264.000 1104.690 264.280 ;
        RECT 1105.530 264.000 1110.670 264.280 ;
        RECT 1111.510 264.000 1116.650 264.280 ;
        RECT 1117.490 264.000 1122.630 264.280 ;
        RECT 1123.470 264.000 1128.610 264.280 ;
        RECT 1129.450 264.000 1134.590 264.280 ;
        RECT 1135.430 264.000 1140.570 264.280 ;
        RECT 1141.410 264.000 1146.550 264.280 ;
        RECT 1147.390 264.000 1152.530 264.280 ;
        RECT 1153.370 264.000 1158.510 264.280 ;
        RECT 1159.350 264.000 1164.490 264.280 ;
        RECT 1165.330 264.000 1170.470 264.280 ;
        RECT 1171.310 264.000 1176.450 264.280 ;
        RECT 1177.290 264.000 1182.430 264.280 ;
        RECT 1183.270 264.000 1188.410 264.280 ;
        RECT 1189.250 264.000 1194.390 264.280 ;
        RECT 1195.230 264.000 1200.370 264.280 ;
        RECT 1201.210 264.000 1206.350 264.280 ;
        RECT 1207.190 264.000 1211.870 264.280 ;
        RECT 1212.710 264.000 1217.850 264.280 ;
        RECT 1218.690 264.000 1223.830 264.280 ;
        RECT 1224.670 264.000 1229.810 264.280 ;
        RECT 1230.650 264.000 1235.790 264.280 ;
        RECT 1236.630 264.000 1241.770 264.280 ;
        RECT 1242.610 264.000 1247.750 264.280 ;
        RECT 1248.590 264.000 1253.730 264.280 ;
        RECT 1254.570 264.000 1259.710 264.280 ;
        RECT 1260.550 264.000 1265.690 264.280 ;
        RECT 1266.530 264.000 1271.670 264.280 ;
        RECT 1272.510 264.000 1277.650 264.280 ;
        RECT 1278.490 264.000 1283.630 264.280 ;
        RECT 1284.470 264.000 1289.610 264.280 ;
        RECT 1290.450 264.000 1295.590 264.280 ;
        RECT 1296.430 264.000 1301.570 264.280 ;
        RECT 1302.410 264.000 1307.550 264.280 ;
        RECT 1308.390 264.000 1313.530 264.280 ;
        RECT 1314.370 264.000 1319.510 264.280 ;
        RECT 1320.350 264.000 1325.490 264.280 ;
        RECT 1326.330 264.000 1331.470 264.280 ;
        RECT 1332.310 264.000 1336.990 264.280 ;
        RECT 1337.830 264.000 1342.970 264.280 ;
        RECT 1343.810 264.000 1348.950 264.280 ;
        RECT 1349.790 264.000 1354.930 264.280 ;
        RECT 1355.770 264.000 1360.910 264.280 ;
        RECT 1361.750 264.000 1366.890 264.280 ;
        RECT 1367.730 264.000 1372.870 264.280 ;
        RECT 1373.710 264.000 1378.850 264.280 ;
        RECT 1379.690 264.000 1384.830 264.280 ;
        RECT 1385.670 264.000 1390.810 264.280 ;
        RECT 1391.650 264.000 1396.790 264.280 ;
        RECT 1397.630 264.000 1402.770 264.280 ;
        RECT 1403.610 264.000 1408.750 264.280 ;
        RECT 1409.590 264.000 1414.730 264.280 ;
        RECT 1415.570 264.000 1420.710 264.280 ;
        RECT 1421.550 264.000 1426.690 264.280 ;
        RECT 1427.530 264.000 1432.670 264.280 ;
        RECT 1433.510 264.000 1438.650 264.280 ;
        RECT 1439.490 264.000 1444.630 264.280 ;
        RECT 1445.470 264.000 1450.610 264.280 ;
        RECT 1451.450 264.000 1456.590 264.280 ;
        RECT 1457.430 264.000 1462.570 264.280 ;
        RECT 1463.410 264.000 1468.090 264.280 ;
        RECT 1468.930 264.000 1474.070 264.280 ;
        RECT 1474.910 264.000 1480.050 264.280 ;
        RECT 1480.890 264.000 1486.030 264.280 ;
        RECT 1486.870 264.000 1492.010 264.280 ;
        RECT 1492.850 264.000 1497.990 264.280 ;
        RECT 1498.830 264.000 1503.970 264.280 ;
        RECT 1504.810 264.000 1509.950 264.280 ;
        RECT 1510.790 264.000 1515.930 264.280 ;
        RECT 1516.770 264.000 1521.910 264.280 ;
        RECT 1522.750 264.000 1527.890 264.280 ;
        RECT 1528.730 264.000 1533.870 264.280 ;
        RECT 1534.710 264.000 1539.850 264.280 ;
        RECT 1540.690 264.000 1545.830 264.280 ;
        RECT 1546.670 264.000 1551.810 264.280 ;
        RECT 1552.650 264.000 1557.790 264.280 ;
        RECT 1558.630 264.000 1563.770 264.280 ;
        RECT 1564.610 264.000 1569.750 264.280 ;
        RECT 1570.590 264.000 1575.730 264.280 ;
        RECT 1576.570 264.000 1581.710 264.280 ;
        RECT 1582.550 264.000 1587.690 264.280 ;
        RECT 1588.530 264.000 1593.210 264.280 ;
        RECT 1594.050 264.000 1599.190 264.280 ;
        RECT 1600.030 264.000 1605.170 264.280 ;
        RECT 1606.010 264.000 1611.150 264.280 ;
        RECT 1611.990 264.000 1617.130 264.280 ;
        RECT 1617.970 264.000 1623.110 264.280 ;
        RECT 1623.950 264.000 1629.090 264.280 ;
        RECT 1629.930 264.000 1635.070 264.280 ;
        RECT 1635.910 264.000 1641.050 264.280 ;
        RECT 1641.890 264.000 1647.030 264.280 ;
        RECT 1647.870 264.000 1653.010 264.280 ;
        RECT 1653.850 264.000 1658.990 264.280 ;
        RECT 1659.830 264.000 1664.970 264.280 ;
        RECT 1665.810 264.000 1670.950 264.280 ;
        RECT 1671.790 264.000 1676.930 264.280 ;
        RECT 1677.770 264.000 1682.910 264.280 ;
        RECT 1683.750 264.000 1688.890 264.280 ;
        RECT 1689.730 264.000 1694.870 264.280 ;
        RECT 1695.710 264.000 1700.850 264.280 ;
        RECT 1701.690 264.000 1706.830 264.280 ;
        RECT 1707.670 264.000 1712.810 264.280 ;
        RECT 1713.650 264.000 1718.330 264.280 ;
        RECT 1719.170 264.000 1724.310 264.280 ;
        RECT 1725.150 264.000 1730.290 264.280 ;
        RECT 1731.130 264.000 1736.270 264.280 ;
        RECT 1737.110 264.000 1742.250 264.280 ;
        RECT 1743.090 264.000 1748.230 264.280 ;
        RECT 1749.070 264.000 1754.210 264.280 ;
        RECT 1755.050 264.000 1760.190 264.280 ;
        RECT 1761.030 264.000 1766.170 264.280 ;
        RECT 1767.010 264.000 1772.150 264.280 ;
        RECT 1772.990 264.000 1778.130 264.280 ;
        RECT 1778.970 264.000 1784.110 264.280 ;
        RECT 1784.950 264.000 1790.090 264.280 ;
        RECT 1790.930 264.000 1796.070 264.280 ;
        RECT 1796.910 264.000 1802.050 264.280 ;
        RECT 1802.890 264.000 1808.030 264.280 ;
        RECT 1808.870 264.000 1814.010 264.280 ;
        RECT 1814.850 264.000 1819.990 264.280 ;
        RECT 1820.830 264.000 1825.970 264.280 ;
        RECT 1826.810 264.000 1831.950 264.280 ;
        RECT 1832.790 264.000 1837.930 264.280 ;
        RECT 1838.770 264.000 1843.910 264.280 ;
        RECT 1844.750 264.000 1849.430 264.280 ;
        RECT 1850.270 264.000 1855.410 264.280 ;
        RECT 1856.250 264.000 1861.390 264.280 ;
        RECT 1862.230 264.000 1867.370 264.280 ;
        RECT 1868.210 264.000 1873.350 264.280 ;
        RECT 1874.190 264.000 1879.330 264.280 ;
        RECT 1880.170 264.000 1885.310 264.280 ;
        RECT 1886.150 264.000 1891.290 264.280 ;
        RECT 1892.130 264.000 1897.270 264.280 ;
        RECT 1898.110 264.000 1903.250 264.280 ;
        RECT 1904.090 264.000 1909.230 264.280 ;
        RECT 1910.070 264.000 1915.210 264.280 ;
        RECT 1916.050 264.000 1921.190 264.280 ;
        RECT 1922.030 264.000 1927.170 264.280 ;
        RECT 1928.010 264.000 1933.150 264.280 ;
        RECT 1933.990 264.000 1939.130 264.280 ;
        RECT 1939.970 264.000 1945.110 264.280 ;
        RECT 1945.950 264.000 1951.090 264.280 ;
        RECT 1951.930 264.000 1957.070 264.280 ;
        RECT 1957.910 264.000 1963.050 264.280 ;
        RECT 1963.890 264.000 1969.030 264.280 ;
        RECT 1969.870 264.000 1974.550 264.280 ;
        RECT 1975.390 264.000 1980.530 264.280 ;
        RECT 1981.370 264.000 1986.510 264.280 ;
        RECT 1987.350 264.000 1992.490 264.280 ;
        RECT 1993.330 264.000 1998.470 264.280 ;
        RECT 1999.310 264.000 2004.450 264.280 ;
        RECT 2005.290 264.000 2010.430 264.280 ;
        RECT 2011.270 264.000 2016.410 264.280 ;
        RECT 2017.250 264.000 2022.390 264.280 ;
        RECT 2023.230 264.000 2028.370 264.280 ;
        RECT 2029.210 264.000 2034.350 264.280 ;
        RECT 2035.190 264.000 2040.330 264.280 ;
        RECT 2041.170 264.000 2046.310 264.280 ;
        RECT 2047.150 264.000 2052.290 264.280 ;
        RECT 2053.130 264.000 2058.270 264.280 ;
        RECT 2059.110 264.000 2064.250 264.280 ;
        RECT 2065.090 264.000 2070.230 264.280 ;
        RECT 2071.070 264.000 2076.210 264.280 ;
        RECT 2077.050 264.000 2082.190 264.280 ;
        RECT 2083.030 264.000 2088.170 264.280 ;
        RECT 2089.010 264.000 2094.150 264.280 ;
        RECT 2094.990 264.000 2100.130 264.280 ;
        RECT 2100.970 264.000 2105.650 264.280 ;
        RECT 2106.490 264.000 2111.630 264.280 ;
        RECT 2112.470 264.000 2117.610 264.280 ;
        RECT 2118.450 264.000 2123.590 264.280 ;
        RECT 2124.430 264.000 2129.570 264.280 ;
        RECT 2130.410 264.000 2135.550 264.280 ;
        RECT 2136.390 264.000 2141.530 264.280 ;
        RECT 2142.370 264.000 2147.510 264.280 ;
        RECT 2148.350 264.000 2153.490 264.280 ;
        RECT 2154.330 264.000 2159.470 264.280 ;
        RECT 2160.310 264.000 2165.450 264.280 ;
        RECT 2166.290 264.000 2171.430 264.280 ;
        RECT 2172.270 264.000 2177.410 264.280 ;
        RECT 2178.250 264.000 2183.390 264.280 ;
        RECT 2184.230 264.000 2189.370 264.280 ;
        RECT 2190.210 264.000 2195.350 264.280 ;
        RECT 2196.190 264.000 2201.330 264.280 ;
        RECT 2202.170 264.000 2207.310 264.280 ;
        RECT 2208.150 264.000 2213.290 264.280 ;
        RECT 2214.130 264.000 2219.270 264.280 ;
        RECT 2220.110 264.000 2225.250 264.280 ;
        RECT 2226.090 264.000 2230.770 264.280 ;
        RECT 2231.610 264.000 2236.750 264.280 ;
        RECT 2237.590 264.000 2242.730 264.280 ;
        RECT 2243.570 264.000 2248.710 264.280 ;
        RECT 2249.550 264.000 2254.690 264.280 ;
        RECT 2255.530 264.000 2260.670 264.280 ;
        RECT 2261.510 264.000 2266.650 264.280 ;
        RECT 2267.490 264.000 2272.630 264.280 ;
        RECT 2273.470 264.000 2278.610 264.280 ;
        RECT 2279.450 264.000 2284.590 264.280 ;
        RECT 2285.430 264.000 2290.570 264.280 ;
        RECT 2291.410 264.000 2296.550 264.280 ;
        RECT 2297.390 264.000 2302.530 264.280 ;
        RECT 2303.370 264.000 2308.510 264.280 ;
        RECT 2309.350 264.000 2314.490 264.280 ;
        RECT 2315.330 264.000 2320.470 264.280 ;
        RECT 2321.310 264.000 2326.450 264.280 ;
        RECT 2327.290 264.000 2332.430 264.280 ;
        RECT 2333.270 264.000 2338.410 264.280 ;
        RECT 2339.250 264.000 2344.390 264.280 ;
        RECT 2345.230 264.000 2350.370 264.280 ;
        RECT 2351.210 264.000 2356.350 264.280 ;
        RECT 2357.190 264.000 2361.870 264.280 ;
        RECT 2362.710 264.000 2367.850 264.280 ;
        RECT 2368.690 264.000 2373.830 264.280 ;
        RECT 2374.670 264.000 2379.810 264.280 ;
        RECT 2380.650 264.000 2385.790 264.280 ;
        RECT 2386.630 264.000 2391.770 264.280 ;
        RECT 2392.610 264.000 2397.750 264.280 ;
        RECT 2398.590 264.000 2403.730 264.280 ;
        RECT 2404.570 264.000 2409.710 264.280 ;
        RECT 2410.550 264.000 2415.690 264.280 ;
        RECT 2416.530 264.000 2421.670 264.280 ;
        RECT 2422.510 264.000 2427.650 264.280 ;
        RECT 2428.490 264.000 2433.630 264.280 ;
        RECT 2434.470 264.000 2439.610 264.280 ;
        RECT 2440.450 264.000 2445.590 264.280 ;
        RECT 2446.430 264.000 2451.570 264.280 ;
        RECT 2452.410 264.000 2457.550 264.280 ;
        RECT 2458.390 264.000 2463.530 264.280 ;
        RECT 2464.370 264.000 2469.510 264.280 ;
        RECT 2470.350 264.000 2475.490 264.280 ;
        RECT 2476.330 264.000 2481.470 264.280 ;
        RECT 2482.310 264.000 2486.990 264.280 ;
        RECT 2487.830 264.000 2492.970 264.280 ;
        RECT 2493.810 264.000 2498.950 264.280 ;
        RECT 2499.790 264.000 2504.930 264.280 ;
        RECT 2505.770 264.000 2510.910 264.280 ;
        RECT 2511.750 264.000 2516.890 264.280 ;
        RECT 2517.730 264.000 2522.870 264.280 ;
        RECT 2523.710 264.000 2528.850 264.280 ;
        RECT 2529.690 264.000 2534.830 264.280 ;
        RECT 2535.670 264.000 2540.810 264.280 ;
        RECT 2541.650 264.000 2546.790 264.280 ;
        RECT 2547.630 264.000 2552.770 264.280 ;
        RECT 2553.610 264.000 2558.750 264.280 ;
        RECT 2559.590 264.000 2564.730 264.280 ;
        RECT 2565.570 264.000 2570.710 264.280 ;
        RECT 2571.550 264.000 2576.690 264.280 ;
        RECT 2577.530 264.000 2582.670 264.280 ;
        RECT 2583.510 264.000 2588.650 264.280 ;
        RECT 2589.490 264.000 2594.630 264.280 ;
        RECT 2595.470 264.000 2600.610 264.280 ;
        RECT 2601.450 264.000 2602.540 264.280 ;
      LAYER met3 ;
        RECT 312.825 3227.200 2606.010 3246.725 ;
        RECT 312.825 3225.800 2605.600 3227.200 ;
        RECT 312.825 3224.480 2606.010 3225.800 ;
        RECT 314.400 3223.080 2606.010 3224.480 ;
        RECT 312.825 3160.560 2606.010 3223.080 ;
        RECT 312.825 3159.160 2605.600 3160.560 ;
        RECT 312.825 3153.080 2606.010 3159.160 ;
        RECT 314.400 3151.680 2606.010 3153.080 ;
        RECT 312.825 3093.920 2606.010 3151.680 ;
        RECT 312.825 3092.520 2605.600 3093.920 ;
        RECT 312.825 3081.680 2606.010 3092.520 ;
        RECT 314.400 3080.280 2606.010 3081.680 ;
        RECT 312.825 3027.280 2606.010 3080.280 ;
        RECT 312.825 3025.880 2605.600 3027.280 ;
        RECT 312.825 3010.280 2606.010 3025.880 ;
        RECT 314.400 3008.880 2606.010 3010.280 ;
        RECT 312.825 2960.640 2606.010 3008.880 ;
        RECT 312.825 2959.240 2605.600 2960.640 ;
        RECT 312.825 2938.880 2606.010 2959.240 ;
        RECT 314.400 2937.480 2606.010 2938.880 ;
        RECT 312.825 2894.000 2606.010 2937.480 ;
        RECT 312.825 2892.600 2605.600 2894.000 ;
        RECT 312.825 2867.480 2606.010 2892.600 ;
        RECT 314.400 2866.080 2606.010 2867.480 ;
        RECT 312.825 2827.360 2606.010 2866.080 ;
        RECT 312.825 2825.960 2605.600 2827.360 ;
        RECT 312.825 2796.080 2606.010 2825.960 ;
        RECT 314.400 2794.680 2606.010 2796.080 ;
        RECT 312.825 2760.720 2606.010 2794.680 ;
        RECT 312.825 2759.320 2605.600 2760.720 ;
        RECT 312.825 2724.680 2606.010 2759.320 ;
        RECT 314.400 2723.280 2606.010 2724.680 ;
        RECT 312.825 2694.080 2606.010 2723.280 ;
        RECT 312.825 2692.680 2605.600 2694.080 ;
        RECT 312.825 2653.280 2606.010 2692.680 ;
        RECT 314.400 2651.880 2606.010 2653.280 ;
        RECT 312.825 2627.440 2606.010 2651.880 ;
        RECT 312.825 2626.040 2605.600 2627.440 ;
        RECT 312.825 2581.880 2606.010 2626.040 ;
        RECT 314.400 2580.480 2606.010 2581.880 ;
        RECT 312.825 2560.800 2606.010 2580.480 ;
        RECT 312.825 2559.400 2605.600 2560.800 ;
        RECT 312.825 2510.480 2606.010 2559.400 ;
        RECT 314.400 2509.080 2606.010 2510.480 ;
        RECT 312.825 2494.160 2606.010 2509.080 ;
        RECT 312.825 2492.760 2605.600 2494.160 ;
        RECT 312.825 2439.080 2606.010 2492.760 ;
        RECT 314.400 2437.680 2606.010 2439.080 ;
        RECT 312.825 2427.520 2606.010 2437.680 ;
        RECT 312.825 2426.120 2605.600 2427.520 ;
        RECT 312.825 2367.680 2606.010 2426.120 ;
        RECT 314.400 2366.280 2606.010 2367.680 ;
        RECT 312.825 2360.880 2606.010 2366.280 ;
        RECT 312.825 2359.480 2605.600 2360.880 ;
        RECT 312.825 2296.280 2606.010 2359.480 ;
        RECT 314.400 2294.880 2606.010 2296.280 ;
        RECT 312.825 2294.240 2606.010 2294.880 ;
        RECT 312.825 2292.840 2605.600 2294.240 ;
        RECT 312.825 2227.600 2606.010 2292.840 ;
        RECT 312.825 2226.200 2605.600 2227.600 ;
        RECT 312.825 2224.880 2606.010 2226.200 ;
        RECT 314.400 2223.480 2606.010 2224.880 ;
        RECT 312.825 2160.960 2606.010 2223.480 ;
        RECT 312.825 2159.560 2605.600 2160.960 ;
        RECT 312.825 2153.480 2606.010 2159.560 ;
        RECT 314.400 2152.080 2606.010 2153.480 ;
        RECT 312.825 2094.320 2606.010 2152.080 ;
        RECT 312.825 2092.920 2605.600 2094.320 ;
        RECT 312.825 2082.080 2606.010 2092.920 ;
        RECT 314.400 2080.680 2606.010 2082.080 ;
        RECT 312.825 2027.680 2606.010 2080.680 ;
        RECT 312.825 2026.280 2605.600 2027.680 ;
        RECT 312.825 2010.680 2606.010 2026.280 ;
        RECT 314.400 2009.280 2606.010 2010.680 ;
        RECT 312.825 1961.040 2606.010 2009.280 ;
        RECT 312.825 1959.640 2605.600 1961.040 ;
        RECT 312.825 1939.280 2606.010 1959.640 ;
        RECT 314.400 1937.880 2606.010 1939.280 ;
        RECT 312.825 1894.400 2606.010 1937.880 ;
        RECT 312.825 1893.000 2605.600 1894.400 ;
        RECT 312.825 1867.880 2606.010 1893.000 ;
        RECT 314.400 1866.480 2606.010 1867.880 ;
        RECT 312.825 1827.760 2606.010 1866.480 ;
        RECT 312.825 1826.360 2605.600 1827.760 ;
        RECT 312.825 1796.480 2606.010 1826.360 ;
        RECT 314.400 1795.080 2606.010 1796.480 ;
        RECT 312.825 1760.440 2606.010 1795.080 ;
        RECT 312.825 1759.040 2605.600 1760.440 ;
        RECT 312.825 1724.400 2606.010 1759.040 ;
        RECT 314.400 1723.000 2606.010 1724.400 ;
        RECT 312.825 1693.800 2606.010 1723.000 ;
        RECT 312.825 1692.400 2605.600 1693.800 ;
        RECT 312.825 1653.000 2606.010 1692.400 ;
        RECT 314.400 1651.600 2606.010 1653.000 ;
        RECT 312.825 1627.160 2606.010 1651.600 ;
        RECT 312.825 1625.760 2605.600 1627.160 ;
        RECT 312.825 1581.600 2606.010 1625.760 ;
        RECT 314.400 1580.200 2606.010 1581.600 ;
        RECT 312.825 1560.520 2606.010 1580.200 ;
        RECT 312.825 1559.120 2605.600 1560.520 ;
        RECT 312.825 1510.200 2606.010 1559.120 ;
        RECT 314.400 1508.800 2606.010 1510.200 ;
        RECT 312.825 1493.880 2606.010 1508.800 ;
        RECT 312.825 1492.480 2605.600 1493.880 ;
        RECT 312.825 1438.800 2606.010 1492.480 ;
        RECT 314.400 1437.400 2606.010 1438.800 ;
        RECT 312.825 1427.240 2606.010 1437.400 ;
        RECT 312.825 1425.840 2605.600 1427.240 ;
        RECT 312.825 1367.400 2606.010 1425.840 ;
        RECT 314.400 1366.000 2606.010 1367.400 ;
        RECT 312.825 1360.600 2606.010 1366.000 ;
        RECT 312.825 1359.200 2605.600 1360.600 ;
        RECT 312.825 1296.000 2606.010 1359.200 ;
        RECT 314.400 1294.600 2606.010 1296.000 ;
        RECT 312.825 1293.960 2606.010 1294.600 ;
        RECT 312.825 1292.560 2605.600 1293.960 ;
        RECT 312.825 1227.320 2606.010 1292.560 ;
        RECT 312.825 1225.920 2605.600 1227.320 ;
        RECT 312.825 1224.600 2606.010 1225.920 ;
        RECT 314.400 1223.200 2606.010 1224.600 ;
        RECT 312.825 1160.680 2606.010 1223.200 ;
        RECT 312.825 1159.280 2605.600 1160.680 ;
        RECT 312.825 1153.200 2606.010 1159.280 ;
        RECT 314.400 1151.800 2606.010 1153.200 ;
        RECT 312.825 1094.040 2606.010 1151.800 ;
        RECT 312.825 1092.640 2605.600 1094.040 ;
        RECT 312.825 1081.800 2606.010 1092.640 ;
        RECT 314.400 1080.400 2606.010 1081.800 ;
        RECT 312.825 1027.400 2606.010 1080.400 ;
        RECT 312.825 1026.000 2605.600 1027.400 ;
        RECT 312.825 1010.400 2606.010 1026.000 ;
        RECT 314.400 1009.000 2606.010 1010.400 ;
        RECT 312.825 960.760 2606.010 1009.000 ;
        RECT 312.825 959.360 2605.600 960.760 ;
        RECT 312.825 939.000 2606.010 959.360 ;
        RECT 314.400 937.600 2606.010 939.000 ;
        RECT 312.825 894.120 2606.010 937.600 ;
        RECT 312.825 892.720 2605.600 894.120 ;
        RECT 312.825 867.600 2606.010 892.720 ;
        RECT 314.400 866.200 2606.010 867.600 ;
        RECT 312.825 827.480 2606.010 866.200 ;
        RECT 312.825 826.080 2605.600 827.480 ;
        RECT 312.825 796.200 2606.010 826.080 ;
        RECT 314.400 794.800 2606.010 796.200 ;
        RECT 312.825 760.840 2606.010 794.800 ;
        RECT 312.825 759.440 2605.600 760.840 ;
        RECT 312.825 724.800 2606.010 759.440 ;
        RECT 314.400 723.400 2606.010 724.800 ;
        RECT 312.825 694.200 2606.010 723.400 ;
        RECT 312.825 692.800 2605.600 694.200 ;
        RECT 312.825 653.400 2606.010 692.800 ;
        RECT 314.400 652.000 2606.010 653.400 ;
        RECT 312.825 627.560 2606.010 652.000 ;
        RECT 312.825 626.160 2605.600 627.560 ;
        RECT 312.825 582.000 2606.010 626.160 ;
        RECT 314.400 580.600 2606.010 582.000 ;
        RECT 312.825 560.920 2606.010 580.600 ;
        RECT 312.825 559.520 2605.600 560.920 ;
        RECT 312.825 510.600 2606.010 559.520 ;
        RECT 314.400 509.200 2606.010 510.600 ;
        RECT 312.825 494.280 2606.010 509.200 ;
        RECT 312.825 492.880 2605.600 494.280 ;
        RECT 312.825 439.200 2606.010 492.880 ;
        RECT 314.400 437.800 2606.010 439.200 ;
        RECT 312.825 427.640 2606.010 437.800 ;
        RECT 312.825 426.240 2605.600 427.640 ;
        RECT 312.825 367.800 2606.010 426.240 ;
        RECT 314.400 366.400 2606.010 367.800 ;
        RECT 312.825 361.000 2606.010 366.400 ;
        RECT 312.825 359.600 2605.600 361.000 ;
        RECT 312.825 296.400 2606.010 359.600 ;
        RECT 314.400 295.000 2606.010 296.400 ;
        RECT 312.825 294.360 2606.010 295.000 ;
        RECT 312.825 292.960 2605.600 294.360 ;
        RECT 312.825 270.715 2606.010 292.960 ;
      LAYER met4 ;
        RECT 326.855 270.640 330.640 3246.800 ;
        RECT 333.040 270.640 407.440 3246.800 ;
        RECT 409.840 270.640 2592.225 3246.800 ;
=======
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 3519.700 97.020 3529.000 ;
        RECT 274.020 3519.700 277.020 3529.000 ;
        RECT 454.020 3519.700 457.020 3529.000 ;
        RECT 634.020 3519.700 637.020 3529.000 ;
        RECT 814.020 3519.700 817.020 3529.000 ;
        RECT 994.020 3519.700 997.020 3529.000 ;
        RECT 1174.020 3519.700 1177.020 3529.000 ;
        RECT 1354.020 3519.700 1357.020 3529.000 ;
        RECT 1534.020 3519.700 1537.020 3529.000 ;
        RECT 1714.020 3519.700 1717.020 3529.000 ;
        RECT 1894.020 3519.700 1897.020 3529.000 ;
        RECT 2074.020 3519.700 2077.020 3529.000 ;
        RECT 2254.020 3519.700 2257.020 3529.000 ;
        RECT 2434.020 3519.700 2437.020 3529.000 ;
        RECT 2614.020 3519.700 2617.020 3529.000 ;
        RECT 2794.020 3519.700 2797.020 3529.000 ;
        RECT 94.020 -9.320 97.020 0.300 ;
        RECT 274.020 -9.320 277.020 0.300 ;
        RECT 454.020 -9.320 457.020 0.300 ;
        RECT 634.020 -9.320 637.020 0.300 ;
        RECT 814.020 -9.320 817.020 0.300 ;
        RECT 994.020 -9.320 997.020 0.300 ;
        RECT 1174.020 -9.320 1177.020 0.300 ;
        RECT 1354.020 -9.320 1357.020 0.300 ;
        RECT 1534.020 -9.320 1537.020 0.300 ;
        RECT 1714.020 -9.320 1717.020 0.300 ;
        RECT 1894.020 -9.320 1897.020 0.300 ;
        RECT 2074.020 -9.320 2077.020 0.300 ;
        RECT 2254.020 -9.320 2257.020 0.300 ;
        RECT 2434.020 -9.320 2437.020 0.300 ;
        RECT 2614.020 -9.320 2617.020 0.300 ;
        RECT 2794.020 -9.320 2797.020 0.300 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3340.850 -12.590 3342.030 ;
        RECT -13.770 3339.250 -12.590 3340.430 ;
        RECT -13.770 3160.850 -12.590 3162.030 ;
        RECT -13.770 3159.250 -12.590 3160.430 ;
        RECT -13.770 2980.850 -12.590 2982.030 ;
        RECT -13.770 2979.250 -12.590 2980.430 ;
        RECT -13.770 2800.850 -12.590 2802.030 ;
        RECT -13.770 2799.250 -12.590 2800.430 ;
        RECT -13.770 2620.850 -12.590 2622.030 ;
        RECT -13.770 2619.250 -12.590 2620.430 ;
        RECT -13.770 2440.850 -12.590 2442.030 ;
        RECT -13.770 2439.250 -12.590 2440.430 ;
        RECT -13.770 2260.850 -12.590 2262.030 ;
        RECT -13.770 2259.250 -12.590 2260.430 ;
        RECT -13.770 2080.850 -12.590 2082.030 ;
        RECT -13.770 2079.250 -12.590 2080.430 ;
        RECT -13.770 1900.850 -12.590 1902.030 ;
        RECT -13.770 1899.250 -12.590 1900.430 ;
        RECT -13.770 1720.850 -12.590 1722.030 ;
        RECT -13.770 1719.250 -12.590 1720.430 ;
        RECT -13.770 1540.850 -12.590 1542.030 ;
        RECT -13.770 1539.250 -12.590 1540.430 ;
        RECT -13.770 1360.850 -12.590 1362.030 ;
        RECT -13.770 1359.250 -12.590 1360.430 ;
        RECT -13.770 1180.850 -12.590 1182.030 ;
        RECT -13.770 1179.250 -12.590 1180.430 ;
        RECT -13.770 1000.850 -12.590 1002.030 ;
        RECT -13.770 999.250 -12.590 1000.430 ;
        RECT -13.770 820.850 -12.590 822.030 ;
        RECT -13.770 819.250 -12.590 820.430 ;
        RECT -13.770 640.850 -12.590 642.030 ;
        RECT -13.770 639.250 -12.590 640.430 ;
        RECT -13.770 460.850 -12.590 462.030 ;
        RECT -13.770 459.250 -12.590 460.430 ;
        RECT -13.770 280.850 -12.590 282.030 ;
        RECT -13.770 279.250 -12.590 280.430 ;
        RECT -13.770 100.850 -12.590 102.030 ;
        RECT -13.770 99.250 -12.590 100.430 ;
        RECT 2932.210 3340.850 2933.390 3342.030 ;
        RECT 2932.210 3339.250 2933.390 3340.430 ;
        RECT 2932.210 3160.850 2933.390 3162.030 ;
        RECT 2932.210 3159.250 2933.390 3160.430 ;
        RECT 2932.210 2980.850 2933.390 2982.030 ;
        RECT 2932.210 2979.250 2933.390 2980.430 ;
        RECT 2932.210 2800.850 2933.390 2802.030 ;
        RECT 2932.210 2799.250 2933.390 2800.430 ;
        RECT 2932.210 2620.850 2933.390 2622.030 ;
        RECT 2932.210 2619.250 2933.390 2620.430 ;
        RECT 2932.210 2440.850 2933.390 2442.030 ;
        RECT 2932.210 2439.250 2933.390 2440.430 ;
        RECT 2932.210 2260.850 2933.390 2262.030 ;
        RECT 2932.210 2259.250 2933.390 2260.430 ;
        RECT 2932.210 2080.850 2933.390 2082.030 ;
        RECT 2932.210 2079.250 2933.390 2080.430 ;
        RECT 2932.210 1900.850 2933.390 1902.030 ;
        RECT 2932.210 1899.250 2933.390 1900.430 ;
        RECT 2932.210 1720.850 2933.390 1722.030 ;
        RECT 2932.210 1719.250 2933.390 1720.430 ;
        RECT 2932.210 1540.850 2933.390 1542.030 ;
        RECT 2932.210 1539.250 2933.390 1540.430 ;
        RECT 2932.210 1360.850 2933.390 1362.030 ;
        RECT 2932.210 1359.250 2933.390 1360.430 ;
        RECT 2932.210 1180.850 2933.390 1182.030 ;
        RECT 2932.210 1179.250 2933.390 1180.430 ;
        RECT 2932.210 1000.850 2933.390 1002.030 ;
        RECT 2932.210 999.250 2933.390 1000.430 ;
        RECT 2932.210 820.850 2933.390 822.030 ;
        RECT 2932.210 819.250 2933.390 820.430 ;
        RECT 2932.210 640.850 2933.390 642.030 ;
        RECT 2932.210 639.250 2933.390 640.430 ;
        RECT 2932.210 460.850 2933.390 462.030 ;
        RECT 2932.210 459.250 2933.390 460.430 ;
        RECT 2932.210 280.850 2933.390 282.030 ;
        RECT 2932.210 279.250 2933.390 280.430 ;
        RECT 2932.210 100.850 2933.390 102.030 ;
        RECT 2932.210 99.250 2933.390 100.430 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.140 -11.680 3342.150 ;
        RECT 2931.300 3342.140 2934.300 3342.150 ;
        RECT -14.680 3339.140 0.300 3342.140 ;
        RECT 2919.700 3339.140 2934.300 3342.140 ;
        RECT -14.680 3339.130 -11.680 3339.140 ;
        RECT 2931.300 3339.130 2934.300 3339.140 ;
        RECT -14.680 3162.140 -11.680 3162.150 ;
        RECT 2931.300 3162.140 2934.300 3162.150 ;
        RECT -14.680 3159.140 0.300 3162.140 ;
        RECT 2919.700 3159.140 2934.300 3162.140 ;
        RECT -14.680 3159.130 -11.680 3159.140 ;
        RECT 2931.300 3159.130 2934.300 3159.140 ;
        RECT -14.680 2982.140 -11.680 2982.150 ;
        RECT 2931.300 2982.140 2934.300 2982.150 ;
        RECT -14.680 2979.140 0.300 2982.140 ;
        RECT 2919.700 2979.140 2934.300 2982.140 ;
        RECT -14.680 2979.130 -11.680 2979.140 ;
        RECT 2931.300 2979.130 2934.300 2979.140 ;
        RECT -14.680 2802.140 -11.680 2802.150 ;
        RECT 2931.300 2802.140 2934.300 2802.150 ;
        RECT -14.680 2799.140 0.300 2802.140 ;
        RECT 2919.700 2799.140 2934.300 2802.140 ;
        RECT -14.680 2799.130 -11.680 2799.140 ;
        RECT 2931.300 2799.130 2934.300 2799.140 ;
        RECT -14.680 2622.140 -11.680 2622.150 ;
        RECT 2931.300 2622.140 2934.300 2622.150 ;
        RECT -14.680 2619.140 0.300 2622.140 ;
        RECT 2919.700 2619.140 2934.300 2622.140 ;
        RECT -14.680 2619.130 -11.680 2619.140 ;
        RECT 2931.300 2619.130 2934.300 2619.140 ;
        RECT -14.680 2442.140 -11.680 2442.150 ;
        RECT 2931.300 2442.140 2934.300 2442.150 ;
        RECT -14.680 2439.140 0.300 2442.140 ;
        RECT 2919.700 2439.140 2934.300 2442.140 ;
        RECT -14.680 2439.130 -11.680 2439.140 ;
        RECT 2931.300 2439.130 2934.300 2439.140 ;
        RECT -14.680 2262.140 -11.680 2262.150 ;
        RECT 2931.300 2262.140 2934.300 2262.150 ;
        RECT -14.680 2259.140 0.300 2262.140 ;
        RECT 2919.700 2259.140 2934.300 2262.140 ;
        RECT -14.680 2259.130 -11.680 2259.140 ;
        RECT 2931.300 2259.130 2934.300 2259.140 ;
        RECT -14.680 2082.140 -11.680 2082.150 ;
        RECT 2931.300 2082.140 2934.300 2082.150 ;
        RECT -14.680 2079.140 0.300 2082.140 ;
        RECT 2919.700 2079.140 2934.300 2082.140 ;
        RECT -14.680 2079.130 -11.680 2079.140 ;
        RECT 2931.300 2079.130 2934.300 2079.140 ;
        RECT -14.680 1902.140 -11.680 1902.150 ;
        RECT 2931.300 1902.140 2934.300 1902.150 ;
        RECT -14.680 1899.140 0.300 1902.140 ;
        RECT 2919.700 1899.140 2934.300 1902.140 ;
        RECT -14.680 1899.130 -11.680 1899.140 ;
        RECT 2931.300 1899.130 2934.300 1899.140 ;
        RECT -14.680 1722.140 -11.680 1722.150 ;
        RECT 2931.300 1722.140 2934.300 1722.150 ;
        RECT -14.680 1719.140 0.300 1722.140 ;
        RECT 2919.700 1719.140 2934.300 1722.140 ;
        RECT -14.680 1719.130 -11.680 1719.140 ;
        RECT 2931.300 1719.130 2934.300 1719.140 ;
        RECT -14.680 1542.140 -11.680 1542.150 ;
        RECT 2931.300 1542.140 2934.300 1542.150 ;
        RECT -14.680 1539.140 0.300 1542.140 ;
        RECT 2919.700 1539.140 2934.300 1542.140 ;
        RECT -14.680 1539.130 -11.680 1539.140 ;
        RECT 2931.300 1539.130 2934.300 1539.140 ;
        RECT -14.680 1362.140 -11.680 1362.150 ;
        RECT 2931.300 1362.140 2934.300 1362.150 ;
        RECT -14.680 1359.140 0.300 1362.140 ;
        RECT 2919.700 1359.140 2934.300 1362.140 ;
        RECT -14.680 1359.130 -11.680 1359.140 ;
        RECT 2931.300 1359.130 2934.300 1359.140 ;
        RECT -14.680 1182.140 -11.680 1182.150 ;
        RECT 2931.300 1182.140 2934.300 1182.150 ;
        RECT -14.680 1179.140 0.300 1182.140 ;
        RECT 2919.700 1179.140 2934.300 1182.140 ;
        RECT -14.680 1179.130 -11.680 1179.140 ;
        RECT 2931.300 1179.130 2934.300 1179.140 ;
        RECT -14.680 1002.140 -11.680 1002.150 ;
        RECT 2931.300 1002.140 2934.300 1002.150 ;
        RECT -14.680 999.140 0.300 1002.140 ;
        RECT 2919.700 999.140 2934.300 1002.140 ;
        RECT -14.680 999.130 -11.680 999.140 ;
        RECT 2931.300 999.130 2934.300 999.140 ;
        RECT -14.680 822.140 -11.680 822.150 ;
        RECT 2931.300 822.140 2934.300 822.150 ;
        RECT -14.680 819.140 0.300 822.140 ;
        RECT 2919.700 819.140 2934.300 822.140 ;
        RECT -14.680 819.130 -11.680 819.140 ;
        RECT 2931.300 819.130 2934.300 819.140 ;
        RECT -14.680 642.140 -11.680 642.150 ;
        RECT 2931.300 642.140 2934.300 642.150 ;
        RECT -14.680 639.140 0.300 642.140 ;
        RECT 2919.700 639.140 2934.300 642.140 ;
        RECT -14.680 639.130 -11.680 639.140 ;
        RECT 2931.300 639.130 2934.300 639.140 ;
        RECT -14.680 462.140 -11.680 462.150 ;
        RECT 2931.300 462.140 2934.300 462.150 ;
        RECT -14.680 459.140 0.300 462.140 ;
        RECT 2919.700 459.140 2934.300 462.140 ;
        RECT -14.680 459.130 -11.680 459.140 ;
        RECT 2931.300 459.130 2934.300 459.140 ;
        RECT -14.680 282.140 -11.680 282.150 ;
        RECT 2931.300 282.140 2934.300 282.150 ;
        RECT -14.680 279.140 0.300 282.140 ;
        RECT 2919.700 279.140 2934.300 282.140 ;
        RECT -14.680 279.130 -11.680 279.140 ;
        RECT 2931.300 279.130 2934.300 279.140 ;
        RECT -14.680 102.140 -11.680 102.150 ;
        RECT 2931.300 102.140 2934.300 102.150 ;
        RECT -14.680 99.140 0.300 102.140 ;
        RECT 2919.700 99.140 2934.300 102.140 ;
        RECT -14.680 99.130 -11.680 99.140 ;
        RECT 2931.300 99.130 2934.300 99.140 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 3519.700 25.020 3538.400 ;
        RECT 202.020 3519.700 205.020 3538.400 ;
        RECT 382.020 3519.700 385.020 3538.400 ;
        RECT 562.020 3519.700 565.020 3538.400 ;
        RECT 742.020 3519.700 745.020 3538.400 ;
        RECT 922.020 3519.700 925.020 3538.400 ;
        RECT 1102.020 3519.700 1105.020 3538.400 ;
        RECT 1282.020 3519.700 1285.020 3538.400 ;
        RECT 1462.020 3519.700 1465.020 3538.400 ;
        RECT 1642.020 3519.700 1645.020 3538.400 ;
        RECT 1822.020 3519.700 1825.020 3538.400 ;
        RECT 2002.020 3519.700 2005.020 3538.400 ;
        RECT 2182.020 3519.700 2185.020 3538.400 ;
        RECT 2362.020 3519.700 2365.020 3538.400 ;
        RECT 2542.020 3519.700 2545.020 3538.400 ;
        RECT 2722.020 3519.700 2725.020 3538.400 ;
        RECT 2902.020 3519.700 2905.020 3538.400 ;
        RECT 22.020 -18.720 25.020 0.300 ;
        RECT 202.020 -18.720 205.020 0.300 ;
        RECT 382.020 -18.720 385.020 0.300 ;
        RECT 562.020 -18.720 565.020 0.300 ;
        RECT 742.020 -18.720 745.020 0.300 ;
        RECT 922.020 -18.720 925.020 0.300 ;
        RECT 1102.020 -18.720 1105.020 0.300 ;
        RECT 1282.020 -18.720 1285.020 0.300 ;
        RECT 1462.020 -18.720 1465.020 0.300 ;
        RECT 1642.020 -18.720 1645.020 0.300 ;
        RECT 1822.020 -18.720 1825.020 0.300 ;
        RECT 2002.020 -18.720 2005.020 0.300 ;
        RECT 2182.020 -18.720 2185.020 0.300 ;
        RECT 2362.020 -18.720 2365.020 0.300 ;
        RECT 2542.020 -18.720 2545.020 0.300 ;
        RECT 2722.020 -18.720 2725.020 0.300 ;
        RECT 2902.020 -18.720 2905.020 0.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 0.300 3450.380 ;
        RECT 2919.700 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 0.300 3270.380 ;
        RECT 2919.700 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 0.300 3090.380 ;
        RECT 2919.700 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 0.300 2910.380 ;
        RECT 2919.700 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 0.300 2730.380 ;
        RECT 2919.700 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 0.300 2550.380 ;
        RECT 2919.700 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 0.300 2370.380 ;
        RECT 2919.700 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 0.300 2190.380 ;
        RECT 2919.700 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 0.300 2010.380 ;
        RECT 2919.700 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 0.300 1830.380 ;
        RECT 2919.700 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 0.300 1650.380 ;
        RECT 2919.700 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 0.300 1470.380 ;
        RECT 2919.700 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 0.300 1290.380 ;
        RECT 2919.700 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 0.300 1110.380 ;
        RECT 2919.700 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 0.300 930.380 ;
        RECT 2919.700 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 0.300 750.380 ;
        RECT 2919.700 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 0.300 570.380 ;
        RECT 2919.700 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 0.300 390.380 ;
        RECT 2919.700 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 0.300 210.380 ;
        RECT 2919.700 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 0.300 30.380 ;
        RECT 2919.700 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 3519.700 115.020 3538.400 ;
        RECT 292.020 3519.700 295.020 3538.400 ;
        RECT 472.020 3519.700 475.020 3538.400 ;
        RECT 652.020 3519.700 655.020 3538.400 ;
        RECT 832.020 3519.700 835.020 3538.400 ;
        RECT 1012.020 3519.700 1015.020 3538.400 ;
        RECT 1192.020 3519.700 1195.020 3538.400 ;
        RECT 1372.020 3519.700 1375.020 3538.400 ;
        RECT 1552.020 3519.700 1555.020 3538.400 ;
        RECT 1732.020 3519.700 1735.020 3538.400 ;
        RECT 1912.020 3519.700 1915.020 3538.400 ;
        RECT 2092.020 3519.700 2095.020 3538.400 ;
        RECT 2272.020 3519.700 2275.020 3538.400 ;
        RECT 2452.020 3519.700 2455.020 3538.400 ;
        RECT 2632.020 3519.700 2635.020 3538.400 ;
        RECT 2812.020 3519.700 2815.020 3538.400 ;
        RECT 112.020 -18.720 115.020 0.300 ;
        RECT 292.020 -18.720 295.020 0.300 ;
        RECT 472.020 -18.720 475.020 0.300 ;
        RECT 652.020 -18.720 655.020 0.300 ;
        RECT 832.020 -18.720 835.020 0.300 ;
        RECT 1012.020 -18.720 1015.020 0.300 ;
        RECT 1192.020 -18.720 1195.020 0.300 ;
        RECT 1372.020 -18.720 1375.020 0.300 ;
        RECT 1552.020 -18.720 1555.020 0.300 ;
        RECT 1732.020 -18.720 1735.020 0.300 ;
        RECT 1912.020 -18.720 1915.020 0.300 ;
        RECT 2092.020 -18.720 2095.020 0.300 ;
        RECT 2272.020 -18.720 2275.020 0.300 ;
        RECT 2452.020 -18.720 2455.020 0.300 ;
        RECT 2632.020 -18.720 2635.020 0.300 ;
        RECT 2812.020 -18.720 2815.020 0.300 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 0.300 3360.380 ;
        RECT 2919.700 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 0.300 3180.380 ;
        RECT 2919.700 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 0.300 3000.380 ;
        RECT 2919.700 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 0.300 2820.380 ;
        RECT 2919.700 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 0.300 2640.380 ;
        RECT 2919.700 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 0.300 2460.380 ;
        RECT 2919.700 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 0.300 2280.380 ;
        RECT 2919.700 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 0.300 2100.380 ;
        RECT 2919.700 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 0.300 1920.380 ;
        RECT 2919.700 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 0.300 1740.380 ;
        RECT 2919.700 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 0.300 1560.380 ;
        RECT 2919.700 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 0.300 1380.380 ;
        RECT 2919.700 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 0.300 1200.380 ;
        RECT 2919.700 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 0.300 1020.380 ;
        RECT 2919.700 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 0.300 840.380 ;
        RECT 2919.700 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 0.300 660.380 ;
        RECT 2919.700 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 0.300 480.380 ;
        RECT 2919.700 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 0.300 300.380 ;
        RECT 2919.700 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 0.300 120.380 ;
        RECT 2919.700 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 3519.700 43.020 3547.800 ;
        RECT 220.020 3519.700 223.020 3547.800 ;
        RECT 400.020 3519.700 403.020 3547.800 ;
        RECT 580.020 3519.700 583.020 3547.800 ;
        RECT 760.020 3519.700 763.020 3547.800 ;
        RECT 940.020 3519.700 943.020 3547.800 ;
        RECT 1120.020 3519.700 1123.020 3547.800 ;
        RECT 1300.020 3519.700 1303.020 3547.800 ;
        RECT 1480.020 3519.700 1483.020 3547.800 ;
        RECT 1660.020 3519.700 1663.020 3547.800 ;
        RECT 1840.020 3519.700 1843.020 3547.800 ;
        RECT 2020.020 3519.700 2023.020 3547.800 ;
        RECT 2200.020 3519.700 2203.020 3547.800 ;
        RECT 2380.020 3519.700 2383.020 3547.800 ;
        RECT 2560.020 3519.700 2563.020 3547.800 ;
        RECT 2740.020 3519.700 2743.020 3547.800 ;
        RECT 40.020 -28.120 43.020 0.300 ;
        RECT 220.020 -28.120 223.020 0.300 ;
        RECT 400.020 -28.120 403.020 0.300 ;
        RECT 580.020 -28.120 583.020 0.300 ;
        RECT 760.020 -28.120 763.020 0.300 ;
        RECT 940.020 -28.120 943.020 0.300 ;
        RECT 1120.020 -28.120 1123.020 0.300 ;
        RECT 1300.020 -28.120 1303.020 0.300 ;
        RECT 1480.020 -28.120 1483.020 0.300 ;
        RECT 1660.020 -28.120 1663.020 0.300 ;
        RECT 1840.020 -28.120 1843.020 0.300 ;
        RECT 2020.020 -28.120 2023.020 0.300 ;
        RECT 2200.020 -28.120 2203.020 0.300 ;
        RECT 2380.020 -28.120 2383.020 0.300 ;
        RECT 2560.020 -28.120 2563.020 0.300 ;
        RECT 2740.020 -28.120 2743.020 0.300 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 0.300 3468.380 ;
        RECT 2919.700 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 0.300 3288.380 ;
        RECT 2919.700 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 0.300 3108.380 ;
        RECT 2919.700 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 0.300 2928.380 ;
        RECT 2919.700 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 0.300 2748.380 ;
        RECT 2919.700 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 0.300 2568.380 ;
        RECT 2919.700 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 0.300 2388.380 ;
        RECT 2919.700 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 0.300 2208.380 ;
        RECT 2919.700 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 0.300 2028.380 ;
        RECT 2919.700 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 0.300 1848.380 ;
        RECT 2919.700 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 0.300 1668.380 ;
        RECT 2919.700 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 0.300 1488.380 ;
        RECT 2919.700 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 0.300 1308.380 ;
        RECT 2919.700 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 0.300 1128.380 ;
        RECT 2919.700 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 0.300 948.380 ;
        RECT 2919.700 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 0.300 768.380 ;
        RECT 2919.700 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 0.300 588.380 ;
        RECT 2919.700 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 0.300 408.380 ;
        RECT 2919.700 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 0.300 228.380 ;
        RECT 2919.700 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 0.300 48.380 ;
        RECT 2919.700 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 3519.700 133.020 3547.800 ;
        RECT 310.020 3519.700 313.020 3547.800 ;
        RECT 490.020 3519.700 493.020 3547.800 ;
        RECT 670.020 3519.700 673.020 3547.800 ;
        RECT 850.020 3519.700 853.020 3547.800 ;
        RECT 1030.020 3519.700 1033.020 3547.800 ;
        RECT 1210.020 3519.700 1213.020 3547.800 ;
        RECT 1390.020 3519.700 1393.020 3547.800 ;
        RECT 1570.020 3519.700 1573.020 3547.800 ;
        RECT 1750.020 3519.700 1753.020 3547.800 ;
        RECT 1930.020 3519.700 1933.020 3547.800 ;
        RECT 2110.020 3519.700 2113.020 3547.800 ;
        RECT 2290.020 3519.700 2293.020 3547.800 ;
        RECT 2470.020 3519.700 2473.020 3547.800 ;
        RECT 2650.020 3519.700 2653.020 3547.800 ;
        RECT 2830.020 3519.700 2833.020 3547.800 ;
        RECT 130.020 -28.120 133.020 0.300 ;
        RECT 310.020 -28.120 313.020 0.300 ;
        RECT 490.020 -28.120 493.020 0.300 ;
        RECT 670.020 -28.120 673.020 0.300 ;
        RECT 850.020 -28.120 853.020 0.300 ;
        RECT 1030.020 -28.120 1033.020 0.300 ;
        RECT 1210.020 -28.120 1213.020 0.300 ;
        RECT 1390.020 -28.120 1393.020 0.300 ;
        RECT 1570.020 -28.120 1573.020 0.300 ;
        RECT 1750.020 -28.120 1753.020 0.300 ;
        RECT 1930.020 -28.120 1933.020 0.300 ;
        RECT 2110.020 -28.120 2113.020 0.300 ;
        RECT 2290.020 -28.120 2293.020 0.300 ;
        RECT 2470.020 -28.120 2473.020 0.300 ;
        RECT 2650.020 -28.120 2653.020 0.300 ;
        RECT 2830.020 -28.120 2833.020 0.300 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 0.300 3378.380 ;
        RECT 2919.700 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 0.300 3198.380 ;
        RECT 2919.700 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 0.300 3018.380 ;
        RECT 2919.700 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 0.300 2838.380 ;
        RECT 2919.700 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 0.300 2658.380 ;
        RECT 2919.700 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 0.300 2478.380 ;
        RECT 2919.700 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 0.300 2298.380 ;
        RECT 2919.700 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 0.300 2118.380 ;
        RECT 2919.700 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 0.300 1938.380 ;
        RECT 2919.700 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 0.300 1758.380 ;
        RECT 2919.700 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 0.300 1578.380 ;
        RECT 2919.700 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 0.300 1398.380 ;
        RECT 2919.700 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 0.300 1218.380 ;
        RECT 2919.700 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 0.300 1038.380 ;
        RECT 2919.700 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 0.300 858.380 ;
        RECT 2919.700 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 0.300 678.380 ;
        RECT 2919.700 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 0.300 498.380 ;
        RECT 2919.700 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 0.300 318.380 ;
        RECT 2919.700 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 0.300 138.380 ;
        RECT 2919.700 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 3519.700 61.020 3557.200 ;
        RECT 238.020 3519.700 241.020 3557.200 ;
        RECT 418.020 3519.700 421.020 3557.200 ;
        RECT 598.020 3519.700 601.020 3557.200 ;
        RECT 778.020 3519.700 781.020 3557.200 ;
        RECT 958.020 3519.700 961.020 3557.200 ;
        RECT 1138.020 3519.700 1141.020 3557.200 ;
        RECT 1318.020 3519.700 1321.020 3557.200 ;
        RECT 1498.020 3519.700 1501.020 3557.200 ;
        RECT 1678.020 3519.700 1681.020 3557.200 ;
        RECT 1858.020 3519.700 1861.020 3557.200 ;
        RECT 2038.020 3519.700 2041.020 3557.200 ;
        RECT 2218.020 3519.700 2221.020 3557.200 ;
        RECT 2398.020 3519.700 2401.020 3557.200 ;
        RECT 2578.020 3519.700 2581.020 3557.200 ;
        RECT 2758.020 3519.700 2761.020 3557.200 ;
        RECT 58.020 -37.520 61.020 0.300 ;
        RECT 238.020 -37.520 241.020 0.300 ;
        RECT 418.020 -37.520 421.020 0.300 ;
        RECT 598.020 -37.520 601.020 0.300 ;
        RECT 778.020 -37.520 781.020 0.300 ;
        RECT 958.020 -37.520 961.020 0.300 ;
        RECT 1138.020 -37.520 1141.020 0.300 ;
        RECT 1318.020 -37.520 1321.020 0.300 ;
        RECT 1498.020 -37.520 1501.020 0.300 ;
        RECT 1678.020 -37.520 1681.020 0.300 ;
        RECT 1858.020 -37.520 1861.020 0.300 ;
        RECT 2038.020 -37.520 2041.020 0.300 ;
        RECT 2218.020 -37.520 2221.020 0.300 ;
        RECT 2398.020 -37.520 2401.020 0.300 ;
        RECT 2578.020 -37.520 2581.020 0.300 ;
        RECT 2758.020 -37.520 2761.020 0.300 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 0.300 3486.380 ;
        RECT 2919.700 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 0.300 3306.380 ;
        RECT 2919.700 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 0.300 3126.380 ;
        RECT 2919.700 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 0.300 2946.380 ;
        RECT 2919.700 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 0.300 2766.380 ;
        RECT 2919.700 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 0.300 2586.380 ;
        RECT 2919.700 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 0.300 2406.380 ;
        RECT 2919.700 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 0.300 2226.380 ;
        RECT 2919.700 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 0.300 2046.380 ;
        RECT 2919.700 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 0.300 1866.380 ;
        RECT 2919.700 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 0.300 1686.380 ;
        RECT 2919.700 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 0.300 1506.380 ;
        RECT 2919.700 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 0.300 1326.380 ;
        RECT 2919.700 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 0.300 1146.380 ;
        RECT 2919.700 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 0.300 966.380 ;
        RECT 2919.700 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 0.300 786.380 ;
        RECT 2919.700 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 0.300 606.380 ;
        RECT 2919.700 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 0.300 426.380 ;
        RECT 2919.700 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 0.300 246.380 ;
        RECT 2919.700 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 0.300 66.380 ;
        RECT 2919.700 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 3519.700 151.020 3557.200 ;
        RECT 328.020 3519.700 331.020 3557.200 ;
        RECT 508.020 3519.700 511.020 3557.200 ;
        RECT 688.020 3519.700 691.020 3557.200 ;
        RECT 868.020 3519.700 871.020 3557.200 ;
        RECT 1048.020 3519.700 1051.020 3557.200 ;
        RECT 1228.020 3519.700 1231.020 3557.200 ;
        RECT 1408.020 3519.700 1411.020 3557.200 ;
        RECT 1588.020 3519.700 1591.020 3557.200 ;
        RECT 1768.020 3519.700 1771.020 3557.200 ;
        RECT 1948.020 3519.700 1951.020 3557.200 ;
        RECT 2128.020 3519.700 2131.020 3557.200 ;
        RECT 2308.020 3519.700 2311.020 3557.200 ;
        RECT 2488.020 3519.700 2491.020 3557.200 ;
        RECT 2668.020 3519.700 2671.020 3557.200 ;
        RECT 2848.020 3519.700 2851.020 3557.200 ;
        RECT 148.020 -37.520 151.020 0.300 ;
        RECT 328.020 -37.520 331.020 0.300 ;
        RECT 508.020 -37.520 511.020 0.300 ;
        RECT 688.020 -37.520 691.020 0.300 ;
        RECT 868.020 -37.520 871.020 0.300 ;
        RECT 1048.020 -37.520 1051.020 0.300 ;
        RECT 1228.020 -37.520 1231.020 0.300 ;
        RECT 1408.020 -37.520 1411.020 0.300 ;
        RECT 1588.020 -37.520 1591.020 0.300 ;
        RECT 1768.020 -37.520 1771.020 0.300 ;
        RECT 1948.020 -37.520 1951.020 0.300 ;
        RECT 2128.020 -37.520 2131.020 0.300 ;
        RECT 2308.020 -37.520 2311.020 0.300 ;
        RECT 2488.020 -37.520 2491.020 0.300 ;
        RECT 2668.020 -37.520 2671.020 0.300 ;
        RECT 2848.020 -37.520 2851.020 0.300 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 0.300 3396.380 ;
        RECT 2919.700 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 0.300 3216.380 ;
        RECT 2919.700 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 0.300 3036.380 ;
        RECT 2919.700 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 0.300 2856.380 ;
        RECT 2919.700 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 0.300 2676.380 ;
        RECT 2919.700 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 0.300 2496.380 ;
        RECT 2919.700 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 0.300 2316.380 ;
        RECT 2919.700 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 0.300 2136.380 ;
        RECT 2919.700 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 0.300 1956.380 ;
        RECT 2919.700 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 0.300 1776.380 ;
        RECT 2919.700 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 0.300 1596.380 ;
        RECT 2919.700 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 0.300 1416.380 ;
        RECT 2919.700 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 0.300 1236.380 ;
        RECT 2919.700 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 0.300 1056.380 ;
        RECT 2919.700 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 0.300 876.380 ;
        RECT 2919.700 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 0.300 696.380 ;
        RECT 2919.700 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 0.300 516.380 ;
        RECT 2919.700 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 0.300 336.380 ;
        RECT 2919.700 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 0.300 156.380 ;
        RECT 2919.700 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 276.145 2.805 2799.415 3477.435 ;
      LAYER met1 ;
        RECT 2.830 2.760 2914.100 3512.160 ;
      LAYER met2 ;
        RECT 2.710 0.300 2917.370 3519.700 ;
      LAYER met3 ;
        RECT 0.300 10.715 2919.700 3508.965 ;
      LAYER met4 ;
        RECT 4.020 0.300 2905.020 3519.700 ;
      LAYER met5 ;
        RECT 0.300 9.130 2919.700 3486.390 ;
>>>>>>> f48448d4736bd6d56fed4dbf7f9cc50552d8745d
  END
END user_project_wrapper
END LIBRARY

